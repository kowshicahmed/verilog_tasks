* NGSPICE file created from program_counter.ext - technology: scmos

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

.subckt program_counter gnd vdd clock opcode[1] opcode[0] pc_in[15] pc_in[14] pc_in[13]
+ pc_in[12] pc_in[11] pc_in[10] pc_in[9] pc_in[8] pc_in[7] pc_in[6] pc_in[5] pc_in[4]
+ pc_in[3] pc_in[2] pc_in[1] pc_in[0] pc_out[15] pc_out[14] pc_out[13] pc_out[12]
+ pc_out[11] pc_out[10] pc_out[9] pc_out[8] pc_out[7] pc_out[6] pc_out[5] pc_out[4]
+ pc_out[3] pc_out[2] pc_out[1] pc_out[0]
X_200_ pc_in[7] _211_/A _214_/C _200_/D gnd _200_/Y vdd AOI22X1
XSFILL7280x2100 gnd vdd FILL
X_131_ _191_/A _131_/B gnd _132_/C vdd NAND2X1
X_277_ _277_/Q _262_/CLK _120_/Y gnd vdd DFFPOSX1
XSFILL17680x10100 gnd vdd FILL
X_114_ _162_/B _134_/B _114_/C gnd _275_/D vdd OAI21X1
XSFILL6320x6100 gnd vdd FILL
X_276_ _276_/Q _284_/CLK _117_/Y gnd vdd DFFPOSX1
X_130_ pc_in[6] gnd _132_/A vdd INVX1
XSFILL18320x100 gnd vdd FILL
XSFILL17360x6100 gnd vdd FILL
X_113_ _162_/C _134_/B gnd _114_/C vdd NAND2X1
X_259_ _243_/A _288_/CLK _259_/D gnd vdd DFFPOSX1
XSFILL7120x2100 gnd vdd FILL
X_258_ _258_/A gnd pc_out[15] vdd BUFX2
X_275_ _162_/C _288_/CLK _275_/D gnd vdd DFFPOSX1
X_189_ pc_in[5] _211_/A _112_/A _188_/Y gnd _189_/Y vdd AOI22X1
XSFILL17840x100 gnd vdd FILL
XSFILL17200x6100 gnd vdd FILL
X_112_ _112_/A _211_/A gnd _112_/Y vdd NOR2X1
XSFILL18160x2100 gnd vdd FILL
X_274_ _258_/A _274_/CLK _242_/Y gnd vdd DFFPOSX1
XSFILL18320x12100 gnd vdd FILL
X_257_ _257_/A gnd pc_out[14] vdd BUFX2
X_111_ opcode[1] _111_/B gnd _211_/A vdd NOR2X1
X_188_ pc_in[5] _186_/Y gnd _188_/Y vdd NAND2X1
XSFILL18000x2100 gnd vdd FILL
X_290_ _158_/A _274_/CLK _290_/D gnd vdd DFFPOSX1
XSFILL16880x6100 gnd vdd FILL
X_256_ _256_/A gnd pc_out[13] vdd BUFX2
XFILL22480x4100 gnd vdd FILL
X_273_ _257_/A _274_/CLK _273_/D gnd vdd DFFPOSX1
X_187_ pc_in[5] _186_/Y gnd _190_/A vdd NOR2X1
X_110_ opcode[0] gnd _111_/B vdd INVX1
X_239_ _238_/A _235_/B gnd _239_/Y vdd NAND2X1
X_272_ _256_/A _274_/CLK _272_/D gnd vdd DFFPOSX1
XSFILL17680x2100 gnd vdd FILL
X_255_ _255_/A gnd pc_out[12] vdd BUFX2
XBUFX2_insert5 _112_/Y gnd _125_/B vdd BUFX2
X_186_ _121_/Y _181_/A _171_/Y gnd _186_/Y vdd NOR3X1
XSFILL7280x10100 gnd vdd FILL
XSFILL6640x8100 gnd vdd FILL
X_169_ _277_/Q _211_/D gnd _169_/Y vdd NAND2X1
X_238_ _238_/A _235_/B gnd _238_/Y vdd NOR2X1
XSFILL6800x12100 gnd vdd FILL
X_254_ _254_/A gnd pc_out[11] vdd BUFX2
X_271_ _255_/A _274_/CLK _228_/Y gnd vdd DFFPOSX1
X_185_ _128_/A _211_/D gnd _185_/Y vdd NAND2X1
XSFILL17680x8100 gnd vdd FILL
XBUFX2_insert6 _112_/Y gnd _117_/B vdd BUFX2
X_237_ _237_/A _237_/B _237_/C gnd _273_/D vdd OAI21X1
X_168_ _168_/A _168_/B _168_/C gnd _168_/Y vdd OAI21X1
X_270_ _254_/A _265_/CLK _221_/Y gnd vdd DFFPOSX1
XSFILL6160x8100 gnd vdd FILL
X_253_ _269_/Q gnd pc_out[10] vdd BUFX2
XSFILL17520x10100 gnd vdd FILL
X_184_ _184_/A _183_/Y gnd _263_/D vdd NAND2X1
XBUFX2_insert7 _112_/Y gnd _147_/B vdd BUFX2
X_219_ _218_/B _217_/Y _219_/C gnd _219_/Y vdd OAI21X1
X_167_ _167_/A _166_/Y pc_in[1] _211_/A gnd _168_/B vdd AOI22X1
X_236_ _211_/A pc_in[14] _289_/Q _211_/D gnd _237_/C vdd AOI22X1
XSFILL17520x8100 gnd vdd FILL
X_252_ _268_/Q gnd pc_out[9] vdd BUFX2
X_166_ pc_in[0] pc_in[1] gnd _166_/Y vdd NAND2X1
X_235_ _219_/C _235_/B gnd _237_/B vdd NAND2X1
X_183_ pc_in[4] _176_/Y _183_/C gnd _183_/Y vdd OAI21X1
XBUFX2_insert8 _112_/Y gnd _131_/B vdd BUFX2
XCLKBUF1_insert0 clock gnd _284_/CLK vdd CLKBUF1
X_218_ _217_/Y _218_/B gnd _221_/A vdd AND2X2
X_149_ _287_/Q _147_/B gnd _149_/Y vdd NAND2X1
X_251_ _267_/Q gnd pc_out[8] vdd BUFX2
XBUFX2_insert9 _112_/Y gnd _134_/B vdd BUFX2
X_182_ _181_/A _204_/B _182_/C gnd _183_/C vdd OAI21X1
XCLKBUF1_insert1 clock gnd _274_/CLK vdd CLKBUF1
X_165_ pc_in[0] pc_in[1] gnd _168_/A vdd NOR2X1
X_217_ pc_in[9] pc_in[10] _208_/B gnd _217_/Y vdd NAND3X1
X_234_ pc_in[13] pc_in[14] _225_/A gnd _235_/B vdd NAND3X1
X_148_ pc_in[12] gnd _224_/B vdd INVX1
X_250_ _266_/Q gnd pc_out[7] vdd BUFX2
X_164_ _276_/Q _211_/D gnd _168_/C vdd NAND2X1
X_233_ _225_/A pc_in[13] pc_in[14] gnd _237_/A vdd AOI21X1
X_181_ _181_/A _178_/D _167_/A gnd _182_/C vdd OAI21X1
X_216_ _213_/Y _214_/Y _215_/Y gnd _216_/Y vdd OAI21X1
XCLKBUF1_insert2 clock gnd _265_/CLK vdd CLKBUF1
X_147_ _218_/B _147_/B _146_/Y gnd _286_/D vdd OAI21X1
XSFILL6480x4100 gnd vdd FILL
XSFILL6800x4100 gnd vdd FILL
XSFILL6960x10100 gnd vdd FILL
XSFILL6000x100 gnd vdd FILL
X_180_ _125_/A _211_/D gnd _184_/A vdd NAND2X1
XSFILL18160x12100 gnd vdd FILL
X_163_ _162_/B _204_/B _163_/C gnd _259_/D vdd OAI21X1
X_232_ _229_/Y _230_/Y _232_/C gnd _272_/D vdd OAI21X1
XSFILL17840x4100 gnd vdd FILL
X_215_ _211_/A pc_in[10] _215_/C _211_/D gnd _215_/Y vdd AOI22X1
X_146_ _220_/C _147_/B gnd _146_/Y vdd NAND2X1
XCLKBUF1_insert3 clock gnd _262_/CLK vdd CLKBUF1
X_129_ _129_/A _125_/B _128_/Y gnd _280_/D vdd OAI21X1
XSFILL6320x4100 gnd vdd FILL
XSFILL7120x10100 gnd vdd FILL
X_162_ _112_/A _162_/B _162_/C _211_/D gnd _163_/C vdd AOI22X1
X_231_ _211_/A pc_in[13] _288_/Q _211_/D gnd _232_/C vdd AOI22X1
X_214_ _142_/Y _214_/B _214_/C gnd _214_/Y vdd OAI21X1
X_145_ pc_in[11] gnd _218_/B vdd INVX2
XCLKBUF1_insert4 clock gnd _288_/CLK vdd CLKBUF1
X_128_ _128_/A _125_/B gnd _128_/Y vdd NAND2X1
X_230_ _153_/A _230_/B _219_/C gnd _230_/Y vdd OAI21X1
X_161_ _108_/Y _111_/B gnd _211_/D vdd NOR2X1
X_213_ _208_/B pc_in[9] pc_in[10] gnd _213_/Y vdd AOI21X1
X_144_ _142_/Y _117_/B _144_/C gnd _144_/Y vdd OAI21X1
X_127_ pc_in[5] gnd _129_/A vdd INVX1
XSFILL6640x12100 gnd vdd FILL
X_212_ _208_/Y _210_/Y _211_/Y gnd _212_/Y vdd OAI21X1
X_143_ _215_/C _117_/B gnd _144_/C vdd NAND2X1
XBUFX2_insert10 _109_/Y gnd _219_/C vdd BUFX2
X_289_ _289_/Q _288_/CLK _156_/Y gnd vdd DFFPOSX1
X_160_ _211_/A gnd _204_/B vdd INVX1
X_126_ _181_/A _125_/B _126_/C gnd _126_/Y vdd OAI21X1
XSFILL17360x10100 gnd vdd FILL
X_109_ opcode[0] _108_/Y gnd _109_/Y vdd NOR2X1
X_288_ _288_/Q _288_/CLK _153_/Y gnd vdd DFFPOSX1
XBUFX2_insert11 _109_/Y gnd _167_/A vdd BUFX2
XSFILL6160x100 gnd vdd FILL
X_125_ _125_/A _125_/B gnd _126_/C vdd NAND2X1
X_211_ _211_/A pc_in[9] _140_/A _211_/D gnd _211_/Y vdd AOI22X1
X_142_ pc_in[10] gnd _142_/Y vdd INVX1
X_108_ opcode[1] gnd _108_/Y vdd INVX1
X_210_ _214_/C _214_/B gnd _210_/Y vdd NAND2X1
X_141_ _141_/A _117_/B _141_/C gnd _141_/Y vdd OAI21X1
XBUFX2_insert12 _109_/Y gnd _112_/A vdd BUFX2
X_287_ _287_/Q _274_/CLK _150_/Y gnd vdd DFFPOSX1
X_124_ pc_in[4] gnd _181_/A vdd INVX2
XFILL22480x8100 gnd vdd FILL
XSFILL6640x6100 gnd vdd FILL
X_107_ pc_in[0] gnd _162_/B vdd INVX1
XBUFX2_insert13 _109_/Y gnd _214_/C vdd BUFX2
X_286_ _220_/C _274_/CLK _286_/D gnd vdd DFFPOSX1
X_269_ _269_/Q _284_/CLK _216_/Y gnd vdd DFFPOSX1
X_140_ _140_/A _117_/B gnd _141_/C vdd NAND2X1
XSFILL18000x12100 gnd vdd FILL
XSFILL6800x10100 gnd vdd FILL
X_123_ _121_/Y _125_/B _123_/C gnd _123_/Y vdd OAI21X1
X_285_ _215_/C _284_/CLK _144_/Y gnd vdd DFFPOSX1
XSFILL6160x6100 gnd vdd FILL
X_268_ _268_/Q _284_/CLK _212_/Y gnd vdd DFFPOSX1
X_199_ _199_/A gnd _200_/D vdd INVX1
X_122_ _174_/A _117_/B gnd _123_/C vdd NAND2X1
X_284_ _140_/A _284_/CLK _141_/Y gnd vdd DFFPOSX1
X_267_ _267_/Q _265_/CLK _267_/D gnd vdd DFFPOSX1
X_198_ _133_/Y _197_/A gnd _199_/A vdd NOR2X1
X_121_ pc_in[3] gnd _121_/Y vdd INVX2
X_283_ _137_/A _265_/CLK _283_/D gnd vdd DFFPOSX1
XSFILL17040x6100 gnd vdd FILL
X_266_ _266_/Q _265_/CLK _201_/Y gnd vdd DFFPOSX1
X_249_ _249_/A gnd pc_out[6] vdd BUFX2
X_197_ _197_/A _133_/Y gnd _197_/Y vdd AND2X2
X_120_ _120_/A _125_/B _120_/C gnd _120_/Y vdd OAI21X1
XSFILL6960x2100 gnd vdd FILL
XSFILL6320x100 gnd vdd FILL
X_265_ _249_/A _265_/CLK _195_/Y gnd vdd DFFPOSX1
X_282_ _282_/Q _265_/CLK _135_/Y gnd vdd DFFPOSX1
X_196_ _282_/Q _211_/D gnd _196_/Y vdd NAND2X1
XSFILL17200x10100 gnd vdd FILL
X_179_ _175_/Y _178_/Y _174_/Y gnd _179_/Y vdd OAI21X1
X_248_ _248_/A gnd pc_out[5] vdd BUFX2
XSFILL6800x2100 gnd vdd FILL
XSFILL6480x12100 gnd vdd FILL
X_281_ _191_/A _288_/CLK _281_/D gnd vdd DFFPOSX1
X_195_ _195_/A _194_/Y _191_/Y gnd _195_/Y vdd OAI21X1
X_247_ _247_/A gnd pc_out[4] vdd BUFX2
X_264_ _248_/A _262_/CLK _190_/Y gnd vdd DFFPOSX1
X_178_ pc_in[3] _211_/A _167_/A _178_/D gnd _178_/Y vdd AOI22X1
XSFILL17840x2100 gnd vdd FILL
XSFILL6480x8100 gnd vdd FILL
X_194_ pc_in[6] _211_/A _112_/A _197_/A gnd _194_/Y vdd AOI22X1
X_280_ _128_/A _288_/CLK _280_/D gnd vdd DFFPOSX1
X_263_ _247_/A _262_/CLK _263_/D gnd vdd DFFPOSX1
X_246_ _262_/Q gnd pc_out[3] vdd BUFX2
X_177_ _176_/Y gnd _178_/D vdd INVX1
X_229_ pc_in[13] _225_/A gnd _229_/Y vdd NOR2X1
XSFILL17840x8100 gnd vdd FILL
X_262_ _262_/Q _262_/CLK _179_/Y gnd vdd DFFPOSX1
X_193_ pc_in[5] pc_in[6] _186_/Y gnd _197_/A vdd NAND3X1
X_245_ _261_/Q gnd pc_out[2] vdd BUFX2
XSFILL6320x8100 gnd vdd FILL
X_228_ _228_/A _228_/B _227_/Y gnd _228_/Y vdd OAI21X1
X_159_ _238_/A _131_/B _158_/Y gnd _290_/D vdd OAI21X1
X_176_ _121_/Y _171_/Y gnd _176_/Y vdd NOR2X1
XSFILL6480x100 gnd vdd FILL
X_261_ _261_/Q _284_/CLK _173_/Y gnd vdd DFFPOSX1
X_192_ _186_/Y pc_in[5] pc_in[6] gnd _195_/A vdd AOI21X1
X_244_ _260_/Q gnd pc_out[1] vdd BUFX2
XSFILL17360x8100 gnd vdd FILL
X_175_ _171_/Y _121_/Y gnd _175_/Y vdd AND2X2
X_158_ _158_/A _131_/B gnd _158_/Y vdd NAND2X1
X_227_ _211_/A pc_in[12] _287_/Q _211_/D gnd _227_/Y vdd AOI22X1
X_260_ _260_/Q _284_/CLK _168_/Y gnd vdd DFFPOSX1
X_191_ _191_/A _211_/D gnd _191_/Y vdd NAND2X1
X_174_ _174_/A _211_/D gnd _174_/Y vdd NAND2X1
X_226_ _219_/C _230_/B gnd _228_/B vdd NAND2X1
X_157_ pc_in[15] gnd _238_/A vdd INVX1
X_243_ _243_/A gnd pc_out[0] vdd BUFX2
X_209_ pc_in[9] _208_/B gnd _214_/B vdd NAND2X1
XSFILL18000x100 gnd vdd FILL
X_173_ _173_/A _172_/Y _169_/Y gnd _173_/Y vdd OAI21X1
X_190_ _190_/A _189_/Y _185_/Y gnd _190_/Y vdd OAI21X1
X_242_ _238_/Y _240_/Y _241_/Y gnd _242_/Y vdd OAI21X1
X_225_ _225_/A gnd _230_/B vdd INVX1
XSFILL18000x4100 gnd vdd FILL
X_156_ _154_/Y _131_/B _156_/C gnd _156_/Y vdd OAI21X1
X_208_ pc_in[9] _208_/B gnd _208_/Y vdd NOR2X1
X_139_ pc_in[9] gnd _141_/A vdd INVX1
XFILL22480x6100 gnd vdd FILL
XSFILL6640x4100 gnd vdd FILL
X_224_ _218_/B _224_/B _217_/Y gnd _225_/A vdd NOR3X1
X_172_ _167_/A _171_/Y pc_in[2] _211_/A gnd _172_/Y vdd AOI22X1
X_241_ _211_/A pc_in[15] _158_/A _211_/D gnd _241_/Y vdd AOI22X1
X_155_ _289_/Q _131_/B gnd _156_/C vdd NAND2X1
XSFILL6320x12100 gnd vdd FILL
XFILL22480x10100 gnd vdd FILL
X_207_ _133_/Y _203_/A _197_/A gnd _208_/B vdd NOR3X1
X_138_ _203_/A _134_/B _137_/Y gnd _283_/D vdd OAI21X1
XSFILL17680x4100 gnd vdd FILL
X_171_ pc_in[0] pc_in[1] pc_in[2] gnd _171_/Y vdd NAND3X1
X_240_ _219_/C _239_/Y gnd _240_/Y vdd NAND2X1
X_223_ _223_/A gnd _228_/A vdd INVX1
X_154_ pc_in[14] gnd _154_/Y vdd INVX1
X_206_ _202_/Y _206_/B gnd _267_/D vdd NAND2X1
X_137_ _137_/A _134_/B gnd _137_/Y vdd NAND2X1
X_170_ pc_in[0] pc_in[1] pc_in[2] gnd _173_/A vdd AOI21X1
XSFILL17520x4100 gnd vdd FILL
X_205_ pc_in[8] _199_/A _205_/C gnd _206_/B vdd OAI21X1
X_136_ pc_in[8] gnd _203_/A vdd INVX2
X_153_ _153_/A _147_/B _153_/C gnd _153_/Y vdd OAI21X1
X_222_ _218_/B _217_/Y _224_/B gnd _223_/A vdd OAI21X1
XSFILL18160x100 gnd vdd FILL
X_119_ _277_/Q _125_/B gnd _120_/C vdd NAND2X1
X_221_ _221_/A _219_/Y _220_/Y gnd _221_/Y vdd OAI21X1
X_152_ _288_/Q _147_/B gnd _153_/C vdd NAND2X1
X_204_ _203_/A _204_/B _204_/C gnd _205_/C vdd OAI21X1
X_135_ _133_/Y _134_/B _135_/C gnd _135_/Y vdd OAI21X1
X_118_ pc_in[2] gnd _120_/A vdd INVX1
XSFILL18480x12100 gnd vdd FILL
X_203_ _203_/A _200_/D _214_/C gnd _204_/C vdd OAI21X1
X_220_ _211_/A pc_in[11] _220_/C _211_/D gnd _220_/Y vdd AOI22X1
X_134_ _282_/Q _134_/B gnd _135_/C vdd NAND2X1
X_151_ pc_in[13] gnd _153_/A vdd INVX1
X_117_ _115_/Y _117_/B _116_/Y gnd _117_/Y vdd OAI21X1
X_279_ _125_/A _262_/CLK _126_/Y gnd vdd DFFPOSX1
X_150_ _224_/B _147_/B _149_/Y gnd _150_/Y vdd OAI21X1
X_133_ pc_in[7] gnd _133_/Y vdd INVX2
X_202_ _137_/A _211_/D gnd _202_/Y vdd NAND2X1
X_116_ _276_/Q _117_/B gnd _116_/Y vdd NAND2X1
X_201_ _197_/Y _200_/Y _196_/Y gnd _201_/Y vdd OAI21X1
X_278_ _174_/A _262_/CLK _123_/Y gnd vdd DFFPOSX1
XSFILL6480x6100 gnd vdd FILL
X_132_ _132_/A _131_/B _132_/C gnd _281_/D vdd OAI21X1
X_115_ pc_in[1] gnd _115_/Y vdd INVX1
.ends

