* NGSPICE file created from map9v3.ext - technology: scmos

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

.subckt map9v3 gnd vdd N[8] N[7] N[6] N[5] N[4] N[3] N[2] N[1] N[0] clock counter[7]
+ counter[6] counter[5] counter[4] counter[3] counter[2] counter[1] counter[0] done
+ dp[8] dp[7] dp[6] dp[5] dp[4] dp[3] dp[2] dp[1] dp[0] reset sr[7] sr[6] sr[5] sr[4]
+ sr[3] sr[2] sr[1] sr[0] start
X_294_ _272_/A _296_/CLK _294_/R vdd _145_/Y gnd vdd DFFSR
X_131_ _131_/A gnd _135_/C vdd INVX1
XSFILL5200x12100 gnd vdd FILL
X_200_ _195_/Y _200_/B gnd _302_/D vdd NAND2X1
X_277_ _158_/A gnd dp[8] vdd BUFX2
XSFILL19600x16100 gnd vdd FILL
X_293_ _271_/A _291_/CLK _304_/R vdd _293_/D gnd vdd DFFSR
X_276_ _155_/A gnd dp[7] vdd BUFX2
X_130_ _256_/A _249_/B _130_/C gnd _130_/Y vdd OAI21X1
XSFILL6800x100 gnd vdd FILL
XSFILL7120x2100 gnd vdd FILL
X_259_ reset gnd _259_/Y vdd INVX8
X_292_ _292_/Q _314_/CLK _314_/R vdd _139_/Y gnd vdd DFFSR
X_275_ _275_/A gnd dp[6] vdd BUFX2
X_189_ _256_/A _260_/A gnd _190_/B vdd AND2X2
X_258_ _258_/A _128_/A gnd _258_/Y vdd AND2X2
XSFILL19920x4100 gnd vdd FILL
X_291_ _161_/A _291_/CLK _304_/R vdd _291_/D gnd vdd DFFSR
XSFILL6640x14100 gnd vdd FILL
XSFILL7120x8100 gnd vdd FILL
X_274_ _296_/Q gnd dp[5] vdd BUFX2
X_257_ _134_/Y _287_/Q gnd _286_/D vdd AND2X2
X_188_ _260_/A _256_/A gnd _188_/Y vdd NOR2X1
X_309_ _255_/A _314_/CLK _314_/R vdd _309_/D gnd vdd DFFSR
X_290_ _131_/A _291_/CLK _304_/R vdd _290_/D gnd vdd DFFSR
X_256_ _256_/A _141_/Y _255_/Y gnd _256_/Y vdd AOI21X1
X_187_ N[1] gnd _187_/Y vdd INVX1
XSFILL6640x2100 gnd vdd FILL
X_273_ _146_/A gnd dp[4] vdd BUFX2
X_239_ _126_/B gnd _239_/Y vdd INVX1
X_308_ _267_/A _302_/CLK _288_/R vdd _250_/Y gnd vdd DFFSR
X_272_ _272_/A gnd dp[3] vdd BUFX2
XSFILL6960x100 gnd vdd FILL
XBUFX2_insert5 _121_/Y gnd _175_/C vdd BUFX2
X_186_ _184_/A _160_/B _186_/C gnd _316_/D vdd AOI21X1
X_255_ _255_/A _177_/B _173_/C gnd _255_/Y vdd OAI21X1
XSFILL7280x10100 gnd vdd FILL
XSFILL6640x8100 gnd vdd FILL
X_169_ _183_/A _160_/B gnd _171_/B vdd NOR2X1
X_307_ _126_/B _302_/CLK _288_/R vdd _307_/D gnd vdd DFFSR
X_238_ N[7] _237_/Y _286_/Q gnd _238_/Y vdd OAI21X1
XSFILL19760x14100 gnd vdd FILL
X_271_ _271_/A gnd dp[2] vdd BUFX2
X_254_ _253_/Y _251_/Y _286_/Q gnd _254_/Y vdd AOI21X1
X_185_ _156_/A _184_/A _175_/C gnd _186_/C vdd OAI21X1
XFILL24560x2100 gnd vdd FILL
X_168_ _285_/A _154_/B gnd _171_/A vdd NOR2X1
XBUFX2_insert6 _121_/Y gnd _216_/A vdd BUFX2
X_237_ _194_/A _218_/Y _236_/Y gnd _237_/Y vdd NAND3X1
X_306_ _306_/Q _302_/CLK _288_/R vdd _306_/D gnd vdd DFFSR
XSFILL7280x16100 gnd vdd FILL
X_270_ _292_/Q gnd dp[1] vdd BUFX2
X_184_ _184_/A _184_/B _183_/Y gnd _315_/D vdd AOI21X1
X_253_ _131_/A _256_/A _253_/C gnd _253_/Y vdd NAND3X1
XBUFX2_insert7 _121_/Y gnd _173_/C vdd BUFX2
X_167_ _165_/Y _167_/B _164_/Y gnd _172_/A vdd OAI21X1
X_219_ _218_/Y _194_/A _219_/C gnd _224_/A vdd AOI21X1
X_305_ _264_/A _302_/CLK _288_/R vdd _305_/D gnd vdd DFFSR
X_236_ N[5] N[6] gnd _236_/Y vdd NOR2X1
XSFILL5040x12100 gnd vdd FILL
X_183_ _183_/A _184_/A _175_/C gnd _183_/Y vdd OAI21X1
X_252_ _290_/D gnd _253_/C vdd INVX1
XBUFX2_insert8 _121_/Y gnd _130_/C vdd BUFX2
X_166_ _166_/A _166_/B gnd _167_/B vdd NOR2X1
X_304_ _304_/Q _291_/CLK _304_/R vdd _216_/Y gnd vdd DFFSR
X_235_ _233_/Y _234_/Y gnd _235_/Y vdd NOR2X1
X_149_ _296_/Q gnd _151_/A vdd INVX1
X_218_ N[3] N[4] gnd _218_/Y vdd NOR2X1
XCLKBUF1_insert0 clock gnd _302_/CLK vdd CLKBUF1
XSFILL20080x4100 gnd vdd FILL
XSFILL19440x16100 gnd vdd FILL
X_251_ _300_/Q gnd _251_/Y vdd INVX1
X_182_ _176_/A _154_/B _181_/Y gnd _314_/D vdd AOI21X1
XBUFX2_insert9 _259_/Y gnd _288_/R vdd BUFX2
XCLKBUF1_insert1 clock gnd _291_/CLK vdd CLKBUF1
X_165_ _181_/A _178_/B gnd _165_/Y vdd NOR2X1
X_234_ _234_/A _211_/A gnd _234_/Y vdd NOR2X1
X_217_ N[5] gnd _219_/C vdd INVX1
X_148_ _146_/Y _178_/B _162_/B gnd _295_/D vdd MUX2X1
X_303_ _212_/B _302_/CLK _288_/R vdd _303_/D gnd vdd DFFSR
XSFILL6960x4100 gnd vdd FILL
XFILL24560x12100 gnd vdd FILL
X_181_ _181_/A _176_/A _175_/C gnd _181_/Y vdd OAI21X1
X_302_ _261_/A _302_/CLK _288_/R vdd _302_/D gnd vdd DFFSR
X_233_ N[7] gnd _233_/Y vdd INVX1
X_250_ _286_/Q _250_/B _248_/Y gnd _250_/Y vdd OAI21X1
X_164_ _183_/A _285_/A gnd _164_/Y vdd XNOR2X1
X_216_ _216_/A _211_/Y _215_/Y gnd _216_/Y vdd OAI21X1
XCLKBUF1_insert2 clock gnd _314_/CLK vdd CLKBUF1
XSFILL6800x4100 gnd vdd FILL
X_147_ _166_/A gnd _178_/B vdd INVX1
XSFILL6480x14100 gnd vdd FILL
XSFILL6960x10100 gnd vdd FILL
X_180_ _177_/B _166_/B _180_/C gnd _313_/D vdd AOI21X1
X_163_ _161_/Y _162_/B _163_/C gnd _291_/D vdd AOI21X1
X_301_ _260_/A _287_/CLK _301_/R vdd _191_/Y gnd vdd DFFSR
X_232_ _216_/A _227_/Y _231_/Y gnd _306_/D vdd OAI21X1
XCLKBUF1_insert3 clock gnd _296_/CLK vdd CLKBUF1
X_215_ _216_/A _214_/Y gnd _215_/Y vdd NAND2X1
X_129_ _129_/A _125_/Y gnd _249_/B vdd NOR2X1
X_146_ _146_/A gnd _146_/Y vdd INVX1
X_162_ N[0] _162_/B gnd _163_/C vdd NOR2X1
X_300_ _300_/Q _287_/CLK _301_/R vdd _254_/Y gnd vdd DFFSR
XSFILL19600x14100 gnd vdd FILL
XSFILL7120x10100 gnd vdd FILL
X_231_ _258_/A _230_/Y _216_/A gnd _231_/Y vdd OAI21X1
XCLKBUF1_insert4 clock gnd _287_/CLK vdd CLKBUF1
X_145_ _145_/A _145_/B _162_/B gnd _145_/Y vdd MUX2X1
X_214_ _221_/B _201_/Y _213_/Y gnd _214_/Y vdd OAI21X1
X_128_ _128_/A _127_/Y gnd _129_/A vdd NAND2X1
X_161_ _161_/A gnd _161_/Y vdd INVX1
X_230_ _230_/A _199_/A _229_/Y gnd _230_/Y vdd AOI21X1
XSFILL7120x16100 gnd vdd FILL
X_144_ _280_/A gnd _145_/B vdd INVX1
X_127_ _261_/A _260_/A gnd _127_/Y vdd NOR2X1
X_213_ _212_/B _201_/Y _304_/Q gnd _213_/Y vdd OAI21X1
XSFILL18640x6100 gnd vdd FILL
XSFILL19280x100 gnd vdd FILL
X_143_ _272_/A gnd _145_/A vdd INVX1
XBUFX2_insert10 _259_/Y gnd _301_/R vdd BUFX2
X_289_ _289_/Q _287_/CLK _301_/R vdd _130_/Y gnd vdd DFFSR
X_212_ _304_/Q _212_/B gnd _221_/B vdd OR2X2
X_160_ _158_/Y _160_/B _162_/B gnd _299_/D vdd MUX2X1
X_126_ _267_/A _126_/B gnd _128_/A vdd NOR2X1
XSFILL19440x2100 gnd vdd FILL
X_288_ _290_/D _302_/CLK _288_/R vdd _258_/Y gnd vdd DFFSR
XBUFX2_insert11 _259_/Y gnd _314_/R vdd BUFX2
X_142_ _140_/Y _141_/Y _162_/B gnd _293_/D vdd MUX2X1
XSFILL19280x10100 gnd vdd FILL
X_211_ _211_/A _211_/B gnd _211_/Y vdd NAND2X1
X_125_ _125_/A _124_/Y gnd _125_/Y vdd NAND2X1
XSFILL19440x8100 gnd vdd FILL
X_287_ _287_/Q _287_/CLK _301_/R vdd _135_/Y gnd vdd DFFSR
XFILL24400x12100 gnd vdd FILL
X_141_ _279_/A gnd _141_/Y vdd INVX1
XBUFX2_insert12 _259_/Y gnd _304_/R vdd BUFX2
X_210_ _203_/Y _210_/B _194_/A gnd _211_/A vdd NAND3X1
XSFILL17840x12100 gnd vdd FILL
X_124_ _306_/Q _264_/A gnd _124_/Y vdd NOR2X1
XSFILL19280x16100 gnd vdd FILL
XSFILL6640x6100 gnd vdd FILL
XBUFX2_insert13 _259_/Y gnd _294_/R vdd BUFX2
X_286_ _286_/Q _287_/CLK vdd _301_/R _286_/D gnd vdd DFFSR
X_269_ _161_/A gnd dp[0] vdd BUFX2
X_140_ _271_/A gnd _140_/Y vdd INVX1
XSFILL18960x2100 gnd vdd FILL
XSFILL18000x12100 gnd vdd FILL
XSFILL6800x10100 gnd vdd FILL
X_123_ _304_/Q _212_/B gnd _125_/A vdd NOR2X1
X_285_ _285_/A gnd sr[7] vdd BUFX2
XBUFX2_insert14 _122_/Y gnd _177_/B vdd BUFX2
X_268_ _300_/Q gnd done vdd BUFX2
X_122_ _289_/Q gnd _122_/Y vdd INVX8
X_199_ _199_/A _199_/B _130_/C gnd _200_/B vdd OAI21X1
XBUFX2_insert15 _122_/Y gnd _256_/A vdd BUFX2
X_284_ _156_/A gnd sr[6] vdd BUFX2
X_198_ _198_/A _188_/Y gnd _199_/B vdd NOR2X1
X_267_ _267_/A gnd counter[7] vdd BUFX2
X_121_ _286_/Q gnd _121_/Y vdd INVX4
XSFILL19440x100 gnd vdd FILL
XSFILL19760x4100 gnd vdd FILL
XSFILL19440x14100 gnd vdd FILL
XBUFX2_insert16 _122_/Y gnd _176_/A vdd BUFX2
X_283_ _183_/A gnd sr[5] vdd BUFX2
X_318_ _134_/A _287_/CLK _301_/R vdd _317_/Q gnd vdd DFFSR
X_197_ _261_/A gnd _198_/A vdd INVX1
X_266_ _126_/B gnd counter[6] vdd BUFX2
X_249_ _289_/Q _249_/B _267_/A _241_/Y gnd _250_/B vdd AOI22X1
XSFILL6960x2100 gnd vdd FILL
XSFILL18960x10100 gnd vdd FILL
XBUFX2_insert17 _122_/Y gnd _184_/A vdd BUFX2
XSFILL5520x12100 gnd vdd FILL
X_196_ _127_/Y _289_/Q gnd _199_/A vdd AND2X2
X_265_ _306_/Q gnd counter[5] vdd BUFX2
X_282_ _181_/A gnd sr[4] vdd BUFX2
X_317_ _317_/Q _291_/CLK _301_/R vdd start gnd vdd DFFSR
X_179_ _166_/A _176_/A _173_/C gnd _180_/C vdd OAI21X1
X_248_ _286_/Q _245_/Y _247_/Y gnd _248_/Y vdd NAND3X1
XSFILL6960x8100 gnd vdd FILL
XSFILL6800x2100 gnd vdd FILL
XSFILL19120x10100 gnd vdd FILL
X_281_ _166_/A gnd sr[3] vdd BUFX2
XFILL24560x16100 gnd vdd FILL
X_195_ _192_/Y _195_/B _286_/Q gnd _195_/Y vdd OAI21X1
X_264_ _264_/A gnd counter[4] vdd BUFX2
X_247_ _233_/Y _246_/Y _234_/Y gnd _247_/Y vdd NAND3X1
X_316_ _285_/A _314_/CLK _314_/R vdd _316_/D gnd vdd DFFSR
X_178_ _177_/B _178_/B _178_/C gnd _312_/D vdd AOI21X1
X_280_ _280_/A gnd sr[2] vdd BUFX2
X_194_ _194_/A gnd _195_/B vdd INVX1
XSFILL6800x8100 gnd vdd FILL
X_263_ _304_/Q gnd counter[3] vdd BUFX2
XSFILL19120x16100 gnd vdd FILL
X_177_ _280_/A _177_/B _175_/C gnd _178_/C vdd OAI21X1
X_315_ _156_/A _296_/CLK _294_/R vdd _315_/D gnd vdd DFFSR
X_246_ N[8] gnd _246_/Y vdd INVX1
XSFILL6960x14100 gnd vdd FILL
X_229_ _306_/Q gnd _229_/Y vdd INVX1
X_193_ N[1] N[2] gnd _194_/A vdd NAND2X1
X_262_ _212_/B gnd counter[2] vdd BUFX2
XSFILL17680x12100 gnd vdd FILL
X_176_ _176_/A _145_/B _175_/Y gnd _176_/Y vdd AOI21X1
X_314_ _183_/A _314_/CLK _314_/R vdd _314_/D gnd vdd DFFSR
X_245_ N[7] _237_/Y N[8] gnd _245_/Y vdd OAI21X1
X_228_ _201_/Y _125_/Y gnd _258_/A vdd NOR2X1
X_159_ _285_/A gnd _160_/B vdd INVX1
X_261_ _261_/A gnd counter[1] vdd BUFX2
X_192_ N[1] N[2] gnd _192_/Y vdd NOR2X1
X_175_ _279_/A _176_/A _175_/C gnd _175_/Y vdd OAI21X1
X_313_ _181_/A _291_/CLK _304_/R vdd _313_/D gnd vdd DFFSR
X_244_ _235_/Y _238_/Y _286_/Q _244_/D gnd _307_/D vdd OAI22X1
XSFILL7120x4100 gnd vdd FILL
X_227_ _211_/A _234_/A _225_/Y gnd _227_/Y vdd OAI21X1
XSFILL19600x100 gnd vdd FILL
X_158_ _158_/A gnd _158_/Y vdd INVX1
X_260_ _260_/A gnd counter[0] vdd BUFX2
X_191_ _130_/C _187_/Y _191_/C gnd _191_/Y vdd OAI21X1
XSFILL20240x4100 gnd vdd FILL
XSFILL7600x16100 gnd vdd FILL
X_157_ _157_/A _184_/B _162_/B gnd _157_/Y vdd MUX2X1
X_226_ N[5] N[6] gnd _234_/A vdd OR2X2
X_243_ _241_/Y _243_/B gnd _244_/D vdd AND2X2
X_174_ _174_/A _289_/Q _173_/Y gnd _309_/D vdd AOI21X1
X_312_ _166_/A _314_/CLK _314_/R vdd _312_/D gnd vdd DFFSR
X_209_ N[4] gnd _210_/B vdd INVX1
X_311_ _280_/A _296_/CLK _294_/R vdd _176_/Y gnd vdd DFFSR
XSFILL18800x10100 gnd vdd FILL
X_190_ _188_/Y _190_/B _130_/C gnd _191_/C vdd OAI21X1
X_242_ _201_/Y _125_/Y _126_/B gnd _243_/B vdd OAI21X1
X_173_ _289_/Q _255_/A _173_/C gnd _173_/Y vdd OAI21X1
X_156_ _156_/A gnd _184_/B vdd INVX1
X_225_ N[5] _211_/A N[6] gnd _225_/Y vdd OAI21X1
X_208_ N[3] _195_/B N[4] gnd _211_/B vdd OAI21X1
X_139_ _139_/A _162_/B _139_/C gnd _139_/Y vdd AOI21X1
XSFILL6640x4100 gnd vdd FILL
X_155_ _155_/A gnd _157_/A vdd INVX1
X_310_ _279_/A _296_/CLK _294_/R vdd _256_/Y gnd vdd DFFSR
X_172_ _172_/A _172_/B gnd _174_/A vdd NAND2X1
X_241_ _239_/Y _199_/A _241_/C gnd _241_/Y vdd NAND3X1
X_224_ _224_/A _220_/Y _286_/Q _224_/D gnd _305_/D vdd OAI22X1
X_207_ _286_/Q _207_/B _207_/C gnd _303_/D vdd OAI21X1
X_138_ _255_/A _162_/B gnd _139_/C vdd NOR2X1
XFILL24400x16100 gnd vdd FILL
XSFILL5360x12100 gnd vdd FILL
X_171_ _171_/A _171_/B _170_/Y gnd _172_/B vdd OAI21X1
X_240_ _125_/A _124_/Y gnd _241_/C vdd AND2X2
X_154_ _152_/Y _154_/B _162_/B gnd _297_/D vdd MUX2X1
XSFILL7120x100 gnd vdd FILL
XSFILL19760x100 gnd vdd FILL
X_223_ _230_/A _199_/A _264_/A _223_/D gnd _224_/D vdd AOI22X1
X_137_ _290_/D _173_/C _177_/B gnd _162_/B vdd NAND3X1
X_206_ _286_/Q _204_/Y _206_/C gnd _207_/C vdd NAND3X1
XSFILL6800x14100 gnd vdd FILL
XSFILL18960x6100 gnd vdd FILL
XFILL24560x4100 gnd vdd FILL
X_170_ _166_/A _181_/A gnd _170_/Y vdd XNOR2X1
X_299_ _158_/A _314_/CLK _314_/R vdd _299_/D gnd vdd DFFSR
X_205_ N[3] _195_/B gnd _206_/C vdd NAND2X1
X_153_ _183_/A gnd _154_/B vdd INVX1
XSFILL6640x100 gnd vdd FILL
X_136_ _292_/Q gnd _139_/A vdd INVX1
XFILL24560x100 gnd vdd FILL
X_222_ _125_/A _199_/A gnd _223_/D vdd NAND2X1
XSFILL17520x12100 gnd vdd FILL
X_152_ _275_/A gnd _152_/Y vdd INVX1
X_298_ _155_/A _296_/CLK _294_/R vdd _157_/Y gnd vdd DFFSR
XSFILL18800x6100 gnd vdd FILL
XSFILL18480x6100 gnd vdd FILL
X_221_ _264_/A _221_/B gnd _230_/A vdd NOR2X1
XFILL24400x4100 gnd vdd FILL
X_135_ _135_/A _134_/Y _135_/C gnd _135_/Y vdd OAI21X1
X_204_ _203_/Y _194_/A gnd _204_/Y vdd NAND2X1
X_297_ _275_/A _291_/CLK _304_/R vdd _297_/D gnd vdd DFFSR
X_151_ _151_/A _166_/B _162_/B gnd _151_/Y vdd MUX2X1
X_134_ _134_/A _134_/B gnd _134_/Y vdd NOR2X1
XSFILL19760x8100 gnd vdd FILL
X_203_ N[3] gnd _203_/Y vdd INVX1
XSFILL19280x2100 gnd vdd FILL
X_220_ N[5] _211_/A _286_/Q gnd _220_/Y vdd OAI21X1
XSFILL19920x14100 gnd vdd FILL
X_296_ _296_/Q _296_/CLK _294_/R vdd _151_/Y gnd vdd DFFSR
X_279_ _279_/A gnd sr[1] vdd BUFX2
X_150_ _181_/A gnd _166_/B vdd INVX1
XSFILL6960x6100 gnd vdd FILL
X_133_ _317_/Q gnd _134_/B vdd INVX1
XSFILL19600x8100 gnd vdd FILL
XSFILL19280x8100 gnd vdd FILL
X_202_ _201_/Y _212_/B gnd _207_/B vdd XOR2X1
XSFILL19120x2100 gnd vdd FILL
XSFILL7440x16100 gnd vdd FILL
X_295_ _146_/A _314_/CLK _314_/R vdd _295_/D gnd vdd DFFSR
X_132_ _287_/Q gnd _135_/A vdd INVX1
X_201_ _289_/Q _127_/Y gnd _201_/Y vdd NAND2X1
XSFILL6800x6100 gnd vdd FILL
XSFILL6480x6100 gnd vdd FILL
X_278_ _255_/A gnd sr[0] vdd BUFX2
.ends

