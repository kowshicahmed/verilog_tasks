/* Verilog module written by vlog2Verilog (qflow) */

module internal_register(
    input clock,
    input [15:0] data_in,
    input enable,
    input [2:0] ra_adrs,
    output [15:0] ra_out,
    input [2:0] rb_adrs,
    output [15:0] rb_out,
    input [2:0] rd_adrs,
    input wr_en
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _588_ ;
wire _168_ ;
wire [15:0] \internal_reg[7]  ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _512_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire rb_adrs_0_bF$buf0 ;
wire rb_adrs_0_bF$buf1 ;
wire rb_adrs_0_bF$buf2 ;
wire rb_adrs_0_bF$buf3 ;
wire rb_adrs_0_bF$buf4 ;
wire rb_adrs_0_bF$buf5 ;
wire rb_adrs_0_bF$buf6 ;
wire rb_adrs_0_bF$buf7 ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire clock ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire [15:0] \internal_reg[2]  ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire _285_ ;
wire [15:0] _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _104__bF$buf0 ;
wire _104__bF$buf1 ;
wire _104__bF$buf2 ;
wire _104__bF$buf3 ;
wire _104__bF$buf4 ;
wire _429_ ;
wire _182_ ;
wire ra_adrs_1_bF$buf0 ;
wire ra_adrs_1_bF$buf1 ;
wire ra_adrs_1_bF$buf2 ;
wire ra_adrs_1_bF$buf3 ;
wire ra_adrs_1_bF$buf4 ;
wire ra_adrs_1_bF$buf5 ;
wire ra_adrs_1_bF$buf6 ;
wire ra_adrs_1_bF$buf7 ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _276_ ;
wire rb_adrs_2_bF$buf0 ;
wire rb_adrs_2_bF$buf1 ;
wire rb_adrs_2_bF$buf2 ;
wire rb_adrs_2_bF$buf3 ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _474__bF$buf0 ;
wire _474__bF$buf1 ;
wire _474__bF$buf2 ;
wire _474__bF$buf3 ;
wire _523_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _273_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire [15:0] \internal_reg[4]  ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _461_ ;
wire _517_ ;
wire _270_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _514_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire [15:0] _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire [15:0] data_in ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _475__bF$buf0 ;
wire _475__bF$buf1 ;
wire _475__bF$buf2 ;
wire _475__bF$buf3 ;
wire _475__bF$buf4 ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _404__bF$buf0 ;
wire _404__bF$buf1 ;
wire _404__bF$buf2 ;
wire _404__bF$buf3 ;
wire _404__bF$buf4 ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire [2:0] ra_adrs ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _423__bF$buf0 ;
wire _423__bF$buf1 ;
wire _423__bF$buf2 ;
wire _423__bF$buf3 ;
wire _423__bF$buf4 ;
wire _9_ ;
wire _505_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [15:0] \internal_reg[6]  ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire enable ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _370__bF$buf0 ;
wire _370__bF$buf1 ;
wire _370__bF$buf2 ;
wire _370__bF$buf3 ;
wire _370__bF$buf4 ;
wire [15:0] rb_out ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire [15:0] _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire [15:0] \internal_reg[1]  ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire clock_bF$buf10 ;
wire clock_bF$buf11 ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _525_ ;
wire _105_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire _525__bF$buf0 ;
wire _525__bF$buf1 ;
wire _525__bF$buf2 ;
wire _525__bF$buf3 ;
wire _525__bF$buf4 ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _272_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _269_ ;
wire _498_ ;
wire _26_ ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire ra_adrs_0_bF$buf0 ;
wire ra_adrs_0_bF$buf1 ;
wire ra_adrs_0_bF$buf2 ;
wire ra_adrs_0_bF$buf3 ;
wire ra_adrs_0_bF$buf4 ;
wire ra_adrs_0_bF$buf5 ;
wire ra_adrs_0_bF$buf6 ;
wire ra_adrs_0_bF$buf7 ;
wire _460_ ;
wire _516_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire rb_adrs_1_bF$buf0 ;
wire rb_adrs_1_bF$buf1 ;
wire rb_adrs_1_bF$buf2 ;
wire rb_adrs_1_bF$buf3 ;
wire rb_adrs_1_bF$buf4 ;
wire rb_adrs_1_bF$buf5 ;
wire rb_adrs_1_bF$buf6 ;
wire rb_adrs_1_bF$buf7 ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _513_ ;
wire [15:0] ra_out ;
wire _322_ ;
wire _94__bF$buf0 ;
wire _94__bF$buf1 ;
wire _94__bF$buf2 ;
wire _94__bF$buf3 ;
wire _94__bF$buf4 ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire [15:0] _683_ ;
wire _263_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire [15:0] \internal_reg[3]  ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _542__bF$buf0 ;
wire _542__bF$buf1 ;
wire _542__bF$buf2 ;
wire _542__bF$buf3 ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire [2:0] rb_adrs ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire [2:0] rd_adrs ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _307_ ;
wire clock_bF$buf0 ;
wire clock_bF$buf1 ;
wire clock_bF$buf2 ;
wire clock_bF$buf3 ;
wire clock_bF$buf4 ;
wire clock_bF$buf5 ;
wire clock_bF$buf6 ;
wire clock_bF$buf7 ;
wire _480_ ;
wire clock_bF$buf8 ;
wire clock_bF$buf9 ;
wire _536_ ;
wire _116_ ;
wire _402__bF$buf0 ;
wire _402__bF$buf1 ;
wire _402__bF$buf2 ;
wire _402__bF$buf3 ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire ra_adrs_2_bF$buf0 ;
wire ra_adrs_2_bF$buf1 ;
wire ra_adrs_2_bF$buf2 ;
wire ra_adrs_2_bF$buf3 ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _304_ ;
wire wr_en_bF$buf0 ;
wire wr_en_bF$buf1 ;
wire wr_en_bF$buf2 ;
wire wr_en_bF$buf3 ;
wire wr_en_bF$buf4 ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire [15:0] \internal_reg[5]  ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _301_ ;
wire _562__bF$buf0 ;
wire _562__bF$buf1 ;
wire _562__bF$buf2 ;
wire _562__bF$buf3 ;
wire _562__bF$buf4 ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire wr_en ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire _34_ ;
wire _116__bF$buf0 ;
wire _116__bF$buf1 ;
wire _116__bF$buf2 ;
wire _116__bF$buf3 ;
wire _116__bF$buf4 ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _524_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _462_ ;
wire _518_ ;
wire [15:0] \internal_reg[0]  ;
wire _271_ ;
wire _327_ ;
wire _422__bF$buf0 ;
wire _422__bF$buf1 ;
wire _422__bF$buf2 ;
wire _422__bF$buf3 ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _268_ ;
wire _497_ ;
wire _441__bF$buf0 ;
wire _441__bF$buf1 ;
wire _441__bF$buf2 ;
wire _441__bF$buf3 ;
wire _441__bF$buf4 ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _515_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert122 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf0)
);

BUFX2 BUFX2_insert121 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf1)
);

BUFX2 BUFX2_insert120 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf2)
);

BUFX2 BUFX2_insert119 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf3)
);

BUFX2 BUFX2_insert118 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf4)
);

BUFX2 BUFX2_insert117 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf5)
);

BUFX2 BUFX2_insert116 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf6)
);

BUFX2 BUFX2_insert115 (
    .A(rb_adrs[1]),
    .Y(rb_adrs_1_bF$buf7)
);

BUFX2 BUFX2_insert114 (
    .A(_562_),
    .Y(_562__bF$buf0)
);

BUFX2 BUFX2_insert113 (
    .A(_562_),
    .Y(_562__bF$buf1)
);

BUFX2 BUFX2_insert112 (
    .A(_562_),
    .Y(_562__bF$buf2)
);

BUFX2 BUFX2_insert111 (
    .A(_562_),
    .Y(_562__bF$buf3)
);

BUFX2 BUFX2_insert110 (
    .A(_562_),
    .Y(_562__bF$buf4)
);

BUFX2 BUFX2_insert109 (
    .A(_104_),
    .Y(_104__bF$buf0)
);

BUFX2 BUFX2_insert108 (
    .A(_104_),
    .Y(_104__bF$buf1)
);

BUFX2 BUFX2_insert107 (
    .A(_104_),
    .Y(_104__bF$buf2)
);

BUFX2 BUFX2_insert106 (
    .A(_104_),
    .Y(_104__bF$buf3)
);

BUFX2 BUFX2_insert105 (
    .A(_104_),
    .Y(_104__bF$buf4)
);

BUFX2 BUFX2_insert104 (
    .A(wr_en),
    .Y(wr_en_bF$buf0)
);

BUFX2 BUFX2_insert103 (
    .A(wr_en),
    .Y(wr_en_bF$buf1)
);

BUFX2 BUFX2_insert102 (
    .A(wr_en),
    .Y(wr_en_bF$buf2)
);

BUFX2 BUFX2_insert101 (
    .A(wr_en),
    .Y(wr_en_bF$buf3)
);

BUFX2 BUFX2_insert100 (
    .A(wr_en),
    .Y(wr_en_bF$buf4)
);

BUFX2 BUFX2_insert99 (
    .A(_474_),
    .Y(_474__bF$buf0)
);

BUFX2 BUFX2_insert98 (
    .A(_474_),
    .Y(_474__bF$buf1)
);

BUFX2 BUFX2_insert97 (
    .A(_474_),
    .Y(_474__bF$buf2)
);

BUFX2 BUFX2_insert96 (
    .A(_474_),
    .Y(_474__bF$buf3)
);

BUFX2 BUFX2_insert95 (
    .A(_116_),
    .Y(_116__bF$buf0)
);

BUFX2 BUFX2_insert94 (
    .A(_116_),
    .Y(_116__bF$buf1)
);

BUFX2 BUFX2_insert93 (
    .A(_116_),
    .Y(_116__bF$buf2)
);

BUFX2 BUFX2_insert92 (
    .A(_116_),
    .Y(_116__bF$buf3)
);

BUFX2 BUFX2_insert91 (
    .A(_116_),
    .Y(_116__bF$buf4)
);

BUFX2 BUFX2_insert90 (
    .A(_404_),
    .Y(_404__bF$buf0)
);

BUFX2 BUFX2_insert89 (
    .A(_404_),
    .Y(_404__bF$buf1)
);

BUFX2 BUFX2_insert88 (
    .A(_404_),
    .Y(_404__bF$buf2)
);

BUFX2 BUFX2_insert87 (
    .A(_404_),
    .Y(_404__bF$buf3)
);

BUFX2 BUFX2_insert86 (
    .A(_404_),
    .Y(_404__bF$buf4)
);

BUFX2 BUFX2_insert85 (
    .A(_542_),
    .Y(_542__bF$buf0)
);

BUFX2 BUFX2_insert84 (
    .A(_542_),
    .Y(_542__bF$buf1)
);

BUFX2 BUFX2_insert83 (
    .A(_542_),
    .Y(_542__bF$buf2)
);

BUFX2 BUFX2_insert82 (
    .A(_542_),
    .Y(_542__bF$buf3)
);

BUFX2 BUFX2_insert81 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf0)
);

BUFX2 BUFX2_insert80 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf1)
);

BUFX2 BUFX2_insert79 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf2)
);

BUFX2 BUFX2_insert78 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf3)
);

BUFX2 BUFX2_insert77 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf4)
);

BUFX2 BUFX2_insert76 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf5)
);

BUFX2 BUFX2_insert75 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf6)
);

BUFX2 BUFX2_insert74 (
    .A(ra_adrs[0]),
    .Y(ra_adrs_0_bF$buf7)
);

BUFX2 BUFX2_insert73 (
    .A(_422_),
    .Y(_422__bF$buf0)
);

BUFX2 BUFX2_insert72 (
    .A(_422_),
    .Y(_422__bF$buf1)
);

BUFX2 BUFX2_insert71 (
    .A(_422_),
    .Y(_422__bF$buf2)
);

BUFX2 BUFX2_insert70 (
    .A(_422_),
    .Y(_422__bF$buf3)
);

BUFX2 BUFX2_insert69 (
    .A(rb_adrs[2]),
    .Y(rb_adrs_2_bF$buf0)
);

BUFX2 BUFX2_insert68 (
    .A(rb_adrs[2]),
    .Y(rb_adrs_2_bF$buf1)
);

BUFX2 BUFX2_insert67 (
    .A(rb_adrs[2]),
    .Y(rb_adrs_2_bF$buf2)
);

BUFX2 BUFX2_insert66 (
    .A(rb_adrs[2]),
    .Y(rb_adrs_2_bF$buf3)
);

BUFX2 BUFX2_insert65 (
    .A(_525_),
    .Y(_525__bF$buf0)
);

BUFX2 BUFX2_insert64 (
    .A(_525_),
    .Y(_525__bF$buf1)
);

BUFX2 BUFX2_insert63 (
    .A(_525_),
    .Y(_525__bF$buf2)
);

BUFX2 BUFX2_insert62 (
    .A(_525_),
    .Y(_525__bF$buf3)
);

BUFX2 BUFX2_insert61 (
    .A(_525_),
    .Y(_525__bF$buf4)
);

BUFX2 BUFX2_insert60 (
    .A(_475_),
    .Y(_475__bF$buf0)
);

BUFX2 BUFX2_insert59 (
    .A(_475_),
    .Y(_475__bF$buf1)
);

BUFX2 BUFX2_insert58 (
    .A(_475_),
    .Y(_475__bF$buf2)
);

BUFX2 BUFX2_insert57 (
    .A(_475_),
    .Y(_475__bF$buf3)
);

BUFX2 BUFX2_insert56 (
    .A(_475_),
    .Y(_475__bF$buf4)
);

BUFX2 BUFX2_insert55 (
    .A(_402_),
    .Y(_402__bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .A(_402_),
    .Y(_402__bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .A(_402_),
    .Y(_402__bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .A(_402_),
    .Y(_402__bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .A(_94_),
    .Y(_94__bF$buf0)
);

BUFX2 BUFX2_insert50 (
    .A(_94_),
    .Y(_94__bF$buf1)
);

BUFX2 BUFX2_insert49 (
    .A(_94_),
    .Y(_94__bF$buf2)
);

BUFX2 BUFX2_insert48 (
    .A(_94_),
    .Y(_94__bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .A(_94_),
    .Y(_94__bF$buf4)
);

BUFX2 BUFX2_insert46 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf0)
);

BUFX2 BUFX2_insert45 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf4)
);

BUFX2 BUFX2_insert41 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf5)
);

BUFX2 BUFX2_insert40 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf6)
);

BUFX2 BUFX2_insert39 (
    .A(ra_adrs[1]),
    .Y(ra_adrs_1_bF$buf7)
);

BUFX2 BUFX2_insert38 (
    .A(_423_),
    .Y(_423__bF$buf0)
);

BUFX2 BUFX2_insert37 (
    .A(_423_),
    .Y(_423__bF$buf1)
);

BUFX2 BUFX2_insert36 (
    .A(_423_),
    .Y(_423__bF$buf2)
);

BUFX2 BUFX2_insert35 (
    .A(_423_),
    .Y(_423__bF$buf3)
);

BUFX2 BUFX2_insert34 (
    .A(_423_),
    .Y(_423__bF$buf4)
);

BUFX2 BUFX2_insert33 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf0)
);

BUFX2 BUFX2_insert32 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf1)
);

BUFX2 BUFX2_insert31 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf2)
);

BUFX2 BUFX2_insert30 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf3)
);

BUFX2 BUFX2_insert29 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf4)
);

BUFX2 BUFX2_insert28 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf5)
);

BUFX2 BUFX2_insert27 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf6)
);

BUFX2 BUFX2_insert26 (
    .A(rb_adrs[0]),
    .Y(rb_adrs_0_bF$buf7)
);

BUFX2 BUFX2_insert25 (
    .A(_370_),
    .Y(_370__bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .A(_370_),
    .Y(_370__bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .A(_370_),
    .Y(_370__bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .A(_370_),
    .Y(_370__bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .A(_370_),
    .Y(_370__bF$buf4)
);

BUFX2 BUFX2_insert20 (
    .A(_441_),
    .Y(_441__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .A(_441_),
    .Y(_441__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .A(_441_),
    .Y(_441__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .A(_441_),
    .Y(_441__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .A(_441_),
    .Y(_441__bF$buf4)
);

CLKBUF1 CLKBUF1_insert15 (
    .A(clock),
    .Y(clock_bF$buf0)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clock),
    .Y(clock_bF$buf1)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clock),
    .Y(clock_bF$buf2)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clock),
    .Y(clock_bF$buf3)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clock),
    .Y(clock_bF$buf4)
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clock),
    .Y(clock_bF$buf5)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clock),
    .Y(clock_bF$buf6)
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clock),
    .Y(clock_bF$buf7)
);

CLKBUF1 CLKBUF1_insert7 (
    .A(clock),
    .Y(clock_bF$buf8)
);

CLKBUF1 CLKBUF1_insert6 (
    .A(clock),
    .Y(clock_bF$buf9)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clock),
    .Y(clock_bF$buf10)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clock),
    .Y(clock_bF$buf11)
);

BUFX2 BUFX2_insert3 (
    .A(ra_adrs[2]),
    .Y(ra_adrs_2_bF$buf0)
);

BUFX2 BUFX2_insert2 (
    .A(ra_adrs[2]),
    .Y(ra_adrs_2_bF$buf1)
);

BUFX2 BUFX2_insert1 (
    .A(ra_adrs[2]),
    .Y(ra_adrs_2_bF$buf2)
);

BUFX2 BUFX2_insert0 (
    .A(ra_adrs[2]),
    .Y(ra_adrs_2_bF$buf3)
);

NAND2X1 _1000_ (
    .A(\internal_reg[2] [14]),
    .B(_423__bF$buf4),
    .Y(_438_)
);

OAI21X1 _1001_ (
    .A(_398_),
    .B(_423__bF$buf3),
    .C(_438_),
    .Y(_117_)
);

NAND2X1 _1002_ (
    .A(\internal_reg[2] [15]),
    .B(_423__bF$buf2),
    .Y(_439_)
);

OAI21X1 _1003_ (
    .A(_400_),
    .B(_423__bF$buf1),
    .C(_439_),
    .Y(_119_)
);

INVX1 _1004_ (
    .A(\internal_reg[3] [0]),
    .Y(_440_)
);

INVX8 _1005_ (
    .A(_404__bF$buf4),
    .Y(_441_)
);

AND2X2 _1006_ (
    .A(_441__bF$buf4),
    .B(_422__bF$buf3),
    .Y(_442_)
);

NAND3X1 _1007_ (
    .A(data_in[0]),
    .B(_422__bF$buf2),
    .C(_441__bF$buf3),
    .Y(_443_)
);

OAI21X1 _1008_ (
    .A(_440_),
    .B(_442_),
    .C(_443_),
    .Y(_123_)
);

INVX1 _1009_ (
    .A(\internal_reg[3] [1]),
    .Y(_444_)
);

NAND3X1 _1010_ (
    .A(data_in[1]),
    .B(_422__bF$buf1),
    .C(_441__bF$buf2),
    .Y(_445_)
);

OAI21X1 _1011_ (
    .A(_444_),
    .B(_442_),
    .C(_445_),
    .Y(_125_)
);

INVX1 _1012_ (
    .A(\internal_reg[3] [2]),
    .Y(_446_)
);

NAND3X1 _1013_ (
    .A(data_in[2]),
    .B(_422__bF$buf0),
    .C(_441__bF$buf1),
    .Y(_447_)
);

OAI21X1 _1014_ (
    .A(_446_),
    .B(_442_),
    .C(_447_),
    .Y(_127_)
);

INVX1 _1015_ (
    .A(\internal_reg[3] [3]),
    .Y(_448_)
);

NAND3X1 _1016_ (
    .A(data_in[3]),
    .B(_422__bF$buf3),
    .C(_441__bF$buf0),
    .Y(_449_)
);

OAI21X1 _1017_ (
    .A(_448_),
    .B(_442_),
    .C(_449_),
    .Y(_129_)
);

INVX1 _1018_ (
    .A(\internal_reg[3] [4]),
    .Y(_450_)
);

NAND3X1 _1019_ (
    .A(data_in[4]),
    .B(_422__bF$buf2),
    .C(_441__bF$buf4),
    .Y(_451_)
);

OAI21X1 _1020_ (
    .A(_450_),
    .B(_442_),
    .C(_451_),
    .Y(_131_)
);

INVX1 _1021_ (
    .A(\internal_reg[3] [5]),
    .Y(_452_)
);

NAND3X1 _1022_ (
    .A(data_in[5]),
    .B(_422__bF$buf1),
    .C(_441__bF$buf3),
    .Y(_453_)
);

OAI21X1 _1023_ (
    .A(_452_),
    .B(_442_),
    .C(_453_),
    .Y(_133_)
);

INVX1 _1024_ (
    .A(\internal_reg[3] [6]),
    .Y(_454_)
);

NAND3X1 _1025_ (
    .A(data_in[6]),
    .B(_422__bF$buf0),
    .C(_441__bF$buf2),
    .Y(_455_)
);

OAI21X1 _1026_ (
    .A(_454_),
    .B(_442_),
    .C(_455_),
    .Y(_135_)
);

INVX1 _1027_ (
    .A(\internal_reg[3] [7]),
    .Y(_456_)
);

NAND3X1 _1028_ (
    .A(data_in[7]),
    .B(_422__bF$buf3),
    .C(_441__bF$buf1),
    .Y(_457_)
);

OAI21X1 _1029_ (
    .A(_456_),
    .B(_442_),
    .C(_457_),
    .Y(_137_)
);

INVX1 _1030_ (
    .A(\internal_reg[3] [8]),
    .Y(_458_)
);

NAND3X1 _1031_ (
    .A(data_in[8]),
    .B(_422__bF$buf2),
    .C(_441__bF$buf0),
    .Y(_459_)
);

OAI21X1 _1032_ (
    .A(_458_),
    .B(_442_),
    .C(_459_),
    .Y(_139_)
);

INVX1 _1033_ (
    .A(\internal_reg[3] [9]),
    .Y(_460_)
);

NAND3X1 _1034_ (
    .A(data_in[9]),
    .B(_422__bF$buf1),
    .C(_441__bF$buf4),
    .Y(_461_)
);

OAI21X1 _1035_ (
    .A(_460_),
    .B(_442_),
    .C(_461_),
    .Y(_140_)
);

INVX1 _1036_ (
    .A(\internal_reg[3] [10]),
    .Y(_462_)
);

NAND3X1 _1037_ (
    .A(data_in[10]),
    .B(_422__bF$buf0),
    .C(_441__bF$buf3),
    .Y(_463_)
);

OAI21X1 _1038_ (
    .A(_462_),
    .B(_442_),
    .C(_463_),
    .Y(_142_)
);

INVX1 _1039_ (
    .A(\internal_reg[3] [11]),
    .Y(_464_)
);

NAND3X1 _1040_ (
    .A(data_in[11]),
    .B(_422__bF$buf3),
    .C(_441__bF$buf2),
    .Y(_465_)
);

OAI21X1 _1041_ (
    .A(_464_),
    .B(_442_),
    .C(_465_),
    .Y(_144_)
);

INVX1 _1042_ (
    .A(\internal_reg[3] [12]),
    .Y(_466_)
);

NAND3X1 _1043_ (
    .A(data_in[12]),
    .B(_422__bF$buf2),
    .C(_441__bF$buf1),
    .Y(_467_)
);

OAI21X1 _1044_ (
    .A(_466_),
    .B(_442_),
    .C(_467_),
    .Y(_146_)
);

INVX1 _1045_ (
    .A(\internal_reg[3] [13]),
    .Y(_468_)
);

NAND3X1 _1046_ (
    .A(data_in[13]),
    .B(_422__bF$buf1),
    .C(_441__bF$buf0),
    .Y(_469_)
);

OAI21X1 _1047_ (
    .A(_468_),
    .B(_442_),
    .C(_469_),
    .Y(_148_)
);

INVX1 _1048_ (
    .A(\internal_reg[3] [14]),
    .Y(_470_)
);

NAND3X1 _1049_ (
    .A(data_in[14]),
    .B(_422__bF$buf0),
    .C(_441__bF$buf4),
    .Y(_471_)
);

OAI21X1 _1050_ (
    .A(_470_),
    .B(_442_),
    .C(_471_),
    .Y(_150_)
);

INVX1 _1051_ (
    .A(\internal_reg[3] [15]),
    .Y(_472_)
);

NAND3X1 _1052_ (
    .A(data_in[15]),
    .B(_422__bF$buf3),
    .C(_441__bF$buf3),
    .Y(_473_)
);

OAI21X1 _1053_ (
    .A(_472_),
    .B(_442_),
    .C(_473_),
    .Y(_152_)
);

NOR2X1 _1054_ (
    .A(rd_adrs[1]),
    .B(_366_),
    .Y(_474_)
);

NAND2X1 _1055_ (
    .A(_474__bF$buf3),
    .B(_369_),
    .Y(_475_)
);

NAND2X1 _1056_ (
    .A(\internal_reg[4] [0]),
    .B(_475__bF$buf4),
    .Y(_476_)
);

OAI21X1 _1057_ (
    .A(_365_),
    .B(_475__bF$buf3),
    .C(_476_),
    .Y(_157_)
);

NAND2X1 _1058_ (
    .A(\internal_reg[4] [1]),
    .B(_475__bF$buf2),
    .Y(_477_)
);

OAI21X1 _1059_ (
    .A(_372_),
    .B(_475__bF$buf1),
    .C(_477_),
    .Y(_159_)
);

NAND2X1 _1060_ (
    .A(\internal_reg[4] [2]),
    .B(_475__bF$buf0),
    .Y(_478_)
);

OAI21X1 _1061_ (
    .A(_374_),
    .B(_475__bF$buf4),
    .C(_478_),
    .Y(_160_)
);

NAND2X1 _1062_ (
    .A(\internal_reg[4] [3]),
    .B(_475__bF$buf3),
    .Y(_479_)
);

OAI21X1 _1063_ (
    .A(_376_),
    .B(_475__bF$buf2),
    .C(_479_),
    .Y(_162_)
);

NAND2X1 _1064_ (
    .A(\internal_reg[4] [4]),
    .B(_475__bF$buf1),
    .Y(_480_)
);

OAI21X1 _1065_ (
    .A(_378_),
    .B(_475__bF$buf0),
    .C(_480_),
    .Y(_164_)
);

NAND2X1 _1066_ (
    .A(\internal_reg[4] [5]),
    .B(_475__bF$buf4),
    .Y(_481_)
);

OAI21X1 _1067_ (
    .A(_380_),
    .B(_475__bF$buf3),
    .C(_481_),
    .Y(_166_)
);

NAND2X1 _1068_ (
    .A(\internal_reg[4] [6]),
    .B(_475__bF$buf2),
    .Y(_482_)
);

OAI21X1 _1069_ (
    .A(_382_),
    .B(_475__bF$buf1),
    .C(_482_),
    .Y(_168_)
);

NAND2X1 _1070_ (
    .A(\internal_reg[4] [7]),
    .B(_475__bF$buf0),
    .Y(_483_)
);

OAI21X1 _1071_ (
    .A(_384_),
    .B(_475__bF$buf4),
    .C(_483_),
    .Y(_170_)
);

NAND2X1 _1072_ (
    .A(\internal_reg[4] [8]),
    .B(_475__bF$buf3),
    .Y(_484_)
);

OAI21X1 _1073_ (
    .A(_386_),
    .B(_475__bF$buf2),
    .C(_484_),
    .Y(_172_)
);

NAND2X1 _1074_ (
    .A(\internal_reg[4] [9]),
    .B(_475__bF$buf1),
    .Y(_485_)
);

OAI21X1 _1075_ (
    .A(_388_),
    .B(_475__bF$buf0),
    .C(_485_),
    .Y(_174_)
);

NAND2X1 _1076_ (
    .A(\internal_reg[4] [10]),
    .B(_475__bF$buf4),
    .Y(_486_)
);

OAI21X1 _1077_ (
    .A(_390_),
    .B(_475__bF$buf3),
    .C(_486_),
    .Y(_176_)
);

NAND2X1 _1078_ (
    .A(\internal_reg[4] [11]),
    .B(_475__bF$buf2),
    .Y(_487_)
);

OAI21X1 _1079_ (
    .A(_392_),
    .B(_475__bF$buf1),
    .C(_487_),
    .Y(_178_)
);

NAND2X1 _1080_ (
    .A(\internal_reg[4] [12]),
    .B(_475__bF$buf0),
    .Y(_488_)
);

OAI21X1 _1081_ (
    .A(_394_),
    .B(_475__bF$buf4),
    .C(_488_),
    .Y(_180_)
);

NAND2X1 _1082_ (
    .A(\internal_reg[4] [13]),
    .B(_475__bF$buf3),
    .Y(_489_)
);

OAI21X1 _1083_ (
    .A(_396_),
    .B(_475__bF$buf2),
    .C(_489_),
    .Y(_182_)
);

NAND2X1 _1084_ (
    .A(\internal_reg[4] [14]),
    .B(_475__bF$buf1),
    .Y(_490_)
);

OAI21X1 _1085_ (
    .A(_398_),
    .B(_475__bF$buf0),
    .C(_490_),
    .Y(_183_)
);

NAND2X1 _1086_ (
    .A(\internal_reg[4] [15]),
    .B(_475__bF$buf4),
    .Y(_491_)
);

OAI21X1 _1087_ (
    .A(_400_),
    .B(_475__bF$buf3),
    .C(_491_),
    .Y(_185_)
);

INVX1 _1088_ (
    .A(\internal_reg[5] [0]),
    .Y(_492_)
);

AND2X2 _1089_ (
    .A(_441__bF$buf2),
    .B(_474__bF$buf2),
    .Y(_493_)
);

NAND3X1 _1090_ (
    .A(data_in[0]),
    .B(_474__bF$buf1),
    .C(_441__bF$buf1),
    .Y(_494_)
);

OAI21X1 _1091_ (
    .A(_492_),
    .B(_493_),
    .C(_494_),
    .Y(_189_)
);

INVX1 _1092_ (
    .A(\internal_reg[5] [1]),
    .Y(_495_)
);

NAND3X1 _1093_ (
    .A(data_in[1]),
    .B(_474__bF$buf0),
    .C(_441__bF$buf0),
    .Y(_496_)
);

OAI21X1 _1094_ (
    .A(_495_),
    .B(_493_),
    .C(_496_),
    .Y(_191_)
);

INVX1 _1095_ (
    .A(\internal_reg[5] [2]),
    .Y(_497_)
);

NAND3X1 _1096_ (
    .A(data_in[2]),
    .B(_474__bF$buf3),
    .C(_441__bF$buf4),
    .Y(_498_)
);

OAI21X1 _1097_ (
    .A(_497_),
    .B(_493_),
    .C(_498_),
    .Y(_193_)
);

INVX1 _1098_ (
    .A(\internal_reg[5] [3]),
    .Y(_499_)
);

NAND3X1 _1099_ (
    .A(data_in[3]),
    .B(_474__bF$buf2),
    .C(_441__bF$buf3),
    .Y(_500_)
);

OAI21X1 _1100_ (
    .A(_499_),
    .B(_493_),
    .C(_500_),
    .Y(_195_)
);

INVX1 _1101_ (
    .A(\internal_reg[5] [4]),
    .Y(_501_)
);

NAND3X1 _1102_ (
    .A(data_in[4]),
    .B(_474__bF$buf1),
    .C(_441__bF$buf2),
    .Y(_502_)
);

OAI21X1 _1103_ (
    .A(_501_),
    .B(_493_),
    .C(_502_),
    .Y(_197_)
);

INVX1 _1104_ (
    .A(\internal_reg[5] [5]),
    .Y(_503_)
);

NAND3X1 _1105_ (
    .A(data_in[5]),
    .B(_474__bF$buf0),
    .C(_441__bF$buf1),
    .Y(_504_)
);

OAI21X1 _1106_ (
    .A(_503_),
    .B(_493_),
    .C(_504_),
    .Y(_199_)
);

INVX1 _1107_ (
    .A(\internal_reg[5] [6]),
    .Y(_505_)
);

NAND3X1 _1108_ (
    .A(data_in[6]),
    .B(_474__bF$buf3),
    .C(_441__bF$buf0),
    .Y(_506_)
);

OAI21X1 _1109_ (
    .A(_505_),
    .B(_493_),
    .C(_506_),
    .Y(_201_)
);

INVX1 _1110_ (
    .A(\internal_reg[5] [7]),
    .Y(_507_)
);

NAND3X1 _1111_ (
    .A(data_in[7]),
    .B(_474__bF$buf2),
    .C(_441__bF$buf4),
    .Y(_508_)
);

OAI21X1 _1112_ (
    .A(_507_),
    .B(_493_),
    .C(_508_),
    .Y(_203_)
);

INVX1 _1113_ (
    .A(\internal_reg[5] [8]),
    .Y(_509_)
);

NAND3X1 _1114_ (
    .A(data_in[8]),
    .B(_474__bF$buf1),
    .C(_441__bF$buf3),
    .Y(_510_)
);

OAI21X1 _1115_ (
    .A(_509_),
    .B(_493_),
    .C(_510_),
    .Y(_204_)
);

INVX1 _1116_ (
    .A(\internal_reg[5] [9]),
    .Y(_511_)
);

NAND3X1 _1117_ (
    .A(data_in[9]),
    .B(_474__bF$buf0),
    .C(_441__bF$buf2),
    .Y(_512_)
);

OAI21X1 _1118_ (
    .A(_511_),
    .B(_493_),
    .C(_512_),
    .Y(_206_)
);

INVX1 _1119_ (
    .A(\internal_reg[5] [10]),
    .Y(_513_)
);

NAND3X1 _1120_ (
    .A(data_in[10]),
    .B(_474__bF$buf3),
    .C(_441__bF$buf1),
    .Y(_514_)
);

OAI21X1 _1121_ (
    .A(_513_),
    .B(_493_),
    .C(_514_),
    .Y(_208_)
);

INVX1 _1122_ (
    .A(\internal_reg[5] [11]),
    .Y(_515_)
);

NAND3X1 _1123_ (
    .A(data_in[11]),
    .B(_474__bF$buf2),
    .C(_441__bF$buf0),
    .Y(_516_)
);

OAI21X1 _1124_ (
    .A(_515_),
    .B(_493_),
    .C(_516_),
    .Y(_210_)
);

INVX1 _1125_ (
    .A(\internal_reg[5] [12]),
    .Y(_517_)
);

NAND3X1 _1126_ (
    .A(data_in[12]),
    .B(_474__bF$buf1),
    .C(_441__bF$buf4),
    .Y(_518_)
);

OAI21X1 _1127_ (
    .A(_517_),
    .B(_493_),
    .C(_518_),
    .Y(_212_)
);

INVX1 _1128_ (
    .A(\internal_reg[5] [13]),
    .Y(_519_)
);

NAND3X1 _1129_ (
    .A(data_in[13]),
    .B(_474__bF$buf0),
    .C(_441__bF$buf3),
    .Y(_520_)
);

OAI21X1 _1130_ (
    .A(_519_),
    .B(_493_),
    .C(_520_),
    .Y(_214_)
);

INVX1 _1131_ (
    .A(\internal_reg[5] [14]),
    .Y(_521_)
);

NAND3X1 _1132_ (
    .A(data_in[14]),
    .B(_474__bF$buf3),
    .C(_441__bF$buf2),
    .Y(_522_)
);

OAI21X1 _1133_ (
    .A(_521_),
    .B(_493_),
    .C(_522_),
    .Y(_216_)
);

INVX1 _1134_ (
    .A(\internal_reg[5] [15]),
    .Y(_523_)
);

NAND3X1 _1135_ (
    .A(data_in[15]),
    .B(_474__bF$buf2),
    .C(_441__bF$buf1),
    .Y(_524_)
);

OAI21X1 _1136_ (
    .A(_523_),
    .B(_493_),
    .C(_524_),
    .Y(_218_)
);

NAND3X1 _1137_ (
    .A(rd_adrs[2]),
    .B(rd_adrs[1]),
    .C(_369_),
    .Y(_525_)
);

NAND2X1 _1138_ (
    .A(\internal_reg[6] [0]),
    .B(_525__bF$buf4),
    .Y(_526_)
);

OAI21X1 _1139_ (
    .A(_365_),
    .B(_525__bF$buf3),
    .C(_526_),
    .Y(_223_)
);

NAND2X1 _1140_ (
    .A(\internal_reg[6] [1]),
    .B(_525__bF$buf2),
    .Y(_527_)
);

OAI21X1 _1141_ (
    .A(_372_),
    .B(_525__bF$buf1),
    .C(_527_),
    .Y(_224_)
);

NAND2X1 _1142_ (
    .A(\internal_reg[6] [2]),
    .B(_525__bF$buf0),
    .Y(_528_)
);

OAI21X1 _1143_ (
    .A(_374_),
    .B(_525__bF$buf4),
    .C(_528_),
    .Y(_226_)
);

NAND2X1 _1144_ (
    .A(\internal_reg[6] [3]),
    .B(_525__bF$buf3),
    .Y(_529_)
);

OAI21X1 _1145_ (
    .A(_376_),
    .B(_525__bF$buf2),
    .C(_529_),
    .Y(_228_)
);

NAND2X1 _1146_ (
    .A(\internal_reg[6] [4]),
    .B(_525__bF$buf1),
    .Y(_530_)
);

OAI21X1 _1147_ (
    .A(_378_),
    .B(_525__bF$buf0),
    .C(_530_),
    .Y(_230_)
);

NAND2X1 _1148_ (
    .A(\internal_reg[6] [5]),
    .B(_525__bF$buf4),
    .Y(_531_)
);

OAI21X1 _1149_ (
    .A(_380_),
    .B(_525__bF$buf3),
    .C(_531_),
    .Y(_232_)
);

NAND2X1 _1150_ (
    .A(\internal_reg[6] [6]),
    .B(_525__bF$buf2),
    .Y(_532_)
);

OAI21X1 _1151_ (
    .A(_382_),
    .B(_525__bF$buf1),
    .C(_532_),
    .Y(_234_)
);

NAND2X1 _1152_ (
    .A(\internal_reg[6] [7]),
    .B(_525__bF$buf0),
    .Y(_533_)
);

OAI21X1 _1153_ (
    .A(_384_),
    .B(_525__bF$buf4),
    .C(_533_),
    .Y(_236_)
);

NAND2X1 _1154_ (
    .A(\internal_reg[6] [8]),
    .B(_525__bF$buf3),
    .Y(_534_)
);

OAI21X1 _1155_ (
    .A(_386_),
    .B(_525__bF$buf2),
    .C(_534_),
    .Y(_238_)
);

NAND2X1 _1156_ (
    .A(\internal_reg[6] [9]),
    .B(_525__bF$buf1),
    .Y(_535_)
);

OAI21X1 _1157_ (
    .A(_388_),
    .B(_525__bF$buf0),
    .C(_535_),
    .Y(_240_)
);

NAND2X1 _1158_ (
    .A(\internal_reg[6] [10]),
    .B(_525__bF$buf4),
    .Y(_536_)
);

OAI21X1 _1159_ (
    .A(_390_),
    .B(_525__bF$buf3),
    .C(_536_),
    .Y(_242_)
);

NAND2X1 _1160_ (
    .A(\internal_reg[6] [11]),
    .B(_525__bF$buf2),
    .Y(_537_)
);

OAI21X1 _1161_ (
    .A(_392_),
    .B(_525__bF$buf1),
    .C(_537_),
    .Y(_244_)
);

NAND2X1 _1162_ (
    .A(\internal_reg[6] [12]),
    .B(_525__bF$buf0),
    .Y(_538_)
);

OAI21X1 _1163_ (
    .A(_394_),
    .B(_525__bF$buf4),
    .C(_538_),
    .Y(_246_)
);

NAND2X1 _1164_ (
    .A(\internal_reg[6] [13]),
    .B(_525__bF$buf3),
    .Y(_539_)
);

OAI21X1 _1165_ (
    .A(_396_),
    .B(_525__bF$buf2),
    .C(_539_),
    .Y(_247_)
);

NAND2X1 _1166_ (
    .A(\internal_reg[6] [14]),
    .B(_525__bF$buf1),
    .Y(_540_)
);

OAI21X1 _1167_ (
    .A(_398_),
    .B(_525__bF$buf0),
    .C(_540_),
    .Y(_249_)
);

NAND2X1 _1168_ (
    .A(\internal_reg[6] [15]),
    .B(_525__bF$buf4),
    .Y(_541_)
);

OAI21X1 _1169_ (
    .A(_400_),
    .B(_525__bF$buf3),
    .C(_541_),
    .Y(_251_)
);

NAND2X1 _1170_ (
    .A(rd_adrs[2]),
    .B(rd_adrs[1]),
    .Y(_542_)
);

OR2X2 _1171_ (
    .A(_404__bF$buf3),
    .B(_542__bF$buf3),
    .Y(_543_)
);

OAI21X1 _1172_ (
    .A(_542__bF$buf2),
    .B(_404__bF$buf2),
    .C(\internal_reg[7] [0]),
    .Y(_544_)
);

OAI21X1 _1173_ (
    .A(_365_),
    .B(_543_),
    .C(_544_),
    .Y(_255_)
);

OAI21X1 _1174_ (
    .A(_542__bF$buf1),
    .B(_404__bF$buf1),
    .C(\internal_reg[7] [1]),
    .Y(_545_)
);

OAI21X1 _1175_ (
    .A(_372_),
    .B(_543_),
    .C(_545_),
    .Y(_257_)
);

OAI21X1 _1176_ (
    .A(_542__bF$buf0),
    .B(_404__bF$buf0),
    .C(\internal_reg[7] [2]),
    .Y(_546_)
);

OAI21X1 _1177_ (
    .A(_374_),
    .B(_543_),
    .C(_546_),
    .Y(_259_)
);

OAI21X1 _1178_ (
    .A(_542__bF$buf3),
    .B(_404__bF$buf4),
    .C(\internal_reg[7] [3]),
    .Y(_547_)
);

OAI21X1 _1179_ (
    .A(_376_),
    .B(_543_),
    .C(_547_),
    .Y(_261_)
);

OAI21X1 _1180_ (
    .A(_542__bF$buf2),
    .B(_404__bF$buf3),
    .C(\internal_reg[7] [4]),
    .Y(_548_)
);

OAI21X1 _1181_ (
    .A(_378_),
    .B(_543_),
    .C(_548_),
    .Y(_263_)
);

OAI21X1 _1182_ (
    .A(_542__bF$buf1),
    .B(_404__bF$buf2),
    .C(\internal_reg[7] [5]),
    .Y(_549_)
);

OAI21X1 _1183_ (
    .A(_380_),
    .B(_543_),
    .C(_549_),
    .Y(_265_)
);

OAI21X1 _1184_ (
    .A(_542__bF$buf0),
    .B(_404__bF$buf1),
    .C(\internal_reg[7] [6]),
    .Y(_550_)
);

OAI21X1 _1185_ (
    .A(_382_),
    .B(_543_),
    .C(_550_),
    .Y(_267_)
);

OAI21X1 _1186_ (
    .A(_542__bF$buf3),
    .B(_404__bF$buf0),
    .C(\internal_reg[7] [7]),
    .Y(_551_)
);

OAI21X1 _1187_ (
    .A(_384_),
    .B(_543_),
    .C(_551_),
    .Y(_268_)
);

OAI21X1 _1188_ (
    .A(_542__bF$buf2),
    .B(_404__bF$buf4),
    .C(\internal_reg[7] [8]),
    .Y(_552_)
);

OAI21X1 _1189_ (
    .A(_386_),
    .B(_543_),
    .C(_552_),
    .Y(_270_)
);

OAI21X1 _1190_ (
    .A(_542__bF$buf1),
    .B(_404__bF$buf3),
    .C(\internal_reg[7] [9]),
    .Y(_553_)
);

OAI21X1 _1191_ (
    .A(_388_),
    .B(_543_),
    .C(_553_),
    .Y(_272_)
);

OAI21X1 _1192_ (
    .A(_542__bF$buf0),
    .B(_404__bF$buf2),
    .C(\internal_reg[7] [10]),
    .Y(_554_)
);

OAI21X1 _1193_ (
    .A(_390_),
    .B(_543_),
    .C(_554_),
    .Y(_274_)
);

OAI21X1 _1194_ (
    .A(_542__bF$buf3),
    .B(_404__bF$buf1),
    .C(\internal_reg[7] [11]),
    .Y(_555_)
);

OAI21X1 _1195_ (
    .A(_392_),
    .B(_543_),
    .C(_555_),
    .Y(_276_)
);

OAI21X1 _1196_ (
    .A(_542__bF$buf2),
    .B(_404__bF$buf0),
    .C(\internal_reg[7] [12]),
    .Y(_556_)
);

OAI21X1 _1197_ (
    .A(_394_),
    .B(_543_),
    .C(_556_),
    .Y(_278_)
);

OAI21X1 _1198_ (
    .A(_542__bF$buf1),
    .B(_404__bF$buf4),
    .C(\internal_reg[7] [13]),
    .Y(_557_)
);

OAI21X1 _1199_ (
    .A(_396_),
    .B(_543_),
    .C(_557_),
    .Y(_280_)
);

OAI21X1 _1200_ (
    .A(_542__bF$buf0),
    .B(_404__bF$buf3),
    .C(\internal_reg[7] [14]),
    .Y(_558_)
);

OAI21X1 _1201_ (
    .A(_398_),
    .B(_543_),
    .C(_558_),
    .Y(_282_)
);

OAI21X1 _1202_ (
    .A(_542__bF$buf3),
    .B(_404__bF$buf2),
    .C(\internal_reg[7] [15]),
    .Y(_559_)
);

OAI21X1 _1203_ (
    .A(_400_),
    .B(_543_),
    .C(_559_),
    .Y(_284_)
);

INVX4 _1204_ (
    .A(rb_adrs_2_bF$buf3),
    .Y(_560_)
);

MUX2X1 _1205_ (
    .A(\internal_reg[5] [0]),
    .B(\internal_reg[4] [0]),
    .S(rb_adrs_0_bF$buf7),
    .Y(_561_)
);

INVX8 _1206_ (
    .A(rb_adrs_0_bF$buf6),
    .Y(_562_)
);

NOR2X1 _1207_ (
    .A(\internal_reg[7] [0]),
    .B(_562__bF$buf4),
    .Y(_563_)
);

OAI21X1 _1208_ (
    .A(\internal_reg[6] [0]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_564_)
);

OAI22X1 _1209_ (
    .A(_564_),
    .B(_563_),
    .C(rb_adrs_1_bF$buf6),
    .D(_561_),
    .Y(_565_)
);

NOR2X1 _1210_ (
    .A(_560_),
    .B(_565_),
    .Y(_566_)
);

OAI21X1 _1211_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_684_[0]),
    .Y(_567_)
);

MUX2X1 _1212_ (
    .A(\internal_reg[1] [0]),
    .B(\internal_reg[0] [0]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_568_)
);

NOR2X1 _1213_ (
    .A(\internal_reg[3] [0]),
    .B(_562__bF$buf3),
    .Y(_569_)
);

OAI21X1 _1214_ (
    .A(\internal_reg[2] [0]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_570_)
);

OAI22X1 _1215_ (
    .A(_570_),
    .B(_569_),
    .C(rb_adrs_1_bF$buf4),
    .D(_568_),
    .Y(_571_)
);

OAI21X1 _1216_ (
    .A(rb_adrs_2_bF$buf2),
    .B(_571_),
    .C(_116__bF$buf4),
    .Y(_572_)
);

OAI21X1 _1217_ (
    .A(_566_),
    .B(_572_),
    .C(_567_),
    .Y(_1_[0])
);

MUX2X1 _1218_ (
    .A(\internal_reg[5] [1]),
    .B(\internal_reg[4] [1]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_573_)
);

NOR2X1 _1219_ (
    .A(\internal_reg[7] [1]),
    .B(_562__bF$buf2),
    .Y(_574_)
);

OAI21X1 _1220_ (
    .A(\internal_reg[6] [1]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_575_)
);

OAI22X1 _1221_ (
    .A(_575_),
    .B(_574_),
    .C(rb_adrs_1_bF$buf2),
    .D(_573_),
    .Y(_576_)
);

NOR2X1 _1222_ (
    .A(_560_),
    .B(_576_),
    .Y(_577_)
);

OAI21X1 _1223_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_684_[1]),
    .Y(_578_)
);

MUX2X1 _1224_ (
    .A(\internal_reg[1] [1]),
    .B(\internal_reg[0] [1]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_579_)
);

NOR2X1 _1225_ (
    .A(\internal_reg[3] [1]),
    .B(_562__bF$buf1),
    .Y(_580_)
);

OAI21X1 _1226_ (
    .A(\internal_reg[2] [1]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_581_)
);

OAI22X1 _1227_ (
    .A(_581_),
    .B(_580_),
    .C(rb_adrs_1_bF$buf0),
    .D(_579_),
    .Y(_582_)
);

OAI21X1 _1228_ (
    .A(rb_adrs_2_bF$buf1),
    .B(_582_),
    .C(_116__bF$buf3),
    .Y(_583_)
);

OAI21X1 _1229_ (
    .A(_577_),
    .B(_583_),
    .C(_578_),
    .Y(_1_[1])
);

MUX2X1 _1230_ (
    .A(\internal_reg[5] [2]),
    .B(\internal_reg[4] [2]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_584_)
);

NOR2X1 _1231_ (
    .A(\internal_reg[7] [2]),
    .B(_562__bF$buf0),
    .Y(_585_)
);

OAI21X1 _1232_ (
    .A(\internal_reg[6] [2]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_586_)
);

OAI22X1 _1233_ (
    .A(_586_),
    .B(_585_),
    .C(rb_adrs_1_bF$buf6),
    .D(_584_),
    .Y(_587_)
);

NOR2X1 _1234_ (
    .A(_560_),
    .B(_587_),
    .Y(_588_)
);

OAI21X1 _1235_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .C(_684_[2]),
    .Y(_589_)
);

MUX2X1 _1236_ (
    .A(\internal_reg[1] [2]),
    .B(\internal_reg[0] [2]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_590_)
);

NOR2X1 _1237_ (
    .A(\internal_reg[3] [2]),
    .B(_562__bF$buf4),
    .Y(_591_)
);

OAI21X1 _1238_ (
    .A(\internal_reg[2] [2]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_592_)
);

OAI22X1 _1239_ (
    .A(_592_),
    .B(_591_),
    .C(rb_adrs_1_bF$buf4),
    .D(_590_),
    .Y(_593_)
);

OAI21X1 _1240_ (
    .A(rb_adrs_2_bF$buf0),
    .B(_593_),
    .C(_116__bF$buf2),
    .Y(_594_)
);

OAI21X1 _1241_ (
    .A(_588_),
    .B(_594_),
    .C(_589_),
    .Y(_1_[2])
);

MUX2X1 _1242_ (
    .A(\internal_reg[5] [3]),
    .B(\internal_reg[4] [3]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_595_)
);

NOR2X1 _1243_ (
    .A(\internal_reg[7] [3]),
    .B(_562__bF$buf3),
    .Y(_596_)
);

OAI21X1 _1244_ (
    .A(\internal_reg[6] [3]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_597_)
);

OAI22X1 _1245_ (
    .A(_597_),
    .B(_596_),
    .C(rb_adrs_1_bF$buf2),
    .D(_595_),
    .Y(_598_)
);

NOR2X1 _1246_ (
    .A(_560_),
    .B(_598_),
    .Y(_599_)
);

OAI21X1 _1247_ (
    .A(wr_en_bF$buf1),
    .B(_104__bF$buf1),
    .C(_684_[3]),
    .Y(_600_)
);

MUX2X1 _1248_ (
    .A(\internal_reg[1] [3]),
    .B(\internal_reg[0] [3]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_601_)
);

NOR2X1 _1249_ (
    .A(\internal_reg[3] [3]),
    .B(_562__bF$buf2),
    .Y(_602_)
);

OAI21X1 _1250_ (
    .A(\internal_reg[2] [3]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_603_)
);

OAI22X1 _1251_ (
    .A(_603_),
    .B(_602_),
    .C(rb_adrs_1_bF$buf0),
    .D(_601_),
    .Y(_604_)
);

OAI21X1 _1252_ (
    .A(rb_adrs_2_bF$buf3),
    .B(_604_),
    .C(_116__bF$buf1),
    .Y(_605_)
);

OAI21X1 _1253_ (
    .A(_599_),
    .B(_605_),
    .C(_600_),
    .Y(_1_[3])
);

MUX2X1 _1254_ (
    .A(\internal_reg[5] [4]),
    .B(\internal_reg[4] [4]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_606_)
);

NOR2X1 _1255_ (
    .A(\internal_reg[7] [4]),
    .B(_562__bF$buf1),
    .Y(_607_)
);

OAI21X1 _1256_ (
    .A(\internal_reg[6] [4]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_608_)
);

OAI22X1 _1257_ (
    .A(_608_),
    .B(_607_),
    .C(rb_adrs_1_bF$buf6),
    .D(_606_),
    .Y(_609_)
);

NOR2X1 _1258_ (
    .A(_560_),
    .B(_609_),
    .Y(_610_)
);

OAI21X1 _1259_ (
    .A(wr_en_bF$buf0),
    .B(_104__bF$buf0),
    .C(_684_[4]),
    .Y(_611_)
);

MUX2X1 _1260_ (
    .A(\internal_reg[1] [4]),
    .B(\internal_reg[0] [4]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_612_)
);

NOR2X1 _1261_ (
    .A(\internal_reg[3] [4]),
    .B(_562__bF$buf0),
    .Y(_613_)
);

OAI21X1 _1262_ (
    .A(\internal_reg[2] [4]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_614_)
);

OAI22X1 _1263_ (
    .A(_614_),
    .B(_613_),
    .C(rb_adrs_1_bF$buf4),
    .D(_612_),
    .Y(_615_)
);

OAI21X1 _1264_ (
    .A(rb_adrs_2_bF$buf2),
    .B(_615_),
    .C(_116__bF$buf0),
    .Y(_616_)
);

OAI21X1 _1265_ (
    .A(_610_),
    .B(_616_),
    .C(_611_),
    .Y(_1_[4])
);

MUX2X1 _1266_ (
    .A(\internal_reg[5] [5]),
    .B(\internal_reg[4] [5]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_617_)
);

NOR2X1 _1267_ (
    .A(\internal_reg[7] [5]),
    .B(_562__bF$buf4),
    .Y(_618_)
);

OAI21X1 _1268_ (
    .A(\internal_reg[6] [5]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_619_)
);

OAI22X1 _1269_ (
    .A(_619_),
    .B(_618_),
    .C(rb_adrs_1_bF$buf2),
    .D(_617_),
    .Y(_620_)
);

NOR2X1 _1270_ (
    .A(_560_),
    .B(_620_),
    .Y(_621_)
);

OAI21X1 _1271_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_684_[5]),
    .Y(_622_)
);

MUX2X1 _1272_ (
    .A(\internal_reg[1] [5]),
    .B(\internal_reg[0] [5]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_623_)
);

NOR2X1 _1273_ (
    .A(\internal_reg[3] [5]),
    .B(_562__bF$buf3),
    .Y(_624_)
);

OAI21X1 _1274_ (
    .A(\internal_reg[2] [5]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_625_)
);

OAI22X1 _1275_ (
    .A(_625_),
    .B(_624_),
    .C(rb_adrs_1_bF$buf0),
    .D(_623_),
    .Y(_626_)
);

OAI21X1 _1276_ (
    .A(rb_adrs_2_bF$buf1),
    .B(_626_),
    .C(_116__bF$buf4),
    .Y(_627_)
);

OAI21X1 _1277_ (
    .A(_621_),
    .B(_627_),
    .C(_622_),
    .Y(_1_[5])
);

MUX2X1 _1278_ (
    .A(\internal_reg[5] [6]),
    .B(\internal_reg[4] [6]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_628_)
);

NOR2X1 _1279_ (
    .A(\internal_reg[7] [6]),
    .B(_562__bF$buf2),
    .Y(_629_)
);

OAI21X1 _1280_ (
    .A(\internal_reg[6] [6]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_630_)
);

OAI22X1 _1281_ (
    .A(_630_),
    .B(_629_),
    .C(rb_adrs_1_bF$buf6),
    .D(_628_),
    .Y(_631_)
);

NOR2X1 _1282_ (
    .A(_560_),
    .B(_631_),
    .Y(_632_)
);

OAI21X1 _1283_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_684_[6]),
    .Y(_633_)
);

MUX2X1 _1284_ (
    .A(\internal_reg[1] [6]),
    .B(\internal_reg[0] [6]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_634_)
);

NOR2X1 _1285_ (
    .A(\internal_reg[3] [6]),
    .B(_562__bF$buf1),
    .Y(_635_)
);

OAI21X1 _1286_ (
    .A(\internal_reg[2] [6]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_636_)
);

OAI22X1 _1287_ (
    .A(_636_),
    .B(_635_),
    .C(rb_adrs_1_bF$buf4),
    .D(_634_),
    .Y(_637_)
);

OAI21X1 _1288_ (
    .A(rb_adrs_2_bF$buf0),
    .B(_637_),
    .C(_116__bF$buf3),
    .Y(_638_)
);

OAI21X1 _1289_ (
    .A(_632_),
    .B(_638_),
    .C(_633_),
    .Y(_1_[6])
);

MUX2X1 _1290_ (
    .A(\internal_reg[5] [7]),
    .B(\internal_reg[4] [7]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_639_)
);

NOR2X1 _1291_ (
    .A(\internal_reg[7] [7]),
    .B(_562__bF$buf0),
    .Y(_640_)
);

OAI21X1 _1292_ (
    .A(\internal_reg[6] [7]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_641_)
);

OAI22X1 _1293_ (
    .A(_641_),
    .B(_640_),
    .C(rb_adrs_1_bF$buf2),
    .D(_639_),
    .Y(_642_)
);

NOR2X1 _1294_ (
    .A(_560_),
    .B(_642_),
    .Y(_643_)
);

OAI21X1 _1295_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .C(_684_[7]),
    .Y(_644_)
);

MUX2X1 _1296_ (
    .A(\internal_reg[1] [7]),
    .B(\internal_reg[0] [7]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_645_)
);

NOR2X1 _1297_ (
    .A(\internal_reg[3] [7]),
    .B(_562__bF$buf4),
    .Y(_646_)
);

OAI21X1 _1298_ (
    .A(\internal_reg[2] [7]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_647_)
);

OAI22X1 _1299_ (
    .A(_647_),
    .B(_646_),
    .C(rb_adrs_1_bF$buf0),
    .D(_645_),
    .Y(_648_)
);

OAI21X1 _1300_ (
    .A(rb_adrs_2_bF$buf3),
    .B(_648_),
    .C(_116__bF$buf2),
    .Y(_649_)
);

OAI21X1 _1301_ (
    .A(_643_),
    .B(_649_),
    .C(_644_),
    .Y(_1_[7])
);

MUX2X1 _1302_ (
    .A(\internal_reg[5] [8]),
    .B(\internal_reg[4] [8]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_650_)
);

NOR2X1 _1303_ (
    .A(\internal_reg[7] [8]),
    .B(_562__bF$buf3),
    .Y(_651_)
);

OAI21X1 _1304_ (
    .A(\internal_reg[6] [8]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_652_)
);

OAI22X1 _1305_ (
    .A(_652_),
    .B(_651_),
    .C(rb_adrs_1_bF$buf6),
    .D(_650_),
    .Y(_653_)
);

NOR2X1 _1306_ (
    .A(_560_),
    .B(_653_),
    .Y(_654_)
);

OAI21X1 _1307_ (
    .A(wr_en_bF$buf1),
    .B(_104__bF$buf1),
    .C(_684_[8]),
    .Y(_655_)
);

MUX2X1 _1308_ (
    .A(\internal_reg[1] [8]),
    .B(\internal_reg[0] [8]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_656_)
);

NOR2X1 _1309_ (
    .A(\internal_reg[3] [8]),
    .B(_562__bF$buf2),
    .Y(_657_)
);

OAI21X1 _1310_ (
    .A(\internal_reg[2] [8]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_658_)
);

OAI22X1 _1311_ (
    .A(_658_),
    .B(_657_),
    .C(rb_adrs_1_bF$buf4),
    .D(_656_),
    .Y(_659_)
);

OAI21X1 _1312_ (
    .A(rb_adrs_2_bF$buf2),
    .B(_659_),
    .C(_116__bF$buf1),
    .Y(_660_)
);

OAI21X1 _1313_ (
    .A(_654_),
    .B(_660_),
    .C(_655_),
    .Y(_1_[8])
);

MUX2X1 _1314_ (
    .A(\internal_reg[5] [9]),
    .B(\internal_reg[4] [9]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_661_)
);

NOR2X1 _1315_ (
    .A(\internal_reg[7] [9]),
    .B(_562__bF$buf1),
    .Y(_662_)
);

OAI21X1 _1316_ (
    .A(\internal_reg[6] [9]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_663_)
);

OAI22X1 _1317_ (
    .A(_663_),
    .B(_662_),
    .C(rb_adrs_1_bF$buf2),
    .D(_661_),
    .Y(_664_)
);

NOR2X1 _1318_ (
    .A(_560_),
    .B(_664_),
    .Y(_665_)
);

OAI21X1 _1319_ (
    .A(wr_en_bF$buf0),
    .B(_104__bF$buf0),
    .C(_684_[9]),
    .Y(_666_)
);

MUX2X1 _1320_ (
    .A(\internal_reg[1] [9]),
    .B(\internal_reg[0] [9]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_667_)
);

NOR2X1 _1321_ (
    .A(\internal_reg[3] [9]),
    .B(_562__bF$buf0),
    .Y(_668_)
);

OAI21X1 _1322_ (
    .A(\internal_reg[2] [9]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_669_)
);

OAI22X1 _1323_ (
    .A(_669_),
    .B(_668_),
    .C(rb_adrs_1_bF$buf0),
    .D(_667_),
    .Y(_670_)
);

OAI21X1 _1324_ (
    .A(rb_adrs_2_bF$buf1),
    .B(_670_),
    .C(_116__bF$buf0),
    .Y(_671_)
);

OAI21X1 _1325_ (
    .A(_665_),
    .B(_671_),
    .C(_666_),
    .Y(_1_[9])
);

MUX2X1 _1326_ (
    .A(\internal_reg[5] [10]),
    .B(\internal_reg[4] [10]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_672_)
);

NOR2X1 _1327_ (
    .A(\internal_reg[7] [10]),
    .B(_562__bF$buf4),
    .Y(_673_)
);

OAI21X1 _1328_ (
    .A(\internal_reg[6] [10]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_674_)
);

OAI22X1 _1329_ (
    .A(_674_),
    .B(_673_),
    .C(rb_adrs_1_bF$buf6),
    .D(_672_),
    .Y(_675_)
);

NOR2X1 _1330_ (
    .A(_560_),
    .B(_675_),
    .Y(_676_)
);

OAI21X1 _1331_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_684_[10]),
    .Y(_677_)
);

MUX2X1 _1332_ (
    .A(\internal_reg[1] [10]),
    .B(\internal_reg[0] [10]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_678_)
);

NOR2X1 _1333_ (
    .A(\internal_reg[3] [10]),
    .B(_562__bF$buf3),
    .Y(_679_)
);

OAI21X1 _1334_ (
    .A(\internal_reg[2] [10]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_680_)
);

OAI22X1 _1335_ (
    .A(_680_),
    .B(_679_),
    .C(rb_adrs_1_bF$buf4),
    .D(_678_),
    .Y(_681_)
);

OAI21X1 _1336_ (
    .A(rb_adrs_2_bF$buf0),
    .B(_681_),
    .C(_116__bF$buf4),
    .Y(_682_)
);

OAI21X1 _1337_ (
    .A(_676_),
    .B(_682_),
    .C(_677_),
    .Y(_1_[10])
);

MUX2X1 _1338_ (
    .A(\internal_reg[5] [11]),
    .B(\internal_reg[4] [11]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_2_)
);

NOR2X1 _1339_ (
    .A(\internal_reg[7] [11]),
    .B(_562__bF$buf2),
    .Y(_3_)
);

OAI21X1 _1340_ (
    .A(\internal_reg[6] [11]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_4_)
);

OAI22X1 _1341_ (
    .A(_4_),
    .B(_3_),
    .C(rb_adrs_1_bF$buf2),
    .D(_2_),
    .Y(_5_)
);

NOR2X1 _1342_ (
    .A(_560_),
    .B(_5_),
    .Y(_6_)
);

OAI21X1 _1343_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_684_[11]),
    .Y(_7_)
);

MUX2X1 _1344_ (
    .A(\internal_reg[1] [11]),
    .B(\internal_reg[0] [11]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_8_)
);

NOR2X1 _1345_ (
    .A(\internal_reg[3] [11]),
    .B(_562__bF$buf1),
    .Y(_9_)
);

OAI21X1 _1346_ (
    .A(\internal_reg[2] [11]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_10_)
);

OAI22X1 _1347_ (
    .A(_10_),
    .B(_9_),
    .C(rb_adrs_1_bF$buf0),
    .D(_8_),
    .Y(_11_)
);

OAI21X1 _1348_ (
    .A(rb_adrs_2_bF$buf3),
    .B(_11_),
    .C(_116__bF$buf3),
    .Y(_12_)
);

OAI21X1 _1349_ (
    .A(_6_),
    .B(_12_),
    .C(_7_),
    .Y(_1_[11])
);

MUX2X1 _1350_ (
    .A(\internal_reg[5] [12]),
    .B(\internal_reg[4] [12]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_13_)
);

NOR2X1 _1351_ (
    .A(\internal_reg[7] [12]),
    .B(_562__bF$buf0),
    .Y(_14_)
);

OAI21X1 _1352_ (
    .A(\internal_reg[6] [12]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_15_)
);

OAI22X1 _1353_ (
    .A(_15_),
    .B(_14_),
    .C(rb_adrs_1_bF$buf6),
    .D(_13_),
    .Y(_16_)
);

NOR2X1 _1354_ (
    .A(_560_),
    .B(_16_),
    .Y(_17_)
);

OAI21X1 _1355_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .C(_684_[12]),
    .Y(_18_)
);

MUX2X1 _1356_ (
    .A(\internal_reg[1] [12]),
    .B(\internal_reg[0] [12]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_19_)
);

NOR2X1 _1357_ (
    .A(\internal_reg[3] [12]),
    .B(_562__bF$buf4),
    .Y(_20_)
);

OAI21X1 _1358_ (
    .A(\internal_reg[2] [12]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_21_)
);

OAI22X1 _1359_ (
    .A(_21_),
    .B(_20_),
    .C(rb_adrs_1_bF$buf4),
    .D(_19_),
    .Y(_22_)
);

OAI21X1 _1360_ (
    .A(rb_adrs_2_bF$buf2),
    .B(_22_),
    .C(_116__bF$buf2),
    .Y(_23_)
);

OAI21X1 _1361_ (
    .A(_17_),
    .B(_23_),
    .C(_18_),
    .Y(_1_[12])
);

MUX2X1 _1362_ (
    .A(\internal_reg[5] [13]),
    .B(\internal_reg[4] [13]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_24_)
);

NOR2X1 _1363_ (
    .A(\internal_reg[7] [13]),
    .B(_562__bF$buf3),
    .Y(_25_)
);

OAI21X1 _1364_ (
    .A(\internal_reg[6] [13]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_26_)
);

OAI22X1 _1365_ (
    .A(_26_),
    .B(_25_),
    .C(rb_adrs_1_bF$buf2),
    .D(_24_),
    .Y(_27_)
);

NOR2X1 _1366_ (
    .A(_560_),
    .B(_27_),
    .Y(_28_)
);

OAI21X1 _1367_ (
    .A(wr_en_bF$buf1),
    .B(_104__bF$buf1),
    .C(_684_[13]),
    .Y(_29_)
);

MUX2X1 _1368_ (
    .A(\internal_reg[1] [13]),
    .B(\internal_reg[0] [13]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_30_)
);

NOR2X1 _1369_ (
    .A(\internal_reg[3] [13]),
    .B(_562__bF$buf2),
    .Y(_31_)
);

OAI21X1 _1370_ (
    .A(\internal_reg[2] [13]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_32_)
);

OAI22X1 _1371_ (
    .A(_32_),
    .B(_31_),
    .C(rb_adrs_1_bF$buf0),
    .D(_30_),
    .Y(_33_)
);

OAI21X1 _1372_ (
    .A(rb_adrs_2_bF$buf1),
    .B(_33_),
    .C(_116__bF$buf1),
    .Y(_34_)
);

OAI21X1 _1373_ (
    .A(_28_),
    .B(_34_),
    .C(_29_),
    .Y(_1_[13])
);

MUX2X1 _1374_ (
    .A(\internal_reg[5] [14]),
    .B(\internal_reg[4] [14]),
    .S(rb_adrs_0_bF$buf6),
    .Y(_35_)
);

NOR2X1 _1375_ (
    .A(\internal_reg[7] [14]),
    .B(_562__bF$buf1),
    .Y(_36_)
);

OAI21X1 _1376_ (
    .A(\internal_reg[6] [14]),
    .B(rb_adrs_0_bF$buf5),
    .C(rb_adrs_1_bF$buf7),
    .Y(_37_)
);

OAI22X1 _1377_ (
    .A(_37_),
    .B(_36_),
    .C(rb_adrs_1_bF$buf6),
    .D(_35_),
    .Y(_38_)
);

NOR2X1 _1378_ (
    .A(_560_),
    .B(_38_),
    .Y(_39_)
);

OAI21X1 _1379_ (
    .A(wr_en_bF$buf0),
    .B(_104__bF$buf0),
    .C(_684_[14]),
    .Y(_40_)
);

MUX2X1 _1380_ (
    .A(\internal_reg[1] [14]),
    .B(\internal_reg[0] [14]),
    .S(rb_adrs_0_bF$buf4),
    .Y(_41_)
);

NOR2X1 _1381_ (
    .A(\internal_reg[3] [14]),
    .B(_562__bF$buf0),
    .Y(_42_)
);

OAI21X1 _1382_ (
    .A(\internal_reg[2] [14]),
    .B(rb_adrs_0_bF$buf3),
    .C(rb_adrs_1_bF$buf5),
    .Y(_43_)
);

OAI22X1 _1383_ (
    .A(_43_),
    .B(_42_),
    .C(rb_adrs_1_bF$buf4),
    .D(_41_),
    .Y(_44_)
);

OAI21X1 _1384_ (
    .A(rb_adrs_2_bF$buf0),
    .B(_44_),
    .C(_116__bF$buf0),
    .Y(_45_)
);

OAI21X1 _1385_ (
    .A(_39_),
    .B(_45_),
    .C(_40_),
    .Y(_1_[14])
);

MUX2X1 _1386_ (
    .A(\internal_reg[5] [15]),
    .B(\internal_reg[4] [15]),
    .S(rb_adrs_0_bF$buf2),
    .Y(_46_)
);

NOR2X1 _1387_ (
    .A(\internal_reg[7] [15]),
    .B(_562__bF$buf4),
    .Y(_47_)
);

OAI21X1 _1388_ (
    .A(\internal_reg[6] [15]),
    .B(rb_adrs_0_bF$buf1),
    .C(rb_adrs_1_bF$buf3),
    .Y(_48_)
);

OAI22X1 _1389_ (
    .A(_48_),
    .B(_47_),
    .C(rb_adrs_1_bF$buf2),
    .D(_46_),
    .Y(_49_)
);

NOR2X1 _1390_ (
    .A(_560_),
    .B(_49_),
    .Y(_50_)
);

OAI21X1 _1391_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_684_[15]),
    .Y(_51_)
);

MUX2X1 _1392_ (
    .A(\internal_reg[1] [15]),
    .B(\internal_reg[0] [15]),
    .S(rb_adrs_0_bF$buf0),
    .Y(_52_)
);

NOR2X1 _1393_ (
    .A(\internal_reg[3] [15]),
    .B(_562__bF$buf3),
    .Y(_53_)
);

OAI21X1 _1394_ (
    .A(\internal_reg[2] [15]),
    .B(rb_adrs_0_bF$buf7),
    .C(rb_adrs_1_bF$buf1),
    .Y(_54_)
);

OAI22X1 _1395_ (
    .A(_54_),
    .B(_53_),
    .C(rb_adrs_1_bF$buf0),
    .D(_52_),
    .Y(_55_)
);

OAI21X1 _1396_ (
    .A(rb_adrs_2_bF$buf3),
    .B(_55_),
    .C(_116__bF$buf4),
    .Y(_56_)
);

OAI21X1 _1397_ (
    .A(_50_),
    .B(_56_),
    .C(_51_),
    .Y(_1_[15])
);

BUFX2 _1398_ (
    .A(_683_[0]),
    .Y(ra_out[0])
);

BUFX2 _1399_ (
    .A(_683_[1]),
    .Y(ra_out[1])
);

BUFX2 _1400_ (
    .A(_683_[2]),
    .Y(ra_out[2])
);

BUFX2 _1401_ (
    .A(_683_[3]),
    .Y(ra_out[3])
);

BUFX2 _1402_ (
    .A(_683_[4]),
    .Y(ra_out[4])
);

BUFX2 _1403_ (
    .A(_683_[5]),
    .Y(ra_out[5])
);

BUFX2 _1404_ (
    .A(_683_[6]),
    .Y(ra_out[6])
);

BUFX2 _1405_ (
    .A(_683_[7]),
    .Y(ra_out[7])
);

BUFX2 _1406_ (
    .A(_683_[8]),
    .Y(ra_out[8])
);

BUFX2 _1407_ (
    .A(_683_[9]),
    .Y(ra_out[9])
);

BUFX2 _1408_ (
    .A(_683_[10]),
    .Y(ra_out[10])
);

BUFX2 _1409_ (
    .A(_683_[11]),
    .Y(ra_out[11])
);

BUFX2 _1410_ (
    .A(_683_[12]),
    .Y(ra_out[12])
);

BUFX2 _1411_ (
    .A(_683_[13]),
    .Y(ra_out[13])
);

BUFX2 _1412_ (
    .A(_683_[14]),
    .Y(ra_out[14])
);

BUFX2 _1413_ (
    .A(_683_[15]),
    .Y(ra_out[15])
);

BUFX2 _1414_ (
    .A(_684_[0]),
    .Y(rb_out[0])
);

BUFX2 _1415_ (
    .A(_684_[1]),
    .Y(rb_out[1])
);

BUFX2 _1416_ (
    .A(_684_[2]),
    .Y(rb_out[2])
);

BUFX2 _1417_ (
    .A(_684_[3]),
    .Y(rb_out[3])
);

BUFX2 _1418_ (
    .A(_684_[4]),
    .Y(rb_out[4])
);

BUFX2 _1419_ (
    .A(_684_[5]),
    .Y(rb_out[5])
);

BUFX2 _1420_ (
    .A(_684_[6]),
    .Y(rb_out[6])
);

BUFX2 _1421_ (
    .A(_684_[7]),
    .Y(rb_out[7])
);

BUFX2 _1422_ (
    .A(_684_[8]),
    .Y(rb_out[8])
);

BUFX2 _1423_ (
    .A(_684_[9]),
    .Y(rb_out[9])
);

BUFX2 _1424_ (
    .A(_684_[10]),
    .Y(rb_out[10])
);

BUFX2 _1425_ (
    .A(_684_[11]),
    .Y(rb_out[11])
);

BUFX2 _1426_ (
    .A(_684_[12]),
    .Y(rb_out[12])
);

BUFX2 _1427_ (
    .A(_684_[13]),
    .Y(rb_out[13])
);

BUFX2 _1428_ (
    .A(_684_[14]),
    .Y(rb_out[14])
);

BUFX2 _1429_ (
    .A(_684_[15]),
    .Y(rb_out[15])
);

DFFPOSX1 _1430_ (
    .CLK(clock_bF$buf11),
    .D(_73_),
    .Q(\internal_reg[1] [0])
);

DFFPOSX1 _1431_ (
    .CLK(clock_bF$buf10),
    .D(_74_),
    .Q(\internal_reg[1] [1])
);

DFFPOSX1 _1432_ (
    .CLK(clock_bF$buf9),
    .D(_75_),
    .Q(\internal_reg[1] [2])
);

DFFPOSX1 _1433_ (
    .CLK(clock_bF$buf8),
    .D(_76_),
    .Q(\internal_reg[1] [3])
);

DFFPOSX1 _1434_ (
    .CLK(clock_bF$buf7),
    .D(_77_),
    .Q(\internal_reg[1] [4])
);

DFFPOSX1 _1435_ (
    .CLK(clock_bF$buf6),
    .D(_78_),
    .Q(\internal_reg[1] [5])
);

DFFPOSX1 _1436_ (
    .CLK(clock_bF$buf5),
    .D(_79_),
    .Q(\internal_reg[1] [6])
);

DFFPOSX1 _1437_ (
    .CLK(clock_bF$buf4),
    .D(_80_),
    .Q(\internal_reg[1] [7])
);

DFFPOSX1 _1438_ (
    .CLK(clock_bF$buf3),
    .D(_81_),
    .Q(\internal_reg[1] [8])
);

DFFPOSX1 _1439_ (
    .CLK(clock_bF$buf2),
    .D(_82_),
    .Q(\internal_reg[1] [9])
);

DFFPOSX1 _1440_ (
    .CLK(clock_bF$buf1),
    .D(_83_),
    .Q(\internal_reg[1] [10])
);

DFFPOSX1 _1441_ (
    .CLK(clock_bF$buf0),
    .D(_84_),
    .Q(\internal_reg[1] [11])
);

DFFPOSX1 _1442_ (
    .CLK(clock_bF$buf11),
    .D(_85_),
    .Q(\internal_reg[1] [12])
);

DFFPOSX1 _1443_ (
    .CLK(clock_bF$buf10),
    .D(_86_),
    .Q(\internal_reg[1] [13])
);

DFFPOSX1 _1444_ (
    .CLK(clock_bF$buf9),
    .D(_87_),
    .Q(\internal_reg[1] [14])
);

DFFPOSX1 _1445_ (
    .CLK(clock_bF$buf8),
    .D(_88_),
    .Q(\internal_reg[1] [15])
);

DFFPOSX1 _1446_ (
    .CLK(clock_bF$buf7),
    .D(_57_),
    .Q(\internal_reg[0] [0])
);

DFFPOSX1 _1447_ (
    .CLK(clock_bF$buf6),
    .D(_58_),
    .Q(\internal_reg[0] [1])
);

DFFPOSX1 _1448_ (
    .CLK(clock_bF$buf5),
    .D(_59_),
    .Q(\internal_reg[0] [2])
);

DFFPOSX1 _1449_ (
    .CLK(clock_bF$buf4),
    .D(_60_),
    .Q(\internal_reg[0] [3])
);

DFFPOSX1 _1450_ (
    .CLK(clock_bF$buf3),
    .D(_61_),
    .Q(\internal_reg[0] [4])
);

DFFPOSX1 _1451_ (
    .CLK(clock_bF$buf2),
    .D(_62_),
    .Q(\internal_reg[0] [5])
);

DFFPOSX1 _1452_ (
    .CLK(clock_bF$buf1),
    .D(_63_),
    .Q(\internal_reg[0] [6])
);

DFFPOSX1 _1453_ (
    .CLK(clock_bF$buf0),
    .D(_64_),
    .Q(\internal_reg[0] [7])
);

DFFPOSX1 _1454_ (
    .CLK(clock_bF$buf11),
    .D(_65_),
    .Q(\internal_reg[0] [8])
);

DFFPOSX1 _1455_ (
    .CLK(clock_bF$buf10),
    .D(_66_),
    .Q(\internal_reg[0] [9])
);

DFFPOSX1 _1456_ (
    .CLK(clock_bF$buf9),
    .D(_67_),
    .Q(\internal_reg[0] [10])
);

DFFPOSX1 _1457_ (
    .CLK(clock_bF$buf8),
    .D(_68_),
    .Q(\internal_reg[0] [11])
);

DFFPOSX1 _1458_ (
    .CLK(clock_bF$buf7),
    .D(_69_),
    .Q(\internal_reg[0] [12])
);

DFFPOSX1 _1459_ (
    .CLK(clock_bF$buf6),
    .D(_70_),
    .Q(\internal_reg[0] [13])
);

DFFPOSX1 _1460_ (
    .CLK(clock_bF$buf5),
    .D(_71_),
    .Q(\internal_reg[0] [14])
);

DFFPOSX1 _1461_ (
    .CLK(clock_bF$buf4),
    .D(_72_),
    .Q(\internal_reg[0] [15])
);

DFFPOSX1 _1462_ (
    .CLK(clock_bF$buf3),
    .D(_255_),
    .Q(\internal_reg[7] [0])
);

DFFPOSX1 _1463_ (
    .CLK(clock_bF$buf2),
    .D(_257_),
    .Q(\internal_reg[7] [1])
);

DFFPOSX1 _1464_ (
    .CLK(clock_bF$buf1),
    .D(_259_),
    .Q(\internal_reg[7] [2])
);

DFFPOSX1 _1465_ (
    .CLK(clock_bF$buf0),
    .D(_261_),
    .Q(\internal_reg[7] [3])
);

DFFPOSX1 _1466_ (
    .CLK(clock_bF$buf11),
    .D(_263_),
    .Q(\internal_reg[7] [4])
);

DFFPOSX1 _1467_ (
    .CLK(clock_bF$buf10),
    .D(_265_),
    .Q(\internal_reg[7] [5])
);

DFFPOSX1 _1468_ (
    .CLK(clock_bF$buf9),
    .D(_267_),
    .Q(\internal_reg[7] [6])
);

DFFPOSX1 _1469_ (
    .CLK(clock_bF$buf8),
    .D(_268_),
    .Q(\internal_reg[7] [7])
);

DFFPOSX1 _1470_ (
    .CLK(clock_bF$buf7),
    .D(_270_),
    .Q(\internal_reg[7] [8])
);

DFFPOSX1 _1471_ (
    .CLK(clock_bF$buf6),
    .D(_272_),
    .Q(\internal_reg[7] [9])
);

DFFPOSX1 _1472_ (
    .CLK(clock_bF$buf5),
    .D(_274_),
    .Q(\internal_reg[7] [10])
);

DFFPOSX1 _1473_ (
    .CLK(clock_bF$buf4),
    .D(_276_),
    .Q(\internal_reg[7] [11])
);

DFFPOSX1 _1474_ (
    .CLK(clock_bF$buf3),
    .D(_278_),
    .Q(\internal_reg[7] [12])
);

DFFPOSX1 _1475_ (
    .CLK(clock_bF$buf2),
    .D(_280_),
    .Q(\internal_reg[7] [13])
);

DFFPOSX1 _1476_ (
    .CLK(clock_bF$buf1),
    .D(_282_),
    .Q(\internal_reg[7] [14])
);

DFFPOSX1 _1477_ (
    .CLK(clock_bF$buf0),
    .D(_284_),
    .Q(\internal_reg[7] [15])
);

DFFPOSX1 _1478_ (
    .CLK(clock_bF$buf11),
    .D(_223_),
    .Q(\internal_reg[6] [0])
);

DFFPOSX1 _1479_ (
    .CLK(clock_bF$buf10),
    .D(_224_),
    .Q(\internal_reg[6] [1])
);

DFFPOSX1 _1480_ (
    .CLK(clock_bF$buf9),
    .D(_226_),
    .Q(\internal_reg[6] [2])
);

DFFPOSX1 _1481_ (
    .CLK(clock_bF$buf8),
    .D(_228_),
    .Q(\internal_reg[6] [3])
);

DFFPOSX1 _1482_ (
    .CLK(clock_bF$buf7),
    .D(_230_),
    .Q(\internal_reg[6] [4])
);

DFFPOSX1 _1483_ (
    .CLK(clock_bF$buf6),
    .D(_232_),
    .Q(\internal_reg[6] [5])
);

DFFPOSX1 _1484_ (
    .CLK(clock_bF$buf5),
    .D(_234_),
    .Q(\internal_reg[6] [6])
);

DFFPOSX1 _1485_ (
    .CLK(clock_bF$buf4),
    .D(_236_),
    .Q(\internal_reg[6] [7])
);

DFFPOSX1 _1486_ (
    .CLK(clock_bF$buf3),
    .D(_238_),
    .Q(\internal_reg[6] [8])
);

DFFPOSX1 _1487_ (
    .CLK(clock_bF$buf2),
    .D(_240_),
    .Q(\internal_reg[6] [9])
);

DFFPOSX1 _1488_ (
    .CLK(clock_bF$buf1),
    .D(_242_),
    .Q(\internal_reg[6] [10])
);

DFFPOSX1 _1489_ (
    .CLK(clock_bF$buf0),
    .D(_244_),
    .Q(\internal_reg[6] [11])
);

DFFPOSX1 _1490_ (
    .CLK(clock_bF$buf11),
    .D(_246_),
    .Q(\internal_reg[6] [12])
);

DFFPOSX1 _1491_ (
    .CLK(clock_bF$buf10),
    .D(_247_),
    .Q(\internal_reg[6] [13])
);

DFFPOSX1 _1492_ (
    .CLK(clock_bF$buf9),
    .D(_249_),
    .Q(\internal_reg[6] [14])
);

DFFPOSX1 _1493_ (
    .CLK(clock_bF$buf8),
    .D(_251_),
    .Q(\internal_reg[6] [15])
);

DFFPOSX1 _1494_ (
    .CLK(clock_bF$buf7),
    .D(_89_),
    .Q(\internal_reg[2] [0])
);

DFFPOSX1 _1495_ (
    .CLK(clock_bF$buf6),
    .D(_91_),
    .Q(\internal_reg[2] [1])
);

DFFPOSX1 _1496_ (
    .CLK(clock_bF$buf5),
    .D(_93_),
    .Q(\internal_reg[2] [2])
);

DFFPOSX1 _1497_ (
    .CLK(clock_bF$buf4),
    .D(_95_),
    .Q(\internal_reg[2] [3])
);

DFFPOSX1 _1498_ (
    .CLK(clock_bF$buf3),
    .D(_97_),
    .Q(\internal_reg[2] [4])
);

DFFPOSX1 _1499_ (
    .CLK(clock_bF$buf2),
    .D(_99_),
    .Q(\internal_reg[2] [5])
);

DFFPOSX1 _1500_ (
    .CLK(clock_bF$buf1),
    .D(_101_),
    .Q(\internal_reg[2] [6])
);

DFFPOSX1 _1501_ (
    .CLK(clock_bF$buf0),
    .D(_103_),
    .Q(\internal_reg[2] [7])
);

DFFPOSX1 _1502_ (
    .CLK(clock_bF$buf11),
    .D(_105_),
    .Q(\internal_reg[2] [8])
);

DFFPOSX1 _1503_ (
    .CLK(clock_bF$buf10),
    .D(_107_),
    .Q(\internal_reg[2] [9])
);

DFFPOSX1 _1504_ (
    .CLK(clock_bF$buf9),
    .D(_109_),
    .Q(\internal_reg[2] [10])
);

DFFPOSX1 _1505_ (
    .CLK(clock_bF$buf8),
    .D(_111_),
    .Q(\internal_reg[2] [11])
);

DFFPOSX1 _1506_ (
    .CLK(clock_bF$buf7),
    .D(_113_),
    .Q(\internal_reg[2] [12])
);

DFFPOSX1 _1507_ (
    .CLK(clock_bF$buf6),
    .D(_115_),
    .Q(\internal_reg[2] [13])
);

DFFPOSX1 _1508_ (
    .CLK(clock_bF$buf5),
    .D(_117_),
    .Q(\internal_reg[2] [14])
);

DFFPOSX1 _1509_ (
    .CLK(clock_bF$buf4),
    .D(_119_),
    .Q(\internal_reg[2] [15])
);

DFFPOSX1 _1510_ (
    .CLK(clock_bF$buf3),
    .D(_189_),
    .Q(\internal_reg[5] [0])
);

DFFPOSX1 _1511_ (
    .CLK(clock_bF$buf2),
    .D(_191_),
    .Q(\internal_reg[5] [1])
);

DFFPOSX1 _1512_ (
    .CLK(clock_bF$buf1),
    .D(_193_),
    .Q(\internal_reg[5] [2])
);

DFFPOSX1 _1513_ (
    .CLK(clock_bF$buf0),
    .D(_195_),
    .Q(\internal_reg[5] [3])
);

DFFPOSX1 _1514_ (
    .CLK(clock_bF$buf11),
    .D(_197_),
    .Q(\internal_reg[5] [4])
);

DFFPOSX1 _1515_ (
    .CLK(clock_bF$buf10),
    .D(_199_),
    .Q(\internal_reg[5] [5])
);

DFFPOSX1 _1516_ (
    .CLK(clock_bF$buf9),
    .D(_201_),
    .Q(\internal_reg[5] [6])
);

DFFPOSX1 _1517_ (
    .CLK(clock_bF$buf8),
    .D(_203_),
    .Q(\internal_reg[5] [7])
);

DFFPOSX1 _1518_ (
    .CLK(clock_bF$buf7),
    .D(_204_),
    .Q(\internal_reg[5] [8])
);

DFFPOSX1 _1519_ (
    .CLK(clock_bF$buf6),
    .D(_206_),
    .Q(\internal_reg[5] [9])
);

DFFPOSX1 _1520_ (
    .CLK(clock_bF$buf5),
    .D(_208_),
    .Q(\internal_reg[5] [10])
);

DFFPOSX1 _1521_ (
    .CLK(clock_bF$buf4),
    .D(_210_),
    .Q(\internal_reg[5] [11])
);

DFFPOSX1 _1522_ (
    .CLK(clock_bF$buf3),
    .D(_212_),
    .Q(\internal_reg[5] [12])
);

DFFPOSX1 _1523_ (
    .CLK(clock_bF$buf2),
    .D(_214_),
    .Q(\internal_reg[5] [13])
);

DFFPOSX1 _1524_ (
    .CLK(clock_bF$buf1),
    .D(_216_),
    .Q(\internal_reg[5] [14])
);

DFFPOSX1 _1525_ (
    .CLK(clock_bF$buf0),
    .D(_218_),
    .Q(\internal_reg[5] [15])
);

DFFPOSX1 _1526_ (
    .CLK(clock_bF$buf11),
    .D(_157_),
    .Q(\internal_reg[4] [0])
);

DFFPOSX1 _1527_ (
    .CLK(clock_bF$buf10),
    .D(_159_),
    .Q(\internal_reg[4] [1])
);

DFFPOSX1 _1528_ (
    .CLK(clock_bF$buf9),
    .D(_160_),
    .Q(\internal_reg[4] [2])
);

DFFPOSX1 _1529_ (
    .CLK(clock_bF$buf8),
    .D(_162_),
    .Q(\internal_reg[4] [3])
);

DFFPOSX1 _1530_ (
    .CLK(clock_bF$buf7),
    .D(_164_),
    .Q(\internal_reg[4] [4])
);

DFFPOSX1 _1531_ (
    .CLK(clock_bF$buf6),
    .D(_166_),
    .Q(\internal_reg[4] [5])
);

DFFPOSX1 _1532_ (
    .CLK(clock_bF$buf5),
    .D(_168_),
    .Q(\internal_reg[4] [6])
);

DFFPOSX1 _1533_ (
    .CLK(clock_bF$buf4),
    .D(_170_),
    .Q(\internal_reg[4] [7])
);

DFFPOSX1 _1534_ (
    .CLK(clock_bF$buf3),
    .D(_172_),
    .Q(\internal_reg[4] [8])
);

DFFPOSX1 _1535_ (
    .CLK(clock_bF$buf2),
    .D(_174_),
    .Q(\internal_reg[4] [9])
);

DFFPOSX1 _1536_ (
    .CLK(clock_bF$buf1),
    .D(_176_),
    .Q(\internal_reg[4] [10])
);

DFFPOSX1 _1537_ (
    .CLK(clock_bF$buf0),
    .D(_178_),
    .Q(\internal_reg[4] [11])
);

DFFPOSX1 _1538_ (
    .CLK(clock_bF$buf11),
    .D(_180_),
    .Q(\internal_reg[4] [12])
);

DFFPOSX1 _1539_ (
    .CLK(clock_bF$buf10),
    .D(_182_),
    .Q(\internal_reg[4] [13])
);

DFFPOSX1 _1540_ (
    .CLK(clock_bF$buf9),
    .D(_183_),
    .Q(\internal_reg[4] [14])
);

DFFPOSX1 _1541_ (
    .CLK(clock_bF$buf8),
    .D(_185_),
    .Q(\internal_reg[4] [15])
);

DFFPOSX1 _1542_ (
    .CLK(clock_bF$buf7),
    .D(_123_),
    .Q(\internal_reg[3] [0])
);

DFFPOSX1 _1543_ (
    .CLK(clock_bF$buf6),
    .D(_125_),
    .Q(\internal_reg[3] [1])
);

DFFPOSX1 _1544_ (
    .CLK(clock_bF$buf5),
    .D(_127_),
    .Q(\internal_reg[3] [2])
);

DFFPOSX1 _1545_ (
    .CLK(clock_bF$buf4),
    .D(_129_),
    .Q(\internal_reg[3] [3])
);

DFFPOSX1 _1546_ (
    .CLK(clock_bF$buf3),
    .D(_131_),
    .Q(\internal_reg[3] [4])
);

DFFPOSX1 _1547_ (
    .CLK(clock_bF$buf2),
    .D(_133_),
    .Q(\internal_reg[3] [5])
);

DFFPOSX1 _1548_ (
    .CLK(clock_bF$buf1),
    .D(_135_),
    .Q(\internal_reg[3] [6])
);

DFFPOSX1 _1549_ (
    .CLK(clock_bF$buf0),
    .D(_137_),
    .Q(\internal_reg[3] [7])
);

DFFPOSX1 _1550_ (
    .CLK(clock_bF$buf11),
    .D(_139_),
    .Q(\internal_reg[3] [8])
);

DFFPOSX1 _1551_ (
    .CLK(clock_bF$buf10),
    .D(_140_),
    .Q(\internal_reg[3] [9])
);

DFFPOSX1 _1552_ (
    .CLK(clock_bF$buf9),
    .D(_142_),
    .Q(\internal_reg[3] [10])
);

DFFPOSX1 _1553_ (
    .CLK(clock_bF$buf8),
    .D(_144_),
    .Q(\internal_reg[3] [11])
);

DFFPOSX1 _1554_ (
    .CLK(clock_bF$buf7),
    .D(_146_),
    .Q(\internal_reg[3] [12])
);

DFFPOSX1 _1555_ (
    .CLK(clock_bF$buf6),
    .D(_148_),
    .Q(\internal_reg[3] [13])
);

DFFPOSX1 _1556_ (
    .CLK(clock_bF$buf5),
    .D(_150_),
    .Q(\internal_reg[3] [14])
);

DFFPOSX1 _1557_ (
    .CLK(clock_bF$buf4),
    .D(_152_),
    .Q(\internal_reg[3] [15])
);

DFFPOSX1 _1558_ (
    .CLK(clock_bF$buf3),
    .D(_1_[0]),
    .Q(_684_[0])
);

DFFPOSX1 _1559_ (
    .CLK(clock_bF$buf2),
    .D(_1_[1]),
    .Q(_684_[1])
);

DFFPOSX1 _1560_ (
    .CLK(clock_bF$buf1),
    .D(_1_[2]),
    .Q(_684_[2])
);

DFFPOSX1 _1561_ (
    .CLK(clock_bF$buf0),
    .D(_1_[3]),
    .Q(_684_[3])
);

DFFPOSX1 _1562_ (
    .CLK(clock_bF$buf11),
    .D(_1_[4]),
    .Q(_684_[4])
);

DFFPOSX1 _1563_ (
    .CLK(clock_bF$buf10),
    .D(_1_[5]),
    .Q(_684_[5])
);

DFFPOSX1 _1564_ (
    .CLK(clock_bF$buf9),
    .D(_1_[6]),
    .Q(_684_[6])
);

DFFPOSX1 _1565_ (
    .CLK(clock_bF$buf8),
    .D(_1_[7]),
    .Q(_684_[7])
);

DFFPOSX1 _1566_ (
    .CLK(clock_bF$buf7),
    .D(_1_[8]),
    .Q(_684_[8])
);

DFFPOSX1 _1567_ (
    .CLK(clock_bF$buf6),
    .D(_1_[9]),
    .Q(_684_[9])
);

DFFPOSX1 _1568_ (
    .CLK(clock_bF$buf5),
    .D(_1_[10]),
    .Q(_684_[10])
);

DFFPOSX1 _1569_ (
    .CLK(clock_bF$buf4),
    .D(_1_[11]),
    .Q(_684_[11])
);

DFFPOSX1 _1570_ (
    .CLK(clock_bF$buf3),
    .D(_1_[12]),
    .Q(_684_[12])
);

DFFPOSX1 _1571_ (
    .CLK(clock_bF$buf2),
    .D(_1_[13]),
    .Q(_684_[13])
);

DFFPOSX1 _1572_ (
    .CLK(clock_bF$buf1),
    .D(_1_[14]),
    .Q(_684_[14])
);

DFFPOSX1 _1573_ (
    .CLK(clock_bF$buf0),
    .D(_1_[15]),
    .Q(_684_[15])
);

DFFPOSX1 _1574_ (
    .CLK(clock_bF$buf11),
    .D(_0_[0]),
    .Q(_683_[0])
);

DFFPOSX1 _1575_ (
    .CLK(clock_bF$buf10),
    .D(_0_[1]),
    .Q(_683_[1])
);

DFFPOSX1 _1576_ (
    .CLK(clock_bF$buf9),
    .D(_0_[2]),
    .Q(_683_[2])
);

DFFPOSX1 _1577_ (
    .CLK(clock_bF$buf8),
    .D(_0_[3]),
    .Q(_683_[3])
);

DFFPOSX1 _1578_ (
    .CLK(clock_bF$buf7),
    .D(_0_[4]),
    .Q(_683_[4])
);

DFFPOSX1 _1579_ (
    .CLK(clock_bF$buf6),
    .D(_0_[5]),
    .Q(_683_[5])
);

DFFPOSX1 _1580_ (
    .CLK(clock_bF$buf5),
    .D(_0_[6]),
    .Q(_683_[6])
);

DFFPOSX1 _1581_ (
    .CLK(clock_bF$buf4),
    .D(_0_[7]),
    .Q(_683_[7])
);

DFFPOSX1 _1582_ (
    .CLK(clock_bF$buf3),
    .D(_0_[8]),
    .Q(_683_[8])
);

DFFPOSX1 _1583_ (
    .CLK(clock_bF$buf2),
    .D(_0_[9]),
    .Q(_683_[9])
);

DFFPOSX1 _1584_ (
    .CLK(clock_bF$buf1),
    .D(_0_[10]),
    .Q(_683_[10])
);

DFFPOSX1 _1585_ (
    .CLK(clock_bF$buf0),
    .D(_0_[11]),
    .Q(_683_[11])
);

DFFPOSX1 _1586_ (
    .CLK(clock_bF$buf11),
    .D(_0_[12]),
    .Q(_683_[12])
);

DFFPOSX1 _1587_ (
    .CLK(clock_bF$buf10),
    .D(_0_[13]),
    .Q(_683_[13])
);

DFFPOSX1 _1588_ (
    .CLK(clock_bF$buf9),
    .D(_0_[14]),
    .Q(_683_[14])
);

DFFPOSX1 _1589_ (
    .CLK(clock_bF$buf8),
    .D(_0_[15]),
    .Q(_683_[15])
);

INVX4 _685_ (
    .A(ra_adrs_2_bF$buf3),
    .Y(_90_)
);

MUX2X1 _686_ (
    .A(\internal_reg[5] [0]),
    .B(\internal_reg[4] [0]),
    .S(ra_adrs_0_bF$buf7),
    .Y(_92_)
);

INVX8 _687_ (
    .A(ra_adrs_0_bF$buf6),
    .Y(_94_)
);

NOR2X1 _688_ (
    .A(\internal_reg[7] [0]),
    .B(_94__bF$buf4),
    .Y(_96_)
);

OAI21X1 _689_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [0]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_98_)
);

OAI22X1 _690_ (
    .A(_98_),
    .B(_96_),
    .C(ra_adrs_1_bF$buf6),
    .D(_92_),
    .Y(_100_)
);

NOR2X1 _691_ (
    .A(_90_),
    .B(_100_),
    .Y(_102_)
);

INVX8 _692_ (
    .A(enable),
    .Y(_104_)
);

OAI21X1 _693_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_683_[0]),
    .Y(_106_)
);

MUX2X1 _694_ (
    .A(\internal_reg[1] [0]),
    .B(\internal_reg[0] [0]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_108_)
);

NOR2X1 _695_ (
    .A(\internal_reg[3] [0]),
    .B(_94__bF$buf3),
    .Y(_110_)
);

OAI21X1 _696_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [0]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_112_)
);

OAI22X1 _697_ (
    .A(_112_),
    .B(_110_),
    .C(ra_adrs_1_bF$buf4),
    .D(_108_),
    .Y(_114_)
);

NOR2X1 _698_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .Y(_116_)
);

OAI21X1 _699_ (
    .A(ra_adrs_2_bF$buf2),
    .B(_114_),
    .C(_116__bF$buf3),
    .Y(_118_)
);

OAI21X1 _700_ (
    .A(_102_),
    .B(_118_),
    .C(_106_),
    .Y(_0_[0])
);

MUX2X1 _701_ (
    .A(\internal_reg[5] [1]),
    .B(\internal_reg[4] [1]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_120_)
);

NOR2X1 _702_ (
    .A(\internal_reg[7] [1]),
    .B(_94__bF$buf2),
    .Y(_121_)
);

OAI21X1 _703_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [1]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_122_)
);

OAI22X1 _704_ (
    .A(_122_),
    .B(_121_),
    .C(ra_adrs_1_bF$buf2),
    .D(_120_),
    .Y(_124_)
);

NOR2X1 _705_ (
    .A(_90_),
    .B(_124_),
    .Y(_126_)
);

OAI21X1 _706_ (
    .A(wr_en_bF$buf1),
    .B(_104__bF$buf1),
    .C(_683_[1]),
    .Y(_128_)
);

MUX2X1 _707_ (
    .A(\internal_reg[1] [1]),
    .B(\internal_reg[0] [1]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_130_)
);

NOR2X1 _708_ (
    .A(\internal_reg[3] [1]),
    .B(_94__bF$buf1),
    .Y(_132_)
);

OAI21X1 _709_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [1]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_134_)
);

OAI22X1 _710_ (
    .A(_134_),
    .B(_132_),
    .C(ra_adrs_1_bF$buf0),
    .D(_130_),
    .Y(_136_)
);

OAI21X1 _711_ (
    .A(ra_adrs_2_bF$buf1),
    .B(_136_),
    .C(_116__bF$buf2),
    .Y(_138_)
);

OAI21X1 _712_ (
    .A(_126_),
    .B(_138_),
    .C(_128_),
    .Y(_0_[1])
);

MUX2X1 _713_ (
    .A(\internal_reg[5] [2]),
    .B(\internal_reg[4] [2]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_141_)
);

NOR2X1 _714_ (
    .A(\internal_reg[7] [2]),
    .B(_94__bF$buf0),
    .Y(_143_)
);

OAI21X1 _715_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [2]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_145_)
);

OAI22X1 _716_ (
    .A(_145_),
    .B(_143_),
    .C(ra_adrs_1_bF$buf6),
    .D(_141_),
    .Y(_147_)
);

NOR2X1 _717_ (
    .A(_90_),
    .B(_147_),
    .Y(_149_)
);

OAI21X1 _718_ (
    .A(wr_en_bF$buf0),
    .B(_104__bF$buf0),
    .C(_683_[2]),
    .Y(_151_)
);

MUX2X1 _719_ (
    .A(\internal_reg[1] [2]),
    .B(\internal_reg[0] [2]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_153_)
);

NOR2X1 _720_ (
    .A(\internal_reg[3] [2]),
    .B(_94__bF$buf4),
    .Y(_154_)
);

OAI21X1 _721_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [2]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_155_)
);

OAI22X1 _722_ (
    .A(_155_),
    .B(_154_),
    .C(ra_adrs_1_bF$buf4),
    .D(_153_),
    .Y(_156_)
);

OAI21X1 _723_ (
    .A(ra_adrs_2_bF$buf0),
    .B(_156_),
    .C(_116__bF$buf1),
    .Y(_158_)
);

OAI21X1 _724_ (
    .A(_149_),
    .B(_158_),
    .C(_151_),
    .Y(_0_[2])
);

MUX2X1 _725_ (
    .A(\internal_reg[5] [3]),
    .B(\internal_reg[4] [3]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_161_)
);

NOR2X1 _726_ (
    .A(\internal_reg[7] [3]),
    .B(_94__bF$buf3),
    .Y(_163_)
);

OAI21X1 _727_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [3]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_165_)
);

OAI22X1 _728_ (
    .A(_165_),
    .B(_163_),
    .C(ra_adrs_1_bF$buf2),
    .D(_161_),
    .Y(_167_)
);

NOR2X1 _729_ (
    .A(_90_),
    .B(_167_),
    .Y(_169_)
);

OAI21X1 _730_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_683_[3]),
    .Y(_171_)
);

MUX2X1 _731_ (
    .A(\internal_reg[1] [3]),
    .B(\internal_reg[0] [3]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_173_)
);

NOR2X1 _732_ (
    .A(\internal_reg[3] [3]),
    .B(_94__bF$buf2),
    .Y(_175_)
);

OAI21X1 _733_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [3]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_177_)
);

OAI22X1 _734_ (
    .A(_177_),
    .B(_175_),
    .C(ra_adrs_1_bF$buf0),
    .D(_173_),
    .Y(_179_)
);

OAI21X1 _735_ (
    .A(ra_adrs_2_bF$buf3),
    .B(_179_),
    .C(_116__bF$buf0),
    .Y(_181_)
);

OAI21X1 _736_ (
    .A(_169_),
    .B(_181_),
    .C(_171_),
    .Y(_0_[3])
);

MUX2X1 _737_ (
    .A(\internal_reg[5] [4]),
    .B(\internal_reg[4] [4]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_184_)
);

NOR2X1 _738_ (
    .A(\internal_reg[7] [4]),
    .B(_94__bF$buf1),
    .Y(_186_)
);

OAI21X1 _739_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [4]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_187_)
);

OAI22X1 _740_ (
    .A(_187_),
    .B(_186_),
    .C(ra_adrs_1_bF$buf6),
    .D(_184_),
    .Y(_188_)
);

NOR2X1 _741_ (
    .A(_90_),
    .B(_188_),
    .Y(_190_)
);

OAI21X1 _742_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_683_[4]),
    .Y(_192_)
);

MUX2X1 _743_ (
    .A(\internal_reg[1] [4]),
    .B(\internal_reg[0] [4]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_194_)
);

NOR2X1 _744_ (
    .A(\internal_reg[3] [4]),
    .B(_94__bF$buf0),
    .Y(_196_)
);

OAI21X1 _745_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [4]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_198_)
);

OAI22X1 _746_ (
    .A(_198_),
    .B(_196_),
    .C(ra_adrs_1_bF$buf4),
    .D(_194_),
    .Y(_200_)
);

OAI21X1 _747_ (
    .A(ra_adrs_2_bF$buf2),
    .B(_200_),
    .C(_116__bF$buf4),
    .Y(_202_)
);

OAI21X1 _748_ (
    .A(_190_),
    .B(_202_),
    .C(_192_),
    .Y(_0_[4])
);

MUX2X1 _749_ (
    .A(\internal_reg[5] [5]),
    .B(\internal_reg[4] [5]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_205_)
);

NOR2X1 _750_ (
    .A(\internal_reg[7] [5]),
    .B(_94__bF$buf4),
    .Y(_207_)
);

OAI21X1 _751_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [5]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_209_)
);

OAI22X1 _752_ (
    .A(_209_),
    .B(_207_),
    .C(ra_adrs_1_bF$buf2),
    .D(_205_),
    .Y(_211_)
);

NOR2X1 _753_ (
    .A(_90_),
    .B(_211_),
    .Y(_213_)
);

OAI21X1 _754_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .C(_683_[5]),
    .Y(_215_)
);

MUX2X1 _755_ (
    .A(\internal_reg[1] [5]),
    .B(\internal_reg[0] [5]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_217_)
);

NOR2X1 _756_ (
    .A(\internal_reg[3] [5]),
    .B(_94__bF$buf3),
    .Y(_219_)
);

OAI21X1 _757_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [5]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_220_)
);

OAI22X1 _758_ (
    .A(_220_),
    .B(_219_),
    .C(ra_adrs_1_bF$buf0),
    .D(_217_),
    .Y(_221_)
);

OAI21X1 _759_ (
    .A(ra_adrs_2_bF$buf1),
    .B(_221_),
    .C(_116__bF$buf3),
    .Y(_222_)
);

OAI21X1 _760_ (
    .A(_213_),
    .B(_222_),
    .C(_215_),
    .Y(_0_[5])
);

MUX2X1 _761_ (
    .A(\internal_reg[5] [6]),
    .B(\internal_reg[4] [6]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_225_)
);

NOR2X1 _762_ (
    .A(\internal_reg[7] [6]),
    .B(_94__bF$buf2),
    .Y(_227_)
);

OAI21X1 _763_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [6]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_229_)
);

OAI22X1 _764_ (
    .A(_229_),
    .B(_227_),
    .C(ra_adrs_1_bF$buf6),
    .D(_225_),
    .Y(_231_)
);

NOR2X1 _765_ (
    .A(_90_),
    .B(_231_),
    .Y(_233_)
);

OAI21X1 _766_ (
    .A(wr_en_bF$buf1),
    .B(_104__bF$buf1),
    .C(_683_[6]),
    .Y(_235_)
);

MUX2X1 _767_ (
    .A(\internal_reg[1] [6]),
    .B(\internal_reg[0] [6]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_237_)
);

NOR2X1 _768_ (
    .A(\internal_reg[3] [6]),
    .B(_94__bF$buf1),
    .Y(_239_)
);

OAI21X1 _769_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [6]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_241_)
);

OAI22X1 _770_ (
    .A(_241_),
    .B(_239_),
    .C(ra_adrs_1_bF$buf4),
    .D(_237_),
    .Y(_243_)
);

OAI21X1 _771_ (
    .A(ra_adrs_2_bF$buf0),
    .B(_243_),
    .C(_116__bF$buf2),
    .Y(_245_)
);

OAI21X1 _772_ (
    .A(_233_),
    .B(_245_),
    .C(_235_),
    .Y(_0_[6])
);

MUX2X1 _773_ (
    .A(\internal_reg[5] [7]),
    .B(\internal_reg[4] [7]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_248_)
);

NOR2X1 _774_ (
    .A(\internal_reg[7] [7]),
    .B(_94__bF$buf0),
    .Y(_250_)
);

OAI21X1 _775_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [7]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_252_)
);

OAI22X1 _776_ (
    .A(_252_),
    .B(_250_),
    .C(ra_adrs_1_bF$buf2),
    .D(_248_),
    .Y(_253_)
);

NOR2X1 _777_ (
    .A(_90_),
    .B(_253_),
    .Y(_254_)
);

OAI21X1 _778_ (
    .A(wr_en_bF$buf0),
    .B(_104__bF$buf0),
    .C(_683_[7]),
    .Y(_256_)
);

MUX2X1 _779_ (
    .A(\internal_reg[1] [7]),
    .B(\internal_reg[0] [7]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_258_)
);

NOR2X1 _780_ (
    .A(\internal_reg[3] [7]),
    .B(_94__bF$buf4),
    .Y(_260_)
);

OAI21X1 _781_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [7]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_262_)
);

OAI22X1 _782_ (
    .A(_262_),
    .B(_260_),
    .C(ra_adrs_1_bF$buf0),
    .D(_258_),
    .Y(_264_)
);

OAI21X1 _783_ (
    .A(ra_adrs_2_bF$buf3),
    .B(_264_),
    .C(_116__bF$buf1),
    .Y(_266_)
);

OAI21X1 _784_ (
    .A(_254_),
    .B(_266_),
    .C(_256_),
    .Y(_0_[7])
);

MUX2X1 _785_ (
    .A(\internal_reg[5] [8]),
    .B(\internal_reg[4] [8]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_269_)
);

NOR2X1 _786_ (
    .A(\internal_reg[7] [8]),
    .B(_94__bF$buf3),
    .Y(_271_)
);

OAI21X1 _787_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [8]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_273_)
);

OAI22X1 _788_ (
    .A(_273_),
    .B(_271_),
    .C(ra_adrs_1_bF$buf6),
    .D(_269_),
    .Y(_275_)
);

NOR2X1 _789_ (
    .A(_90_),
    .B(_275_),
    .Y(_277_)
);

OAI21X1 _790_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_683_[8]),
    .Y(_279_)
);

MUX2X1 _791_ (
    .A(\internal_reg[1] [8]),
    .B(\internal_reg[0] [8]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_281_)
);

NOR2X1 _792_ (
    .A(\internal_reg[3] [8]),
    .B(_94__bF$buf2),
    .Y(_283_)
);

OAI21X1 _793_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [8]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_285_)
);

OAI22X1 _794_ (
    .A(_285_),
    .B(_283_),
    .C(ra_adrs_1_bF$buf4),
    .D(_281_),
    .Y(_286_)
);

OAI21X1 _795_ (
    .A(ra_adrs_2_bF$buf2),
    .B(_286_),
    .C(_116__bF$buf0),
    .Y(_287_)
);

OAI21X1 _796_ (
    .A(_277_),
    .B(_287_),
    .C(_279_),
    .Y(_0_[8])
);

MUX2X1 _797_ (
    .A(\internal_reg[5] [9]),
    .B(\internal_reg[4] [9]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_288_)
);

NOR2X1 _798_ (
    .A(\internal_reg[7] [9]),
    .B(_94__bF$buf1),
    .Y(_289_)
);

OAI21X1 _799_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [9]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_290_)
);

OAI22X1 _800_ (
    .A(_290_),
    .B(_289_),
    .C(ra_adrs_1_bF$buf2),
    .D(_288_),
    .Y(_291_)
);

NOR2X1 _801_ (
    .A(_90_),
    .B(_291_),
    .Y(_292_)
);

OAI21X1 _802_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_683_[9]),
    .Y(_293_)
);

MUX2X1 _803_ (
    .A(\internal_reg[1] [9]),
    .B(\internal_reg[0] [9]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_294_)
);

NOR2X1 _804_ (
    .A(\internal_reg[3] [9]),
    .B(_94__bF$buf0),
    .Y(_295_)
);

OAI21X1 _805_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [9]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_296_)
);

OAI22X1 _806_ (
    .A(_296_),
    .B(_295_),
    .C(ra_adrs_1_bF$buf0),
    .D(_294_),
    .Y(_297_)
);

OAI21X1 _807_ (
    .A(ra_adrs_2_bF$buf1),
    .B(_297_),
    .C(_116__bF$buf4),
    .Y(_298_)
);

OAI21X1 _808_ (
    .A(_292_),
    .B(_298_),
    .C(_293_),
    .Y(_0_[9])
);

MUX2X1 _809_ (
    .A(\internal_reg[5] [10]),
    .B(\internal_reg[4] [10]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_299_)
);

NOR2X1 _810_ (
    .A(\internal_reg[7] [10]),
    .B(_94__bF$buf4),
    .Y(_300_)
);

OAI21X1 _811_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [10]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_301_)
);

OAI22X1 _812_ (
    .A(_301_),
    .B(_300_),
    .C(ra_adrs_1_bF$buf6),
    .D(_299_),
    .Y(_302_)
);

NOR2X1 _813_ (
    .A(_90_),
    .B(_302_),
    .Y(_303_)
);

OAI21X1 _814_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .C(_683_[10]),
    .Y(_304_)
);

MUX2X1 _815_ (
    .A(\internal_reg[1] [10]),
    .B(\internal_reg[0] [10]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_305_)
);

NOR2X1 _816_ (
    .A(\internal_reg[3] [10]),
    .B(_94__bF$buf3),
    .Y(_306_)
);

OAI21X1 _817_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [10]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_307_)
);

OAI22X1 _818_ (
    .A(_307_),
    .B(_306_),
    .C(ra_adrs_1_bF$buf4),
    .D(_305_),
    .Y(_308_)
);

OAI21X1 _819_ (
    .A(ra_adrs_2_bF$buf0),
    .B(_308_),
    .C(_116__bF$buf3),
    .Y(_309_)
);

OAI21X1 _820_ (
    .A(_303_),
    .B(_309_),
    .C(_304_),
    .Y(_0_[10])
);

MUX2X1 _821_ (
    .A(\internal_reg[5] [11]),
    .B(\internal_reg[4] [11]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_310_)
);

NOR2X1 _822_ (
    .A(\internal_reg[7] [11]),
    .B(_94__bF$buf2),
    .Y(_311_)
);

OAI21X1 _823_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [11]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_312_)
);

OAI22X1 _824_ (
    .A(_312_),
    .B(_311_),
    .C(ra_adrs_1_bF$buf2),
    .D(_310_),
    .Y(_313_)
);

NOR2X1 _825_ (
    .A(_90_),
    .B(_313_),
    .Y(_314_)
);

OAI21X1 _826_ (
    .A(wr_en_bF$buf1),
    .B(_104__bF$buf1),
    .C(_683_[11]),
    .Y(_315_)
);

MUX2X1 _827_ (
    .A(\internal_reg[1] [11]),
    .B(\internal_reg[0] [11]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_316_)
);

NOR2X1 _828_ (
    .A(\internal_reg[3] [11]),
    .B(_94__bF$buf1),
    .Y(_317_)
);

OAI21X1 _829_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [11]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_318_)
);

OAI22X1 _830_ (
    .A(_318_),
    .B(_317_),
    .C(ra_adrs_1_bF$buf0),
    .D(_316_),
    .Y(_319_)
);

OAI21X1 _831_ (
    .A(ra_adrs_2_bF$buf3),
    .B(_319_),
    .C(_116__bF$buf2),
    .Y(_320_)
);

OAI21X1 _832_ (
    .A(_314_),
    .B(_320_),
    .C(_315_),
    .Y(_0_[11])
);

MUX2X1 _833_ (
    .A(\internal_reg[5] [12]),
    .B(\internal_reg[4] [12]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_321_)
);

NOR2X1 _834_ (
    .A(\internal_reg[7] [12]),
    .B(_94__bF$buf0),
    .Y(_322_)
);

OAI21X1 _835_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [12]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_323_)
);

OAI22X1 _836_ (
    .A(_323_),
    .B(_322_),
    .C(ra_adrs_1_bF$buf6),
    .D(_321_),
    .Y(_324_)
);

NOR2X1 _837_ (
    .A(_90_),
    .B(_324_),
    .Y(_325_)
);

OAI21X1 _838_ (
    .A(wr_en_bF$buf0),
    .B(_104__bF$buf0),
    .C(_683_[12]),
    .Y(_326_)
);

MUX2X1 _839_ (
    .A(\internal_reg[1] [12]),
    .B(\internal_reg[0] [12]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_327_)
);

NOR2X1 _840_ (
    .A(\internal_reg[3] [12]),
    .B(_94__bF$buf4),
    .Y(_328_)
);

OAI21X1 _841_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [12]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_329_)
);

OAI22X1 _842_ (
    .A(_329_),
    .B(_328_),
    .C(ra_adrs_1_bF$buf4),
    .D(_327_),
    .Y(_330_)
);

OAI21X1 _843_ (
    .A(ra_adrs_2_bF$buf2),
    .B(_330_),
    .C(_116__bF$buf1),
    .Y(_331_)
);

OAI21X1 _844_ (
    .A(_325_),
    .B(_331_),
    .C(_326_),
    .Y(_0_[12])
);

MUX2X1 _845_ (
    .A(\internal_reg[5] [13]),
    .B(\internal_reg[4] [13]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_332_)
);

NOR2X1 _846_ (
    .A(\internal_reg[7] [13]),
    .B(_94__bF$buf3),
    .Y(_333_)
);

OAI21X1 _847_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [13]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_334_)
);

OAI22X1 _848_ (
    .A(_334_),
    .B(_333_),
    .C(ra_adrs_1_bF$buf2),
    .D(_332_),
    .Y(_335_)
);

NOR2X1 _849_ (
    .A(_90_),
    .B(_335_),
    .Y(_336_)
);

OAI21X1 _850_ (
    .A(wr_en_bF$buf4),
    .B(_104__bF$buf4),
    .C(_683_[13]),
    .Y(_337_)
);

MUX2X1 _851_ (
    .A(\internal_reg[1] [13]),
    .B(\internal_reg[0] [13]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_338_)
);

NOR2X1 _852_ (
    .A(\internal_reg[3] [13]),
    .B(_94__bF$buf2),
    .Y(_339_)
);

OAI21X1 _853_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [13]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_340_)
);

OAI22X1 _854_ (
    .A(_340_),
    .B(_339_),
    .C(ra_adrs_1_bF$buf0),
    .D(_338_),
    .Y(_341_)
);

OAI21X1 _855_ (
    .A(ra_adrs_2_bF$buf1),
    .B(_341_),
    .C(_116__bF$buf0),
    .Y(_342_)
);

OAI21X1 _856_ (
    .A(_336_),
    .B(_342_),
    .C(_337_),
    .Y(_0_[13])
);

MUX2X1 _857_ (
    .A(\internal_reg[5] [14]),
    .B(\internal_reg[4] [14]),
    .S(ra_adrs_0_bF$buf6),
    .Y(_343_)
);

NOR2X1 _858_ (
    .A(\internal_reg[7] [14]),
    .B(_94__bF$buf1),
    .Y(_344_)
);

OAI21X1 _859_ (
    .A(ra_adrs_0_bF$buf5),
    .B(\internal_reg[6] [14]),
    .C(ra_adrs_1_bF$buf7),
    .Y(_345_)
);

OAI22X1 _860_ (
    .A(_345_),
    .B(_344_),
    .C(ra_adrs_1_bF$buf6),
    .D(_343_),
    .Y(_346_)
);

NOR2X1 _861_ (
    .A(_90_),
    .B(_346_),
    .Y(_347_)
);

OAI21X1 _862_ (
    .A(wr_en_bF$buf3),
    .B(_104__bF$buf3),
    .C(_683_[14]),
    .Y(_348_)
);

MUX2X1 _863_ (
    .A(\internal_reg[1] [14]),
    .B(\internal_reg[0] [14]),
    .S(ra_adrs_0_bF$buf4),
    .Y(_349_)
);

NOR2X1 _864_ (
    .A(\internal_reg[3] [14]),
    .B(_94__bF$buf0),
    .Y(_350_)
);

OAI21X1 _865_ (
    .A(ra_adrs_0_bF$buf3),
    .B(\internal_reg[2] [14]),
    .C(ra_adrs_1_bF$buf5),
    .Y(_351_)
);

OAI22X1 _866_ (
    .A(_351_),
    .B(_350_),
    .C(ra_adrs_1_bF$buf4),
    .D(_349_),
    .Y(_352_)
);

OAI21X1 _867_ (
    .A(ra_adrs_2_bF$buf0),
    .B(_352_),
    .C(_116__bF$buf4),
    .Y(_353_)
);

OAI21X1 _868_ (
    .A(_347_),
    .B(_353_),
    .C(_348_),
    .Y(_0_[14])
);

MUX2X1 _869_ (
    .A(\internal_reg[5] [15]),
    .B(\internal_reg[4] [15]),
    .S(ra_adrs_0_bF$buf2),
    .Y(_354_)
);

NOR2X1 _870_ (
    .A(\internal_reg[7] [15]),
    .B(_94__bF$buf4),
    .Y(_355_)
);

OAI21X1 _871_ (
    .A(ra_adrs_0_bF$buf1),
    .B(\internal_reg[6] [15]),
    .C(ra_adrs_1_bF$buf3),
    .Y(_356_)
);

OAI22X1 _872_ (
    .A(_356_),
    .B(_355_),
    .C(ra_adrs_1_bF$buf2),
    .D(_354_),
    .Y(_357_)
);

NOR2X1 _873_ (
    .A(_90_),
    .B(_357_),
    .Y(_358_)
);

OAI21X1 _874_ (
    .A(wr_en_bF$buf2),
    .B(_104__bF$buf2),
    .C(_683_[15]),
    .Y(_359_)
);

MUX2X1 _875_ (
    .A(\internal_reg[1] [15]),
    .B(\internal_reg[0] [15]),
    .S(ra_adrs_0_bF$buf0),
    .Y(_360_)
);

NOR2X1 _876_ (
    .A(\internal_reg[3] [15]),
    .B(_94__bF$buf3),
    .Y(_361_)
);

OAI21X1 _877_ (
    .A(ra_adrs_0_bF$buf7),
    .B(\internal_reg[2] [15]),
    .C(ra_adrs_1_bF$buf1),
    .Y(_362_)
);

OAI22X1 _878_ (
    .A(_362_),
    .B(_361_),
    .C(ra_adrs_1_bF$buf0),
    .D(_360_),
    .Y(_363_)
);

OAI21X1 _879_ (
    .A(ra_adrs_2_bF$buf3),
    .B(_363_),
    .C(_116__bF$buf3),
    .Y(_364_)
);

OAI21X1 _880_ (
    .A(_358_),
    .B(_364_),
    .C(_359_),
    .Y(_0_[15])
);

INVX2 _881_ (
    .A(data_in[0]),
    .Y(_365_)
);

INVX1 _882_ (
    .A(rd_adrs[2]),
    .Y(_366_)
);

INVX1 _883_ (
    .A(rd_adrs[1]),
    .Y(_367_)
);

NAND2X1 _884_ (
    .A(wr_en_bF$buf1),
    .B(enable),
    .Y(_368_)
);

NOR2X1 _885_ (
    .A(rd_adrs[0]),
    .B(_368_),
    .Y(_369_)
);

NAND3X1 _886_ (
    .A(_366_),
    .B(_367_),
    .C(_369_),
    .Y(_370_)
);

NAND2X1 _887_ (
    .A(\internal_reg[0] [0]),
    .B(_370__bF$buf4),
    .Y(_371_)
);

OAI21X1 _888_ (
    .A(_365_),
    .B(_370__bF$buf3),
    .C(_371_),
    .Y(_57_)
);

INVX2 _889_ (
    .A(data_in[1]),
    .Y(_372_)
);

NAND2X1 _890_ (
    .A(\internal_reg[0] [1]),
    .B(_370__bF$buf2),
    .Y(_373_)
);

OAI21X1 _891_ (
    .A(_372_),
    .B(_370__bF$buf1),
    .C(_373_),
    .Y(_58_)
);

INVX2 _892_ (
    .A(data_in[2]),
    .Y(_374_)
);

NAND2X1 _893_ (
    .A(\internal_reg[0] [2]),
    .B(_370__bF$buf0),
    .Y(_375_)
);

OAI21X1 _894_ (
    .A(_374_),
    .B(_370__bF$buf4),
    .C(_375_),
    .Y(_59_)
);

INVX2 _895_ (
    .A(data_in[3]),
    .Y(_376_)
);

NAND2X1 _896_ (
    .A(\internal_reg[0] [3]),
    .B(_370__bF$buf3),
    .Y(_377_)
);

OAI21X1 _897_ (
    .A(_376_),
    .B(_370__bF$buf2),
    .C(_377_),
    .Y(_60_)
);

INVX2 _898_ (
    .A(data_in[4]),
    .Y(_378_)
);

NAND2X1 _899_ (
    .A(\internal_reg[0] [4]),
    .B(_370__bF$buf1),
    .Y(_379_)
);

OAI21X1 _900_ (
    .A(_378_),
    .B(_370__bF$buf0),
    .C(_379_),
    .Y(_61_)
);

INVX2 _901_ (
    .A(data_in[5]),
    .Y(_380_)
);

NAND2X1 _902_ (
    .A(\internal_reg[0] [5]),
    .B(_370__bF$buf4),
    .Y(_381_)
);

OAI21X1 _903_ (
    .A(_380_),
    .B(_370__bF$buf3),
    .C(_381_),
    .Y(_62_)
);

INVX2 _904_ (
    .A(data_in[6]),
    .Y(_382_)
);

NAND2X1 _905_ (
    .A(\internal_reg[0] [6]),
    .B(_370__bF$buf2),
    .Y(_383_)
);

OAI21X1 _906_ (
    .A(_382_),
    .B(_370__bF$buf1),
    .C(_383_),
    .Y(_63_)
);

INVX2 _907_ (
    .A(data_in[7]),
    .Y(_384_)
);

NAND2X1 _908_ (
    .A(\internal_reg[0] [7]),
    .B(_370__bF$buf0),
    .Y(_385_)
);

OAI21X1 _909_ (
    .A(_384_),
    .B(_370__bF$buf4),
    .C(_385_),
    .Y(_64_)
);

INVX2 _910_ (
    .A(data_in[8]),
    .Y(_386_)
);

NAND2X1 _911_ (
    .A(\internal_reg[0] [8]),
    .B(_370__bF$buf3),
    .Y(_387_)
);

OAI21X1 _912_ (
    .A(_386_),
    .B(_370__bF$buf2),
    .C(_387_),
    .Y(_65_)
);

INVX2 _913_ (
    .A(data_in[9]),
    .Y(_388_)
);

NAND2X1 _914_ (
    .A(\internal_reg[0] [9]),
    .B(_370__bF$buf1),
    .Y(_389_)
);

OAI21X1 _915_ (
    .A(_388_),
    .B(_370__bF$buf0),
    .C(_389_),
    .Y(_66_)
);

INVX2 _916_ (
    .A(data_in[10]),
    .Y(_390_)
);

NAND2X1 _917_ (
    .A(\internal_reg[0] [10]),
    .B(_370__bF$buf4),
    .Y(_391_)
);

OAI21X1 _918_ (
    .A(_390_),
    .B(_370__bF$buf3),
    .C(_391_),
    .Y(_67_)
);

INVX2 _919_ (
    .A(data_in[11]),
    .Y(_392_)
);

NAND2X1 _920_ (
    .A(\internal_reg[0] [11]),
    .B(_370__bF$buf2),
    .Y(_393_)
);

OAI21X1 _921_ (
    .A(_392_),
    .B(_370__bF$buf1),
    .C(_393_),
    .Y(_68_)
);

INVX2 _922_ (
    .A(data_in[12]),
    .Y(_394_)
);

NAND2X1 _923_ (
    .A(\internal_reg[0] [12]),
    .B(_370__bF$buf0),
    .Y(_395_)
);

OAI21X1 _924_ (
    .A(_394_),
    .B(_370__bF$buf4),
    .C(_395_),
    .Y(_69_)
);

INVX2 _925_ (
    .A(data_in[13]),
    .Y(_396_)
);

NAND2X1 _926_ (
    .A(\internal_reg[0] [13]),
    .B(_370__bF$buf3),
    .Y(_397_)
);

OAI21X1 _927_ (
    .A(_396_),
    .B(_370__bF$buf2),
    .C(_397_),
    .Y(_70_)
);

INVX2 _928_ (
    .A(data_in[14]),
    .Y(_398_)
);

NAND2X1 _929_ (
    .A(\internal_reg[0] [14]),
    .B(_370__bF$buf1),
    .Y(_399_)
);

OAI21X1 _930_ (
    .A(_398_),
    .B(_370__bF$buf0),
    .C(_399_),
    .Y(_71_)
);

INVX2 _931_ (
    .A(data_in[15]),
    .Y(_400_)
);

NAND2X1 _932_ (
    .A(\internal_reg[0] [15]),
    .B(_370__bF$buf4),
    .Y(_401_)
);

OAI21X1 _933_ (
    .A(_400_),
    .B(_370__bF$buf3),
    .C(_401_),
    .Y(_72_)
);

NAND2X1 _934_ (
    .A(_366_),
    .B(_367_),
    .Y(_402_)
);

AND2X2 _935_ (
    .A(wr_en_bF$buf0),
    .B(enable),
    .Y(_403_)
);

NAND2X1 _936_ (
    .A(rd_adrs[0]),
    .B(_403_),
    .Y(_404_)
);

OR2X2 _937_ (
    .A(_404__bF$buf1),
    .B(_402__bF$buf3),
    .Y(_405_)
);

OAI21X1 _938_ (
    .A(_402__bF$buf2),
    .B(_404__bF$buf0),
    .C(\internal_reg[1] [0]),
    .Y(_406_)
);

OAI21X1 _939_ (
    .A(_365_),
    .B(_405_),
    .C(_406_),
    .Y(_73_)
);

OAI21X1 _940_ (
    .A(_402__bF$buf1),
    .B(_404__bF$buf4),
    .C(\internal_reg[1] [1]),
    .Y(_407_)
);

OAI21X1 _941_ (
    .A(_372_),
    .B(_405_),
    .C(_407_),
    .Y(_74_)
);

OAI21X1 _942_ (
    .A(_402__bF$buf0),
    .B(_404__bF$buf3),
    .C(\internal_reg[1] [2]),
    .Y(_408_)
);

OAI21X1 _943_ (
    .A(_374_),
    .B(_405_),
    .C(_408_),
    .Y(_75_)
);

OAI21X1 _944_ (
    .A(_402__bF$buf3),
    .B(_404__bF$buf2),
    .C(\internal_reg[1] [3]),
    .Y(_409_)
);

OAI21X1 _945_ (
    .A(_376_),
    .B(_405_),
    .C(_409_),
    .Y(_76_)
);

OAI21X1 _946_ (
    .A(_402__bF$buf2),
    .B(_404__bF$buf1),
    .C(\internal_reg[1] [4]),
    .Y(_410_)
);

OAI21X1 _947_ (
    .A(_378_),
    .B(_405_),
    .C(_410_),
    .Y(_77_)
);

OAI21X1 _948_ (
    .A(_402__bF$buf1),
    .B(_404__bF$buf0),
    .C(\internal_reg[1] [5]),
    .Y(_411_)
);

OAI21X1 _949_ (
    .A(_380_),
    .B(_405_),
    .C(_411_),
    .Y(_78_)
);

OAI21X1 _950_ (
    .A(_402__bF$buf0),
    .B(_404__bF$buf4),
    .C(\internal_reg[1] [6]),
    .Y(_412_)
);

OAI21X1 _951_ (
    .A(_382_),
    .B(_405_),
    .C(_412_),
    .Y(_79_)
);

OAI21X1 _952_ (
    .A(_402__bF$buf3),
    .B(_404__bF$buf3),
    .C(\internal_reg[1] [7]),
    .Y(_413_)
);

OAI21X1 _953_ (
    .A(_384_),
    .B(_405_),
    .C(_413_),
    .Y(_80_)
);

OAI21X1 _954_ (
    .A(_402__bF$buf2),
    .B(_404__bF$buf2),
    .C(\internal_reg[1] [8]),
    .Y(_414_)
);

OAI21X1 _955_ (
    .A(_386_),
    .B(_405_),
    .C(_414_),
    .Y(_81_)
);

OAI21X1 _956_ (
    .A(_402__bF$buf1),
    .B(_404__bF$buf1),
    .C(\internal_reg[1] [9]),
    .Y(_415_)
);

OAI21X1 _957_ (
    .A(_388_),
    .B(_405_),
    .C(_415_),
    .Y(_82_)
);

OAI21X1 _958_ (
    .A(_402__bF$buf0),
    .B(_404__bF$buf0),
    .C(\internal_reg[1] [10]),
    .Y(_416_)
);

OAI21X1 _959_ (
    .A(_390_),
    .B(_405_),
    .C(_416_),
    .Y(_83_)
);

OAI21X1 _960_ (
    .A(_402__bF$buf3),
    .B(_404__bF$buf4),
    .C(\internal_reg[1] [11]),
    .Y(_417_)
);

OAI21X1 _961_ (
    .A(_392_),
    .B(_405_),
    .C(_417_),
    .Y(_84_)
);

OAI21X1 _962_ (
    .A(_402__bF$buf2),
    .B(_404__bF$buf3),
    .C(\internal_reg[1] [12]),
    .Y(_418_)
);

OAI21X1 _963_ (
    .A(_394_),
    .B(_405_),
    .C(_418_),
    .Y(_85_)
);

OAI21X1 _964_ (
    .A(_402__bF$buf1),
    .B(_404__bF$buf2),
    .C(\internal_reg[1] [13]),
    .Y(_419_)
);

OAI21X1 _965_ (
    .A(_396_),
    .B(_405_),
    .C(_419_),
    .Y(_86_)
);

OAI21X1 _966_ (
    .A(_402__bF$buf0),
    .B(_404__bF$buf1),
    .C(\internal_reg[1] [14]),
    .Y(_420_)
);

OAI21X1 _967_ (
    .A(_398_),
    .B(_405_),
    .C(_420_),
    .Y(_87_)
);

OAI21X1 _968_ (
    .A(_402__bF$buf3),
    .B(_404__bF$buf0),
    .C(\internal_reg[1] [15]),
    .Y(_421_)
);

OAI21X1 _969_ (
    .A(_400_),
    .B(_405_),
    .C(_421_),
    .Y(_88_)
);

NOR2X1 _970_ (
    .A(rd_adrs[2]),
    .B(_367_),
    .Y(_422_)
);

NAND2X1 _971_ (
    .A(_422__bF$buf2),
    .B(_369_),
    .Y(_423_)
);

NAND2X1 _972_ (
    .A(\internal_reg[2] [0]),
    .B(_423__bF$buf0),
    .Y(_424_)
);

OAI21X1 _973_ (
    .A(_365_),
    .B(_423__bF$buf4),
    .C(_424_),
    .Y(_89_)
);

NAND2X1 _974_ (
    .A(\internal_reg[2] [1]),
    .B(_423__bF$buf3),
    .Y(_425_)
);

OAI21X1 _975_ (
    .A(_372_),
    .B(_423__bF$buf2),
    .C(_425_),
    .Y(_91_)
);

NAND2X1 _976_ (
    .A(\internal_reg[2] [2]),
    .B(_423__bF$buf1),
    .Y(_426_)
);

OAI21X1 _977_ (
    .A(_374_),
    .B(_423__bF$buf0),
    .C(_426_),
    .Y(_93_)
);

NAND2X1 _978_ (
    .A(\internal_reg[2] [3]),
    .B(_423__bF$buf4),
    .Y(_427_)
);

OAI21X1 _979_ (
    .A(_376_),
    .B(_423__bF$buf3),
    .C(_427_),
    .Y(_95_)
);

NAND2X1 _980_ (
    .A(\internal_reg[2] [4]),
    .B(_423__bF$buf2),
    .Y(_428_)
);

OAI21X1 _981_ (
    .A(_378_),
    .B(_423__bF$buf1),
    .C(_428_),
    .Y(_97_)
);

NAND2X1 _982_ (
    .A(\internal_reg[2] [5]),
    .B(_423__bF$buf0),
    .Y(_429_)
);

OAI21X1 _983_ (
    .A(_380_),
    .B(_423__bF$buf4),
    .C(_429_),
    .Y(_99_)
);

NAND2X1 _984_ (
    .A(\internal_reg[2] [6]),
    .B(_423__bF$buf3),
    .Y(_430_)
);

OAI21X1 _985_ (
    .A(_382_),
    .B(_423__bF$buf2),
    .C(_430_),
    .Y(_101_)
);

NAND2X1 _986_ (
    .A(\internal_reg[2] [7]),
    .B(_423__bF$buf1),
    .Y(_431_)
);

OAI21X1 _987_ (
    .A(_384_),
    .B(_423__bF$buf0),
    .C(_431_),
    .Y(_103_)
);

NAND2X1 _988_ (
    .A(\internal_reg[2] [8]),
    .B(_423__bF$buf4),
    .Y(_432_)
);

OAI21X1 _989_ (
    .A(_386_),
    .B(_423__bF$buf3),
    .C(_432_),
    .Y(_105_)
);

NAND2X1 _990_ (
    .A(\internal_reg[2] [9]),
    .B(_423__bF$buf2),
    .Y(_433_)
);

OAI21X1 _991_ (
    .A(_388_),
    .B(_423__bF$buf1),
    .C(_433_),
    .Y(_107_)
);

NAND2X1 _992_ (
    .A(\internal_reg[2] [10]),
    .B(_423__bF$buf0),
    .Y(_434_)
);

OAI21X1 _993_ (
    .A(_390_),
    .B(_423__bF$buf4),
    .C(_434_),
    .Y(_109_)
);

NAND2X1 _994_ (
    .A(\internal_reg[2] [11]),
    .B(_423__bF$buf3),
    .Y(_435_)
);

OAI21X1 _995_ (
    .A(_392_),
    .B(_423__bF$buf2),
    .C(_435_),
    .Y(_111_)
);

NAND2X1 _996_ (
    .A(\internal_reg[2] [12]),
    .B(_423__bF$buf1),
    .Y(_436_)
);

OAI21X1 _997_ (
    .A(_394_),
    .B(_423__bF$buf0),
    .C(_436_),
    .Y(_113_)
);

NAND2X1 _998_ (
    .A(\internal_reg[2] [13]),
    .B(_423__bF$buf4),
    .Y(_437_)
);

OAI21X1 _999_ (
    .A(_396_),
    .B(_423__bF$buf3),
    .C(_437_),
    .Y(_115_)
);

endmodule
