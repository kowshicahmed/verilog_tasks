magic
tech scmos
magscale 1 2
timestamp 1594572398
<< metal1 >>
rect 762 614 774 616
rect 747 606 749 614
rect 757 606 759 614
rect 767 606 769 614
rect 777 606 779 614
rect 787 606 789 614
rect 762 604 774 606
rect 749 557 812 563
rect 596 537 611 543
rect 1053 537 1068 543
rect 637 517 675 523
rect 733 517 796 523
rect 820 517 835 523
rect 605 497 627 503
rect 298 414 310 416
rect 283 406 285 414
rect 293 406 295 414
rect 303 406 305 414
rect 313 406 315 414
rect 323 406 325 414
rect 298 404 310 406
rect 205 377 252 383
rect 506 376 508 384
rect 109 297 131 303
rect 708 297 739 303
rect 228 277 292 283
rect 589 277 627 283
rect 701 277 723 283
rect 717 264 723 277
rect 989 277 1004 283
rect 1005 257 1020 263
rect 205 237 236 243
rect 762 214 774 216
rect 747 206 749 214
rect 757 206 759 214
rect 767 206 769 214
rect 777 206 779 214
rect 787 206 789 214
rect 762 204 774 206
rect 740 177 803 183
rect 1028 176 1030 184
rect 188 157 211 163
rect 188 154 196 157
rect 221 117 236 123
rect 605 117 627 123
rect 669 117 691 123
rect 836 97 851 103
rect 893 97 915 103
rect 948 97 963 103
rect 956 84 964 88
rect 269 77 332 83
rect 298 14 310 16
rect 283 6 285 14
rect 293 6 295 14
rect 303 6 305 14
rect 313 6 315 14
rect 323 6 325 14
rect 298 4 310 6
<< m2contact >>
rect 739 606 747 614
rect 749 606 757 614
rect 759 606 767 614
rect 769 606 777 614
rect 779 606 787 614
rect 789 606 797 614
rect 572 576 580 584
rect 700 576 708 584
rect 860 576 868 584
rect 908 576 916 584
rect 956 576 964 584
rect 284 556 292 564
rect 364 556 372 564
rect 588 556 596 564
rect 812 556 820 564
rect 988 558 996 566
rect 1036 558 1044 566
rect 220 536 228 544
rect 412 536 420 544
rect 588 536 596 544
rect 652 536 660 544
rect 1068 536 1076 544
rect 44 516 52 524
rect 188 518 196 526
rect 252 516 260 524
rect 268 516 276 524
rect 380 516 388 524
rect 444 518 452 526
rect 716 516 724 524
rect 796 516 804 524
rect 812 516 820 524
rect 876 516 884 524
rect 924 516 932 524
rect 972 516 980 524
rect 1020 516 1028 524
rect 12 476 20 484
rect 1004 476 1012 484
rect 60 456 68 464
rect 275 406 283 414
rect 285 406 293 414
rect 295 406 303 414
rect 305 406 313 414
rect 315 406 323 414
rect 325 406 333 414
rect 252 376 260 384
rect 460 376 468 384
rect 508 376 516 384
rect 860 376 868 384
rect 76 356 84 364
rect 476 316 484 324
rect 652 316 660 324
rect 28 296 36 304
rect 332 294 340 302
rect 508 296 516 304
rect 572 296 580 304
rect 636 296 644 304
rect 684 296 692 304
rect 700 296 708 304
rect 748 296 756 304
rect 860 296 868 304
rect 892 296 900 304
rect 908 296 916 304
rect 924 296 932 304
rect 12 276 20 284
rect 156 280 164 288
rect 172 276 180 284
rect 220 276 228 284
rect 396 276 404 284
rect 524 276 532 284
rect 876 276 884 284
rect 940 276 948 284
rect 1004 276 1012 284
rect 188 256 196 264
rect 604 256 612 264
rect 716 256 724 264
rect 828 256 836 264
rect 956 256 964 264
rect 1020 256 1028 264
rect 60 236 68 244
rect 236 236 244 244
rect 540 236 548 244
rect 652 236 660 244
rect 1036 236 1044 244
rect 739 206 747 214
rect 749 206 757 214
rect 759 206 767 214
rect 769 206 777 214
rect 779 206 787 214
rect 789 206 797 214
rect 188 176 196 184
rect 524 176 532 184
rect 732 176 740 184
rect 908 176 916 184
rect 956 176 964 184
rect 1020 176 1028 184
rect 236 156 244 164
rect 396 156 404 164
rect 588 156 596 164
rect 668 156 676 164
rect 860 156 868 164
rect 876 156 884 164
rect 92 136 100 144
rect 636 136 644 144
rect 828 136 836 144
rect 940 136 948 144
rect 988 136 996 144
rect 1004 136 1012 144
rect 60 118 68 126
rect 236 116 244 124
rect 268 116 276 124
rect 396 118 404 126
rect 540 116 548 124
rect 796 96 804 104
rect 828 96 836 104
rect 940 96 948 104
rect 1036 96 1044 104
rect 332 76 340 84
rect 956 76 964 84
rect 572 36 580 44
rect 716 36 724 44
rect 275 6 283 14
rect 285 6 293 14
rect 295 6 303 14
rect 305 6 313 14
rect 315 6 323 14
rect 325 6 333 14
<< metal2 >>
rect 685 657 707 663
rect 845 657 867 663
rect 893 657 915 663
rect 941 657 963 663
rect 701 584 707 657
rect 762 614 774 616
rect 747 606 749 614
rect 757 606 759 614
rect 767 606 769 614
rect 777 606 779 614
rect 787 606 789 614
rect 762 604 774 606
rect 861 584 867 657
rect 909 584 915 657
rect 957 584 963 657
rect 573 563 579 576
rect 573 557 588 563
rect 973 558 988 563
rect 1021 558 1036 563
rect 973 557 995 558
rect 1021 557 1043 558
rect 285 544 291 556
rect 13 484 19 496
rect 45 463 51 516
rect 29 457 60 463
rect 29 304 35 457
rect 221 284 227 536
rect 253 384 259 516
rect 413 483 419 536
rect 397 477 419 483
rect 298 414 310 416
rect 283 406 285 414
rect 293 406 295 414
rect 303 406 305 414
rect 313 406 315 414
rect 323 406 325 414
rect 298 404 310 406
rect 61 126 67 236
rect 157 184 163 280
rect 173 264 179 276
rect 189 264 195 276
rect 221 144 227 276
rect 237 244 243 296
rect 397 284 403 477
rect 509 384 515 556
rect 653 384 659 536
rect 717 524 723 536
rect 813 524 819 556
rect 973 524 979 557
rect 1021 524 1027 557
rect 925 504 931 516
rect 861 384 867 496
rect 1005 484 1011 496
rect 477 284 483 316
rect 237 164 243 236
rect 397 164 403 276
rect 509 183 515 296
rect 525 284 531 376
rect 653 304 659 316
rect 509 177 524 183
rect 541 124 547 236
rect 589 164 595 296
rect 605 264 611 276
rect 637 184 643 296
rect 669 164 675 296
rect 685 184 691 296
rect 701 264 707 296
rect 749 284 755 296
rect 829 244 835 256
rect 893 244 899 296
rect 762 214 774 216
rect 747 206 749 214
rect 757 206 759 214
rect 767 206 769 214
rect 777 206 779 214
rect 787 206 789 214
rect 762 204 774 206
rect 909 184 915 276
rect 925 224 931 296
rect 957 184 963 216
rect 829 144 835 156
rect 861 144 867 156
rect 989 144 995 156
rect 1005 144 1011 276
rect 1021 264 1027 296
rect 1021 184 1027 236
rect 637 124 643 136
rect 397 104 403 118
rect 941 104 947 136
rect 1005 124 1011 136
rect 1037 104 1043 236
rect 333 84 339 96
rect 298 14 310 16
rect 283 6 285 14
rect 293 6 295 14
rect 303 6 305 14
rect 313 6 315 14
rect 323 6 325 14
rect 298 4 310 6
rect 573 -17 579 36
rect 717 -17 723 36
rect 557 -23 579 -17
rect 701 -23 723 -17
rect 957 -23 963 76
<< m3contact >>
rect 739 606 747 614
rect 749 606 757 614
rect 759 606 767 614
rect 769 606 777 614
rect 779 606 787 614
rect 789 606 797 614
rect 364 556 372 564
rect 508 556 516 564
rect 588 556 596 564
rect 812 556 820 564
rect 284 536 292 544
rect 188 518 196 524
rect 188 516 196 518
rect 12 496 20 504
rect 76 356 84 364
rect 12 276 20 284
rect 268 516 276 524
rect 380 516 388 524
rect 444 518 452 524
rect 444 516 452 518
rect 275 406 283 414
rect 285 406 293 414
rect 295 406 303 414
rect 305 406 313 414
rect 315 406 323 414
rect 325 406 333 414
rect 236 296 244 304
rect 332 302 340 304
rect 332 296 340 302
rect 188 276 196 284
rect 172 256 180 264
rect 156 176 164 184
rect 188 176 196 184
rect 588 536 596 544
rect 652 536 660 544
rect 716 536 724 544
rect 1068 536 1076 544
rect 796 516 804 524
rect 876 516 884 524
rect 860 496 868 504
rect 924 496 932 504
rect 1004 496 1012 504
rect 460 376 468 384
rect 524 376 532 384
rect 652 376 660 384
rect 508 296 516 304
rect 476 276 484 284
rect 572 296 580 304
rect 588 296 596 304
rect 652 296 660 304
rect 668 296 676 304
rect 860 296 868 304
rect 908 296 916 304
rect 1020 296 1028 304
rect 92 136 100 144
rect 220 136 228 144
rect 236 116 244 124
rect 268 116 276 124
rect 604 276 612 284
rect 652 236 660 244
rect 636 176 644 184
rect 748 276 756 284
rect 876 276 884 284
rect 700 256 708 264
rect 716 256 724 264
rect 908 276 916 284
rect 828 236 836 244
rect 892 236 900 244
rect 739 206 747 214
rect 749 206 757 214
rect 759 206 767 214
rect 769 206 777 214
rect 779 206 787 214
rect 789 206 797 214
rect 940 276 948 284
rect 1004 276 1012 284
rect 956 256 964 264
rect 924 216 932 224
rect 956 216 964 224
rect 684 176 692 184
rect 732 176 740 184
rect 828 156 836 164
rect 876 156 884 164
rect 988 156 996 164
rect 1020 236 1028 244
rect 860 136 868 144
rect 940 136 948 144
rect 636 116 644 124
rect 1004 116 1012 124
rect 332 96 340 104
rect 396 96 404 104
rect 796 96 804 104
rect 828 96 836 104
rect 275 6 283 14
rect 285 6 293 14
rect 295 6 303 14
rect 305 6 313 14
rect 315 6 323 14
rect 325 6 333 14
<< metal3 >>
rect 738 614 798 616
rect 738 606 739 614
rect 748 606 749 614
rect 787 606 788 614
rect 797 606 798 614
rect 738 604 798 606
rect 372 557 508 563
rect 596 557 812 563
rect 292 537 588 543
rect 660 537 716 543
rect 1076 537 1107 543
rect 196 517 268 523
rect 388 517 444 523
rect 804 517 876 523
rect -35 497 12 503
rect 868 497 924 503
rect 1012 497 1107 503
rect 274 414 334 416
rect 274 406 275 414
rect 284 406 285 414
rect 323 406 324 414
rect 333 406 334 414
rect 274 404 334 406
rect 468 377 524 383
rect 532 377 652 383
rect -35 357 76 363
rect -35 317 -29 323
rect 244 297 332 303
rect 516 297 572 303
rect 580 297 588 303
rect 596 297 652 303
rect 676 297 860 303
rect 868 297 908 303
rect 1028 297 1107 303
rect -35 277 12 283
rect 20 277 188 283
rect 196 277 476 283
rect 612 277 723 283
rect 717 264 723 277
rect 756 277 876 283
rect 884 277 908 283
rect 948 277 1004 283
rect 180 257 700 263
rect 724 257 956 263
rect 660 237 828 243
rect 900 237 1020 243
rect 932 217 956 223
rect 738 214 798 216
rect 738 206 739 214
rect 748 206 749 214
rect 787 206 788 214
rect 797 206 798 214
rect 738 204 798 206
rect 164 177 188 183
rect 644 177 684 183
rect 692 177 732 183
rect 836 157 876 163
rect 884 157 988 163
rect 996 157 1107 163
rect -35 137 92 143
rect 100 137 220 143
rect 868 137 940 143
rect 244 117 268 123
rect 276 117 636 123
rect 1012 117 1107 123
rect 340 97 396 103
rect 804 97 828 103
rect 274 14 334 16
rect 274 6 275 14
rect 284 6 285 14
rect 323 6 324 14
rect 333 6 334 14
rect 274 4 334 6
<< m4contact >>
rect 740 606 747 614
rect 747 606 748 614
rect 752 606 757 614
rect 757 606 759 614
rect 759 606 760 614
rect 764 606 767 614
rect 767 606 769 614
rect 769 606 772 614
rect 776 606 777 614
rect 777 606 779 614
rect 779 606 784 614
rect 788 606 789 614
rect 789 606 796 614
rect 276 406 283 414
rect 283 406 284 414
rect 288 406 293 414
rect 293 406 295 414
rect 295 406 296 414
rect 300 406 303 414
rect 303 406 305 414
rect 305 406 308 414
rect 312 406 313 414
rect 313 406 315 414
rect 315 406 320 414
rect 324 406 325 414
rect 325 406 332 414
rect 740 206 747 214
rect 747 206 748 214
rect 752 206 757 214
rect 757 206 759 214
rect 759 206 760 214
rect 764 206 767 214
rect 767 206 769 214
rect 769 206 772 214
rect 776 206 777 214
rect 777 206 779 214
rect 779 206 784 214
rect 788 206 789 214
rect 789 206 796 214
rect 276 6 283 14
rect 283 6 284 14
rect 288 6 293 14
rect 293 6 295 14
rect 295 6 296 14
rect 300 6 303 14
rect 303 6 305 14
rect 305 6 308 14
rect 312 6 313 14
rect 313 6 315 14
rect 315 6 320 14
rect 324 6 325 14
rect 325 6 332 14
<< metal4 >>
rect 272 414 336 616
rect 272 406 276 414
rect 284 406 288 414
rect 296 406 300 414
rect 308 406 312 414
rect 320 406 324 414
rect 332 406 336 414
rect 272 14 336 406
rect 272 6 276 14
rect 284 6 288 14
rect 296 6 300 14
rect 308 6 312 14
rect 320 6 324 14
rect 332 6 336 14
rect 272 -10 336 6
rect 736 614 800 616
rect 736 606 740 614
rect 748 606 752 614
rect 760 606 764 614
rect 772 606 776 614
rect 784 606 788 614
rect 796 606 800 614
rect 736 214 800 606
rect 736 206 740 214
rect 748 206 752 214
rect 760 206 764 214
rect 772 206 776 214
rect 784 206 788 214
rect 796 206 800 214
rect 736 -10 800 206
use DFFPOSX1  _66_
timestamp 1594572398
transform 1 0 8 0 -1 210
box -4 -6 196 206
use INVX1  _51_
timestamp 1594572398
transform 1 0 200 0 -1 210
box -4 -6 36 206
use AND2X2  _54_
timestamp 1594572398
transform 1 0 8 0 1 210
box -4 -6 68 206
use BUFX2  _59_
timestamp 1594572398
transform -1 0 120 0 1 210
box -4 -6 52 206
use AND2X2  _41_
timestamp 1594572398
transform -1 0 184 0 1 210
box -4 -6 68 206
use INVX1  _31_
timestamp 1594572398
transform 1 0 184 0 1 210
box -4 -6 36 206
use FILL  SFILL2640x2100
timestamp 1594572398
transform 1 0 264 0 1 210
box -4 -6 20 206
use FILL  SFILL2480x2100
timestamp 1594572398
transform 1 0 248 0 1 210
box -4 -6 20 206
use FILL  SFILL2320x2100
timestamp 1594572398
transform 1 0 232 0 1 210
box -4 -6 20 206
use FILL  SFILL2160x2100
timestamp 1594572398
transform 1 0 216 0 1 210
box -4 -6 20 206
use FILL  SFILL2960x100
timestamp 1594572398
transform -1 0 312 0 -1 210
box -4 -6 20 206
use FILL  SFILL2800x100
timestamp 1594572398
transform -1 0 296 0 -1 210
box -4 -6 20 206
use NOR2X1  _53_
timestamp 1594572398
transform 1 0 232 0 -1 210
box -4 -6 52 206
use FILL  SFILL3280x100
timestamp 1594572398
transform -1 0 344 0 -1 210
box -4 -6 20 206
use FILL  SFILL3120x100
timestamp 1594572398
transform -1 0 328 0 -1 210
box -4 -6 20 206
use DFFPOSX1  _65_
timestamp 1594572398
transform 1 0 280 0 1 210
box -4 -6 196 206
use DFFPOSX1  _67_
timestamp 1594572398
transform 1 0 344 0 -1 210
box -4 -6 196 206
use BUFX2  _60_
timestamp 1594572398
transform 1 0 536 0 -1 210
box -4 -6 52 206
use INVX1  _50_
timestamp 1594572398
transform 1 0 584 0 -1 210
box -4 -6 36 206
use OAI21X1  _48_
timestamp 1594572398
transform -1 0 536 0 1 210
box -4 -6 68 206
use AND2X2  _37_
timestamp 1594572398
transform -1 0 600 0 1 210
box -4 -6 68 206
use NOR2X1  _36_
timestamp 1594572398
transform 1 0 600 0 1 210
box -4 -6 52 206
use OAI21X1  _46_
timestamp 1594572398
transform -1 0 712 0 1 210
box -4 -6 68 206
use BUFX2  _64_
timestamp 1594572398
transform 1 0 680 0 -1 210
box -4 -6 52 206
use AOI21X1  _52_
timestamp 1594572398
transform 1 0 616 0 -1 210
box -4 -6 68 206
use FILL  SFILL7440x100
timestamp 1594572398
transform -1 0 760 0 -1 210
box -4 -6 20 206
use FILL  SFILL7280x100
timestamp 1594572398
transform -1 0 744 0 -1 210
box -4 -6 20 206
use NOR2X1  _40_
timestamp 1594572398
transform 1 0 712 0 1 210
box -4 -6 52 206
use FILL  SFILL8080x2100
timestamp 1594572398
transform 1 0 808 0 1 210
box -4 -6 20 206
use FILL  SFILL7920x2100
timestamp 1594572398
transform 1 0 792 0 1 210
box -4 -6 20 206
use FILL  SFILL7760x2100
timestamp 1594572398
transform 1 0 776 0 1 210
box -4 -6 20 206
use FILL  SFILL7600x2100
timestamp 1594572398
transform 1 0 760 0 1 210
box -4 -6 20 206
use FILL  SFILL7760x100
timestamp 1594572398
transform -1 0 792 0 -1 210
box -4 -6 20 206
use FILL  SFILL7600x100
timestamp 1594572398
transform -1 0 776 0 -1 210
box -4 -6 20 206
use NAND2X1  _35_
timestamp 1594572398
transform -1 0 840 0 -1 210
box -4 -6 52 206
use INVX1  _34_
timestamp 1594572398
transform -1 0 872 0 -1 210
box -4 -6 36 206
use INVX1  _38_
timestamp 1594572398
transform 1 0 872 0 -1 210
box -4 -6 36 206
use NAND2X1  _39_
timestamp 1594572398
transform -1 0 952 0 -1 210
box -4 -6 52 206
use NAND2X1  _44_
timestamp 1594572398
transform -1 0 1000 0 -1 210
box -4 -6 52 206
use NAND2X1  _43_
timestamp 1594572398
transform 1 0 1000 0 -1 210
box -4 -6 52 206
use NOR2X1  _47_
timestamp 1594572398
transform 1 0 824 0 1 210
box -4 -6 52 206
use OAI22X1  _45_
timestamp 1594572398
transform -1 0 952 0 1 210
box -4 -6 84 206
use OR2X2  _33_
timestamp 1594572398
transform -1 0 1016 0 1 210
box -4 -6 68 206
use INVX1  _42_
timestamp 1594572398
transform 1 0 1016 0 1 210
box -4 -6 36 206
use FILL  FILL9200x100
timestamp 1594572398
transform -1 0 1064 0 -1 210
box -4 -6 20 206
use FILL  FILL9200x2100
timestamp 1594572398
transform 1 0 1048 0 1 210
box -4 -6 20 206
use BUFX2  _56_
timestamp 1594572398
transform -1 0 56 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _69_
timestamp 1594572398
transform -1 0 248 0 -1 610
box -4 -6 196 206
use NOR2X1  _32_
timestamp 1594572398
transform -1 0 296 0 -1 610
box -4 -6 52 206
use INVX1  _49_
timestamp 1594572398
transform 1 0 360 0 -1 610
box -4 -6 36 206
use DFFPOSX1  _68_
timestamp 1594572398
transform 1 0 392 0 -1 610
box -4 -6 196 206
use FILL  SFILL2960x4100
timestamp 1594572398
transform -1 0 312 0 -1 610
box -4 -6 20 206
use FILL  SFILL3120x4100
timestamp 1594572398
transform -1 0 328 0 -1 610
box -4 -6 20 206
use FILL  SFILL3280x4100
timestamp 1594572398
transform -1 0 344 0 -1 610
box -4 -6 20 206
use FILL  SFILL3440x4100
timestamp 1594572398
transform -1 0 360 0 -1 610
box -4 -6 20 206
use INVX1  _29_
timestamp 1594572398
transform 1 0 584 0 -1 610
box -4 -6 36 206
use NAND2X1  _30_
timestamp 1594572398
transform -1 0 664 0 -1 610
box -4 -6 52 206
use BUFX2  _62_
timestamp 1594572398
transform 1 0 664 0 -1 610
box -4 -6 52 206
use NOR2X1  _28_
timestamp 1594572398
transform -1 0 760 0 -1 610
box -4 -6 52 206
use FILL  SFILL7600x4100
timestamp 1594572398
transform -1 0 776 0 -1 610
box -4 -6 20 206
use FILL  SFILL7760x4100
timestamp 1594572398
transform -1 0 792 0 -1 610
box -4 -6 20 206
use FILL  SFILL7920x4100
timestamp 1594572398
transform -1 0 808 0 -1 610
box -4 -6 20 206
use FILL  SFILL8080x4100
timestamp 1594572398
transform -1 0 824 0 -1 610
box -4 -6 20 206
use BUFX2  _58_
timestamp 1594572398
transform 1 0 824 0 -1 610
box -4 -6 52 206
use BUFX2  _61_
timestamp 1594572398
transform 1 0 872 0 -1 610
box -4 -6 52 206
use BUFX2  _63_
timestamp 1594572398
transform 1 0 920 0 -1 610
box -4 -6 52 206
use BUFX2  _57_
timestamp 1594572398
transform 1 0 968 0 -1 610
box -4 -6 52 206
use BUFX2  _55_
timestamp 1594572398
transform 1 0 1016 0 -1 610
box -4 -6 52 206
<< labels >>
flabel metal4 s 736 -10 800 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 272 -10 336 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal3 s 1101 537 1107 543 3 FreeSans 24 0 0 0 adrs_ctrl
port 2 nsew
flabel metal3 s -35 137 -29 143 7 FreeSans 24 0 0 0 clock
port 3 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 decoder_en
port 4 nsew
flabel metal3 s -35 317 -29 323 7 FreeSans 24 0 0 0 flag
port 5 nsew
flabel metal3 s 1101 497 1107 503 3 FreeSans 24 0 0 0 imm_en
port 6 nsew
flabel metal2 s 845 657 851 663 3 FreeSans 24 90 0 0 inst_wr
port 7 nsew
flabel metal3 s -35 357 -29 363 7 FreeSans 24 0 0 0 mem_rd
port 8 nsew
flabel metal2 s 557 -23 563 -17 7 FreeSans 24 270 0 0 mem_wr
port 9 nsew
flabel metal3 s 1101 297 1107 303 3 FreeSans 24 0 0 0 opcode[3]
port 10 nsew
flabel metal3 s 1101 117 1107 123 3 FreeSans 24 0 0 0 opcode[2]
port 11 nsew
flabel metal3 s 1101 157 1107 163 3 FreeSans 24 0 0 0 opcode[1]
port 12 nsew
flabel metal2 s 957 -23 963 -17 7 FreeSans 24 270 0 0 opcode[0]
port 13 nsew
flabel metal2 s 685 657 691 663 3 FreeSans 24 90 0 0 pc_op[1]
port 14 nsew
flabel metal2 s 893 657 899 663 3 FreeSans 24 90 0 0 pc_op[0]
port 15 nsew
flabel metal2 s 941 657 947 663 3 FreeSans 24 90 0 0 rD_wr
port 16 nsew
flabel metal2 s 701 -23 707 -17 7 FreeSans 24 270 0 0 reg_en
port 17 nsew
flabel metal3 s -35 277 -29 283 7 FreeSans 24 0 0 0 reset
port 18 nsew
<< end >>
