magic
tech scmos
magscale 1 2
timestamp 1596991774
<< metal1 >>
rect 2938 5414 2950 5416
rect 5946 5414 5958 5416
rect 2923 5406 2925 5414
rect 2933 5406 2935 5414
rect 2943 5406 2945 5414
rect 2953 5406 2955 5414
rect 2963 5406 2965 5414
rect 5931 5406 5933 5414
rect 5941 5406 5943 5414
rect 5951 5406 5953 5414
rect 5961 5406 5963 5414
rect 5971 5406 5973 5414
rect 2938 5404 2950 5406
rect 5946 5404 5958 5406
rect 2884 5377 2931 5383
rect 2157 5357 2195 5363
rect 2461 5357 2499 5363
rect 180 5337 195 5343
rect 676 5337 691 5343
rect 781 5337 796 5343
rect 829 5337 844 5343
rect 1101 5337 1116 5343
rect 1789 5337 1804 5343
rect 2845 5337 2892 5343
rect 3100 5337 3124 5343
rect 3741 5343 3747 5363
rect 5165 5357 5203 5363
rect 3741 5337 3779 5343
rect 4036 5337 4051 5343
rect 4861 5337 4876 5343
rect 5469 5343 5475 5363
rect 5437 5337 5475 5343
rect 340 5317 355 5323
rect 1053 5317 1068 5323
rect 1133 5317 1171 5323
rect 2621 5317 2668 5323
rect 2733 5317 2748 5323
rect 2765 5317 2803 5323
rect 2829 5317 2908 5323
rect 781 5297 803 5303
rect 861 5297 876 5303
rect 2797 5297 2803 5317
rect 3181 5317 3196 5323
rect 4013 5317 4051 5323
rect 2820 5296 2828 5304
rect 4045 5297 4051 5317
rect 4333 5317 4396 5323
rect 4861 5317 4899 5323
rect 4269 5297 4307 5303
rect 4861 5297 4867 5317
rect 5940 5297 6003 5303
rect 1194 5276 1196 5284
rect 2086 5276 2092 5284
rect 2390 5276 2396 5284
rect 5062 5276 5068 5284
rect 314 5236 316 5244
rect 2596 5236 2598 5244
rect 2698 5236 2700 5244
rect 1434 5214 1446 5216
rect 4442 5214 4454 5216
rect 1419 5206 1421 5214
rect 1429 5206 1431 5214
rect 1439 5206 1441 5214
rect 1449 5206 1451 5214
rect 1459 5206 1461 5214
rect 4427 5206 4429 5214
rect 4437 5206 4439 5214
rect 4447 5206 4449 5214
rect 4457 5206 4459 5214
rect 4467 5206 4469 5214
rect 1434 5204 1446 5206
rect 4442 5204 4454 5206
rect 4100 5176 4102 5184
rect 4298 5176 4300 5184
rect 122 5136 124 5144
rect 1588 5137 1619 5143
rect 2989 5137 3004 5143
rect 5492 5136 5494 5144
rect 5812 5136 5814 5144
rect 13 5097 67 5103
rect 77 5097 108 5103
rect 189 5097 204 5103
rect 381 5103 387 5123
rect 372 5097 387 5103
rect 413 5097 460 5103
rect 516 5097 531 5103
rect 669 5103 675 5123
rect 820 5116 828 5124
rect 1044 5116 1052 5124
rect 1373 5117 1388 5123
rect 1533 5117 1555 5123
rect 1613 5117 1635 5123
rect 669 5097 707 5103
rect 1005 5097 1036 5103
rect 1261 5097 1299 5103
rect 1677 5097 1692 5103
rect 1933 5097 1964 5103
rect 2173 5097 2188 5103
rect 3117 5103 3123 5123
rect 3085 5097 3123 5103
rect 3252 5097 3299 5103
rect 3517 5097 3571 5103
rect 3581 5097 3596 5103
rect 3812 5097 3843 5103
rect 3853 5097 3900 5103
rect 4125 5103 4131 5123
rect 4228 5116 4236 5124
rect 4125 5097 4163 5103
rect 4397 5097 4508 5103
rect 4653 5103 4659 5123
rect 5876 5116 5884 5124
rect 4621 5097 4659 5103
rect 5277 5097 5292 5103
rect 6100 5097 6115 5103
rect 6180 5097 6195 5103
rect 6356 5097 6371 5103
rect 6436 5097 6483 5103
rect 7076 5097 7091 5103
rect 7268 5097 7283 5103
rect 205 5077 220 5083
rect 429 5077 444 5083
rect 1156 5077 1176 5083
rect 1556 5077 1571 5083
rect 1581 5077 1603 5083
rect 1597 5064 1603 5077
rect 1693 5077 1708 5083
rect 1869 5077 1907 5083
rect 1917 5077 1948 5083
rect 1869 5057 1875 5077
rect 2372 5077 2387 5083
rect 2796 5077 2820 5083
rect 3012 5077 3075 5083
rect 3245 5077 3276 5083
rect 3933 5077 3955 5083
rect 4036 5077 4051 5083
rect 4420 5077 4515 5083
rect 5316 5076 5318 5084
rect 5388 5077 5411 5083
rect 5453 5077 5475 5083
rect 5533 5077 5548 5083
rect 5388 5072 5396 5077
rect 6084 5077 6099 5083
rect 6573 5077 6611 5083
rect 2045 5057 2060 5063
rect 2349 5057 2371 5063
rect 3322 5056 3324 5064
rect 5596 5063 5604 5066
rect 5117 5057 5155 5063
rect 5581 5057 5604 5063
rect 6605 5057 6611 5077
rect 234 5036 236 5044
rect 1642 5036 1644 5044
rect 3764 5036 3766 5044
rect 4372 5036 4374 5044
rect 6404 5036 6406 5044
rect 2938 5014 2950 5016
rect 5946 5014 5958 5016
rect 2923 5006 2925 5014
rect 2933 5006 2935 5014
rect 2943 5006 2945 5014
rect 2953 5006 2955 5014
rect 2963 5006 2965 5014
rect 5931 5006 5933 5014
rect 5941 5006 5943 5014
rect 5951 5006 5953 5014
rect 5961 5006 5963 5014
rect 5971 5006 5973 5014
rect 2938 5004 2950 5006
rect 5946 5004 5958 5006
rect 474 4976 476 4984
rect 1412 4977 1475 4983
rect 1674 4976 1676 4984
rect 2228 4976 2230 4984
rect 244 4957 259 4963
rect 1261 4957 1276 4963
rect 1805 4944 1811 4963
rect 1837 4957 1859 4963
rect 2157 4957 2172 4963
rect 2925 4957 3011 4963
rect 4717 4957 4732 4963
rect 5389 4957 5427 4963
rect 5533 4957 5571 4963
rect 5748 4957 5763 4963
rect 6388 4957 6403 4963
rect 6772 4956 6774 4964
rect 7261 4957 7276 4963
rect 7309 4957 7324 4963
rect 61 4923 67 4943
rect 996 4937 1011 4943
rect 1293 4937 1331 4943
rect 1501 4937 1523 4943
rect 1517 4924 1523 4937
rect 3565 4937 3587 4943
rect 3636 4937 3651 4943
rect 3748 4937 3779 4943
rect 3917 4937 3932 4943
rect 3972 4937 3987 4943
rect 4877 4937 4892 4943
rect 5581 4943 5587 4956
rect 5581 4937 5603 4943
rect 5645 4937 5667 4943
rect 5773 4943 5779 4956
rect 5773 4937 5795 4943
rect 5805 4937 5836 4943
rect 6893 4937 6908 4943
rect 7197 4937 7235 4943
rect 52 4917 67 4923
rect 109 4917 124 4923
rect 189 4917 227 4923
rect 365 4917 403 4923
rect 813 4917 851 4923
rect 909 4917 931 4923
rect 973 4917 988 4923
rect 1885 4917 1900 4923
rect 2189 4917 2211 4923
rect 2269 4917 2291 4923
rect 2397 4917 2451 4923
rect 2884 4917 2899 4923
rect 3053 4917 3068 4923
rect 3396 4917 3411 4923
rect 3428 4917 3459 4923
rect 93 4897 115 4903
rect 770 4896 780 4904
rect 1389 4897 1468 4903
rect 3453 4897 3459 4917
rect 3901 4917 3955 4923
rect 4013 4917 4060 4923
rect 4205 4917 4220 4923
rect 4301 4917 4316 4923
rect 4500 4917 4515 4923
rect 4836 4917 4851 4923
rect 4884 4917 4899 4923
rect 5149 4917 5164 4923
rect 7197 4924 7203 4937
rect 5940 4917 5996 4923
rect 6013 4917 6067 4923
rect 6189 4917 6220 4923
rect 6276 4917 6307 4923
rect 6365 4917 6396 4923
rect 6452 4917 6467 4923
rect 6557 4917 6588 4923
rect 6797 4917 6812 4923
rect 7060 4917 7091 4923
rect 3876 4896 3886 4904
rect 4516 4896 4524 4904
rect 4541 4897 4579 4903
rect 1844 4877 1859 4883
rect 5684 4876 5686 4884
rect 6468 4876 6470 4884
rect 1732 4856 1734 4864
rect 1194 4836 1196 4844
rect 1242 4836 1244 4844
rect 1604 4836 1606 4844
rect 2372 4836 2374 4844
rect 3546 4836 3548 4844
rect 4068 4836 4070 4844
rect 4180 4836 4182 4844
rect 4772 4836 4774 4844
rect 6164 4836 6166 4844
rect 1434 4814 1446 4816
rect 4442 4814 4454 4816
rect 1419 4806 1421 4814
rect 1429 4806 1431 4814
rect 1439 4806 1441 4814
rect 1449 4806 1451 4814
rect 1459 4806 1461 4814
rect 4427 4806 4429 4814
rect 4437 4806 4439 4814
rect 4447 4806 4449 4814
rect 4457 4806 4459 4814
rect 4467 4806 4469 4814
rect 1434 4804 1446 4806
rect 4442 4804 4454 4806
rect 900 4776 902 4784
rect 2932 4777 2995 4783
rect 3716 4776 3718 4784
rect 5236 4776 5238 4784
rect 5933 4777 5980 4783
rect 5140 4756 5142 4764
rect 212 4737 227 4743
rect 2088 4736 2092 4744
rect 3430 4736 3436 4744
rect 4100 4737 4115 4743
rect 5066 4736 5068 4744
rect 6650 4736 6652 4744
rect 45 4717 67 4723
rect 141 4717 179 4723
rect 1101 4717 1123 4723
rect 1405 4717 1491 4723
rect 1860 4717 1875 4723
rect 125 4697 147 4703
rect 420 4697 435 4703
rect 701 4697 723 4703
rect 788 4697 803 4703
rect 925 4697 963 4703
rect 1101 4697 1116 4703
rect 1149 4697 1171 4703
rect 1229 4697 1251 4703
rect 1149 4684 1155 4697
rect 2244 4697 2259 4703
rect 3492 4697 3507 4703
rect 3629 4703 3635 4723
rect 3597 4697 3635 4703
rect 3741 4697 3795 4703
rect 4045 4703 4051 4723
rect 4045 4697 4083 4703
rect 4196 4697 4227 4703
rect 5037 4703 5043 4723
rect 5005 4697 5043 4703
rect 5188 4697 5203 4703
rect 5261 4697 5276 4703
rect 5837 4703 5843 4723
rect 5805 4697 5843 4703
rect 6317 4703 6323 4723
rect 6589 4717 6627 4723
rect 6285 4697 6323 4703
rect 7149 4697 7164 4703
rect 724 4677 739 4683
rect 861 4677 883 4683
rect 1261 4677 1283 4683
rect 1261 4664 1267 4677
rect 1565 4677 1580 4683
rect 1725 4677 1740 4683
rect 2893 4677 2940 4683
rect 3757 4677 3772 4683
rect 3812 4677 3827 4683
rect 3869 4677 3891 4683
rect 3885 4664 3891 4677
rect 4045 4677 4060 4683
rect 4284 4677 4308 4683
rect 5284 4677 5299 4683
rect 5828 4677 5843 4683
rect 6556 4677 6572 4683
rect 109 4657 124 4663
rect 1604 4656 1612 4664
rect 3901 4657 3939 4663
rect 36 4636 38 4644
rect 186 4636 188 4644
rect 1188 4636 1190 4644
rect 1316 4636 1320 4644
rect 1428 4637 1491 4643
rect 1546 4636 1548 4644
rect 1796 4636 1798 4644
rect 2938 4614 2950 4616
rect 5946 4614 5958 4616
rect 2923 4606 2925 4614
rect 2933 4606 2935 4614
rect 2943 4606 2945 4614
rect 2953 4606 2955 4614
rect 2963 4606 2965 4614
rect 5931 4606 5933 4614
rect 5941 4606 5943 4614
rect 5951 4606 5953 4614
rect 5961 4606 5963 4614
rect 5971 4606 5973 4614
rect 2938 4604 2950 4606
rect 5946 4604 5958 4606
rect 954 4576 956 4584
rect 2196 4576 2200 4584
rect 6740 4576 6742 4584
rect 285 4557 300 4563
rect 461 4543 467 4563
rect 573 4557 588 4563
rect 1556 4556 1564 4564
rect 4221 4557 4259 4563
rect 429 4537 467 4543
rect 980 4537 1011 4543
rect 1517 4537 1532 4543
rect 1604 4537 1635 4543
rect 1933 4537 1971 4543
rect 1988 4537 2003 4543
rect 2765 4537 2780 4543
rect 3836 4543 3844 4548
rect 3821 4537 3844 4543
rect 5101 4543 5107 4563
rect 5213 4543 5219 4563
rect 6052 4557 6067 4563
rect 5101 4537 5139 4543
rect 5181 4537 5219 4543
rect 5380 4536 5382 4544
rect 5949 4537 6035 4543
rect 84 4517 99 4523
rect 173 4517 211 4523
rect 877 4517 915 4523
rect 1229 4517 1244 4523
rect 1597 4517 1612 4523
rect 1652 4517 1667 4523
rect 1684 4517 1715 4523
rect 2077 4517 2108 4523
rect 2884 4517 2915 4523
rect 3693 4517 3747 4523
rect 4349 4517 4364 4523
rect 4372 4517 4403 4523
rect 4573 4517 4611 4523
rect 269 4497 284 4503
rect 541 4497 563 4503
rect 605 4497 627 4503
rect 1373 4497 1420 4503
rect 3309 4497 3347 4503
rect 4605 4497 4611 4517
rect 4756 4517 4787 4523
rect 4925 4517 4940 4523
rect 5156 4517 5171 4523
rect 5501 4517 5516 4523
rect 5581 4517 5596 4523
rect 5773 4517 5788 4523
rect 5868 4523 5876 4528
rect 5853 4517 5876 4523
rect 5853 4497 5859 4517
rect 5949 4523 5955 4537
rect 6269 4537 6291 4543
rect 7085 4543 7091 4563
rect 7085 4537 7123 4543
rect 7197 4543 7203 4563
rect 7140 4537 7171 4543
rect 7197 4537 7235 4543
rect 7341 4537 7404 4543
rect 5917 4517 5955 4523
rect 6004 4517 6019 4523
rect 6157 4517 6195 4523
rect 6205 4517 6220 4523
rect 6157 4497 6163 4517
rect 6317 4517 6355 4523
rect 6381 4517 6396 4523
rect 6349 4497 6355 4517
rect 6372 4496 6380 4504
rect 173 4477 188 4483
rect 516 4477 531 4483
rect 5892 4476 5894 4484
rect 6452 4476 6458 4484
rect 5828 4456 5830 4464
rect 6980 4456 6982 4464
rect 100 4436 102 4444
rect 314 4436 316 4444
rect 378 4436 380 4444
rect 5498 4436 5500 4444
rect 5556 4436 5558 4444
rect 6084 4436 6086 4444
rect 6884 4436 6886 4444
rect 1434 4414 1446 4416
rect 4442 4414 4454 4416
rect 1419 4406 1421 4414
rect 1429 4406 1431 4414
rect 1439 4406 1441 4414
rect 1449 4406 1451 4414
rect 1459 4406 1461 4414
rect 4427 4406 4429 4414
rect 4437 4406 4439 4414
rect 4447 4406 4449 4414
rect 4457 4406 4459 4414
rect 4467 4406 4469 4414
rect 1434 4404 1446 4406
rect 4442 4404 4454 4406
rect 4989 4337 5004 4343
rect 6884 4337 6899 4343
rect 852 4316 860 4324
rect 1165 4317 1187 4323
rect 1885 4317 1907 4323
rect 2253 4317 2275 4323
rect 2356 4317 2387 4323
rect 2397 4317 2419 4323
rect 4164 4316 4172 4324
rect 404 4297 419 4303
rect 493 4297 556 4303
rect 861 4297 876 4303
rect 1037 4297 1075 4303
rect 1684 4297 1699 4303
rect 1892 4297 1907 4303
rect 2061 4297 2076 4303
rect 2436 4297 2483 4303
rect 2621 4297 2636 4303
rect 2852 4297 2867 4303
rect 3533 4297 3548 4303
rect 3693 4297 3708 4303
rect 4173 4297 4188 4303
rect 4269 4297 4323 4303
rect 4877 4297 4892 4303
rect 5053 4303 5059 4323
rect 5812 4316 5820 4324
rect 5021 4297 5059 4303
rect 5421 4297 5436 4303
rect 5485 4297 5500 4303
rect 5821 4297 5836 4303
rect 5997 4303 6003 4323
rect 5916 4297 6003 4303
rect 6029 4297 6044 4303
rect 5916 4292 5924 4297
rect 6573 4303 6579 4323
rect 6541 4297 6579 4303
rect 6829 4303 6835 4323
rect 6829 4297 6867 4303
rect 7133 4303 7139 4323
rect 7156 4316 7164 4324
rect 6980 4297 7011 4303
rect 7101 4297 7139 4303
rect 7261 4297 7276 4303
rect 125 4277 147 4283
rect 157 4277 179 4283
rect 157 4264 163 4277
rect 212 4277 227 4283
rect 1172 4277 1187 4283
rect 1389 4277 1475 4283
rect 1389 4264 1395 4277
rect 1869 4277 1884 4283
rect 2029 4277 2067 4283
rect 2077 4277 2092 4283
rect 436 4256 444 4264
rect 1940 4256 1944 4264
rect 2077 4257 2083 4277
rect 2109 4277 2124 4283
rect 2349 4277 2371 4283
rect 2349 4264 2355 4277
rect 3322 4276 3324 4284
rect 3485 4277 3523 4283
rect 2324 4257 2339 4263
rect 3485 4257 3491 4277
rect 3709 4277 3731 4283
rect 3796 4277 3811 4283
rect 4189 4277 4211 4283
rect 4468 4277 4547 4283
rect 4596 4277 4611 4283
rect 5044 4277 5059 4283
rect 6180 4277 6211 4283
rect 6829 4277 6844 4283
rect 4956 4264 4964 4272
rect 196 4236 198 4244
rect 280 4236 284 4244
rect 584 4236 588 4244
rect 676 4236 680 4244
rect 1528 4236 1532 4244
rect 2996 4237 3011 4243
rect 5940 4237 5980 4243
rect 2938 4214 2950 4216
rect 5946 4214 5958 4216
rect 2923 4206 2925 4214
rect 2933 4206 2935 4214
rect 2943 4206 2945 4214
rect 2953 4206 2955 4214
rect 2963 4206 2965 4214
rect 5931 4206 5933 4214
rect 5941 4206 5943 4214
rect 5951 4206 5953 4214
rect 5961 4206 5963 4214
rect 5971 4206 5973 4214
rect 2938 4204 2950 4206
rect 5946 4204 5958 4206
rect 1604 4176 1608 4184
rect 2234 4176 2236 4184
rect 157 4157 172 4163
rect 2813 4157 2835 4163
rect 2941 4157 3027 4163
rect 4996 4157 5011 4163
rect 5252 4157 5267 4163
rect 5892 4157 5907 4163
rect 6941 4157 6979 4163
rect 109 4143 115 4156
rect 93 4137 115 4143
rect 212 4137 227 4143
rect 317 4137 348 4143
rect 381 4137 403 4143
rect 557 4137 588 4143
rect 660 4137 675 4143
rect 797 4137 812 4143
rect 1172 4137 1187 4143
rect 1348 4137 1363 4143
rect 1501 4137 1516 4143
rect 1924 4137 1939 4143
rect 2109 4137 2147 4143
rect 2637 4137 2652 4143
rect 2685 4137 2716 4143
rect 3117 4137 3148 4143
rect 3428 4137 3443 4143
rect 3565 4137 3596 4143
rect 3908 4137 3923 4143
rect 4221 4137 4236 4143
rect 4588 4143 4596 4148
rect 4445 4137 4531 4143
rect 4573 4137 4596 4143
rect 4973 4137 4988 4143
rect 5028 4137 5043 4143
rect 5085 4137 5100 4143
rect 5149 4137 5171 4143
rect 5229 4137 5244 4143
rect 5284 4137 5315 4143
rect 5676 4143 5684 4148
rect 5676 4137 5699 4143
rect 6173 4137 6188 4143
rect 6349 4137 6371 4143
rect 301 4117 316 4123
rect 781 4117 796 4123
rect 804 4117 835 4123
rect 845 4117 883 4123
rect 893 4117 908 4123
rect 1156 4117 1171 4123
rect 1389 4117 1404 4123
rect 29 4097 51 4103
rect 1165 4097 1171 4117
rect 1533 4117 1564 4123
rect 1725 4117 1740 4123
rect 1773 4117 1811 4123
rect 1805 4097 1811 4117
rect 1917 4117 1955 4123
rect 2205 4117 2227 4123
rect 2221 4104 2227 4117
rect 2260 4117 2275 4123
rect 3405 4117 3443 4123
rect 1997 4097 2019 4103
rect 2941 4097 2988 4103
rect 3437 4097 3443 4117
rect 3789 4117 3843 4123
rect 3924 4117 3939 4123
rect 4045 4117 4060 4123
rect 4317 4117 4332 4123
rect 4957 4117 4972 4123
rect 5405 4117 5443 4123
rect 5437 4097 5443 4117
rect 5773 4117 5827 4123
rect 6013 4117 6067 4123
rect 7028 4117 7043 4123
rect 5460 4096 5468 4104
rect 74 4076 76 4084
rect 596 4077 611 4083
rect 2029 4077 2044 4083
rect 4020 4076 4026 4084
rect 4628 4076 4634 4084
rect 6445 4077 6460 4083
rect 6516 4076 6522 4084
rect 5188 4056 5190 4064
rect 6234 4056 6236 4064
rect 186 4036 188 4044
rect 244 4036 246 4044
rect 1140 4036 1142 4044
rect 1284 4036 1288 4044
rect 3764 4036 3766 4044
rect 5828 4036 5830 4044
rect 6068 4036 6070 4044
rect 6308 4036 6310 4044
rect 1434 4014 1446 4016
rect 4442 4014 4454 4016
rect 1419 4006 1421 4014
rect 1429 4006 1431 4014
rect 1439 4006 1441 4014
rect 1449 4006 1451 4014
rect 1459 4006 1461 4014
rect 4427 4006 4429 4014
rect 4437 4006 4439 4014
rect 4447 4006 4449 4014
rect 4457 4006 4459 4014
rect 4467 4006 4469 4014
rect 1434 4004 1446 4006
rect 4442 4004 4454 4006
rect 3434 3976 3436 3984
rect 3530 3976 3532 3984
rect 3780 3976 3782 3984
rect 5933 3977 5996 3983
rect 4922 3956 4924 3964
rect 1588 3936 1590 3944
rect 4052 3936 4054 3944
rect 237 3883 243 3903
rect 308 3897 323 3903
rect 429 3897 444 3903
rect 580 3897 595 3903
rect 772 3897 787 3903
rect 989 3903 995 3923
rect 1076 3917 1091 3923
rect 2068 3917 2083 3923
rect 957 3897 995 3903
rect 2173 3903 2179 3923
rect 2173 3897 2211 3903
rect 2260 3897 2275 3903
rect 3133 3903 3139 3923
rect 3101 3897 3139 3903
rect 3261 3897 3292 3903
rect 3492 3897 3507 3903
rect 3572 3897 3603 3903
rect 4077 3903 4083 3923
rect 4077 3897 4115 3903
rect 4125 3897 4140 3903
rect 5069 3897 5084 3903
rect 5508 3897 5523 3903
rect 6804 3897 6819 3903
rect 7012 3897 7043 3903
rect 180 3877 195 3883
rect 205 3877 243 3883
rect 189 3857 195 3877
rect 276 3877 291 3883
rect 340 3877 371 3883
rect 557 3877 579 3883
rect 573 3864 579 3877
rect 813 3877 828 3883
rect 1101 3877 1116 3883
rect 228 3857 259 3863
rect 1101 3857 1107 3877
rect 1165 3877 1180 3883
rect 1373 3877 1388 3883
rect 1373 3857 1379 3877
rect 1556 3877 1571 3883
rect 1965 3877 1987 3883
rect 1997 3877 2019 3883
rect 1981 3864 1987 3877
rect 2120 3877 2147 3883
rect 3028 3877 3091 3883
rect 3124 3877 3139 3883
rect 4506 3876 4508 3884
rect 5021 3877 5043 3883
rect 5085 3877 5108 3883
rect 5100 3872 5108 3877
rect 5332 3877 5363 3883
rect 5677 3877 5692 3883
rect 6317 3877 6355 3883
rect 6381 3877 6396 3883
rect 3677 3857 3692 3863
rect 5309 3857 5347 3863
rect 5613 3857 5651 3863
rect 6349 3857 6355 3877
rect 6685 3877 6700 3883
rect 6861 3877 6899 3883
rect 6717 3857 6755 3863
rect 6861 3857 6867 3877
rect 7149 3877 7187 3883
rect 7357 3877 7388 3883
rect 72 3836 76 3844
rect 1002 3836 1004 3844
rect 1928 3836 1932 3844
rect 2356 3836 2360 3844
rect 2536 3836 2540 3844
rect 3005 3837 3020 3843
rect 2938 3814 2950 3816
rect 5946 3814 5958 3816
rect 2923 3806 2925 3814
rect 2933 3806 2935 3814
rect 2943 3806 2945 3814
rect 2953 3806 2955 3814
rect 2963 3806 2965 3814
rect 5931 3806 5933 3814
rect 5941 3806 5943 3814
rect 5951 3806 5953 3814
rect 5961 3806 5963 3814
rect 5971 3806 5973 3814
rect 2938 3804 2950 3806
rect 5946 3804 5958 3806
rect 968 3776 972 3784
rect 2116 3776 2120 3784
rect 5268 3776 5270 3784
rect 6596 3776 6598 3784
rect 125 3757 156 3763
rect 557 3757 579 3763
rect 1421 3757 1436 3763
rect 3325 3757 3363 3763
rect 3530 3756 3532 3764
rect 4221 3757 4236 3763
rect 260 3737 291 3743
rect 1005 3737 1020 3743
rect 1204 3737 1235 3743
rect 1661 3737 1699 3743
rect 2052 3737 2083 3743
rect 2900 3737 2980 3743
rect 5149 3737 5171 3743
rect 5316 3737 5347 3743
rect 5517 3743 5523 3763
rect 5517 3737 5555 3743
rect 5940 3737 6003 3743
rect 6468 3737 6483 3743
rect 6893 3743 6899 3763
rect 6861 3737 6899 3743
rect 7197 3743 7203 3763
rect 7197 3737 7235 3743
rect 845 3717 876 3723
rect 1444 3717 1507 3723
rect 1517 3717 1532 3723
rect 1581 3717 1596 3723
rect 1604 3717 1612 3723
rect 1748 3717 1763 3723
rect 2285 3717 2300 3723
rect 3213 3717 3251 3723
rect 205 3697 220 3703
rect 1572 3696 1580 3704
rect 3188 3696 3196 3704
rect 3213 3697 3219 3717
rect 3588 3717 3603 3723
rect 3741 3717 3779 3723
rect 3773 3697 3779 3717
rect 4157 3717 4172 3723
rect 4749 3717 4787 3723
rect 4781 3697 4787 3717
rect 4932 3717 4963 3723
rect 5197 3717 5212 3723
rect 5293 3717 5340 3723
rect 6093 3717 6147 3723
rect 6285 3717 6339 3723
rect 6380 3723 6388 3728
rect 6380 3717 6403 3723
rect 6397 3697 6403 3717
rect 6468 3717 6483 3723
rect 429 3677 444 3683
rect 2189 3677 2204 3683
rect 3802 3676 3804 3684
rect 4052 3676 4054 3684
rect 4634 3676 4636 3684
rect 6426 3676 6428 3684
rect 6340 3656 6342 3664
rect 346 3636 348 3644
rect 1160 3636 1164 3644
rect 1300 3636 1304 3644
rect 1642 3636 1644 3644
rect 1722 3636 1724 3644
rect 2340 3636 2344 3644
rect 3434 3636 3436 3644
rect 3604 3636 3606 3644
rect 3668 3636 3670 3644
rect 4154 3636 4156 3644
rect 5860 3636 5862 3644
rect 1434 3614 1446 3616
rect 4442 3614 4454 3616
rect 1419 3606 1421 3614
rect 1429 3606 1431 3614
rect 1439 3606 1441 3614
rect 1449 3606 1451 3614
rect 1459 3606 1461 3614
rect 4427 3606 4429 3614
rect 4437 3606 4439 3614
rect 4447 3606 4449 3614
rect 4457 3606 4459 3614
rect 4467 3606 4469 3614
rect 1434 3604 1446 3606
rect 4442 3604 4454 3606
rect 2900 3577 2931 3583
rect 3940 3576 3942 3584
rect 4036 3576 4038 3584
rect 4858 3576 4860 3584
rect 244 3556 246 3564
rect 541 3537 556 3543
rect 1764 3536 1766 3544
rect 2468 3537 2483 3543
rect 3466 3536 3468 3544
rect 3700 3536 3702 3544
rect 4564 3536 4566 3544
rect 29 3517 51 3523
rect 852 3516 860 3524
rect 1412 3517 1491 3523
rect 436 3497 451 3503
rect 637 3497 684 3503
rect 813 3497 828 3503
rect 2372 3497 2387 3503
rect 2813 3503 2819 3523
rect 2765 3497 2819 3503
rect 93 3477 108 3483
rect 164 3477 179 3483
rect 205 3477 227 3483
rect 573 3477 595 3483
rect 733 3477 755 3483
rect 893 3477 915 3483
rect 957 3477 979 3483
rect 1341 3477 1363 3483
rect 1517 3477 1532 3483
rect 1661 3477 1699 3483
rect 1725 3477 1740 3483
rect 148 3457 163 3463
rect 797 3457 812 3463
rect 1405 3457 1436 3463
rect 1725 3457 1731 3477
rect 1837 3477 1864 3483
rect 2061 3483 2067 3496
rect 3220 3497 3235 3503
rect 3412 3497 3443 3503
rect 6100 3497 6115 3503
rect 6461 3497 6476 3503
rect 6692 3497 6707 3503
rect 2045 3477 2067 3483
rect 2125 3477 2147 3483
rect 2349 3477 2371 3483
rect 2429 3477 2451 3483
rect 2685 3477 2700 3483
rect 3100 3477 3124 3483
rect 3805 3477 3843 3483
rect 3869 3477 3884 3483
rect 2020 3456 2028 3464
rect 2317 3457 2339 3463
rect 3357 3457 3395 3463
rect 3837 3457 3843 3477
rect 4605 3477 4627 3483
rect 5412 3477 5427 3483
rect 5437 3477 5452 3483
rect 5741 3477 5779 3483
rect 4436 3457 4499 3463
rect 4989 3457 5027 3463
rect 5261 3457 5299 3463
rect 5373 3457 5411 3463
rect 5773 3457 5779 3477
rect 6012 3477 6099 3483
rect 6012 3472 6020 3477
rect 6532 3477 6563 3483
rect 6708 3477 6723 3483
rect 6765 3483 6771 3503
rect 6756 3477 6771 3483
rect 7181 3483 7187 3503
rect 7284 3497 7299 3503
rect 7165 3477 7187 3483
rect 7197 3477 7235 3483
rect 6509 3457 6547 3463
rect 6749 3457 6787 3463
rect 7229 3457 7235 3477
rect 7341 3457 7379 3463
rect 1498 3436 1500 3444
rect 1572 3436 1576 3444
rect 1818 3436 1820 3444
rect 2564 3436 2568 3444
rect 2826 3436 2828 3444
rect 4772 3436 4774 3444
rect 6196 3436 6198 3444
rect 2938 3414 2950 3416
rect 5946 3414 5958 3416
rect 2923 3406 2925 3414
rect 2933 3406 2935 3414
rect 2943 3406 2945 3414
rect 2953 3406 2955 3414
rect 2963 3406 2965 3414
rect 5931 3406 5933 3414
rect 5941 3406 5943 3414
rect 5951 3406 5953 3414
rect 5961 3406 5963 3414
rect 5971 3406 5973 3414
rect 2938 3404 2950 3406
rect 5946 3404 5958 3406
rect 116 3376 118 3384
rect 1444 3377 1507 3383
rect 1674 3376 1676 3384
rect 3005 3377 3027 3383
rect 212 3356 220 3364
rect 397 3357 435 3363
rect 61 3337 99 3343
rect 253 3343 259 3356
rect 237 3337 259 3343
rect 452 3337 467 3343
rect 605 3337 627 3343
rect 813 3337 835 3343
rect 925 3337 963 3343
rect 1133 3337 1155 3343
rect 1565 3337 1603 3343
rect 1885 3343 1891 3363
rect 2173 3357 2195 3363
rect 2237 3357 2252 3363
rect 2269 3357 2307 3363
rect 3021 3363 3027 3377
rect 5044 3376 5046 3384
rect 3021 3357 3084 3363
rect 3101 3357 3139 3363
rect 3629 3357 3667 3363
rect 4868 3357 4883 3363
rect 5228 3348 5236 3356
rect 1853 3337 1891 3343
rect 2292 3337 2323 3343
rect 4813 3337 4828 3343
rect 4916 3337 4931 3343
rect 5092 3337 5123 3343
rect 5885 3337 5964 3343
rect 6221 3337 6243 3343
rect 29 3317 51 3323
rect 300 3323 308 3328
rect 189 3317 227 3323
rect 285 3317 308 3323
rect 189 3297 195 3317
rect 349 3317 371 3323
rect 733 3317 748 3323
rect 868 3317 883 3323
rect 1028 3317 1043 3323
rect 1053 3317 1068 3323
rect 1629 3317 1667 3323
rect 772 3296 780 3304
rect 1092 3296 1100 3304
rect 1661 3297 1667 3317
rect 1917 3317 1939 3323
rect 2084 3317 2099 3323
rect 2333 3317 2355 3323
rect 2893 3317 2908 3323
rect 3261 3317 3276 3323
rect 3300 3317 3315 3323
rect 3469 3317 3484 3323
rect 4317 3317 4355 3323
rect 4317 3297 4323 3317
rect 4388 3317 4403 3323
rect 4413 3317 4531 3323
rect 4572 3323 4580 3328
rect 4572 3317 4595 3323
rect 4589 3297 4595 3317
rect 4797 3317 4812 3323
rect 5069 3317 5116 3323
rect 6653 3317 6668 3323
rect 6861 3317 6876 3323
rect 7268 3317 7299 3323
rect 6701 3297 6739 3303
rect 6756 3296 6764 3304
rect 532 3277 563 3283
rect 573 3277 588 3283
rect 1364 3277 1379 3283
rect 4970 3276 4972 3284
rect 58 3236 60 3244
rect 164 3236 166 3244
rect 3434 3236 3436 3244
rect 6004 3236 6006 3244
rect 6100 3236 6102 3244
rect 6628 3236 6630 3244
rect 1434 3214 1446 3216
rect 4442 3214 4454 3216
rect 1419 3206 1421 3214
rect 1429 3206 1431 3214
rect 1439 3206 1441 3214
rect 1449 3206 1451 3214
rect 1459 3206 1461 3214
rect 4427 3206 4429 3214
rect 4437 3206 4439 3214
rect 4447 3206 4449 3214
rect 4457 3206 4459 3214
rect 4467 3206 4469 3214
rect 1434 3204 1446 3206
rect 4442 3204 4454 3206
rect 36 3176 38 3184
rect 1101 3143 1107 3163
rect 1101 3137 1139 3143
rect 61 3103 67 3123
rect 685 3117 700 3123
rect 1133 3117 1139 3137
rect 1908 3137 1955 3143
rect 3300 3136 3306 3144
rect 5060 3137 5075 3143
rect 6916 3136 6918 3144
rect 2370 3116 2380 3124
rect 61 3097 99 3103
rect 132 3097 147 3103
rect 820 3097 835 3103
rect 1005 3097 1027 3103
rect 164 3077 179 3083
rect 1021 3077 1027 3097
rect 1117 3077 1123 3108
rect 1757 3097 1772 3103
rect 2100 3097 2115 3103
rect 2253 3097 2275 3103
rect 1245 3077 1260 3083
rect 1284 3077 1299 3083
rect 1565 3077 1587 3083
rect 1789 3077 1811 3083
rect 1869 3077 1891 3083
rect 2253 3077 2259 3097
rect 2877 3097 2892 3103
rect 2909 3097 2988 3103
rect 3053 3097 3075 3103
rect 3501 3097 3516 3103
rect 3741 3103 3747 3123
rect 3709 3097 3747 3103
rect 4205 3103 4211 3123
rect 4444 3103 4452 3106
rect 4205 3097 4243 3103
rect 4444 3097 4547 3103
rect 5005 3103 5011 3123
rect 5005 3097 5043 3103
rect 5268 3097 5283 3103
rect 5732 3097 5747 3103
rect 6269 3103 6275 3123
rect 6237 3097 6275 3103
rect 6925 3097 6940 3103
rect 6973 3097 7027 3103
rect 2397 3077 2419 3083
rect 2637 3077 2652 3083
rect 765 3057 780 3063
rect 1741 3057 1756 3063
rect 1901 3057 1923 3063
rect 1988 3056 1996 3064
rect 2429 3057 2451 3063
rect 232 3036 236 3044
rect 468 3037 483 3043
rect 532 3037 547 3043
rect 884 3036 886 3044
rect 1338 3036 1340 3044
rect 1421 3037 1484 3043
rect 2045 3037 2060 3043
rect 2445 3037 2451 3057
rect 2637 3057 2643 3077
rect 2781 3077 2819 3083
rect 2932 3077 3027 3083
rect 3076 3077 3091 3083
rect 3117 3077 3155 3083
rect 3517 3077 3539 3083
rect 3869 3077 3907 3083
rect 2836 3057 2851 3063
rect 2980 3057 3011 3063
rect 3901 3057 3907 3077
rect 3956 3077 3971 3083
rect 4205 3077 4220 3083
rect 5405 3077 5443 3083
rect 5405 3057 5411 3077
rect 5476 3077 5491 3083
rect 6068 3077 6083 3083
rect 7101 3083 7107 3103
rect 7101 3077 7132 3083
rect 5901 3057 5980 3063
rect 7085 3057 7100 3063
rect 2552 3036 2556 3044
rect 3114 3036 3116 3044
rect 2938 3014 2950 3016
rect 5946 3014 5958 3016
rect 2923 3006 2925 3014
rect 2933 3006 2935 3014
rect 2943 3006 2945 3014
rect 2953 3006 2955 3014
rect 2963 3006 2965 3014
rect 5931 3006 5933 3014
rect 5941 3006 5943 3014
rect 5951 3006 5953 3014
rect 5961 3006 5963 3014
rect 5971 3006 5973 3014
rect 2938 3004 2950 3006
rect 5946 3004 5958 3006
rect 3258 2976 3260 2984
rect 52 2957 67 2963
rect 125 2957 163 2963
rect 109 2937 124 2943
rect 237 2943 243 2963
rect 1524 2956 1532 2964
rect 2868 2957 2883 2963
rect 3341 2957 3363 2963
rect 3469 2957 3491 2963
rect 3693 2957 3731 2963
rect 4156 2957 4179 2963
rect 4189 2957 4227 2963
rect 4156 2954 4164 2957
rect 6141 2957 6164 2963
rect 6156 2954 6164 2957
rect 6980 2957 6995 2963
rect 7005 2957 7027 2963
rect 4924 2944 4932 2948
rect 5452 2944 5460 2948
rect 205 2937 243 2943
rect 573 2937 595 2943
rect 45 2917 67 2923
rect 180 2917 195 2923
rect 548 2917 563 2923
rect 701 2912 707 2943
rect 829 2912 835 2943
rect 1021 2937 1036 2943
rect 1117 2912 1123 2943
rect 1277 2937 1292 2943
rect 1357 2912 1363 2943
rect 1549 2937 1564 2943
rect 2068 2937 2083 2943
rect 2125 2937 2147 2943
rect 1709 2917 1724 2923
rect 2125 2917 2131 2937
rect 2429 2937 2444 2943
rect 2525 2937 2547 2943
rect 2189 2917 2204 2923
rect 2468 2917 2483 2923
rect 2605 2923 2611 2943
rect 2669 2937 2684 2943
rect 3964 2937 3988 2943
rect 4228 2937 4243 2943
rect 4996 2937 5011 2943
rect 5668 2937 5683 2943
rect 6388 2937 6403 2943
rect 6436 2937 6451 2943
rect 6957 2937 6995 2943
rect 7293 2943 7299 2963
rect 7284 2937 7299 2943
rect 2605 2917 2627 2923
rect 2749 2917 2780 2923
rect 2845 2917 2915 2923
rect 3284 2917 3315 2923
rect 3348 2917 3363 2923
rect 4829 2917 4844 2923
rect 4973 2917 5011 2923
rect 285 2883 291 2903
rect 580 2897 595 2903
rect 269 2877 291 2883
rect 596 2877 627 2883
rect 669 2877 700 2883
rect 845 2883 851 2903
rect 813 2877 851 2883
rect 813 2857 819 2877
rect 1101 2883 1107 2903
rect 1101 2877 1139 2883
rect 1133 2857 1139 2877
rect 1373 2883 1379 2903
rect 1981 2897 1996 2903
rect 2484 2896 2492 2904
rect 4724 2896 4732 2904
rect 5005 2897 5011 2917
rect 5133 2917 5187 2923
rect 5309 2917 5324 2923
rect 5645 2917 5683 2923
rect 5677 2897 5683 2917
rect 6381 2917 6396 2923
rect 6413 2917 6451 2923
rect 6445 2897 6451 2917
rect 6756 2917 6787 2923
rect 7124 2917 7139 2923
rect 6573 2897 6611 2903
rect 6628 2896 6636 2904
rect 1341 2877 1379 2883
rect 1341 2857 1347 2877
rect 1844 2877 1907 2883
rect 3828 2876 3834 2884
rect 4330 2876 4332 2884
rect 4941 2877 4956 2883
rect 5188 2876 5190 2884
rect 6004 2877 6067 2883
rect 7069 2877 7084 2883
rect 7236 2877 7251 2883
rect 7373 2877 7404 2883
rect 3044 2837 3059 2843
rect 5818 2836 5820 2844
rect 6122 2836 6124 2844
rect 1434 2814 1446 2816
rect 4442 2814 4454 2816
rect 1419 2806 1421 2814
rect 1429 2806 1431 2814
rect 1439 2806 1441 2814
rect 1449 2806 1451 2814
rect 1459 2806 1461 2814
rect 4427 2806 4429 2814
rect 4437 2806 4439 2814
rect 4447 2806 4449 2814
rect 4457 2806 4459 2814
rect 4467 2806 4469 2814
rect 1434 2804 1446 2806
rect 4442 2804 4454 2806
rect 154 2776 156 2784
rect 4324 2776 4326 2784
rect 4516 2776 4518 2784
rect 5242 2776 5244 2784
rect 5428 2776 5430 2784
rect 1322 2756 1324 2764
rect 445 2737 460 2743
rect 1101 2737 1148 2743
rect 1380 2737 1395 2743
rect 1805 2737 1820 2743
rect 3085 2737 3116 2743
rect 3981 2737 3996 2743
rect 4250 2736 4252 2744
rect 6836 2736 6842 2744
rect 1245 2717 1260 2723
rect 2861 2717 2963 2723
rect 3172 2716 3176 2724
rect 205 2697 220 2703
rect 365 2677 371 2708
rect 388 2677 404 2683
rect 477 2677 483 2708
rect 541 2677 547 2708
rect 628 2697 643 2703
rect 396 2676 404 2677
rect 941 2677 956 2683
rect 1100 2677 1116 2683
rect 1100 2676 1108 2677
rect 1357 2677 1363 2708
rect 1581 2677 1587 2708
rect 1645 2677 1651 2708
rect 1709 2677 1715 2708
rect 2141 2677 2147 2708
rect 2269 2677 2275 2708
rect 2317 2697 2332 2703
rect 2484 2697 2499 2703
rect 2564 2697 2579 2703
rect 2589 2697 2659 2703
rect 3005 2697 3075 2703
rect 4045 2703 4051 2723
rect 4578 2716 4588 2724
rect 5796 2716 5804 2724
rect 6180 2716 6188 2724
rect 4013 2697 4051 2703
rect 4077 2697 4092 2703
rect 4189 2697 4204 2703
rect 4525 2697 4540 2703
rect 4669 2697 4691 2703
rect 4532 2677 4547 2683
rect 4669 2683 4675 2697
rect 4861 2697 4876 2703
rect 4957 2697 4972 2703
rect 4996 2697 5011 2703
rect 5101 2697 5155 2703
rect 5252 2697 5276 2703
rect 6148 2697 6179 2703
rect 4660 2677 4675 2683
rect 4804 2677 4819 2683
rect 4980 2677 5011 2683
rect 6141 2677 6163 2683
rect 6253 2677 6268 2683
rect 6733 2677 6771 2683
rect 573 2657 588 2663
rect 685 2657 700 2663
rect 1613 2657 1628 2663
rect 1933 2657 1948 2663
rect 2324 2657 2339 2663
rect 3037 2657 3052 2663
rect 3293 2657 3315 2663
rect 3421 2657 3443 2663
rect 3709 2657 3747 2663
rect 4388 2657 4403 2663
rect 4420 2657 4499 2663
rect 5293 2657 5331 2663
rect 6733 2657 6739 2677
rect 6796 2663 6804 2666
rect 6788 2657 6804 2663
rect 6828 2663 6836 2672
rect 6828 2657 6860 2663
rect 72 2636 76 2644
rect 280 2636 284 2644
rect 1288 2636 1292 2644
rect 2173 2637 2188 2643
rect 2420 2636 2424 2644
rect 2756 2636 2760 2644
rect 2861 2637 2876 2643
rect 5524 2636 5526 2644
rect 2938 2614 2950 2616
rect 5946 2614 5958 2616
rect 2923 2606 2925 2614
rect 2933 2606 2935 2614
rect 2943 2606 2945 2614
rect 2953 2606 2955 2614
rect 2963 2606 2965 2614
rect 5931 2606 5933 2614
rect 5941 2606 5943 2614
rect 5951 2606 5953 2614
rect 5961 2606 5963 2614
rect 5971 2606 5973 2614
rect 2938 2604 2950 2606
rect 5946 2604 5958 2606
rect 109 2557 147 2563
rect 781 2557 796 2563
rect 1053 2563 1059 2583
rect 1213 2563 1219 2583
rect 2488 2576 2492 2584
rect 2600 2576 2604 2584
rect 2925 2577 2988 2583
rect 3096 2576 3100 2584
rect 4445 2577 4508 2583
rect 1053 2557 1075 2563
rect 1197 2557 1219 2563
rect 4013 2557 4051 2563
rect 6269 2557 6307 2563
rect 5276 2548 5284 2556
rect 164 2537 179 2543
rect 893 2537 915 2543
rect 973 2537 995 2543
rect 1037 2537 1052 2543
rect 1085 2537 1107 2543
rect 1165 2537 1187 2543
rect 1220 2537 1235 2543
rect 1277 2537 1299 2543
rect 1341 2537 1356 2543
rect 1581 2537 1603 2543
rect 1661 2537 1683 2543
rect 1949 2537 1971 2543
rect 541 2517 556 2523
rect 573 2517 588 2523
rect 797 2517 812 2523
rect 1300 2517 1315 2523
rect 1341 2517 1379 2523
rect 836 2496 844 2504
rect 1341 2497 1347 2517
rect 2141 2512 2147 2543
rect 2228 2517 2243 2523
rect 2893 2523 2899 2543
rect 4381 2537 4396 2543
rect 5780 2537 5795 2543
rect 6148 2537 6163 2543
rect 6317 2543 6323 2556
rect 6317 2537 6339 2543
rect 6381 2537 6403 2543
rect 7133 2537 7155 2543
rect 2884 2517 2899 2523
rect 3565 2517 3580 2523
rect 3716 2517 3731 2523
rect 4093 2517 4108 2523
rect 4365 2517 4380 2523
rect 4828 2523 4836 2528
rect 4813 2517 4836 2523
rect 1933 2497 1971 2503
rect 4356 2496 4364 2504
rect 4445 2497 4524 2503
rect 4628 2496 4636 2504
rect 4813 2497 4819 2517
rect 5060 2517 5091 2523
rect 5156 2517 5171 2523
rect 5309 2517 5324 2523
rect 5348 2517 5363 2523
rect 7133 2524 7139 2537
rect 5757 2517 5795 2523
rect 5821 2517 5884 2523
rect 4868 2496 4876 2504
rect 5460 2496 5468 2504
rect 5789 2497 5795 2517
rect 5981 2517 5996 2523
rect 6125 2517 6163 2523
rect 6157 2497 6163 2517
rect 6340 2517 6355 2523
rect 6388 2517 6419 2523
rect 6628 2517 6659 2523
rect 6765 2517 6780 2523
rect 7341 2517 7372 2523
rect 6596 2496 6604 2504
rect 7236 2496 7244 2504
rect 7309 2497 7324 2503
rect 1844 2476 1846 2484
rect 2840 2476 2844 2484
rect 6093 2477 6108 2483
rect 4186 2436 4188 2444
rect 4708 2436 4710 2444
rect 5012 2436 5014 2444
rect 6420 2436 6422 2444
rect 1434 2414 1446 2416
rect 4442 2414 4454 2416
rect 1419 2406 1421 2414
rect 1429 2406 1431 2414
rect 1439 2406 1441 2414
rect 1449 2406 1451 2414
rect 1459 2406 1461 2414
rect 4427 2406 4429 2414
rect 4437 2406 4439 2414
rect 4447 2406 4449 2414
rect 4457 2406 4459 2414
rect 4467 2406 4469 2414
rect 1434 2404 1446 2406
rect 4442 2404 4454 2406
rect 1060 2376 1062 2384
rect 1940 2376 1942 2384
rect 2744 2376 2748 2384
rect 4932 2356 4934 2364
rect 554 2336 556 2344
rect 1178 2336 1180 2344
rect 2612 2337 2627 2343
rect 4589 2337 4604 2343
rect 5258 2336 5260 2344
rect 5610 2336 5612 2344
rect 61 2303 67 2323
rect 141 2317 163 2323
rect 381 2317 396 2323
rect 852 2316 860 2324
rect 52 2297 67 2303
rect 285 2297 316 2303
rect 29 2277 60 2283
rect 125 2277 140 2283
rect 461 2277 467 2308
rect 484 2277 500 2283
rect 492 2276 500 2277
rect 589 2277 595 2308
rect 756 2297 771 2303
rect 877 2303 883 2323
rect 4100 2316 4108 2324
rect 877 2297 915 2303
rect 1437 2297 1523 2303
rect 1581 2297 1619 2303
rect 813 2277 835 2283
rect 952 2277 972 2283
rect 1021 2277 1043 2283
rect 1197 2277 1219 2283
rect 1261 2277 1283 2283
rect 1357 2277 1379 2283
rect 1437 2277 1443 2297
rect 1949 2297 2012 2303
rect 3380 2297 3395 2303
rect 4125 2303 4131 2323
rect 4125 2297 4163 2303
rect 4653 2303 4659 2323
rect 4621 2297 4659 2303
rect 4916 2297 4931 2303
rect 1645 2277 1667 2283
rect 1741 2277 1756 2283
rect 1933 2277 1964 2283
rect 2036 2276 2040 2284
rect 2093 2277 2131 2283
rect 781 2257 803 2263
rect 989 2257 1011 2263
rect 781 2237 787 2257
rect 1108 2257 1123 2263
rect 1565 2257 1580 2263
rect 1956 2257 1971 2263
rect 2093 2257 2099 2277
rect 2461 2277 2483 2283
rect 2676 2277 2691 2283
rect 3620 2277 3651 2283
rect 4644 2277 4659 2283
rect 5277 2277 5292 2283
rect 5373 2283 5379 2303
rect 5508 2297 5523 2303
rect 5764 2297 5779 2303
rect 6020 2297 6035 2303
rect 6413 2297 6428 2303
rect 6941 2297 6956 2303
rect 5373 2277 5388 2283
rect 5396 2277 5411 2283
rect 5549 2277 5571 2283
rect 5933 2277 6019 2283
rect 6340 2277 6355 2283
rect 7341 2277 7372 2283
rect 3373 2257 3395 2263
rect 3565 2257 3587 2263
rect 4285 2257 4323 2263
rect 4333 2257 4396 2263
rect 4989 2257 5027 2263
rect 5652 2257 5667 2263
rect 6292 2257 6307 2263
rect 6532 2257 6547 2263
rect 6589 2257 6627 2263
rect 2938 2214 2950 2216
rect 5946 2214 5958 2216
rect 2923 2206 2925 2214
rect 2933 2206 2935 2214
rect 2943 2206 2945 2214
rect 2953 2206 2955 2214
rect 2963 2206 2965 2214
rect 5931 2206 5933 2214
rect 5941 2206 5943 2214
rect 5951 2206 5953 2214
rect 5961 2206 5963 2214
rect 5971 2206 5973 2214
rect 2938 2204 2950 2206
rect 5946 2204 5958 2206
rect 1348 2176 1350 2184
rect 1732 2177 1747 2183
rect 1956 2176 1958 2184
rect 2356 2176 2358 2184
rect 2724 2176 2728 2184
rect 2836 2176 2840 2184
rect 4842 2176 4844 2184
rect 5112 2176 5116 2184
rect 5498 2176 5500 2184
rect 6772 2176 6774 2184
rect 356 2156 364 2164
rect 2189 2157 2204 2163
rect 2228 2156 2236 2164
rect 2461 2157 2483 2163
rect 6388 2156 6390 2164
rect 7261 2157 7276 2163
rect 301 2137 339 2143
rect 436 2137 467 2143
rect 109 2117 124 2123
rect 276 2117 291 2123
rect 509 2117 548 2123
rect 540 2112 548 2117
rect 717 2112 723 2143
rect 733 2112 739 2143
rect 845 2112 851 2143
rect 925 2137 947 2143
rect 1005 2137 1027 2143
rect 1197 2137 1219 2143
rect 1277 2137 1299 2143
rect 1597 2137 1612 2143
rect 1821 2137 1836 2143
rect 1677 2117 1692 2123
rect 1933 2123 1939 2143
rect 2317 2137 2339 2143
rect 1924 2117 1939 2123
rect 2317 2112 2323 2137
rect 2333 2117 2339 2137
rect 2381 2137 2396 2143
rect 2493 2137 2508 2143
rect 2548 2137 2563 2143
rect 4236 2137 4260 2143
rect 4660 2137 4668 2143
rect 6196 2137 6211 2143
rect 6253 2137 6275 2143
rect 6493 2137 6515 2143
rect 6580 2137 6595 2143
rect 6644 2137 6659 2143
rect 6852 2137 6867 2143
rect 6909 2137 6924 2143
rect 7220 2137 7235 2143
rect 7268 2137 7299 2143
rect 7309 2137 7363 2143
rect 2669 2117 2684 2123
rect 3597 2117 3620 2123
rect 3612 2114 3620 2117
rect 4644 2117 4691 2123
rect 4868 2117 4884 2123
rect 4876 2114 4884 2117
rect 6100 2117 6115 2123
rect 6452 2117 6467 2123
rect 6909 2117 6947 2123
rect 232 2096 236 2104
rect 1364 2097 1372 2103
rect 1652 2098 1656 2106
rect 2580 2096 2590 2104
rect 4468 2097 4515 2103
rect 5357 2097 5379 2103
rect 6292 2096 6300 2104
rect 6532 2096 6540 2104
rect 6909 2097 6915 2117
rect 7076 2117 7091 2123
rect 7181 2117 7219 2123
rect 564 2077 579 2083
rect 612 2077 636 2083
rect 692 2077 771 2083
rect 1165 2077 1180 2083
rect 2285 2077 2316 2083
rect 4538 2076 4540 2084
rect 5229 2077 5244 2083
rect 5229 2057 5235 2077
rect 1428 2037 1491 2043
rect 2196 2036 2198 2044
rect 2916 2037 2979 2043
rect 4634 2036 4636 2044
rect 5620 2036 5622 2044
rect 5914 2036 5916 2044
rect 6052 2036 6054 2044
rect 6148 2036 6150 2044
rect 1434 2014 1446 2016
rect 4442 2014 4454 2016
rect 1419 2006 1421 2014
rect 1429 2006 1431 2014
rect 1439 2006 1441 2014
rect 1449 2006 1451 2014
rect 1459 2006 1461 2014
rect 4427 2006 4429 2014
rect 4437 2006 4439 2014
rect 4447 2006 4449 2014
rect 4457 2006 4459 2014
rect 4467 2006 4469 2014
rect 1434 2004 1446 2006
rect 4442 2004 4454 2006
rect 148 1976 150 1984
rect 436 1976 438 1984
rect 1722 1976 1724 1984
rect 3028 1976 3032 1984
rect 3220 1976 3224 1984
rect 3364 1976 3366 1984
rect 360 1936 364 1944
rect 520 1936 524 1944
rect 1117 1943 1123 1963
rect 1556 1956 1558 1964
rect 1117 1937 1155 1943
rect 20 1897 35 1903
rect 109 1903 115 1923
rect 1149 1917 1155 1937
rect 1357 1937 1388 1943
rect 1652 1937 1683 1943
rect 1981 1937 1996 1943
rect 6804 1937 6819 1943
rect 1964 1932 1972 1936
rect 1421 1917 1484 1923
rect 1853 1917 1891 1923
rect 1949 1917 1971 1923
rect 6100 1916 6108 1924
rect 109 1897 131 1903
rect 125 1884 131 1897
rect 445 1897 460 1903
rect 52 1877 67 1883
rect 221 1877 236 1883
rect 244 1877 259 1883
rect 269 1877 307 1883
rect 452 1877 467 1883
rect 616 1876 620 1884
rect 925 1877 940 1883
rect 1021 1877 1036 1883
rect 1133 1877 1139 1908
rect 1220 1897 1235 1903
rect 1844 1897 1859 1903
rect 1876 1897 1939 1903
rect 1309 1877 1324 1883
rect 1517 1877 1539 1883
rect 1796 1877 1827 1883
rect 1284 1856 1292 1864
rect 1933 1857 1939 1897
rect 2156 1903 2164 1908
rect 2156 1897 2179 1903
rect 2173 1877 2179 1897
rect 2285 1884 2291 1903
rect 2484 1897 2499 1903
rect 3284 1897 3299 1903
rect 3309 1897 3324 1903
rect 4173 1897 4195 1903
rect 4413 1897 4476 1903
rect 6020 1897 6035 1903
rect 6125 1903 6131 1923
rect 6084 1897 6099 1903
rect 6125 1897 6163 1903
rect 6253 1897 6284 1903
rect 6749 1903 6755 1923
rect 6749 1897 6787 1903
rect 6916 1897 6931 1903
rect 7053 1897 7068 1903
rect 7101 1897 7139 1903
rect 2269 1877 2284 1883
rect 2340 1877 2371 1883
rect 2893 1877 2908 1883
rect 3277 1877 3292 1883
rect 3405 1877 3443 1883
rect 3693 1877 3715 1883
rect 3869 1877 3884 1883
rect 5069 1877 5092 1883
rect 5084 1872 5092 1877
rect 5708 1877 5732 1883
rect 5924 1877 6003 1883
rect 6493 1877 6531 1883
rect 2333 1857 2348 1863
rect 2845 1857 2867 1863
rect 2909 1857 2924 1863
rect 3156 1856 3164 1864
rect 3581 1857 3603 1863
rect 3821 1857 3843 1863
rect 4349 1857 4371 1863
rect 4797 1857 4819 1863
rect 6525 1857 6531 1877
rect 6685 1883 6691 1896
rect 6685 1877 6707 1883
rect 6749 1877 6764 1883
rect 6605 1857 6643 1863
rect 1684 1836 1686 1844
rect 2212 1836 2216 1844
rect 2938 1814 2950 1816
rect 5946 1814 5958 1816
rect 2923 1806 2925 1814
rect 2933 1806 2935 1814
rect 2943 1806 2945 1814
rect 2953 1806 2955 1814
rect 2963 1806 2965 1814
rect 5931 1806 5933 1814
rect 5941 1806 5943 1814
rect 5951 1806 5953 1814
rect 5961 1806 5963 1814
rect 5971 1806 5973 1814
rect 2938 1804 2950 1806
rect 5946 1804 5958 1806
rect 532 1776 536 1784
rect 3252 1776 3254 1784
rect 4778 1776 4780 1784
rect 5620 1776 5622 1784
rect 5668 1776 5670 1784
rect 5716 1776 5718 1784
rect 6234 1776 6236 1784
rect 317 1757 332 1763
rect 45 1737 83 1743
rect 253 1737 284 1743
rect 253 1724 259 1737
rect 365 1743 371 1763
rect 2516 1756 2524 1764
rect 2829 1757 2860 1763
rect 365 1737 403 1743
rect 1037 1737 1059 1743
rect 157 1717 172 1723
rect 733 1717 748 1723
rect 900 1717 915 1723
rect 1012 1717 1027 1723
rect 1053 1712 1059 1737
rect 1172 1737 1187 1743
rect 1357 1737 1379 1743
rect 1357 1712 1363 1737
rect 1373 1717 1379 1737
rect 1421 1737 1436 1743
rect 1437 1717 1484 1723
rect 1725 1712 1731 1743
rect 1789 1712 1795 1743
rect 1853 1712 1859 1743
rect 2116 1717 2147 1723
rect 2221 1712 2227 1743
rect 2429 1737 2444 1743
rect 2653 1737 2668 1743
rect 2740 1737 2755 1743
rect 2909 1743 2915 1763
rect 2909 1737 3004 1743
rect 3037 1737 3052 1743
rect 3268 1737 3283 1743
rect 3501 1743 3507 1763
rect 4157 1757 4179 1763
rect 5245 1757 5260 1763
rect 3501 1737 3539 1743
rect 5588 1737 5603 1743
rect 5901 1737 6003 1743
rect 2836 1717 2867 1723
rect 3117 1717 3155 1723
rect 3549 1717 3587 1723
rect 3604 1717 3619 1723
rect 3876 1717 3907 1723
rect 4269 1717 4291 1723
rect 4404 1717 4483 1723
rect 5165 1717 5203 1723
rect 5901 1717 5907 1737
rect 6541 1717 6579 1723
rect 3581 1697 3603 1703
rect 4941 1697 4963 1703
rect 6260 1697 6275 1703
rect 5548 1684 5556 1688
rect 2228 1677 2259 1683
rect 2301 1677 2316 1683
rect 2596 1676 2600 1684
rect 2788 1677 2803 1683
rect 3828 1676 3834 1684
rect 4077 1677 4092 1683
rect 5628 1683 5636 1688
rect 5628 1677 5644 1683
rect 5676 1683 5684 1688
rect 5724 1684 5732 1688
rect 5676 1677 5692 1683
rect 7126 1676 7132 1684
rect 3316 1636 3320 1644
rect 4260 1636 4262 1644
rect 7373 1637 7388 1643
rect 1434 1614 1446 1616
rect 4442 1614 4454 1616
rect 1419 1606 1421 1614
rect 1429 1606 1431 1614
rect 1439 1606 1441 1614
rect 1449 1606 1451 1614
rect 1459 1606 1461 1614
rect 4427 1606 4429 1614
rect 4437 1606 4439 1614
rect 4447 1606 4449 1614
rect 4457 1606 4459 1614
rect 4467 1606 4469 1614
rect 1434 1604 1446 1606
rect 4442 1604 4454 1606
rect 440 1576 444 1584
rect 1754 1576 1756 1584
rect 618 1556 620 1564
rect 2180 1537 2211 1543
rect 2381 1543 2387 1563
rect 2381 1537 2419 1543
rect 701 1517 707 1536
rect 2413 1517 2419 1537
rect 4612 1537 4627 1543
rect 5124 1537 5155 1543
rect 5668 1537 5683 1543
rect 20 1497 35 1503
rect 301 1497 316 1503
rect 589 1497 611 1503
rect 1117 1497 1132 1503
rect 1165 1497 1187 1503
rect 228 1477 259 1483
rect 365 1477 387 1483
rect 365 1464 371 1477
rect 952 1477 972 1483
rect 1101 1477 1116 1483
rect 1293 1477 1299 1508
rect 1501 1477 1523 1483
rect 1693 1477 1715 1483
rect 1773 1477 1795 1483
rect 2397 1477 2403 1508
rect 2548 1497 2563 1503
rect 2653 1497 2668 1503
rect 2733 1497 2755 1503
rect 2877 1503 2883 1523
rect 4573 1517 4595 1523
rect 5101 1517 5123 1523
rect 5357 1517 5372 1523
rect 5940 1517 6019 1523
rect 2877 1497 2892 1503
rect 3325 1497 3379 1503
rect 2525 1477 2556 1483
rect 2564 1477 2579 1483
rect 2829 1477 2844 1483
rect 52 1457 83 1463
rect 317 1457 355 1463
rect 1604 1456 1612 1464
rect 2216 1456 2220 1464
rect 2781 1457 2819 1463
rect 2829 1457 2835 1477
rect 3373 1477 3379 1497
rect 4372 1497 4387 1503
rect 5613 1497 5651 1503
rect 6429 1503 6435 1523
rect 6429 1497 6467 1503
rect 6557 1497 6572 1503
rect 6845 1497 6860 1503
rect 7261 1497 7276 1503
rect 3732 1477 3747 1483
rect 3812 1477 3827 1483
rect 5188 1477 5203 1483
rect 6317 1477 6332 1483
rect 6484 1477 6499 1483
rect 7220 1477 7235 1483
rect 2925 1457 2988 1463
rect 3661 1457 3683 1463
rect 3789 1457 3811 1463
rect 4413 1457 4499 1463
rect 4749 1457 4771 1463
rect 5933 1457 5996 1463
rect 2008 1436 2012 1444
rect 2868 1436 2870 1444
rect 6244 1436 6246 1444
rect 6516 1436 6518 1444
rect 2938 1414 2950 1416
rect 5946 1414 5958 1416
rect 2923 1406 2925 1414
rect 2933 1406 2935 1414
rect 2943 1406 2945 1414
rect 2953 1406 2955 1414
rect 2963 1406 2965 1414
rect 5931 1406 5933 1414
rect 5941 1406 5943 1414
rect 5951 1406 5953 1414
rect 5961 1406 5963 1414
rect 5971 1406 5973 1414
rect 2938 1404 2950 1406
rect 5946 1404 5958 1406
rect 74 1376 76 1384
rect 1162 1376 1164 1384
rect 2090 1376 2092 1384
rect 2164 1376 2168 1384
rect 2394 1376 2396 1384
rect 3412 1376 3416 1384
rect 3956 1376 3958 1384
rect 4468 1377 4531 1383
rect 4765 1377 4780 1383
rect 4970 1376 4972 1384
rect 5018 1376 5020 1384
rect 5066 1376 5068 1384
rect 5908 1376 5910 1384
rect 6196 1376 6198 1384
rect 1928 1356 1932 1364
rect 2308 1356 2316 1364
rect 701 1337 723 1343
rect 781 1323 787 1343
rect 845 1337 867 1343
rect 909 1337 924 1343
rect 765 1317 787 1323
rect 909 1317 947 1323
rect 909 1297 915 1317
rect 1053 1317 1068 1323
rect 1181 1323 1187 1343
rect 1960 1336 1964 1344
rect 2685 1343 2691 1363
rect 3092 1357 3107 1363
rect 5940 1357 6003 1363
rect 6813 1357 6835 1363
rect 2685 1337 2700 1343
rect 2932 1337 3011 1343
rect 4941 1337 4956 1343
rect 5092 1337 5107 1343
rect 5492 1337 5507 1343
rect 5581 1337 5596 1343
rect 1181 1317 1203 1323
rect 1325 1317 1363 1323
rect 1741 1317 1756 1323
rect 1853 1317 1868 1323
rect 2452 1317 2467 1323
rect 2804 1317 2835 1323
rect 3133 1317 3148 1323
rect 3908 1317 3955 1323
rect 4100 1317 4131 1323
rect 4292 1317 4323 1323
rect 5245 1317 5267 1323
rect 5540 1317 5555 1323
rect 5885 1323 5891 1343
rect 6125 1323 6131 1343
rect 6548 1337 6563 1343
rect 6676 1337 6707 1343
rect 6925 1337 6947 1343
rect 5853 1317 5891 1323
rect 6013 1317 6035 1323
rect 6045 1317 6083 1323
rect 6093 1317 6131 1323
rect 1988 1297 2003 1303
rect 2052 1297 2067 1303
rect 3965 1297 3987 1303
rect 4509 1297 4531 1303
rect 1965 1277 1996 1283
rect 2036 1277 2060 1283
rect 2429 1277 2444 1283
rect 2644 1277 2659 1283
rect 3224 1276 3228 1284
rect 4509 1283 4515 1297
rect 4685 1297 4707 1303
rect 4861 1297 4883 1303
rect 6077 1297 6083 1317
rect 6365 1317 6380 1323
rect 6461 1317 6499 1323
rect 6861 1317 6876 1323
rect 7172 1317 7187 1323
rect 5308 1284 5316 1288
rect 4429 1277 4515 1283
rect 4429 1257 4435 1277
rect 5356 1284 5364 1288
rect 5404 1283 5412 1288
rect 5396 1277 5412 1283
rect 5596 1284 5604 1288
rect 6204 1284 6212 1288
rect 6765 1277 6780 1283
rect 1524 1236 1526 1244
rect 1434 1214 1446 1216
rect 4442 1214 4454 1216
rect 1419 1206 1421 1214
rect 1429 1206 1431 1214
rect 1439 1206 1441 1214
rect 1449 1206 1451 1214
rect 1459 1206 1461 1214
rect 4427 1206 4429 1214
rect 4437 1206 4439 1214
rect 4447 1206 4449 1214
rect 4457 1206 4459 1214
rect 4467 1206 4469 1214
rect 1434 1204 1446 1206
rect 4442 1204 4454 1206
rect 266 1176 268 1184
rect 1754 1176 1756 1184
rect 6474 1176 6476 1184
rect 6858 1176 6860 1184
rect 1117 1137 1132 1143
rect 2621 1137 2636 1143
rect 4077 1137 4092 1143
rect 4205 1137 4236 1143
rect 4436 1137 4531 1143
rect 4676 1137 4691 1143
rect 7261 1137 7276 1143
rect 125 1117 147 1123
rect 468 1116 476 1124
rect 1325 1117 1340 1123
rect 93 1097 108 1103
rect 541 1103 547 1116
rect 541 1097 579 1103
rect 781 1097 819 1103
rect 829 1097 844 1103
rect 1229 1097 1251 1103
rect 1517 1103 1523 1123
rect 2232 1114 2236 1122
rect 3005 1117 3027 1123
rect 3981 1117 3996 1123
rect 4109 1117 4131 1123
rect 4237 1117 4259 1123
rect 4445 1117 4492 1123
rect 4605 1117 4627 1123
rect 1517 1097 1532 1103
rect 1629 1097 1667 1103
rect 1965 1097 1987 1103
rect 2141 1097 2156 1103
rect 2461 1097 2476 1103
rect 2509 1097 2524 1103
rect 2676 1097 2691 1103
rect 2893 1097 2956 1103
rect 3044 1097 3059 1103
rect 3213 1097 3228 1103
rect 3373 1097 3395 1103
rect 173 1077 195 1083
rect 381 1077 396 1083
rect 413 1077 435 1083
rect 685 1077 716 1083
rect 1149 1077 1187 1083
rect 1213 1077 1228 1083
rect 1245 1077 1283 1083
rect 1549 1077 1587 1083
rect 1508 1057 1532 1063
rect 1581 1057 1587 1077
rect 1933 1083 1939 1096
rect 3389 1084 3395 1097
rect 3741 1097 3756 1103
rect 5117 1097 5132 1103
rect 5229 1097 5251 1103
rect 5469 1103 5475 1123
rect 5469 1097 5507 1103
rect 5549 1097 5580 1103
rect 5661 1097 5699 1103
rect 6285 1097 6300 1103
rect 6333 1097 6371 1103
rect 6669 1097 6700 1103
rect 6861 1097 6915 1103
rect 6925 1097 6972 1103
rect 7149 1097 7164 1103
rect 7293 1097 7331 1103
rect 1908 1077 1923 1083
rect 1933 1077 1948 1083
rect 2100 1077 2131 1083
rect 2525 1077 2547 1083
rect 2557 1077 2588 1083
rect 2004 1056 2012 1064
rect 2189 1057 2204 1063
rect 2260 1057 2291 1063
rect 2557 1057 2563 1077
rect 2653 1077 2707 1083
rect 2756 1077 2787 1083
rect 3261 1077 3276 1083
rect 3181 1057 3196 1063
rect 3261 1057 3267 1077
rect 3293 1077 3324 1083
rect 3357 1077 3372 1083
rect 4941 1077 4963 1083
rect 5037 1077 5052 1083
rect 5405 1077 5420 1083
rect 5572 1077 5587 1083
rect 5757 1077 5772 1083
rect 6269 1077 6284 1083
rect 3804 1063 3812 1072
rect 7228 1064 7236 1072
rect 3804 1057 3836 1063
rect 5837 1057 5852 1063
rect 6797 1057 6812 1063
rect 6989 1057 7004 1063
rect 154 1036 156 1044
rect 1405 1037 1468 1043
rect 2708 1036 2710 1044
rect 2826 1036 2828 1044
rect 5738 1036 5740 1044
rect 5786 1036 5788 1044
rect 2938 1014 2950 1016
rect 5946 1014 5958 1016
rect 2923 1006 2925 1014
rect 2933 1006 2935 1014
rect 2943 1006 2945 1014
rect 2953 1006 2955 1014
rect 2963 1006 2965 1014
rect 5931 1006 5933 1014
rect 5941 1006 5943 1014
rect 5951 1006 5953 1014
rect 5961 1006 5963 1014
rect 5971 1006 5973 1014
rect 2938 1004 2950 1006
rect 5946 1004 5958 1006
rect 564 976 566 984
rect 2029 977 2051 983
rect 189 943 195 963
rect 692 957 707 963
rect 925 957 940 963
rect 189 937 227 943
rect 317 937 339 943
rect 77 917 92 923
rect 109 917 147 923
rect 244 917 259 923
rect 317 917 323 937
rect 868 937 899 943
rect 1252 937 1267 943
rect 1325 943 1331 963
rect 2029 963 2035 977
rect 2301 977 2316 983
rect 2932 977 2995 983
rect 3940 977 3955 983
rect 5076 976 5078 984
rect 2013 957 2035 963
rect 2749 957 2764 963
rect 2781 957 2796 963
rect 1300 937 1331 943
rect 1508 937 1523 943
rect 1613 937 1628 943
rect 1837 937 1891 943
rect 1981 937 2003 943
rect 2349 937 2387 943
rect 2509 937 2547 943
rect 525 917 547 923
rect 605 917 627 923
rect 941 917 963 923
rect 1069 917 1091 923
rect 1156 917 1171 923
rect 1229 917 1251 923
rect 1364 917 1379 923
rect 2452 917 2467 923
rect 2605 923 2611 943
rect 2669 937 2707 943
rect 2868 937 2883 943
rect 3101 943 3107 963
rect 3101 937 3139 943
rect 3156 937 3187 943
rect 3277 937 3299 943
rect 5044 937 5059 943
rect 5293 943 5299 963
rect 7028 956 7036 964
rect 7332 957 7347 963
rect 5261 937 5299 943
rect 5629 937 5644 943
rect 5700 937 5715 943
rect 5940 937 6035 943
rect 6061 937 6076 943
rect 6884 937 6899 943
rect 6996 937 7011 943
rect 2605 917 2620 923
rect 2724 917 2739 923
rect 3156 917 3171 923
rect 2420 896 2428 904
rect 2948 897 2995 903
rect 3165 897 3171 917
rect 3204 917 3219 923
rect 3485 917 3500 923
rect 3508 917 3571 923
rect 4013 917 4092 923
rect 4189 917 4227 923
rect 4381 917 4396 923
rect 4532 917 4579 923
rect 4621 917 4659 923
rect 5181 917 5219 923
rect 5565 917 5603 923
rect 5780 917 5795 923
rect 5828 917 5843 923
rect 6212 917 6227 923
rect 6333 917 6371 923
rect 7181 917 7196 923
rect 3380 897 3411 903
rect 3444 897 3459 903
rect 3592 898 3596 906
rect 4276 896 4284 904
rect 4740 897 4755 903
rect 4797 897 4819 903
rect 5341 897 5379 903
rect 6669 897 6691 903
rect 6749 897 6764 903
rect 6813 897 6828 903
rect 7092 896 7100 904
rect 749 877 764 883
rect 980 877 995 883
rect 1108 877 1123 883
rect 2301 877 2332 883
rect 3924 877 3955 883
rect 4717 877 4764 883
rect 1940 856 1942 864
rect 3818 856 3820 864
rect 4717 857 4723 877
rect 5084 883 5092 888
rect 5084 877 5100 883
rect 3482 836 3484 844
rect 3882 836 3884 844
rect 1434 814 1446 816
rect 4442 814 4454 816
rect 1419 806 1421 814
rect 1429 806 1431 814
rect 1439 806 1441 814
rect 1449 806 1451 814
rect 1459 806 1461 814
rect 4427 806 4429 814
rect 4437 806 4439 814
rect 4447 806 4449 814
rect 4457 806 4459 814
rect 4467 806 4469 814
rect 1434 804 1446 806
rect 4442 804 4454 806
rect 314 776 316 784
rect 820 776 822 784
rect 1764 776 1766 784
rect 1994 776 1996 784
rect 3402 776 3404 784
rect 4477 777 4492 783
rect 6906 776 6908 784
rect 660 737 675 743
rect 2426 736 2428 744
rect 2653 737 2684 743
rect 4109 737 4140 743
rect 7284 736 7286 744
rect 477 717 492 723
rect 573 717 595 723
rect 1092 717 1107 723
rect 1405 717 1452 723
rect 13 697 44 703
rect 13 684 19 697
rect 157 697 179 703
rect 221 697 243 703
rect 349 697 396 703
rect 605 697 620 703
rect 829 697 844 703
rect 1309 697 1331 703
rect 1389 697 1468 703
rect 1677 697 1708 703
rect 2020 697 2051 703
rect 2269 697 2284 703
rect 2333 703 2339 723
rect 4669 717 4691 723
rect 4765 717 4787 723
rect 4884 717 4899 723
rect 5469 717 5484 723
rect 5812 717 5827 723
rect 7144 714 7148 722
rect 7309 717 7331 723
rect 2324 697 2339 703
rect 2525 697 2563 703
rect 2781 697 2796 703
rect 3277 697 3299 703
rect 3581 697 3603 703
rect 3924 697 3939 703
rect 3981 697 4019 703
rect 4157 697 4172 703
rect 4852 697 4867 703
rect 4989 697 5027 703
rect 5357 697 5379 703
rect 6388 697 6403 703
rect 6868 697 6899 703
rect 6932 697 6947 703
rect 7053 697 7068 703
rect 493 677 515 683
rect 564 677 579 683
rect 861 677 883 683
rect 941 677 956 683
rect 973 677 995 683
rect 1053 677 1075 683
rect 1229 677 1267 683
rect 1325 677 1363 683
rect 1629 677 1651 683
rect 1725 677 1747 683
rect 1821 677 1843 683
rect 1901 677 1923 683
rect 2212 677 2227 683
rect 2365 677 2380 683
rect 2925 677 3043 683
rect 3060 677 3075 683
rect 3316 677 3331 683
rect 4052 677 4067 683
rect 4221 677 4275 683
rect 5485 677 5500 683
rect 6980 677 7011 683
rect 829 657 851 663
rect 72 636 76 644
rect 829 637 835 657
rect 1085 657 1107 663
rect 1197 657 1219 663
rect 1965 657 1987 663
rect 1981 637 1987 657
rect 2861 657 2899 663
rect 3604 657 3619 663
rect 4477 637 4508 643
rect 5636 636 5638 644
rect 5748 636 5750 644
rect 7034 636 7036 644
rect 2938 614 2950 616
rect 5946 614 5958 616
rect 2923 606 2925 614
rect 2933 606 2935 614
rect 2943 606 2945 614
rect 2953 606 2955 614
rect 2963 606 2965 614
rect 5931 606 5933 614
rect 5941 606 5943 614
rect 5951 606 5953 614
rect 5961 606 5963 614
rect 5971 606 5973 614
rect 2938 604 2950 606
rect 5946 604 5958 606
rect 660 576 662 584
rect 1005 563 1011 583
rect 1373 577 1420 583
rect 1556 576 1558 584
rect 2634 576 2636 584
rect 3044 576 3046 584
rect 3348 576 3350 584
rect 6013 577 6028 583
rect 6074 576 6076 584
rect 989 557 1011 563
rect 1597 557 1612 563
rect 1661 557 1683 563
rect 2381 557 2403 563
rect 3140 556 3148 564
rect 173 537 195 543
rect 285 537 323 543
rect 173 524 179 537
rect 621 537 659 543
rect 845 537 867 543
rect 957 537 979 543
rect 1181 537 1203 543
rect 1380 537 1459 543
rect 1524 537 1539 543
rect 1821 537 1843 543
rect 1917 537 1939 543
rect 1997 537 2035 543
rect 2205 537 2227 543
rect 2269 537 2291 543
rect 2452 537 2467 543
rect 2573 537 2604 543
rect 2637 537 2675 543
rect 2989 537 3004 543
rect 3165 537 3180 543
rect 3220 537 3235 543
rect 3453 537 3484 543
rect 3501 537 3539 543
rect 3533 524 3539 537
rect 3812 537 3827 543
rect 589 517 604 523
rect 701 517 723 523
rect 788 517 803 523
rect 1325 517 1340 523
rect 1572 517 1587 523
rect 1844 517 1859 523
rect 1869 517 1900 523
rect 2669 517 2707 523
rect 2877 517 2979 523
rect 3261 517 3276 523
rect 3389 517 3404 523
rect 1245 497 1283 503
rect 1476 496 1486 504
rect 1565 497 1587 503
rect 3821 497 3827 537
rect 4044 537 4068 543
rect 4420 537 4436 543
rect 4653 537 4668 543
rect 5085 543 5091 563
rect 4733 537 4787 543
rect 5085 537 5100 543
rect 5236 537 5251 543
rect 5549 537 5564 543
rect 5700 537 5715 543
rect 5885 537 5948 543
rect 6253 537 6268 543
rect 6989 537 7004 543
rect 7085 537 7100 543
rect 5037 517 5059 523
rect 5117 517 5155 523
rect 5149 497 5155 517
rect 5181 517 5219 523
rect 5341 517 5356 523
rect 5437 517 5468 523
rect 5485 517 5500 523
rect 6044 517 6060 523
rect 6044 512 6052 517
rect 6484 517 6499 523
rect 5789 497 5804 503
rect 5821 497 5843 503
rect 7148 492 7156 496
rect 3820 484 3828 488
rect 4566 476 4572 484
rect 5866 476 5868 484
rect 5940 477 5980 483
rect 6301 477 6355 483
rect 7124 477 7155 483
rect 52 436 56 444
rect 452 436 456 444
rect 3732 436 3734 444
rect 6132 436 6134 444
rect 1434 414 1446 416
rect 4442 414 4454 416
rect 1419 406 1421 414
rect 1429 406 1431 414
rect 1439 406 1441 414
rect 1449 406 1451 414
rect 1459 406 1461 414
rect 4427 406 4429 414
rect 4437 406 4439 414
rect 4447 406 4449 414
rect 4457 406 4459 414
rect 4467 406 4469 414
rect 1434 404 1446 406
rect 4442 404 4454 406
rect 132 376 134 384
rect 186 376 188 384
rect 3930 376 3932 384
rect 4250 376 4252 384
rect 4308 376 4310 384
rect 3668 356 3670 364
rect 1293 337 1315 343
rect 237 317 259 323
rect 356 316 364 324
rect 317 297 348 303
rect 637 303 643 323
rect 1309 317 1315 337
rect 1332 337 1347 343
rect 1869 337 1884 343
rect 3485 337 3500 343
rect 6684 337 6739 343
rect 6749 337 6780 343
rect 6684 332 6692 337
rect 6858 336 6860 344
rect 7044 337 7091 343
rect 637 297 675 303
rect 692 297 739 303
rect 893 297 908 303
rect 1012 297 1027 303
rect 1565 303 1571 323
rect 1588 316 1596 324
rect 1533 297 1571 303
rect 1597 297 1612 303
rect 1757 303 1763 323
rect 1780 316 1788 324
rect 1652 297 1667 303
rect 1725 297 1763 303
rect 1789 297 1804 303
rect 1892 297 1907 303
rect 1917 297 1948 303
rect 2132 297 2147 303
rect 2180 297 2195 303
rect 2452 297 2504 303
rect 3005 297 3027 303
rect 3188 297 3203 303
rect 3229 297 3251 303
rect 3309 297 3331 303
rect 3357 297 3395 303
rect 3789 303 3795 323
rect 4205 317 4227 323
rect 3652 297 3667 303
rect 3709 297 3747 303
rect 3757 297 3795 303
rect 3933 297 3948 303
rect 29 277 60 283
rect 285 277 307 283
rect 301 264 307 277
rect 413 277 444 283
rect 541 277 595 283
rect 685 277 691 296
rect 4253 297 4300 303
rect 4813 297 4851 303
rect 5213 303 5219 323
rect 6461 317 6476 323
rect 6605 317 6643 323
rect 5181 297 5219 303
rect 6861 297 6876 303
rect 6884 297 6947 303
rect 7101 297 7116 303
rect 7124 297 7139 303
rect 7149 297 7187 303
rect 829 277 851 283
rect 909 277 931 283
rect 1613 277 1635 283
rect 1805 277 1827 283
rect 1965 277 1987 283
rect 2237 277 2275 283
rect 2765 277 2803 283
rect 3069 277 3107 283
rect 3101 264 3107 277
rect 3293 277 3308 283
rect 3613 277 3651 283
rect 4372 277 4387 283
rect 4541 277 4556 283
rect 4573 277 4627 283
rect 4733 277 4764 283
rect 5149 277 5164 283
rect 5396 277 5411 283
rect 5444 277 5459 283
rect 5492 277 5507 283
rect 5597 277 5619 283
rect 6036 277 6067 283
rect 6285 277 6307 283
rect 6349 277 6380 283
rect 6285 264 6291 277
rect 6884 277 6915 283
rect 452 256 460 264
rect 1133 257 1155 263
rect 1645 257 1667 263
rect 266 236 268 244
rect 1236 236 1238 244
rect 1661 237 1667 257
rect 2909 257 2972 263
rect 3572 256 3580 264
rect 3892 257 3907 263
rect 6237 257 6275 263
rect 6909 257 6915 277
rect 2356 236 2360 244
rect 2376 236 2380 244
rect 2708 236 2712 244
rect 2794 236 2796 244
rect 4900 236 4902 244
rect 5524 236 5526 244
rect 5882 236 5884 244
rect 6676 236 6678 244
rect 2938 214 2950 216
rect 5946 214 5958 216
rect 2923 206 2925 214
rect 2933 206 2935 214
rect 2943 206 2945 214
rect 2953 206 2955 214
rect 2963 206 2965 214
rect 5931 206 5933 214
rect 5941 206 5943 214
rect 5951 206 5953 214
rect 5961 206 5963 214
rect 5971 206 5973 214
rect 2938 204 2950 206
rect 5946 204 5958 206
rect 100 176 104 184
rect 212 176 216 184
rect 392 176 396 184
rect 776 176 780 184
rect 888 176 892 184
rect 980 176 984 184
rect 1533 163 1539 183
rect 2212 176 2216 184
rect 3012 177 3027 183
rect 1437 157 1507 163
rect 1517 157 1539 163
rect 157 137 172 143
rect 541 137 556 143
rect 637 137 668 143
rect 1069 137 1091 143
rect 1149 137 1171 143
rect 1213 137 1235 143
rect 1293 137 1315 143
rect 1437 143 1443 157
rect 2349 157 2387 163
rect 3245 157 3260 163
rect 4221 157 4243 163
rect 1421 137 1443 143
rect 1597 137 1619 143
rect 1677 137 1699 143
rect 1789 137 1827 143
rect 1885 137 1907 143
rect 1949 137 1971 143
rect 2029 137 2067 143
rect 2157 137 2172 143
rect 2269 137 2284 143
rect 2413 137 2467 143
rect 2644 137 2675 143
rect 3181 143 3187 156
rect 3140 137 3155 143
rect 3165 137 3187 143
rect 3252 137 3283 143
rect 4781 137 4796 143
rect 5476 137 5491 143
rect 6756 137 6771 143
rect 6813 137 6828 143
rect 61 123 67 136
rect 7037 137 7059 143
rect 7101 137 7139 143
rect 45 117 67 123
rect 232 117 284 123
rect 589 117 620 123
rect 1405 117 1484 123
rect 1828 117 1843 123
rect 2276 117 2307 123
rect 2685 117 2707 123
rect 2724 117 2771 123
rect 3076 117 3091 123
rect 3172 117 3203 123
rect 3220 117 3235 123
rect 3293 117 3315 123
rect 3309 104 3315 117
rect 3757 117 3779 123
rect 3837 117 3852 123
rect 4173 117 4188 123
rect 4260 117 4275 123
rect 4621 117 4636 123
rect 4877 117 4915 123
rect 5012 117 5027 123
rect 5101 117 5139 123
rect 5149 117 5187 123
rect 5293 117 5331 123
rect 6861 117 6876 123
rect 7085 117 7100 123
rect 2484 97 2499 103
rect 3060 97 3075 103
rect 3364 97 3379 103
rect 3901 97 3939 103
rect 6436 77 6451 83
rect 1434 14 1446 16
rect 4442 14 4454 16
rect 1419 6 1421 14
rect 1429 6 1431 14
rect 1439 6 1441 14
rect 1449 6 1451 14
rect 1459 6 1461 14
rect 4427 6 4429 14
rect 4437 6 4439 14
rect 4447 6 4449 14
rect 4457 6 4459 14
rect 4467 6 4469 14
rect 1434 4 1446 6
rect 4442 4 4454 6
<< m2contact >>
rect 2915 5406 2923 5414
rect 2925 5406 2933 5414
rect 2935 5406 2943 5414
rect 2945 5406 2953 5414
rect 2955 5406 2963 5414
rect 2965 5406 2973 5414
rect 5923 5406 5931 5414
rect 5933 5406 5941 5414
rect 5943 5406 5951 5414
rect 5953 5406 5961 5414
rect 5963 5406 5971 5414
rect 5973 5406 5981 5414
rect 412 5376 420 5384
rect 556 5376 564 5384
rect 796 5376 804 5384
rect 924 5376 932 5384
rect 972 5376 980 5384
rect 1228 5376 1236 5384
rect 1548 5376 1556 5384
rect 2124 5376 2132 5384
rect 2428 5376 2436 5384
rect 2876 5376 2884 5384
rect 3676 5376 3684 5384
rect 3804 5376 3812 5384
rect 4604 5376 4612 5384
rect 5100 5376 5108 5384
rect 5404 5376 5412 5384
rect 6252 5376 6260 5384
rect 364 5356 372 5364
rect 524 5356 532 5364
rect 764 5356 772 5364
rect 844 5356 852 5364
rect 1116 5356 1124 5364
rect 1532 5356 1540 5364
rect 2140 5356 2148 5364
rect 2204 5356 2212 5364
rect 2444 5356 2452 5364
rect 2508 5356 2516 5364
rect 12 5336 20 5344
rect 60 5336 68 5344
rect 172 5336 180 5344
rect 204 5336 212 5344
rect 252 5336 260 5344
rect 268 5336 276 5344
rect 332 5336 340 5344
rect 476 5336 484 5344
rect 508 5336 516 5344
rect 636 5336 644 5344
rect 668 5336 676 5344
rect 700 5336 708 5344
rect 748 5336 756 5344
rect 796 5336 804 5344
rect 844 5336 852 5344
rect 876 5336 884 5344
rect 1020 5336 1028 5344
rect 1116 5336 1124 5344
rect 1148 5336 1156 5344
rect 1212 5336 1220 5344
rect 1436 5336 1444 5344
rect 1564 5336 1572 5344
rect 1596 5336 1604 5344
rect 1628 5336 1636 5344
rect 1804 5336 1812 5344
rect 1932 5336 1940 5344
rect 1964 5336 1972 5344
rect 2220 5336 2228 5344
rect 2268 5336 2276 5344
rect 2524 5336 2532 5344
rect 2748 5336 2756 5344
rect 2892 5336 2900 5344
rect 3228 5336 3236 5344
rect 3324 5336 3332 5344
rect 3516 5336 3524 5344
rect 3708 5336 3716 5344
rect 3756 5356 3764 5364
rect 5212 5356 5220 5364
rect 5452 5356 5460 5364
rect 3964 5336 3972 5344
rect 3996 5336 4004 5344
rect 4028 5336 4036 5344
rect 4092 5336 4100 5344
rect 4236 5336 4244 5344
rect 4284 5336 4292 5344
rect 4348 5336 4356 5344
rect 4444 5336 4452 5344
rect 4636 5336 4644 5344
rect 4812 5336 4820 5344
rect 4876 5336 4884 5344
rect 4908 5336 4916 5344
rect 4940 5336 4948 5344
rect 5132 5336 5140 5344
rect 5308 5336 5316 5344
rect 5868 5356 5876 5364
rect 6012 5356 6020 5364
rect 5484 5336 5492 5344
rect 5500 5336 5508 5344
rect 5852 5336 5860 5344
rect 5900 5336 5908 5344
rect 6060 5336 6068 5344
rect 6428 5336 6436 5344
rect 6620 5336 6628 5344
rect 6812 5336 6820 5344
rect 7228 5336 7236 5344
rect 7356 5336 7364 5344
rect 44 5316 52 5324
rect 92 5316 100 5324
rect 140 5316 148 5324
rect 284 5316 292 5324
rect 316 5316 324 5324
rect 332 5316 340 5324
rect 380 5316 388 5324
rect 492 5316 500 5324
rect 588 5316 596 5324
rect 620 5316 628 5324
rect 956 5316 964 5324
rect 1004 5316 1012 5324
rect 1068 5316 1076 5324
rect 1196 5316 1204 5324
rect 1260 5316 1268 5324
rect 1404 5318 1412 5326
rect 1580 5316 1588 5324
rect 1612 5316 1620 5324
rect 1660 5316 1668 5324
rect 2012 5316 2020 5324
rect 2172 5316 2180 5324
rect 2236 5316 2244 5324
rect 2316 5316 2324 5324
rect 2476 5316 2484 5324
rect 2540 5316 2548 5324
rect 2556 5316 2564 5324
rect 2572 5316 2580 5324
rect 2668 5316 2676 5324
rect 2716 5316 2724 5324
rect 2748 5316 2756 5324
rect 156 5296 164 5304
rect 172 5296 180 5304
rect 220 5296 228 5304
rect 236 5296 244 5304
rect 604 5296 612 5304
rect 668 5296 676 5304
rect 716 5296 724 5304
rect 876 5296 884 5304
rect 908 5296 916 5304
rect 1644 5296 1652 5304
rect 2780 5296 2788 5304
rect 2908 5316 2916 5324
rect 2988 5316 2996 5324
rect 3036 5316 3044 5324
rect 3196 5316 3204 5324
rect 3372 5316 3380 5324
rect 3564 5316 3572 5324
rect 3692 5316 3700 5324
rect 3724 5316 3732 5324
rect 3788 5316 3796 5324
rect 3932 5318 3940 5326
rect 2828 5296 2836 5304
rect 4028 5296 4036 5304
rect 4076 5316 4084 5324
rect 4108 5316 4116 5324
rect 4316 5316 4324 5324
rect 4396 5316 4404 5324
rect 4476 5318 4484 5326
rect 4684 5316 4692 5324
rect 4828 5316 4836 5324
rect 4972 5318 4980 5326
rect 4252 5296 4260 5304
rect 5116 5316 5124 5324
rect 5164 5316 5172 5324
rect 5180 5316 5188 5324
rect 5292 5316 5300 5324
rect 5420 5316 5428 5324
rect 5516 5316 5524 5324
rect 5580 5318 5588 5326
rect 5644 5316 5652 5324
rect 5724 5316 5732 5324
rect 5916 5316 5924 5324
rect 6140 5316 6148 5324
rect 6188 5316 6196 5324
rect 6396 5318 6404 5326
rect 6588 5318 6596 5326
rect 6780 5318 6788 5326
rect 6908 5316 6916 5324
rect 6972 5318 6980 5326
rect 7100 5316 7108 5324
rect 7164 5318 7172 5326
rect 4876 5296 4884 5304
rect 5932 5296 5940 5304
rect 6028 5296 6036 5304
rect 124 5276 132 5284
rect 636 5276 644 5284
rect 732 5276 740 5284
rect 1196 5276 1204 5284
rect 2092 5276 2100 5284
rect 2396 5276 2404 5284
rect 5068 5276 5076 5284
rect 140 5236 148 5244
rect 316 5236 324 5244
rect 892 5236 900 5244
rect 1132 5236 1140 5244
rect 1276 5236 1284 5244
rect 2588 5236 2596 5244
rect 2700 5236 2708 5244
rect 3292 5236 3300 5244
rect 3484 5236 3492 5244
rect 4796 5236 4804 5244
rect 5708 5236 5716 5244
rect 5868 5236 5876 5244
rect 6044 5236 6052 5244
rect 6268 5236 6276 5244
rect 6460 5236 6468 5244
rect 6652 5236 6660 5244
rect 6844 5236 6852 5244
rect 7036 5236 7044 5244
rect 1411 5206 1419 5214
rect 1421 5206 1429 5214
rect 1431 5206 1439 5214
rect 1441 5206 1449 5214
rect 1451 5206 1459 5214
rect 1461 5206 1469 5214
rect 4419 5206 4427 5214
rect 4429 5206 4437 5214
rect 4439 5206 4447 5214
rect 4449 5206 4457 5214
rect 4459 5206 4467 5214
rect 4469 5206 4477 5214
rect 588 5176 596 5184
rect 1404 5176 1412 5184
rect 3404 5176 3412 5184
rect 4092 5176 4100 5184
rect 4300 5176 4308 5184
rect 4892 5176 4900 5184
rect 2620 5156 2628 5164
rect 6492 5156 6500 5164
rect 124 5136 132 5144
rect 1164 5136 1172 5144
rect 1420 5136 1428 5144
rect 1580 5136 1588 5144
rect 3004 5136 3012 5144
rect 4140 5136 4148 5144
rect 4204 5136 4212 5144
rect 4636 5136 4644 5144
rect 4908 5136 4916 5144
rect 5484 5136 5492 5144
rect 5548 5136 5556 5144
rect 5804 5136 5812 5144
rect 6076 5136 6084 5144
rect 92 5116 100 5124
rect 156 5116 164 5124
rect 220 5116 228 5124
rect 316 5116 324 5124
rect 108 5096 116 5104
rect 204 5096 212 5104
rect 284 5096 292 5104
rect 332 5096 340 5104
rect 364 5096 372 5104
rect 492 5116 500 5124
rect 460 5096 468 5104
rect 508 5096 516 5104
rect 540 5096 548 5104
rect 636 5096 644 5104
rect 684 5116 692 5124
rect 812 5116 820 5124
rect 972 5116 980 5124
rect 1036 5116 1044 5124
rect 1068 5116 1076 5124
rect 1132 5116 1140 5124
rect 1276 5116 1284 5124
rect 1388 5116 1396 5124
rect 2348 5116 2356 5124
rect 3100 5116 3108 5124
rect 716 5096 724 5104
rect 780 5096 788 5104
rect 812 5096 820 5104
rect 844 5096 852 5104
rect 876 5096 884 5104
rect 1036 5096 1044 5104
rect 1116 5096 1124 5104
rect 1148 5096 1156 5104
rect 1196 5096 1204 5104
rect 1228 5096 1236 5104
rect 1340 5096 1348 5104
rect 1404 5096 1412 5104
rect 1692 5096 1700 5104
rect 1708 5096 1716 5104
rect 1772 5096 1780 5104
rect 1788 5096 1796 5104
rect 1820 5096 1828 5104
rect 1964 5096 1972 5104
rect 1996 5096 2004 5104
rect 2060 5096 2068 5104
rect 2076 5096 2084 5104
rect 2188 5096 2196 5104
rect 2236 5094 2244 5102
rect 2316 5096 2324 5104
rect 2412 5096 2420 5104
rect 2492 5096 2500 5104
rect 2556 5094 2564 5102
rect 2684 5096 2692 5104
rect 2732 5096 2740 5104
rect 2876 5096 2884 5104
rect 3820 5116 3828 5124
rect 3932 5116 3940 5124
rect 3148 5096 3156 5104
rect 3180 5096 3188 5104
rect 3196 5096 3204 5104
rect 3244 5096 3252 5104
rect 3340 5096 3348 5104
rect 3356 5096 3364 5104
rect 3388 5096 3396 5104
rect 3436 5096 3444 5104
rect 3452 5096 3460 5104
rect 3484 5096 3492 5104
rect 3596 5096 3604 5104
rect 3660 5096 3668 5104
rect 3692 5096 3700 5104
rect 3724 5096 3732 5104
rect 3740 5096 3748 5104
rect 3788 5096 3796 5104
rect 3804 5096 3812 5104
rect 3900 5096 3908 5104
rect 3964 5096 3972 5104
rect 3996 5096 4004 5104
rect 4028 5096 4036 5104
rect 4092 5096 4100 5104
rect 4236 5116 4244 5124
rect 4268 5116 4276 5124
rect 4172 5096 4180 5104
rect 4236 5096 4244 5104
rect 4300 5096 4308 5104
rect 4332 5096 4340 5104
rect 4348 5096 4356 5104
rect 4508 5096 4516 5104
rect 4556 5096 4564 5104
rect 4572 5096 4580 5104
rect 4604 5096 4612 5104
rect 5452 5116 5460 5124
rect 5836 5116 5844 5124
rect 5868 5116 5876 5124
rect 5900 5116 5908 5124
rect 6028 5116 6036 5124
rect 6204 5116 6212 5124
rect 4668 5096 4676 5104
rect 4684 5096 4692 5104
rect 4764 5094 4772 5102
rect 5036 5094 5044 5102
rect 5132 5096 5140 5104
rect 5148 5096 5156 5104
rect 5196 5096 5204 5104
rect 5292 5096 5300 5104
rect 5420 5096 5428 5104
rect 5484 5096 5492 5104
rect 5516 5096 5524 5104
rect 5548 5096 5556 5104
rect 5660 5096 5668 5104
rect 5724 5094 5732 5102
rect 5804 5096 5812 5104
rect 5868 5096 5876 5104
rect 5996 5096 6004 5104
rect 6012 5096 6020 5104
rect 6076 5096 6084 5104
rect 6092 5096 6100 5104
rect 6140 5096 6148 5104
rect 6172 5096 6180 5104
rect 6236 5096 6244 5104
rect 6252 5096 6260 5104
rect 6284 5096 6292 5104
rect 6332 5096 6340 5104
rect 6348 5096 6356 5104
rect 6380 5096 6388 5104
rect 6428 5096 6436 5104
rect 6524 5096 6532 5104
rect 6540 5096 6548 5104
rect 6556 5096 6564 5104
rect 6620 5096 6628 5104
rect 6652 5096 6660 5104
rect 6716 5094 6724 5102
rect 6860 5096 6868 5104
rect 6908 5096 6916 5104
rect 7068 5096 7076 5104
rect 7228 5096 7236 5104
rect 7260 5096 7268 5104
rect 44 5076 52 5084
rect 172 5076 180 5084
rect 220 5076 228 5084
rect 252 5076 260 5084
rect 268 5076 276 5084
rect 300 5076 308 5084
rect 380 5076 388 5084
rect 444 5076 452 5084
rect 476 5076 484 5084
rect 620 5076 628 5084
rect 668 5076 676 5084
rect 732 5076 740 5084
rect 796 5076 804 5084
rect 860 5076 868 5084
rect 892 5076 900 5084
rect 940 5076 948 5084
rect 1020 5076 1028 5084
rect 1148 5076 1156 5084
rect 1212 5076 1220 5084
rect 1244 5076 1252 5084
rect 1308 5076 1316 5084
rect 1324 5076 1332 5084
rect 1356 5076 1364 5084
rect 1548 5076 1556 5084
rect 1660 5076 1668 5084
rect 1708 5076 1716 5084
rect 1724 5076 1732 5084
rect 1756 5076 1764 5084
rect 1836 5076 1844 5084
rect 28 5056 36 5064
rect 140 5056 148 5064
rect 348 5056 356 5064
rect 364 5056 372 5064
rect 508 5056 516 5064
rect 604 5056 612 5064
rect 748 5056 756 5064
rect 924 5056 932 5064
rect 988 5056 996 5064
rect 1084 5056 1092 5064
rect 1516 5056 1524 5064
rect 1596 5056 1604 5064
rect 1804 5056 1812 5064
rect 1948 5076 1956 5084
rect 2012 5076 2020 5084
rect 2300 5076 2308 5084
rect 2364 5076 2372 5084
rect 2396 5076 2404 5084
rect 2540 5076 2548 5084
rect 3004 5076 3012 5084
rect 3116 5076 3124 5084
rect 3164 5076 3172 5084
rect 3276 5076 3284 5084
rect 3468 5076 3476 5084
rect 3500 5076 3508 5084
rect 3532 5076 3540 5084
rect 3644 5076 3652 5084
rect 3708 5076 3716 5084
rect 3868 5076 3876 5084
rect 3884 5076 3892 5084
rect 3980 5076 3988 5084
rect 4012 5076 4020 5084
rect 4028 5076 4036 5084
rect 4076 5076 4084 5084
rect 4188 5076 4196 5084
rect 4252 5076 4260 5084
rect 4316 5076 4324 5084
rect 4412 5076 4420 5084
rect 4588 5076 4596 5084
rect 4700 5076 4708 5084
rect 4780 5076 4788 5084
rect 5068 5076 5076 5084
rect 5180 5076 5188 5084
rect 5228 5076 5236 5084
rect 5308 5076 5316 5084
rect 5548 5076 5556 5084
rect 5788 5076 5796 5084
rect 5852 5076 5860 5084
rect 5980 5076 5988 5084
rect 6076 5076 6084 5084
rect 6156 5076 6164 5084
rect 1884 5056 1892 5064
rect 1996 5056 2004 5064
rect 2028 5056 2036 5064
rect 2060 5056 2068 5064
rect 2092 5056 2100 5064
rect 3324 5056 3332 5064
rect 3548 5056 3556 5064
rect 3612 5056 3620 5064
rect 3628 5056 3636 5064
rect 4060 5056 4068 5064
rect 5100 5056 5108 5064
rect 6044 5056 6052 5064
rect 6588 5056 6596 5064
rect 6636 5076 6644 5084
rect 6684 5076 6692 5084
rect 6924 5076 6932 5084
rect 7084 5076 7092 5084
rect 7100 5076 7108 5084
rect 6892 5056 6900 5064
rect 6956 5056 6964 5064
rect 236 5036 244 5044
rect 572 5036 580 5044
rect 764 5036 772 5044
rect 908 5036 916 5044
rect 972 5036 980 5044
rect 1100 5036 1108 5044
rect 1644 5036 1652 5044
rect 1740 5036 1748 5044
rect 1852 5036 1860 5044
rect 2108 5036 2116 5044
rect 2428 5036 2436 5044
rect 2620 5036 2628 5044
rect 3660 5036 3668 5044
rect 3756 5036 3764 5044
rect 4364 5036 4372 5044
rect 5388 5036 5396 5044
rect 5596 5036 5604 5044
rect 6140 5036 6148 5044
rect 6300 5036 6308 5044
rect 6396 5036 6404 5044
rect 6844 5036 6852 5044
rect 6876 5036 6884 5044
rect 6940 5036 6948 5044
rect 6972 5036 6980 5044
rect 7164 5036 7172 5044
rect 2915 5006 2923 5014
rect 2925 5006 2933 5014
rect 2935 5006 2943 5014
rect 2945 5006 2953 5014
rect 2955 5006 2963 5014
rect 2965 5006 2973 5014
rect 5923 5006 5931 5014
rect 5933 5006 5941 5014
rect 5943 5006 5951 5014
rect 5953 5006 5961 5014
rect 5963 5006 5971 5014
rect 5973 5006 5981 5014
rect 92 4976 100 4984
rect 156 4976 164 4984
rect 220 4976 228 4984
rect 284 4976 292 4984
rect 476 4976 484 4984
rect 508 4976 516 4984
rect 684 4976 692 4984
rect 812 4976 820 4984
rect 876 4976 884 4984
rect 924 4976 932 4984
rect 1084 4976 1092 4984
rect 1148 4976 1156 4984
rect 1404 4976 1412 4984
rect 1548 4976 1556 4984
rect 1676 4976 1684 4984
rect 1820 4976 1828 4984
rect 2220 4976 2228 4984
rect 2556 4976 2564 4984
rect 3020 4976 3028 4984
rect 3148 4976 3156 4984
rect 3372 4976 3380 4984
rect 4236 4976 4244 4984
rect 5180 4976 5188 4984
rect 5516 4976 5524 4984
rect 6220 4976 6228 4984
rect 6668 4976 6676 4984
rect 6940 4976 6948 4984
rect 7244 4976 7252 4984
rect 124 4956 132 4964
rect 236 4956 244 4964
rect 332 4956 340 4964
rect 348 4956 356 4964
rect 604 4956 612 4964
rect 700 4956 708 4964
rect 828 4956 836 4964
rect 940 4956 948 4964
rect 988 4956 996 4964
rect 1276 4956 1284 4964
rect 1356 4956 1364 4964
rect 1372 4956 1380 4964
rect 1564 4956 1572 4964
rect 1964 4956 1972 4964
rect 1980 4956 1988 4964
rect 2172 4956 2180 4964
rect 2300 4956 2308 4964
rect 2316 4956 2324 4964
rect 2428 4956 2436 4964
rect 2492 4956 2500 4964
rect 2812 4956 2820 4964
rect 3132 4956 3140 4964
rect 3740 4956 3748 4964
rect 3932 4956 3940 4964
rect 4108 4956 4116 4964
rect 4700 4956 4708 4964
rect 4732 4956 4740 4964
rect 4924 4956 4932 4964
rect 5116 4956 5124 4964
rect 5308 4956 5316 4964
rect 5372 4956 5380 4964
rect 5580 4956 5588 4964
rect 5740 4956 5748 4964
rect 5772 4956 5780 4964
rect 6028 4956 6036 4964
rect 6380 4956 6388 4964
rect 6524 4956 6532 4964
rect 6764 4956 6772 4964
rect 6956 4956 6964 4964
rect 7164 4956 7172 4964
rect 7276 4956 7284 4964
rect 7324 4956 7332 4964
rect 7340 4956 7348 4964
rect 7356 4956 7364 4964
rect 44 4916 52 4924
rect 140 4936 148 4944
rect 204 4936 212 4944
rect 316 4936 324 4944
rect 380 4936 388 4944
rect 412 4936 420 4944
rect 444 4936 452 4944
rect 492 4936 500 4944
rect 636 4936 644 4944
rect 732 4936 740 4944
rect 796 4936 804 4944
rect 860 4936 868 4944
rect 892 4936 900 4944
rect 988 4936 996 4944
rect 1052 4936 1060 4944
rect 1100 4936 1108 4944
rect 1212 4936 1220 4944
rect 1532 4936 1540 4944
rect 1580 4936 1588 4944
rect 1644 4936 1652 4944
rect 1692 4936 1700 4944
rect 1708 4936 1716 4944
rect 1772 4936 1780 4944
rect 1804 4936 1812 4944
rect 1948 4936 1956 4944
rect 2108 4936 2116 4944
rect 2220 4936 2228 4944
rect 2252 4936 2260 4944
rect 2332 4936 2340 4944
rect 2348 4936 2356 4944
rect 2412 4936 2420 4944
rect 2508 4936 2516 4944
rect 2844 4936 2852 4944
rect 2876 4936 2884 4944
rect 3036 4936 3044 4944
rect 3084 4936 3092 4944
rect 3116 4936 3124 4944
rect 3164 4936 3172 4944
rect 3212 4936 3220 4944
rect 3436 4936 3444 4944
rect 3484 4936 3492 4944
rect 3500 4936 3508 4944
rect 3628 4936 3636 4944
rect 3740 4936 3748 4944
rect 3852 4936 3860 4944
rect 3932 4936 3940 4944
rect 3964 4936 3972 4944
rect 4028 4936 4036 4944
rect 4044 4936 4052 4944
rect 4156 4936 4164 4944
rect 4220 4936 4228 4944
rect 4492 4936 4500 4944
rect 4556 4936 4564 4944
rect 4748 4936 4756 4944
rect 4812 4936 4820 4944
rect 4892 4936 4900 4944
rect 5036 4936 5044 4944
rect 5100 4936 5108 4944
rect 5164 4936 5172 4944
rect 5452 4936 5460 4944
rect 5500 4936 5508 4944
rect 5724 4936 5732 4944
rect 5836 4936 5844 4944
rect 6044 4936 6052 4944
rect 6108 4936 6116 4944
rect 6268 4936 6276 4944
rect 6332 4936 6340 4944
rect 6444 4936 6452 4944
rect 6508 4936 6516 4944
rect 6572 4936 6580 4944
rect 6588 4936 6596 4944
rect 6620 4936 6628 4944
rect 6652 4936 6660 4944
rect 6716 4936 6724 4944
rect 6908 4936 6916 4944
rect 7084 4936 7092 4944
rect 124 4916 132 4924
rect 156 4916 164 4924
rect 268 4916 276 4924
rect 428 4916 436 4924
rect 540 4916 548 4924
rect 588 4916 596 4924
rect 652 4916 660 4924
rect 716 4916 724 4924
rect 748 4916 756 4924
rect 780 4916 788 4924
rect 956 4916 964 4924
rect 988 4916 996 4924
rect 1036 4916 1044 4924
rect 1116 4916 1124 4924
rect 1196 4916 1204 4924
rect 1228 4916 1236 4924
rect 1308 4916 1316 4924
rect 1516 4916 1524 4924
rect 1596 4916 1604 4924
rect 1628 4916 1636 4924
rect 1724 4916 1732 4924
rect 1756 4916 1764 4924
rect 1900 4916 1908 4924
rect 1916 4916 1924 4924
rect 1932 4916 1940 4924
rect 2012 4916 2020 4924
rect 2076 4916 2084 4924
rect 2092 4916 2100 4924
rect 2124 4916 2132 4924
rect 2364 4916 2372 4924
rect 2460 4916 2468 4924
rect 2524 4916 2532 4924
rect 2604 4916 2612 4924
rect 2684 4916 2692 4924
rect 2748 4918 2756 4926
rect 2812 4916 2820 4924
rect 2860 4916 2868 4924
rect 2876 4916 2884 4924
rect 3068 4916 3076 4924
rect 3100 4916 3108 4924
rect 3180 4916 3188 4924
rect 3260 4916 3268 4924
rect 3388 4916 3396 4924
rect 3420 4916 3428 4924
rect 460 4896 468 4904
rect 684 4896 692 4904
rect 780 4896 788 4904
rect 1084 4896 1092 4904
rect 1164 4896 1172 4904
rect 1468 4896 1476 4904
rect 1660 4896 1668 4904
rect 1788 4896 1796 4904
rect 1900 4896 1908 4904
rect 1996 4896 2004 4904
rect 2060 4896 2068 4904
rect 2556 4896 2564 4904
rect 2924 4896 2932 4904
rect 3068 4896 3076 4904
rect 3388 4896 3396 4904
rect 3468 4916 3476 4924
rect 3516 4916 3524 4924
rect 3548 4916 3556 4924
rect 3612 4916 3620 4924
rect 3660 4916 3668 4924
rect 3676 4916 3684 4924
rect 3708 4916 3716 4924
rect 3772 4916 3780 4924
rect 3820 4916 3828 4924
rect 3836 4916 3844 4924
rect 3868 4916 3876 4924
rect 3964 4916 3972 4924
rect 4060 4916 4068 4924
rect 4140 4916 4148 4924
rect 4172 4916 4180 4924
rect 4220 4916 4228 4924
rect 4316 4916 4324 4924
rect 4364 4918 4372 4926
rect 4492 4916 4500 4924
rect 4620 4916 4628 4924
rect 4668 4916 4676 4924
rect 4684 4916 4692 4924
rect 4732 4916 4740 4924
rect 4764 4916 4772 4924
rect 4796 4916 4804 4924
rect 4828 4916 4836 4924
rect 4860 4916 4868 4924
rect 4876 4916 4884 4924
rect 4956 4916 4964 4924
rect 5004 4916 5012 4924
rect 5020 4916 5028 4924
rect 5052 4916 5060 4924
rect 5084 4916 5092 4924
rect 5164 4916 5172 4924
rect 5308 4918 5316 4926
rect 5404 4916 5412 4924
rect 5468 4916 5476 4924
rect 5484 4916 5492 4924
rect 5548 4916 5556 4924
rect 5612 4916 5620 4924
rect 5676 4916 5684 4924
rect 5708 4916 5716 4924
rect 5740 4916 5748 4924
rect 5852 4916 5860 4924
rect 5900 4916 5908 4924
rect 5916 4916 5924 4924
rect 5932 4916 5940 4924
rect 5996 4916 6004 4924
rect 6076 4916 6084 4924
rect 6092 4916 6100 4924
rect 6124 4916 6132 4924
rect 6140 4916 6148 4924
rect 6220 4916 6228 4924
rect 6252 4916 6260 4924
rect 6268 4916 6276 4924
rect 6316 4916 6324 4924
rect 6348 4916 6356 4924
rect 6396 4916 6404 4924
rect 6428 4916 6436 4924
rect 6444 4916 6452 4924
rect 6492 4916 6500 4924
rect 6588 4916 6596 4924
rect 6604 4916 6612 4924
rect 6636 4916 6644 4924
rect 6700 4916 6708 4924
rect 6732 4916 6740 4924
rect 6748 4916 6756 4924
rect 6812 4916 6820 4924
rect 6828 4916 6836 4924
rect 6844 4916 6852 4924
rect 6892 4916 6900 4924
rect 6924 4916 6932 4924
rect 7052 4916 7060 4924
rect 7196 4916 7204 4924
rect 7212 4916 7220 4924
rect 7276 4916 7284 4924
rect 7324 4916 7332 4924
rect 3580 4896 3588 4904
rect 3692 4896 3700 4904
rect 3868 4896 3876 4904
rect 3980 4896 3988 4904
rect 4092 4896 4100 4904
rect 4508 4896 4516 4904
rect 4588 4896 4596 4904
rect 4828 4896 4836 4904
rect 4908 4896 4916 4904
rect 5068 4896 5076 4904
rect 5116 4896 5124 4904
rect 5644 4896 5652 4904
rect 5820 4896 5828 4904
rect 6220 4896 6228 4904
rect 6284 4896 6292 4904
rect 6524 4896 6532 4904
rect 6668 4896 6676 4904
rect 12 4876 20 4884
rect 1836 4876 1844 4884
rect 2028 4876 2036 4884
rect 2572 4876 2580 4884
rect 4140 4876 4148 4884
rect 5420 4876 5428 4884
rect 5676 4876 5684 4884
rect 6460 4876 6468 4884
rect 6972 4876 6980 4884
rect 1724 4856 1732 4864
rect 3708 4856 3716 4864
rect 6428 4856 6436 4864
rect 556 4836 564 4844
rect 620 4836 628 4844
rect 1004 4836 1012 4844
rect 1196 4836 1204 4844
rect 1244 4836 1252 4844
rect 1356 4836 1364 4844
rect 1596 4836 1604 4844
rect 2012 4836 2020 4844
rect 2364 4836 2372 4844
rect 2620 4836 2628 4844
rect 3548 4836 3556 4844
rect 4060 4836 4068 4844
rect 4172 4836 4180 4844
rect 4636 4836 4644 4844
rect 4764 4836 4772 4844
rect 4972 4836 4980 4844
rect 5868 4836 5876 4844
rect 6156 4836 6164 4844
rect 7196 4836 7204 4844
rect 7276 4836 7284 4844
rect 1411 4806 1419 4814
rect 1421 4806 1429 4814
rect 1431 4806 1439 4814
rect 1441 4806 1449 4814
rect 1451 4806 1459 4814
rect 1461 4806 1469 4814
rect 4419 4806 4427 4814
rect 4429 4806 4437 4814
rect 4439 4806 4447 4814
rect 4449 4806 4457 4814
rect 4459 4806 4467 4814
rect 4469 4806 4477 4814
rect 460 4776 468 4784
rect 892 4776 900 4784
rect 1036 4776 1044 4784
rect 1948 4776 1956 4784
rect 2012 4776 2020 4784
rect 2332 4776 2340 4784
rect 2924 4776 2932 4784
rect 3036 4776 3044 4784
rect 3708 4776 3716 4784
rect 4108 4776 4116 4784
rect 4556 4776 4564 4784
rect 4748 4776 4756 4784
rect 4796 4776 4804 4784
rect 5228 4776 5236 4784
rect 5980 4776 5988 4784
rect 6236 4776 6244 4784
rect 6380 4776 6388 4784
rect 5132 4756 5140 4764
rect 6908 4756 6916 4764
rect 7180 4756 7188 4764
rect 204 4736 212 4744
rect 1756 4736 1764 4744
rect 2092 4736 2100 4744
rect 2380 4736 2388 4744
rect 2636 4736 2644 4744
rect 3436 4736 3444 4744
rect 4092 4736 4100 4744
rect 5068 4736 5076 4744
rect 6300 4736 6308 4744
rect 6652 4736 6660 4744
rect 636 4716 644 4724
rect 1532 4716 1540 4724
rect 1804 4716 1812 4724
rect 1820 4716 1828 4724
rect 1852 4716 1860 4724
rect 2140 4716 2148 4724
rect 2284 4716 2292 4724
rect 2732 4716 2740 4724
rect 2844 4716 2852 4724
rect 3612 4716 3620 4724
rect 252 4696 260 4704
rect 300 4696 308 4704
rect 412 4696 420 4704
rect 524 4696 532 4704
rect 572 4696 580 4704
rect 588 4696 596 4704
rect 780 4696 788 4704
rect 892 4696 900 4704
rect 988 4696 996 4704
rect 1068 4696 1076 4704
rect 1116 4696 1124 4704
rect 12 4676 20 4684
rect 204 4676 212 4684
rect 268 4676 276 4684
rect 348 4680 356 4688
rect 1580 4696 1588 4704
rect 1644 4696 1652 4704
rect 1676 4696 1684 4704
rect 1708 4696 1716 4704
rect 1932 4696 1940 4704
rect 1980 4696 1988 4704
rect 2188 4696 2196 4704
rect 2236 4696 2244 4704
rect 2364 4696 2372 4704
rect 2508 4694 2516 4702
rect 2572 4696 2580 4704
rect 2620 4696 2628 4704
rect 2668 4696 2676 4704
rect 2700 4696 2708 4704
rect 2780 4696 2788 4704
rect 2812 4696 2820 4704
rect 2908 4696 2916 4704
rect 3020 4696 3028 4704
rect 3164 4694 3172 4702
rect 3228 4696 3236 4704
rect 3276 4696 3284 4704
rect 3356 4696 3364 4704
rect 3484 4696 3492 4704
rect 3548 4696 3556 4704
rect 3564 4696 3572 4704
rect 3820 4716 3828 4724
rect 3660 4696 3668 4704
rect 3708 4696 3716 4704
rect 3804 4696 3812 4704
rect 3852 4696 3860 4704
rect 3916 4696 3924 4704
rect 3980 4696 3988 4704
rect 4012 4696 4020 4704
rect 4060 4716 4068 4724
rect 5020 4716 5028 4724
rect 4172 4696 4180 4704
rect 4188 4696 4196 4704
rect 4348 4694 4356 4702
rect 4588 4696 4596 4704
rect 4620 4696 4628 4704
rect 4780 4696 4788 4704
rect 4860 4696 4868 4704
rect 5340 4716 5348 4724
rect 5548 4716 5556 4724
rect 5564 4716 5572 4724
rect 5820 4716 5828 4724
rect 4924 4694 4932 4702
rect 5068 4696 5076 4704
rect 5100 4696 5108 4704
rect 5116 4696 5124 4704
rect 5164 4696 5172 4704
rect 5180 4696 5188 4704
rect 5212 4696 5220 4704
rect 5276 4696 5284 4704
rect 5308 4696 5316 4704
rect 5404 4694 5412 4702
rect 5660 4696 5668 4704
rect 5724 4694 5732 4702
rect 5868 4696 5876 4704
rect 5900 4696 5908 4704
rect 6140 4694 6148 4702
rect 6204 4696 6212 4704
rect 6268 4696 6276 4704
rect 6572 4716 6580 4724
rect 7164 4716 7172 4724
rect 6332 4696 6340 4704
rect 6348 4696 6356 4704
rect 6444 4696 6452 4704
rect 6492 4696 6500 4704
rect 6652 4696 6660 4704
rect 6716 4696 6724 4704
rect 6796 4696 6804 4704
rect 6988 4696 6996 4704
rect 7052 4694 7060 4702
rect 7132 4696 7140 4704
rect 7164 4696 7172 4704
rect 7244 4696 7252 4704
rect 7292 4696 7300 4704
rect 364 4676 372 4684
rect 540 4676 548 4684
rect 620 4676 628 4684
rect 668 4676 676 4684
rect 716 4676 724 4684
rect 764 4676 772 4684
rect 940 4676 948 4684
rect 1148 4676 1156 4684
rect 1180 4676 1188 4684
rect 1212 4676 1220 4684
rect 1372 4676 1380 4684
rect 1516 4676 1524 4684
rect 1580 4676 1588 4684
rect 1596 4676 1604 4684
rect 1628 4676 1636 4684
rect 1660 4676 1668 4684
rect 1692 4676 1700 4684
rect 1740 4676 1748 4684
rect 1772 4676 1780 4684
rect 1852 4676 1860 4684
rect 2028 4676 2036 4684
rect 2124 4676 2132 4684
rect 2172 4676 2180 4684
rect 2220 4676 2228 4684
rect 2236 4676 2244 4684
rect 2300 4676 2308 4684
rect 2476 4676 2484 4684
rect 2540 4676 2548 4684
rect 2604 4676 2612 4684
rect 2684 4676 2692 4684
rect 2748 4676 2756 4684
rect 2796 4676 2804 4684
rect 2940 4676 2948 4684
rect 3132 4676 3140 4684
rect 3196 4676 3204 4684
rect 3260 4676 3268 4684
rect 3308 4676 3316 4684
rect 3404 4676 3412 4684
rect 3500 4676 3508 4684
rect 3580 4676 3588 4684
rect 3628 4676 3636 4684
rect 3676 4676 3684 4684
rect 3692 4676 3700 4684
rect 3772 4676 3780 4684
rect 3804 4676 3812 4684
rect 3964 4676 3972 4684
rect 3996 4676 4004 4684
rect 4060 4676 4068 4684
rect 4092 4676 4100 4684
rect 4316 4676 4324 4684
rect 4412 4676 4420 4684
rect 4732 4676 4740 4684
rect 4988 4676 4996 4684
rect 5084 4676 5092 4684
rect 5276 4676 5284 4684
rect 5340 4676 5348 4684
rect 5372 4676 5380 4684
rect 5580 4676 5588 4684
rect 5788 4676 5796 4684
rect 5820 4676 5828 4684
rect 5884 4676 5892 4684
rect 6172 4676 6180 4684
rect 6252 4676 6260 4684
rect 6364 4676 6372 4684
rect 6572 4676 6580 4684
rect 6604 4676 6612 4684
rect 6668 4676 6676 4684
rect 6748 4676 6756 4684
rect 7084 4676 7092 4684
rect 7116 4676 7124 4684
rect 76 4656 84 4664
rect 92 4656 100 4664
rect 124 4656 132 4664
rect 156 4656 164 4664
rect 380 4656 388 4664
rect 444 4656 452 4664
rect 476 4656 484 4664
rect 556 4656 564 4664
rect 652 4656 660 4664
rect 684 4656 692 4664
rect 828 4656 836 4664
rect 844 4656 852 4664
rect 972 4656 980 4664
rect 1020 4656 1028 4664
rect 1036 4656 1044 4664
rect 1084 4656 1092 4664
rect 1260 4656 1268 4664
rect 1388 4656 1396 4664
rect 1596 4656 1604 4664
rect 1740 4656 1748 4664
rect 1884 4656 1892 4664
rect 1996 4656 2004 4664
rect 2316 4656 2324 4664
rect 2572 4656 2580 4664
rect 2844 4656 2852 4664
rect 2860 4656 2868 4664
rect 3228 4656 3236 4664
rect 3772 4656 3780 4664
rect 3884 4656 3892 4664
rect 4924 4656 4932 4664
rect 6684 4656 6692 4664
rect 28 4636 36 4644
rect 60 4636 68 4644
rect 188 4636 196 4644
rect 316 4636 324 4644
rect 396 4636 404 4644
rect 492 4636 500 4644
rect 748 4636 756 4644
rect 812 4636 820 4644
rect 1116 4636 1124 4644
rect 1180 4636 1188 4644
rect 1308 4636 1316 4644
rect 1420 4636 1428 4644
rect 1548 4636 1556 4644
rect 1788 4636 1796 4644
rect 1820 4636 1828 4644
rect 1900 4636 1908 4644
rect 2140 4636 2148 4644
rect 2284 4636 2292 4644
rect 2732 4636 2740 4644
rect 2876 4636 2884 4644
rect 3468 4636 3476 4644
rect 3948 4636 3956 4644
rect 4476 4636 4484 4644
rect 5532 4636 5540 4644
rect 5596 4636 5604 4644
rect 6012 4636 6020 4644
rect 6924 4636 6932 4644
rect 2915 4606 2923 4614
rect 2925 4606 2933 4614
rect 2935 4606 2943 4614
rect 2945 4606 2953 4614
rect 2955 4606 2963 4614
rect 2965 4606 2973 4614
rect 5923 4606 5931 4614
rect 5933 4606 5941 4614
rect 5943 4606 5951 4614
rect 5953 4606 5961 4614
rect 5963 4606 5971 4614
rect 5973 4606 5981 4614
rect 732 4576 740 4584
rect 828 4576 836 4584
rect 956 4576 964 4584
rect 2044 4576 2052 4584
rect 2188 4576 2196 4584
rect 2268 4576 2276 4584
rect 2316 4576 2324 4584
rect 2652 4576 2660 4584
rect 3244 4576 3252 4584
rect 3580 4576 3588 4584
rect 3660 4576 3668 4584
rect 3836 4576 3844 4584
rect 4204 4576 4212 4584
rect 5036 4576 5044 4584
rect 5452 4576 5460 4584
rect 5756 4576 5764 4584
rect 6156 4576 6164 4584
rect 6268 4576 6276 4584
rect 6604 4576 6612 4584
rect 6684 4576 6692 4584
rect 6732 4576 6740 4584
rect 7068 4576 7076 4584
rect 7180 4576 7188 4584
rect 60 4556 68 4564
rect 140 4556 148 4564
rect 188 4556 196 4564
rect 220 4556 228 4564
rect 300 4556 308 4564
rect 332 4556 340 4564
rect 444 4556 452 4564
rect 44 4536 52 4544
rect 76 4536 84 4544
rect 396 4536 404 4544
rect 588 4556 596 4564
rect 812 4556 820 4564
rect 892 4556 900 4564
rect 988 4556 996 4564
rect 1116 4556 1124 4564
rect 1548 4556 1556 4564
rect 1644 4556 1652 4564
rect 1676 4556 1684 4564
rect 1868 4556 1876 4564
rect 1980 4556 1988 4564
rect 2140 4556 2148 4564
rect 2732 4556 2740 4564
rect 2748 4556 2756 4564
rect 3724 4556 3732 4564
rect 4060 4556 4068 4564
rect 4268 4556 4276 4564
rect 4796 4556 4804 4564
rect 508 4536 516 4544
rect 652 4536 660 4544
rect 924 4536 932 4544
rect 956 4536 964 4544
rect 972 4536 980 4544
rect 1164 4536 1172 4544
rect 1212 4536 1220 4544
rect 1340 4536 1348 4544
rect 1452 4536 1460 4544
rect 1484 4536 1492 4544
rect 1532 4536 1540 4544
rect 1548 4536 1556 4544
rect 1580 4536 1588 4544
rect 1596 4536 1604 4544
rect 1740 4536 1748 4544
rect 1836 4536 1844 4544
rect 1900 4536 1908 4544
rect 1980 4536 1988 4544
rect 2092 4536 2100 4544
rect 2156 4536 2164 4544
rect 2252 4536 2260 4544
rect 2476 4536 2484 4544
rect 2556 4536 2564 4544
rect 2588 4536 2596 4544
rect 2684 4536 2692 4544
rect 2716 4536 2724 4544
rect 2780 4536 2788 4544
rect 3212 4536 3220 4544
rect 3324 4536 3332 4544
rect 3388 4536 3396 4544
rect 3420 4536 3428 4544
rect 3644 4536 3652 4544
rect 3708 4536 3716 4544
rect 3772 4536 3780 4544
rect 3932 4536 3940 4544
rect 4076 4536 4084 4544
rect 4124 4536 4132 4544
rect 4188 4536 4196 4544
rect 4348 4536 4356 4544
rect 4540 4536 4548 4544
rect 4652 4536 4660 4544
rect 4876 4536 4884 4544
rect 5068 4536 5076 4544
rect 5084 4536 5092 4544
rect 5116 4556 5124 4564
rect 5196 4556 5204 4564
rect 5324 4556 5332 4564
rect 6044 4556 6052 4564
rect 6828 4556 6836 4564
rect 5244 4536 5252 4544
rect 5372 4536 5380 4544
rect 5516 4536 5524 4544
rect 5532 4536 5540 4544
rect 5596 4536 5604 4544
rect 5804 4536 5812 4544
rect 5868 4536 5876 4544
rect 5932 4536 5940 4544
rect 76 4516 84 4524
rect 252 4516 260 4524
rect 300 4516 308 4524
rect 380 4516 388 4524
rect 412 4516 420 4524
rect 492 4516 500 4524
rect 636 4516 644 4524
rect 684 4516 692 4524
rect 764 4516 772 4524
rect 780 4516 788 4524
rect 860 4516 868 4524
rect 972 4516 980 4524
rect 1084 4516 1092 4524
rect 1148 4516 1156 4524
rect 1196 4516 1204 4524
rect 1244 4516 1252 4524
rect 1276 4516 1284 4524
rect 1356 4516 1364 4524
rect 1468 4516 1476 4524
rect 1500 4516 1508 4524
rect 1532 4516 1540 4524
rect 1612 4516 1620 4524
rect 1644 4516 1652 4524
rect 1676 4516 1684 4524
rect 1724 4516 1732 4524
rect 1788 4516 1796 4524
rect 1820 4516 1828 4524
rect 1884 4516 1892 4524
rect 1916 4516 1924 4524
rect 1948 4516 1956 4524
rect 2028 4516 2036 4524
rect 2108 4516 2116 4524
rect 2300 4516 2308 4524
rect 2348 4516 2356 4524
rect 2492 4518 2500 4526
rect 2572 4516 2580 4524
rect 2620 4516 2628 4524
rect 2700 4516 2708 4524
rect 2780 4516 2788 4524
rect 2860 4516 2868 4524
rect 2876 4516 2884 4524
rect 3164 4516 3172 4524
rect 3276 4516 3284 4524
rect 3356 4516 3364 4524
rect 3372 4516 3380 4524
rect 3452 4518 3460 4526
rect 3628 4516 3636 4524
rect 3660 4516 3668 4524
rect 3756 4516 3764 4524
rect 3804 4516 3812 4524
rect 3948 4516 3956 4524
rect 4028 4516 4036 4524
rect 4108 4516 4116 4524
rect 4156 4516 4164 4524
rect 4172 4516 4180 4524
rect 4236 4516 4244 4524
rect 4284 4516 4292 4524
rect 4300 4516 4308 4524
rect 4364 4516 4372 4524
rect 4444 4516 4452 4524
rect 4460 4516 4468 4524
rect 4556 4516 4564 4524
rect 124 4496 132 4504
rect 284 4496 292 4504
rect 348 4496 356 4504
rect 668 4496 676 4504
rect 1100 4496 1108 4504
rect 1244 4496 1252 4504
rect 1260 4496 1268 4504
rect 1420 4496 1428 4504
rect 1692 4496 1700 4504
rect 1804 4496 1812 4504
rect 2044 4496 2052 4504
rect 2604 4496 2612 4504
rect 2668 4496 2676 4504
rect 3292 4496 3300 4504
rect 3772 4496 3780 4504
rect 4620 4516 4628 4524
rect 4636 4516 4644 4524
rect 4748 4516 4756 4524
rect 4940 4516 4948 4524
rect 5052 4516 5060 4524
rect 5148 4516 5156 4524
rect 5228 4516 5236 4524
rect 5260 4516 5268 4524
rect 5324 4518 5332 4526
rect 5516 4516 5524 4524
rect 5548 4516 5556 4524
rect 5596 4516 5604 4524
rect 5612 4516 5620 4524
rect 5628 4516 5636 4524
rect 5660 4516 5668 4524
rect 5676 4516 5684 4524
rect 5708 4516 5716 4524
rect 5724 4516 5732 4524
rect 5788 4516 5796 4524
rect 5820 4516 5828 4524
rect 5468 4496 5476 4504
rect 5884 4516 5892 4524
rect 6108 4536 6116 4544
rect 6220 4536 6228 4544
rect 6396 4536 6404 4544
rect 7052 4536 7060 4544
rect 7100 4556 7108 4564
rect 7132 4536 7140 4544
rect 7212 4556 7220 4564
rect 7404 4536 7412 4544
rect 5996 4516 6004 4524
rect 6092 4516 6100 4524
rect 6124 4516 6132 4524
rect 6220 4516 6228 4524
rect 6236 4516 6244 4524
rect 6300 4516 6308 4524
rect 6172 4496 6180 4504
rect 6396 4516 6404 4524
rect 6476 4516 6484 4524
rect 6524 4516 6532 4524
rect 6636 4516 6644 4524
rect 6652 4516 6660 4524
rect 6700 4516 6708 4524
rect 6716 4516 6724 4524
rect 6764 4516 6772 4524
rect 6796 4516 6804 4524
rect 6844 4516 6852 4524
rect 6860 4516 6868 4524
rect 6908 4516 6916 4524
rect 6940 4516 6948 4524
rect 6956 4516 6964 4524
rect 7004 4516 7012 4524
rect 7036 4516 7044 4524
rect 7132 4516 7140 4524
rect 7148 4516 7156 4524
rect 7244 4516 7252 4524
rect 7260 4516 7268 4524
rect 7308 4516 7316 4524
rect 6380 4496 6388 4504
rect 188 4476 196 4484
rect 508 4476 516 4484
rect 700 4476 708 4484
rect 1036 4476 1044 4484
rect 1068 4476 1076 4484
rect 1292 4476 1300 4484
rect 1340 4476 1348 4484
rect 1772 4476 1780 4484
rect 4588 4476 4596 4484
rect 4668 4476 4676 4484
rect 5884 4476 5892 4484
rect 6332 4476 6340 4484
rect 6412 4476 6420 4484
rect 6444 4476 6452 4484
rect 7292 4476 7300 4484
rect 2108 4456 2116 4464
rect 3052 4456 3060 4464
rect 5452 4456 5460 4464
rect 5820 4456 5828 4464
rect 6972 4456 6980 4464
rect 12 4436 20 4444
rect 92 4436 100 4444
rect 316 4436 324 4444
rect 380 4436 388 4444
rect 492 4436 500 4444
rect 684 4436 692 4444
rect 828 4436 836 4444
rect 1084 4436 1092 4444
rect 1276 4436 1284 4444
rect 1756 4436 1764 4444
rect 1868 4436 1876 4444
rect 2364 4436 2372 4444
rect 2652 4436 2660 4444
rect 2796 4436 2804 4444
rect 3596 4436 3604 4444
rect 4412 4436 4420 4444
rect 5500 4436 5508 4444
rect 5548 4436 5556 4444
rect 6076 4436 6084 4444
rect 6604 4436 6612 4444
rect 6876 4436 6884 4444
rect 1411 4406 1419 4414
rect 1421 4406 1429 4414
rect 1431 4406 1439 4414
rect 1441 4406 1449 4414
rect 1451 4406 1459 4414
rect 1461 4406 1469 4414
rect 4419 4406 4427 4414
rect 4429 4406 4437 4414
rect 4439 4406 4447 4414
rect 4449 4406 4457 4414
rect 4459 4406 4467 4414
rect 4469 4406 4477 4414
rect 988 4376 996 4384
rect 1372 4376 1380 4384
rect 2172 4376 2180 4384
rect 2204 4376 2212 4384
rect 2556 4376 2564 4384
rect 4204 4376 4212 4384
rect 4620 4376 4628 4384
rect 4764 4376 4772 4384
rect 5148 4376 5156 4384
rect 5196 4376 5204 4384
rect 5244 4376 5252 4384
rect 5260 4376 5268 4384
rect 5596 4376 5604 4384
rect 5772 4376 5780 4384
rect 892 4356 900 4364
rect 6092 4356 6100 4364
rect 6732 4356 6740 4364
rect 7196 4356 7204 4364
rect 940 4336 948 4344
rect 1948 4336 1956 4344
rect 2220 4336 2228 4344
rect 4684 4336 4692 4344
rect 5004 4336 5012 4344
rect 5548 4336 5556 4344
rect 6636 4336 6644 4344
rect 6876 4336 6884 4344
rect 76 4316 84 4324
rect 204 4316 212 4324
rect 428 4316 436 4324
rect 476 4316 484 4324
rect 860 4316 868 4324
rect 1292 4316 1300 4324
rect 1724 4316 1732 4324
rect 1740 4316 1748 4324
rect 1980 4316 1988 4324
rect 2348 4316 2356 4324
rect 3580 4316 3588 4324
rect 3724 4316 3732 4324
rect 3884 4316 3892 4324
rect 4140 4316 4148 4324
rect 4172 4316 4180 4324
rect 4540 4316 4548 4324
rect 4636 4316 4644 4324
rect 4700 4316 4708 4324
rect 5036 4316 5044 4324
rect 28 4296 36 4304
rect 108 4296 116 4304
rect 332 4296 340 4304
rect 396 4296 404 4304
rect 556 4296 564 4304
rect 780 4296 788 4304
rect 828 4296 836 4304
rect 876 4296 884 4304
rect 924 4296 932 4304
rect 972 4296 980 4304
rect 1100 4296 1108 4304
rect 1212 4296 1220 4304
rect 1276 4296 1284 4304
rect 1324 4296 1332 4304
rect 1580 4296 1588 4304
rect 1660 4296 1668 4304
rect 1676 4296 1684 4304
rect 1708 4296 1716 4304
rect 1788 4296 1796 4304
rect 1820 4296 1828 4304
rect 1884 4296 1892 4304
rect 1964 4296 1972 4304
rect 2012 4296 2020 4304
rect 2044 4296 2052 4304
rect 2076 4296 2084 4304
rect 2124 4296 2132 4304
rect 2188 4296 2196 4304
rect 2236 4296 2244 4304
rect 2428 4296 2436 4304
rect 2636 4296 2644 4304
rect 2668 4296 2676 4304
rect 2812 4296 2820 4304
rect 2844 4296 2852 4304
rect 3036 4296 3044 4304
rect 3100 4294 3108 4302
rect 3372 4294 3380 4302
rect 3436 4296 3444 4304
rect 3468 4296 3476 4304
rect 3548 4296 3556 4304
rect 3564 4296 3572 4304
rect 3612 4296 3620 4304
rect 3628 4296 3636 4304
rect 3660 4296 3668 4304
rect 3708 4296 3716 4304
rect 3756 4296 3764 4304
rect 3788 4296 3796 4304
rect 3852 4296 3860 4304
rect 4012 4296 4020 4304
rect 4124 4296 4132 4304
rect 4188 4296 4196 4304
rect 4236 4296 4244 4304
rect 4252 4296 4260 4304
rect 4348 4296 4356 4304
rect 4380 4296 4388 4304
rect 4396 4296 4404 4304
rect 4428 4296 4436 4304
rect 4444 4296 4452 4304
rect 4572 4296 4580 4304
rect 4652 4296 4660 4304
rect 4732 4296 4740 4304
rect 4796 4296 4804 4304
rect 4892 4296 4900 4304
rect 4924 4296 4932 4304
rect 5500 4316 5508 4324
rect 5788 4316 5796 4324
rect 5820 4316 5828 4324
rect 5084 4296 5092 4304
rect 5116 4296 5124 4304
rect 5164 4296 5172 4304
rect 5212 4296 5220 4304
rect 5292 4296 5300 4304
rect 5324 4296 5332 4304
rect 5372 4296 5380 4304
rect 5388 4296 5396 4304
rect 5436 4296 5444 4304
rect 5468 4296 5476 4304
rect 5500 4296 5508 4304
rect 5516 4296 5524 4304
rect 5564 4296 5572 4304
rect 5628 4296 5636 4304
rect 5660 4296 5668 4304
rect 5692 4296 5700 4304
rect 5708 4296 5716 4304
rect 5740 4296 5748 4304
rect 5836 4296 5844 4304
rect 5868 4296 5876 4304
rect 5900 4296 5908 4304
rect 6556 4316 6564 4324
rect 6044 4296 6052 4304
rect 6076 4296 6084 4304
rect 6108 4296 6116 4304
rect 6140 4296 6148 4304
rect 6204 4296 6212 4304
rect 6252 4296 6260 4304
rect 6268 4296 6276 4304
rect 6284 4296 6292 4304
rect 6460 4294 6468 4302
rect 6604 4296 6612 4304
rect 6668 4296 6676 4304
rect 6684 4296 6692 4304
rect 6700 4296 6708 4304
rect 6748 4296 6756 4304
rect 6796 4296 6804 4304
rect 6844 4316 6852 4324
rect 7116 4316 7124 4324
rect 6972 4296 6980 4304
rect 7164 4316 7172 4324
rect 7164 4296 7172 4304
rect 7276 4296 7284 4304
rect 7308 4296 7316 4304
rect 12 4276 20 4284
rect 92 4276 100 4284
rect 204 4276 212 4284
rect 316 4276 324 4284
rect 348 4276 356 4284
rect 460 4276 468 4284
rect 508 4276 516 4284
rect 524 4276 532 4284
rect 620 4276 628 4284
rect 636 4276 644 4284
rect 796 4276 804 4284
rect 812 4276 820 4284
rect 876 4276 884 4284
rect 1052 4276 1060 4284
rect 1116 4276 1124 4284
rect 1132 4276 1140 4284
rect 1164 4276 1172 4284
rect 1228 4276 1236 4284
rect 1564 4276 1572 4284
rect 1612 4276 1620 4284
rect 1676 4276 1684 4284
rect 1772 4276 1780 4284
rect 1804 4276 1812 4284
rect 1852 4276 1860 4284
rect 1884 4276 1892 4284
rect 156 4256 164 4264
rect 380 4256 388 4264
rect 396 4256 404 4264
rect 428 4256 436 4264
rect 1004 4256 1012 4264
rect 1020 4256 1028 4264
rect 1148 4256 1156 4264
rect 1196 4256 1204 4264
rect 1260 4256 1268 4264
rect 1308 4256 1316 4264
rect 1356 4256 1364 4264
rect 1388 4256 1396 4264
rect 1628 4256 1636 4264
rect 1836 4256 1844 4264
rect 1916 4256 1924 4264
rect 1932 4256 1940 4264
rect 1996 4256 2004 4264
rect 2092 4276 2100 4284
rect 2124 4276 2132 4284
rect 2140 4276 2148 4284
rect 2172 4276 2180 4284
rect 2300 4276 2308 4284
rect 2444 4276 2452 4284
rect 2540 4276 2548 4284
rect 2860 4276 2868 4284
rect 3068 4276 3076 4284
rect 3132 4276 3140 4284
rect 3324 4276 3332 4284
rect 3404 4276 3412 4284
rect 3452 4276 3460 4284
rect 2092 4256 2100 4264
rect 2316 4256 2324 4264
rect 2348 4256 2356 4264
rect 2428 4256 2436 4264
rect 3644 4276 3652 4284
rect 3772 4276 3780 4284
rect 3788 4276 3796 4284
rect 3836 4276 3844 4284
rect 3884 4276 3892 4284
rect 4060 4276 4068 4284
rect 4300 4276 4308 4284
rect 4364 4276 4372 4284
rect 4460 4276 4468 4284
rect 4588 4276 4596 4284
rect 4748 4276 4756 4284
rect 4828 4276 4836 4284
rect 5004 4276 5012 4284
rect 5036 4276 5044 4284
rect 5100 4276 5108 4284
rect 5404 4276 5412 4284
rect 5452 4276 5460 4284
rect 5612 4276 5620 4284
rect 5676 4276 5684 4284
rect 5836 4276 5844 4284
rect 5852 4276 5860 4284
rect 5916 4276 5924 4284
rect 6012 4276 6020 4284
rect 6044 4276 6052 4284
rect 6060 4276 6068 4284
rect 6124 4276 6132 4284
rect 6172 4276 6180 4284
rect 6444 4276 6452 4284
rect 6524 4276 6532 4284
rect 6572 4276 6580 4284
rect 6620 4276 6628 4284
rect 6780 4276 6788 4284
rect 6844 4276 6852 4284
rect 6876 4276 6884 4284
rect 7020 4276 7028 4284
rect 7084 4276 7092 4284
rect 7180 4276 7188 4284
rect 3500 4256 3508 4264
rect 3820 4256 3828 4264
rect 4284 4256 4292 4264
rect 4956 4256 4964 4264
rect 5724 4256 5732 4264
rect 6172 4256 6180 4264
rect 6316 4256 6324 4264
rect 60 4236 68 4244
rect 188 4236 196 4244
rect 284 4236 292 4244
rect 364 4236 372 4244
rect 588 4236 596 4244
rect 668 4236 676 4244
rect 748 4236 756 4244
rect 1100 4236 1108 4244
rect 1244 4236 1252 4244
rect 1532 4236 1540 4244
rect 1644 4236 1652 4244
rect 1740 4236 1748 4244
rect 2556 4236 2564 4244
rect 2748 4236 2756 4244
rect 2988 4236 2996 4244
rect 3228 4236 3236 4244
rect 3244 4236 3252 4244
rect 3660 4236 3668 4244
rect 3900 4236 3908 4244
rect 4092 4236 4100 4244
rect 4348 4236 4356 4244
rect 4700 4236 4708 4244
rect 5260 4236 5268 4244
rect 5340 4236 5348 4244
rect 5660 4236 5668 4244
rect 5900 4236 5908 4244
rect 5932 4236 5940 4244
rect 5980 4236 5988 4244
rect 6156 4236 6164 4244
rect 6300 4236 6308 4244
rect 6332 4236 6340 4244
rect 2915 4206 2923 4214
rect 2925 4206 2933 4214
rect 2935 4206 2943 4214
rect 2945 4206 2953 4214
rect 2955 4206 2963 4214
rect 2965 4206 2973 4214
rect 5923 4206 5931 4214
rect 5933 4206 5941 4214
rect 5943 4206 5951 4214
rect 5953 4206 5961 4214
rect 5963 4206 5971 4214
rect 5973 4206 5981 4214
rect 1596 4176 1604 4184
rect 1692 4176 1700 4184
rect 2060 4176 2068 4184
rect 2236 4176 2244 4184
rect 2396 4176 2404 4184
rect 2444 4176 2452 4184
rect 2588 4176 2596 4184
rect 2668 4176 2676 4184
rect 2844 4176 2852 4184
rect 3036 4176 3044 4184
rect 3100 4176 3108 4184
rect 3692 4176 3700 4184
rect 3868 4176 3876 4184
rect 3980 4176 3988 4184
rect 4268 4176 4276 4184
rect 4588 4176 4596 4184
rect 4876 4176 4884 4184
rect 4924 4176 4932 4184
rect 5676 4176 5684 4184
rect 5740 4176 5748 4184
rect 6476 4176 6484 4184
rect 6732 4176 6740 4184
rect 7100 4176 7108 4184
rect 12 4156 20 4164
rect 108 4156 116 4164
rect 172 4156 180 4164
rect 204 4156 212 4164
rect 332 4156 340 4164
rect 460 4156 468 4164
rect 572 4156 580 4164
rect 588 4156 596 4164
rect 620 4156 628 4164
rect 716 4156 724 4164
rect 748 4156 756 4164
rect 908 4156 916 4164
rect 1116 4156 1124 4164
rect 1228 4156 1236 4164
rect 1548 4156 1556 4164
rect 1676 4156 1684 4164
rect 1708 4156 1716 4164
rect 1820 4156 1828 4164
rect 1980 4156 1988 4164
rect 2156 4156 2164 4164
rect 2172 4156 2180 4164
rect 2188 4156 2196 4164
rect 2284 4156 2292 4164
rect 2524 4156 2532 4164
rect 2652 4156 2660 4164
rect 3084 4156 3092 4164
rect 3164 4156 3172 4164
rect 3180 4156 3188 4164
rect 3324 4156 3332 4164
rect 3820 4156 3828 4164
rect 4332 4156 4340 4164
rect 4348 4156 4356 4164
rect 4396 4156 4404 4164
rect 4716 4156 4724 4164
rect 4988 4156 4996 4164
rect 5020 4156 5028 4164
rect 5244 4156 5252 4164
rect 5276 4156 5284 4164
rect 5788 4156 5796 4164
rect 5884 4156 5892 4164
rect 5916 4156 5924 4164
rect 6028 4156 6036 4164
rect 6924 4156 6932 4164
rect 7084 4156 7092 4164
rect 124 4136 132 4144
rect 204 4136 212 4144
rect 348 4136 356 4144
rect 588 4136 596 4144
rect 652 4136 660 4144
rect 732 4136 740 4144
rect 812 4136 820 4144
rect 988 4136 996 4144
rect 1164 4136 1172 4144
rect 1196 4136 1204 4144
rect 1212 4136 1220 4144
rect 1244 4136 1252 4144
rect 1340 4136 1348 4144
rect 1516 4136 1524 4144
rect 1564 4136 1572 4144
rect 1660 4136 1668 4144
rect 1740 4136 1748 4144
rect 1836 4136 1844 4144
rect 1868 4136 1876 4144
rect 1900 4136 1908 4144
rect 1916 4136 1924 4144
rect 2044 4136 2052 4144
rect 2252 4136 2260 4144
rect 2540 4136 2548 4144
rect 2652 4136 2660 4144
rect 2716 4136 2724 4144
rect 2764 4136 2772 4144
rect 2860 4136 2868 4144
rect 2892 4136 2900 4144
rect 3052 4136 3060 4144
rect 3148 4136 3156 4144
rect 3388 4136 3396 4144
rect 3420 4136 3428 4144
rect 3484 4136 3492 4144
rect 3596 4136 3604 4144
rect 3612 4136 3620 4144
rect 3740 4136 3748 4144
rect 3804 4136 3812 4144
rect 3900 4136 3908 4144
rect 3948 4136 3956 4144
rect 4188 4136 4196 4144
rect 4236 4136 4244 4144
rect 4380 4136 4388 4144
rect 4892 4136 4900 4144
rect 4908 4136 4916 4144
rect 4988 4136 4996 4144
rect 5020 4136 5028 4144
rect 5100 4136 5108 4144
rect 5244 4136 5252 4144
rect 5276 4136 5284 4144
rect 5388 4136 5396 4144
rect 5484 4136 5492 4144
rect 5516 4136 5524 4144
rect 5804 4136 5812 4144
rect 5868 4136 5876 4144
rect 6044 4136 6052 4144
rect 6108 4136 6116 4144
rect 6124 4136 6132 4144
rect 6188 4136 6196 4144
rect 6284 4136 6292 4144
rect 6412 4136 6420 4144
rect 6460 4136 6468 4144
rect 6636 4136 6644 4144
rect 6684 4136 6692 4144
rect 6716 4136 6724 4144
rect 6828 4136 6836 4144
rect 7004 4136 7012 4144
rect 7052 4136 7060 4144
rect 7228 4136 7236 4144
rect 76 4116 84 4124
rect 172 4116 180 4124
rect 236 4116 244 4124
rect 316 4116 324 4124
rect 412 4116 420 4124
rect 524 4116 532 4124
rect 540 4116 548 4124
rect 652 4116 660 4124
rect 700 4116 708 4124
rect 796 4116 804 4124
rect 908 4116 916 4124
rect 940 4116 948 4124
rect 1004 4116 1012 4124
rect 1036 4116 1044 4124
rect 1068 4116 1076 4124
rect 1148 4116 1156 4124
rect 268 4096 276 4104
rect 284 4096 292 4104
rect 748 4096 756 4104
rect 860 4096 868 4104
rect 924 4096 932 4104
rect 1052 4096 1060 4104
rect 1404 4116 1412 4124
rect 1468 4116 1476 4124
rect 1516 4116 1524 4124
rect 1564 4116 1572 4124
rect 1740 4116 1748 4124
rect 1756 4116 1764 4124
rect 1788 4096 1796 4104
rect 1852 4116 1860 4124
rect 2092 4116 2100 4124
rect 2124 4116 2132 4124
rect 2252 4116 2260 4124
rect 2300 4116 2308 4124
rect 2380 4116 2388 4124
rect 2428 4116 2436 4124
rect 2476 4116 2484 4124
rect 2492 4116 2500 4124
rect 2556 4116 2564 4124
rect 2604 4116 2612 4124
rect 2700 4116 2708 4124
rect 2748 4116 2756 4124
rect 2780 4116 2788 4124
rect 2876 4116 2884 4124
rect 2908 4116 2916 4124
rect 3068 4116 3076 4124
rect 3132 4116 3140 4124
rect 3148 4116 3156 4124
rect 3324 4118 3332 4126
rect 1948 4096 1956 4104
rect 1964 4096 1972 4104
rect 2060 4096 2068 4104
rect 2220 4096 2228 4104
rect 2588 4096 2596 4104
rect 2812 4096 2820 4104
rect 2988 4096 2996 4104
rect 3420 4096 3428 4104
rect 3468 4116 3476 4124
rect 3500 4116 3508 4124
rect 3516 4116 3524 4124
rect 3564 4116 3572 4124
rect 3612 4116 3620 4124
rect 3660 4116 3668 4124
rect 3676 4116 3684 4124
rect 3724 4116 3732 4124
rect 3756 4116 3764 4124
rect 3852 4116 3860 4124
rect 3916 4116 3924 4124
rect 4060 4116 4068 4124
rect 4108 4118 4116 4126
rect 4204 4116 4212 4124
rect 4252 4116 4260 4124
rect 4300 4116 4308 4124
rect 4332 4116 4340 4124
rect 4364 4116 4372 4124
rect 4396 4116 4404 4124
rect 4428 4116 4436 4124
rect 4556 4116 4564 4124
rect 4700 4116 4708 4124
rect 4812 4116 4820 4124
rect 4844 4116 4852 4124
rect 4924 4116 4932 4124
rect 4972 4116 4980 4124
rect 4988 4116 4996 4124
rect 5068 4116 5076 4124
rect 5116 4116 5124 4124
rect 5180 4116 5188 4124
rect 5212 4116 5220 4124
rect 5244 4116 5252 4124
rect 5308 4116 5316 4124
rect 5356 4116 5364 4124
rect 5372 4116 5380 4124
rect 3868 4096 3876 4104
rect 3964 4096 3972 4104
rect 4172 4096 4180 4104
rect 4524 4096 4532 4104
rect 5036 4096 5044 4104
rect 5148 4096 5156 4104
rect 5420 4096 5428 4104
rect 5468 4116 5476 4124
rect 5548 4118 5556 4126
rect 5612 4116 5620 4124
rect 5708 4116 5716 4124
rect 5756 4116 5764 4124
rect 5852 4116 5860 4124
rect 5884 4116 5892 4124
rect 5996 4116 6004 4124
rect 6092 4116 6100 4124
rect 6156 4116 6164 4124
rect 6204 4116 6212 4124
rect 6252 4116 6260 4124
rect 6268 4116 6276 4124
rect 6300 4116 6308 4124
rect 6332 4116 6340 4124
rect 6396 4116 6404 4124
rect 6588 4116 6596 4124
rect 6700 4116 6708 4124
rect 6860 4118 6868 4126
rect 6956 4116 6964 4124
rect 6972 4116 6980 4124
rect 7020 4116 7028 4124
rect 7084 4116 7092 4124
rect 7212 4116 7220 4124
rect 7308 4116 7316 4124
rect 5468 4096 5476 4104
rect 5740 4096 5748 4104
rect 6124 4096 6132 4104
rect 6364 4096 6372 4104
rect 6428 4096 6436 4104
rect 6668 4096 6676 4104
rect 7292 4096 7300 4104
rect 76 4076 84 4084
rect 588 4076 596 4084
rect 956 4076 964 4084
rect 1084 4076 1092 4084
rect 2044 4076 2052 4084
rect 3196 4076 3204 4084
rect 4012 4076 4020 4084
rect 4620 4076 4628 4084
rect 6460 4076 6468 4084
rect 6508 4076 6516 4084
rect 7324 4076 7332 4084
rect 5180 4056 5188 4064
rect 6236 4056 6244 4064
rect 7100 4056 7108 4064
rect 188 4036 196 4044
rect 236 4036 244 4044
rect 444 4036 452 4044
rect 476 4036 484 4044
rect 492 4036 500 4044
rect 652 4036 660 4044
rect 668 4036 676 4044
rect 940 4036 948 4044
rect 1068 4036 1076 4044
rect 1132 4036 1140 4044
rect 1276 4036 1284 4044
rect 1356 4036 1364 4044
rect 1900 4036 1908 4044
rect 2332 4036 2340 4044
rect 2348 4036 2356 4044
rect 3756 4036 3764 4044
rect 4780 4036 4788 4044
rect 5820 4036 5828 4044
rect 6060 4036 6068 4044
rect 6300 4036 6308 4044
rect 7308 4036 7316 4044
rect 1411 4006 1419 4014
rect 1421 4006 1429 4014
rect 1431 4006 1439 4014
rect 1441 4006 1449 4014
rect 1451 4006 1459 4014
rect 1461 4006 1469 4014
rect 4419 4006 4427 4014
rect 4429 4006 4437 4014
rect 4439 4006 4447 4014
rect 4449 4006 4457 4014
rect 4459 4006 4467 4014
rect 4469 4006 4477 4014
rect 844 3976 852 3984
rect 2236 3976 2244 3984
rect 3436 3976 3444 3984
rect 3532 3976 3540 3984
rect 3772 3976 3780 3984
rect 4220 3976 4228 3984
rect 4620 3976 4628 3984
rect 4748 3976 4756 3984
rect 4764 3976 4772 3984
rect 4828 3976 4836 3984
rect 4892 3976 4900 3984
rect 5708 3976 5716 3984
rect 5996 3976 6004 3984
rect 6012 3976 6020 3984
rect 6188 3976 6196 3984
rect 6252 3976 6260 3984
rect 6412 3976 6420 3984
rect 7148 3976 7156 3984
rect 7212 3976 7220 3984
rect 4316 3956 4324 3964
rect 4700 3956 4708 3964
rect 4924 3956 4932 3964
rect 460 3936 468 3944
rect 1580 3936 1588 3944
rect 2108 3936 2116 3944
rect 3372 3936 3380 3944
rect 3836 3936 3844 3944
rect 4044 3936 4052 3944
rect 5644 3936 5652 3944
rect 6924 3936 6932 3944
rect 124 3916 132 3924
rect 396 3916 404 3924
rect 508 3916 516 3924
rect 972 3916 980 3924
rect 156 3896 164 3904
rect 220 3896 228 3904
rect 12 3876 20 3884
rect 108 3876 116 3884
rect 172 3876 180 3884
rect 300 3896 308 3904
rect 380 3896 388 3904
rect 412 3896 420 3904
rect 444 3896 452 3904
rect 460 3896 468 3904
rect 540 3896 548 3904
rect 572 3896 580 3904
rect 604 3896 612 3904
rect 764 3896 772 3904
rect 940 3896 948 3904
rect 1036 3916 1044 3924
rect 1068 3916 1076 3924
rect 1164 3916 1172 3924
rect 1228 3916 1236 3924
rect 1308 3916 1316 3924
rect 1612 3916 1620 3924
rect 2060 3916 2068 3924
rect 1132 3896 1140 3904
rect 1180 3896 1188 3904
rect 1244 3896 1252 3904
rect 1404 3896 1412 3904
rect 1516 3896 1524 3904
rect 1580 3896 1588 3904
rect 1692 3896 1700 3904
rect 1804 3896 1812 3904
rect 1852 3896 1860 3904
rect 2028 3896 2036 3904
rect 2092 3896 2100 3904
rect 2188 3916 2196 3924
rect 2636 3916 2644 3924
rect 2812 3916 2820 3924
rect 3116 3916 3124 3924
rect 2252 3896 2260 3904
rect 2460 3896 2468 3904
rect 2588 3896 2596 3904
rect 2668 3896 2676 3904
rect 2748 3896 2756 3904
rect 2780 3896 2788 3904
rect 2892 3896 2900 3904
rect 3628 3916 3636 3924
rect 3164 3896 3172 3904
rect 3292 3896 3300 3904
rect 3404 3896 3412 3904
rect 3452 3896 3460 3904
rect 3468 3896 3476 3904
rect 3484 3896 3492 3904
rect 3548 3896 3556 3904
rect 3564 3896 3572 3904
rect 3644 3896 3652 3904
rect 3724 3896 3732 3904
rect 3740 3896 3748 3904
rect 3756 3896 3764 3904
rect 3804 3896 3812 3904
rect 3948 3896 3956 3904
rect 4044 3896 4052 3904
rect 4092 3916 4100 3924
rect 4252 3916 4260 3924
rect 5036 3916 5044 3924
rect 4140 3896 4148 3904
rect 4156 3896 4164 3904
rect 4284 3896 4292 3904
rect 4348 3896 4356 3904
rect 4556 3894 4564 3902
rect 4652 3896 4660 3904
rect 4668 3896 4676 3904
rect 4716 3896 4724 3904
rect 4796 3896 4804 3904
rect 4860 3896 4868 3904
rect 4908 3896 4916 3904
rect 4972 3896 4980 3904
rect 5004 3896 5012 3904
rect 5084 3896 5092 3904
rect 5164 3896 5172 3904
rect 5228 3894 5236 3902
rect 5324 3896 5332 3904
rect 5388 3896 5396 3904
rect 5500 3896 5508 3904
rect 5628 3896 5636 3904
rect 5692 3896 5700 3904
rect 5772 3896 5780 3904
rect 5820 3896 5828 3904
rect 5900 3896 5908 3904
rect 6044 3896 6052 3904
rect 6076 3896 6084 3904
rect 6124 3896 6132 3904
rect 6140 3896 6148 3904
rect 6172 3896 6180 3904
rect 6220 3896 6228 3904
rect 6236 3896 6244 3904
rect 6284 3896 6292 3904
rect 6300 3896 6308 3904
rect 6364 3896 6372 3904
rect 6396 3896 6404 3904
rect 6524 3896 6532 3904
rect 6636 3896 6644 3904
rect 6652 3896 6660 3904
rect 6732 3896 6740 3904
rect 6796 3896 6804 3904
rect 6860 3896 6868 3904
rect 6908 3896 6916 3904
rect 7004 3896 7012 3904
rect 7116 3896 7124 3904
rect 7164 3896 7172 3904
rect 7228 3896 7236 3904
rect 268 3876 276 3884
rect 332 3876 340 3884
rect 444 3876 452 3884
rect 620 3876 628 3884
rect 636 3880 644 3888
rect 700 3876 708 3884
rect 828 3876 836 3884
rect 892 3876 900 3884
rect 924 3876 932 3884
rect 1020 3876 1028 3884
rect 1068 3876 1076 3884
rect 220 3856 228 3864
rect 268 3856 276 3864
rect 300 3856 308 3864
rect 332 3856 340 3864
rect 348 3856 356 3864
rect 492 3856 500 3864
rect 572 3856 580 3864
rect 684 3856 692 3864
rect 764 3856 772 3864
rect 828 3856 836 3864
rect 908 3856 916 3864
rect 1116 3876 1124 3884
rect 1180 3876 1188 3884
rect 1196 3876 1204 3884
rect 1276 3876 1284 3884
rect 1340 3876 1348 3884
rect 1228 3856 1236 3864
rect 1292 3856 1300 3864
rect 1356 3856 1364 3864
rect 1388 3876 1396 3884
rect 1548 3876 1556 3884
rect 1724 3876 1732 3884
rect 1772 3876 1780 3884
rect 1868 3876 1876 3884
rect 2060 3876 2068 3884
rect 2220 3876 2228 3884
rect 2316 3876 2324 3884
rect 2412 3876 2420 3884
rect 2428 3876 2436 3884
rect 2476 3876 2484 3884
rect 2572 3876 2580 3884
rect 2684 3876 2692 3884
rect 2732 3876 2740 3884
rect 2764 3876 2772 3884
rect 2892 3876 2900 3884
rect 3020 3876 3028 3884
rect 3116 3876 3124 3884
rect 3180 3876 3188 3884
rect 3212 3876 3220 3884
rect 3580 3876 3588 3884
rect 3996 3876 4004 3884
rect 4028 3876 4036 3884
rect 4140 3876 4148 3884
rect 4236 3876 4244 3884
rect 4300 3876 4308 3884
rect 4508 3876 4516 3884
rect 4588 3876 4596 3884
rect 4844 3876 4852 3884
rect 4956 3876 4964 3884
rect 5324 3876 5332 3884
rect 5372 3876 5380 3884
rect 5516 3876 5524 3884
rect 5692 3876 5700 3884
rect 1548 3856 1556 3864
rect 1628 3856 1636 3864
rect 1708 3856 1716 3864
rect 1980 3856 1988 3864
rect 2252 3856 2260 3864
rect 2620 3856 2628 3864
rect 2700 3856 2708 3864
rect 3692 3856 3700 3864
rect 4940 3856 4948 3864
rect 5292 3856 5300 3864
rect 5596 3856 5604 3864
rect 6332 3856 6340 3864
rect 6396 3876 6404 3884
rect 6508 3876 6516 3884
rect 6604 3876 6612 3884
rect 6700 3876 6708 3884
rect 6780 3876 6788 3884
rect 6828 3876 6836 3884
rect 6700 3856 6708 3864
rect 7084 3876 7092 3884
rect 7388 3876 7396 3884
rect 6876 3856 6884 3864
rect 7212 3856 7220 3864
rect 76 3836 84 3844
rect 124 3836 132 3844
rect 668 3836 676 3844
rect 732 3836 740 3844
rect 748 3836 756 3844
rect 860 3836 868 3844
rect 1004 3836 1012 3844
rect 1036 3836 1044 3844
rect 1308 3836 1316 3844
rect 1436 3836 1444 3844
rect 1532 3836 1540 3844
rect 1644 3836 1652 3844
rect 1660 3836 1668 3844
rect 1756 3836 1764 3844
rect 1820 3836 1828 3844
rect 1932 3836 1940 3844
rect 2172 3836 2180 3844
rect 2300 3836 2308 3844
rect 2348 3836 2356 3844
rect 2540 3836 2548 3844
rect 2636 3836 2644 3844
rect 2716 3836 2724 3844
rect 2812 3836 2820 3844
rect 3020 3836 3028 3844
rect 3628 3836 3636 3844
rect 3660 3836 3668 3844
rect 3708 3836 3716 3844
rect 4188 3836 4196 3844
rect 4252 3836 4260 3844
rect 4428 3836 4436 3844
rect 4972 3836 4980 3844
rect 5100 3836 5108 3844
rect 5404 3836 5412 3844
rect 6092 3836 6100 3844
rect 6684 3836 6692 3844
rect 6764 3836 6772 3844
rect 2915 3806 2923 3814
rect 2925 3806 2933 3814
rect 2935 3806 2943 3814
rect 2945 3806 2953 3814
rect 2955 3806 2963 3814
rect 2965 3806 2973 3814
rect 5923 3806 5931 3814
rect 5933 3806 5941 3814
rect 5943 3806 5951 3814
rect 5953 3806 5961 3814
rect 5963 3806 5971 3814
rect 5973 3806 5981 3814
rect 700 3776 708 3784
rect 796 3776 804 3784
rect 972 3776 980 3784
rect 2108 3776 2116 3784
rect 2460 3776 2468 3784
rect 2652 3776 2660 3784
rect 3148 3776 3156 3784
rect 3308 3776 3316 3784
rect 3836 3776 3844 3784
rect 4252 3776 4260 3784
rect 4780 3776 4788 3784
rect 5100 3776 5108 3784
rect 5260 3776 5268 3784
rect 5500 3776 5508 3784
rect 5628 3776 5636 3784
rect 5708 3776 5716 3784
rect 5756 3776 5764 3784
rect 6588 3776 6596 3784
rect 6652 3776 6660 3784
rect 6908 3776 6916 3784
rect 6956 3776 6964 3784
rect 7180 3776 7188 3784
rect 60 3756 68 3764
rect 76 3756 84 3764
rect 188 3756 196 3764
rect 300 3756 308 3764
rect 444 3756 452 3764
rect 508 3756 516 3764
rect 716 3756 724 3764
rect 732 3756 740 3764
rect 876 3756 884 3764
rect 1036 3756 1044 3764
rect 1052 3756 1060 3764
rect 1068 3756 1076 3764
rect 1404 3756 1412 3764
rect 1436 3756 1444 3764
rect 1532 3756 1540 3764
rect 1676 3756 1684 3764
rect 1740 3756 1748 3764
rect 1836 3756 1844 3764
rect 1852 3756 1860 3764
rect 2060 3756 2068 3764
rect 2204 3756 2212 3764
rect 2220 3756 2228 3764
rect 2844 3756 2852 3764
rect 3372 3756 3380 3764
rect 3532 3756 3540 3764
rect 4236 3756 4244 3764
rect 4284 3756 4292 3764
rect 4668 3756 4676 3764
rect 4972 3756 4980 3764
rect 5036 3756 5044 3764
rect 28 3736 36 3744
rect 172 3736 180 3744
rect 220 3736 228 3744
rect 252 3736 260 3744
rect 364 3736 372 3744
rect 524 3736 532 3744
rect 604 3736 612 3744
rect 684 3736 692 3744
rect 812 3736 820 3744
rect 908 3736 916 3744
rect 1020 3736 1028 3744
rect 1100 3736 1108 3744
rect 1196 3736 1204 3744
rect 1244 3736 1252 3744
rect 1260 3736 1268 3744
rect 1356 3736 1364 3744
rect 1388 3736 1396 3744
rect 1596 3736 1604 3744
rect 1804 3736 1812 3744
rect 1948 3736 1956 3744
rect 2044 3736 2052 3744
rect 2172 3736 2180 3744
rect 2300 3736 2308 3744
rect 2396 3736 2404 3744
rect 2620 3736 2628 3744
rect 2812 3736 2820 3744
rect 2876 3736 2884 3744
rect 2892 3736 2900 3744
rect 3164 3736 3172 3744
rect 3260 3736 3268 3744
rect 3292 3736 3300 3744
rect 3580 3736 3588 3744
rect 3644 3736 3652 3744
rect 3708 3736 3716 3744
rect 3724 3736 3732 3744
rect 3820 3736 3828 3744
rect 3948 3736 3956 3744
rect 4028 3736 4036 3744
rect 4092 3736 4100 3744
rect 4108 3736 4116 3744
rect 4172 3736 4180 3744
rect 4332 3736 4340 3744
rect 4508 3736 4516 3744
rect 4652 3736 4660 3744
rect 4716 3736 4724 3744
rect 4732 3736 4740 3744
rect 4828 3736 4836 3744
rect 5052 3736 5060 3744
rect 5084 3736 5092 3744
rect 5212 3736 5220 3744
rect 5308 3736 5316 3744
rect 5420 3736 5428 3744
rect 5484 3736 5492 3744
rect 5532 3756 5540 3764
rect 6108 3756 6116 3764
rect 6300 3756 6308 3764
rect 6876 3756 6884 3764
rect 5932 3736 5940 3744
rect 6124 3736 6132 3744
rect 6156 3736 6164 3744
rect 6188 3736 6196 3744
rect 6252 3736 6260 3744
rect 6316 3736 6324 3744
rect 6380 3736 6388 3744
rect 6444 3736 6452 3744
rect 6460 3736 6468 3744
rect 6812 3736 6820 3744
rect 7084 3756 7092 3764
rect 6924 3736 6932 3744
rect 7164 3736 7172 3744
rect 7212 3756 7220 3764
rect 7388 3736 7396 3744
rect 12 3716 20 3724
rect 108 3716 116 3724
rect 268 3716 276 3724
rect 348 3716 356 3724
rect 380 3716 388 3724
rect 492 3716 500 3724
rect 620 3716 628 3724
rect 652 3716 660 3724
rect 668 3716 676 3724
rect 764 3716 772 3724
rect 828 3716 836 3724
rect 876 3716 884 3724
rect 1020 3716 1028 3724
rect 1372 3716 1380 3724
rect 1436 3716 1444 3724
rect 1532 3716 1540 3724
rect 1596 3716 1604 3724
rect 1612 3716 1620 3724
rect 1644 3716 1652 3724
rect 1708 3716 1716 3724
rect 1740 3716 1748 3724
rect 1788 3716 1796 3724
rect 1820 3716 1828 3724
rect 1868 3716 1876 3724
rect 1916 3716 1924 3724
rect 1964 3716 1972 3724
rect 2300 3716 2308 3724
rect 2444 3716 2452 3724
rect 2588 3718 2596 3726
rect 2780 3718 2788 3726
rect 2844 3716 2852 3724
rect 2892 3716 2900 3724
rect 3036 3716 3044 3724
rect 3084 3716 3092 3724
rect 3180 3716 3188 3724
rect 140 3696 148 3704
rect 220 3696 228 3704
rect 252 3696 260 3704
rect 316 3696 324 3704
rect 860 3696 868 3704
rect 1212 3696 1220 3704
rect 1548 3696 1556 3704
rect 1580 3696 1588 3704
rect 1612 3696 1620 3704
rect 3180 3696 3188 3704
rect 3276 3716 3284 3724
rect 3340 3716 3348 3724
rect 3404 3716 3412 3724
rect 3452 3716 3460 3724
rect 3468 3716 3476 3724
rect 3500 3716 3508 3724
rect 3548 3716 3556 3724
rect 3564 3716 3572 3724
rect 3580 3716 3588 3724
rect 3660 3716 3668 3724
rect 3692 3716 3700 3724
rect 3228 3696 3236 3704
rect 3628 3696 3636 3704
rect 3756 3696 3764 3704
rect 3804 3716 3812 3724
rect 3948 3716 3956 3724
rect 4044 3716 4052 3724
rect 4076 3716 4084 3724
rect 4124 3716 4132 3724
rect 4172 3716 4180 3724
rect 4188 3716 4196 3724
rect 4268 3716 4276 3724
rect 4316 3716 4324 3724
rect 4540 3718 4548 3726
rect 4636 3716 4644 3724
rect 4700 3716 4708 3724
rect 4284 3696 4292 3704
rect 4604 3696 4612 3704
rect 4668 3696 4676 3704
rect 4764 3696 4772 3704
rect 4812 3716 4820 3724
rect 4924 3716 4932 3724
rect 5068 3716 5076 3724
rect 5100 3716 5108 3724
rect 5132 3716 5140 3724
rect 5212 3716 5220 3724
rect 5228 3716 5236 3724
rect 5244 3716 5252 3724
rect 5340 3716 5348 3724
rect 5388 3716 5396 3724
rect 5404 3716 5412 3724
rect 5452 3716 5460 3724
rect 5468 3716 5476 3724
rect 5564 3716 5572 3724
rect 5580 3716 5588 3724
rect 5660 3716 5668 3724
rect 5676 3716 5684 3724
rect 5724 3716 5732 3724
rect 5804 3716 5812 3724
rect 5820 3716 5828 3724
rect 5836 3716 5844 3724
rect 5884 3716 5892 3724
rect 5996 3716 6004 3724
rect 6044 3716 6052 3724
rect 6060 3716 6068 3724
rect 6076 3716 6084 3724
rect 6172 3716 6180 3724
rect 6220 3716 6228 3724
rect 6236 3716 6244 3724
rect 6268 3716 6276 3724
rect 6364 3716 6372 3724
rect 5164 3696 5172 3704
rect 6204 3696 6212 3704
rect 6428 3716 6436 3724
rect 6460 3716 6468 3724
rect 6524 3716 6532 3724
rect 6540 3716 6548 3724
rect 6556 3716 6564 3724
rect 6572 3716 6580 3724
rect 6620 3716 6628 3724
rect 6764 3716 6772 3724
rect 6844 3716 6852 3724
rect 6940 3716 6948 3724
rect 7068 3716 7076 3724
rect 7148 3716 7156 3724
rect 7244 3716 7252 3724
rect 444 3676 452 3684
rect 2204 3676 2212 3684
rect 3804 3676 3812 3684
rect 4044 3676 4052 3684
rect 4188 3676 4196 3684
rect 4412 3676 4420 3684
rect 4636 3676 4644 3684
rect 6428 3676 6436 3684
rect 6332 3656 6340 3664
rect 60 3636 68 3644
rect 92 3636 100 3644
rect 156 3636 164 3644
rect 236 3636 244 3644
rect 348 3636 356 3644
rect 412 3636 420 3644
rect 460 3636 468 3644
rect 588 3636 596 3644
rect 748 3636 756 3644
rect 796 3636 804 3644
rect 892 3636 900 3644
rect 1084 3636 1092 3644
rect 1164 3636 1172 3644
rect 1292 3636 1300 3644
rect 1644 3636 1652 3644
rect 1724 3636 1732 3644
rect 1900 3636 1908 3644
rect 1996 3636 2004 3644
rect 2012 3636 2020 3644
rect 2236 3636 2244 3644
rect 2252 3636 2260 3644
rect 2332 3636 2340 3644
rect 2412 3636 2420 3644
rect 3436 3636 3444 3644
rect 3596 3636 3604 3644
rect 3660 3636 3668 3644
rect 4156 3636 4164 3644
rect 4844 3636 4852 3644
rect 5612 3636 5620 3644
rect 5628 3636 5636 3644
rect 5772 3636 5780 3644
rect 5852 3636 5860 3644
rect 7276 3636 7284 3644
rect 1411 3606 1419 3614
rect 1421 3606 1429 3614
rect 1431 3606 1439 3614
rect 1441 3606 1449 3614
rect 1451 3606 1459 3614
rect 1461 3606 1469 3614
rect 4419 3606 4427 3614
rect 4429 3606 4437 3614
rect 4439 3606 4447 3614
rect 4449 3606 4457 3614
rect 4459 3606 4467 3614
rect 4469 3606 4477 3614
rect 284 3576 292 3584
rect 1388 3576 1396 3584
rect 2636 3576 2644 3584
rect 2892 3576 2900 3584
rect 3932 3576 3940 3584
rect 4028 3576 4036 3584
rect 4140 3576 4148 3584
rect 4364 3576 4372 3584
rect 4684 3576 4692 3584
rect 4860 3576 4868 3584
rect 4988 3576 4996 3584
rect 5228 3576 5236 3584
rect 6284 3576 6292 3584
rect 7004 3576 7012 3584
rect 7164 3576 7172 3584
rect 7340 3576 7348 3584
rect 236 3556 244 3564
rect 4092 3556 4100 3564
rect 556 3536 564 3544
rect 1756 3536 1764 3544
rect 1868 3536 1876 3544
rect 2460 3536 2468 3544
rect 3468 3536 3476 3544
rect 3692 3536 3700 3544
rect 4556 3536 4564 3544
rect 5468 3536 5476 3544
rect 6012 3536 6020 3544
rect 6332 3536 6340 3544
rect 6748 3536 6756 3544
rect 268 3516 276 3524
rect 380 3516 388 3524
rect 844 3516 852 3524
rect 1404 3516 1412 3524
rect 1788 3516 1796 3524
rect 1804 3516 1812 3524
rect 1900 3516 1908 3524
rect 2012 3516 2020 3524
rect 76 3496 84 3504
rect 108 3496 116 3504
rect 236 3496 244 3504
rect 316 3496 324 3504
rect 396 3496 404 3504
rect 428 3496 436 3504
rect 492 3496 500 3504
rect 604 3496 612 3504
rect 684 3496 692 3504
rect 716 3496 724 3504
rect 828 3496 836 3504
rect 844 3496 852 3504
rect 876 3496 884 3504
rect 988 3496 996 3504
rect 1020 3496 1028 3504
rect 1164 3496 1172 3504
rect 1196 3496 1204 3504
rect 1260 3496 1268 3504
rect 1292 3496 1300 3504
rect 1324 3496 1332 3504
rect 1676 3496 1684 3504
rect 1756 3496 1764 3504
rect 1884 3496 1892 3504
rect 1916 3496 1924 3504
rect 2060 3496 2068 3504
rect 2156 3496 2164 3504
rect 2188 3496 2196 3504
rect 2252 3496 2260 3504
rect 2364 3496 2372 3504
rect 2412 3496 2420 3504
rect 2508 3496 2516 3504
rect 2668 3496 2676 3504
rect 3724 3516 3732 3524
rect 4508 3516 4516 3524
rect 4620 3516 4628 3524
rect 4828 3516 4836 3524
rect 5660 3516 5668 3524
rect 6140 3516 6148 3524
rect 6428 3516 6436 3524
rect 6652 3516 6660 3524
rect 7116 3516 7124 3524
rect 60 3476 68 3484
rect 108 3476 116 3484
rect 156 3476 164 3484
rect 332 3476 340 3484
rect 348 3476 356 3484
rect 508 3476 516 3484
rect 652 3476 660 3484
rect 668 3476 676 3484
rect 828 3476 836 3484
rect 1036 3476 1044 3484
rect 1068 3476 1076 3484
rect 1148 3476 1156 3484
rect 1212 3476 1220 3484
rect 1276 3476 1284 3484
rect 1308 3476 1316 3484
rect 1532 3476 1540 3484
rect 1628 3476 1636 3484
rect 12 3456 20 3464
rect 140 3456 148 3464
rect 412 3456 420 3464
rect 428 3456 436 3464
rect 476 3456 484 3464
rect 540 3456 548 3464
rect 556 3456 564 3464
rect 716 3456 724 3464
rect 764 3456 772 3464
rect 780 3456 788 3464
rect 812 3456 820 3464
rect 924 3456 932 3464
rect 940 3456 948 3464
rect 1052 3456 1060 3464
rect 1100 3456 1108 3464
rect 1132 3456 1140 3464
rect 1196 3456 1204 3464
rect 1228 3456 1236 3464
rect 1372 3456 1380 3464
rect 1436 3456 1444 3464
rect 1644 3456 1652 3464
rect 1740 3476 1748 3484
rect 1948 3476 1956 3484
rect 1964 3480 1972 3488
rect 3052 3494 3060 3502
rect 3180 3496 3188 3504
rect 3212 3496 3220 3504
rect 3308 3496 3316 3504
rect 3340 3496 3348 3504
rect 3372 3496 3380 3504
rect 3404 3496 3412 3504
rect 3484 3496 3492 3504
rect 3500 3496 3508 3504
rect 3532 3496 3540 3504
rect 3564 3496 3572 3504
rect 3612 3496 3620 3504
rect 3644 3496 3652 3504
rect 3692 3496 3700 3504
rect 3772 3496 3780 3504
rect 3788 3496 3796 3504
rect 3852 3496 3860 3504
rect 3884 3496 3892 3504
rect 3900 3496 3908 3504
rect 3916 3496 3924 3504
rect 3964 3496 3972 3504
rect 3996 3496 4004 3504
rect 4012 3496 4020 3504
rect 4060 3496 4068 3504
rect 4124 3496 4132 3504
rect 4204 3496 4212 3504
rect 4252 3496 4260 3504
rect 4348 3496 4356 3504
rect 4396 3496 4404 3504
rect 4412 3496 4420 3504
rect 4524 3496 4532 3504
rect 4556 3496 4564 3504
rect 4588 3496 4596 3504
rect 4652 3496 4660 3504
rect 4716 3496 4724 3504
rect 4732 3496 4740 3504
rect 4748 3496 4756 3504
rect 4796 3496 4804 3504
rect 4860 3496 4868 3504
rect 4924 3496 4932 3504
rect 4940 3496 4948 3504
rect 5004 3496 5012 3504
rect 5116 3496 5124 3504
rect 5276 3496 5284 3504
rect 5340 3496 5348 3504
rect 5388 3496 5396 3504
rect 5452 3496 5460 3504
rect 5580 3496 5588 3504
rect 5692 3496 5700 3504
rect 5724 3496 5732 3504
rect 5820 3496 5828 3504
rect 5900 3496 5908 3504
rect 6092 3496 6100 3504
rect 6156 3496 6164 3504
rect 6172 3496 6180 3504
rect 6220 3496 6228 3504
rect 6252 3496 6260 3504
rect 6300 3496 6308 3504
rect 6364 3496 6372 3504
rect 6380 3496 6388 3504
rect 6396 3496 6404 3504
rect 6476 3496 6484 3504
rect 6524 3496 6532 3504
rect 6588 3496 6596 3504
rect 6604 3496 6612 3504
rect 6620 3496 6628 3504
rect 6668 3496 6676 3504
rect 6684 3496 6692 3504
rect 2172 3476 2180 3484
rect 2204 3476 2212 3484
rect 2284 3476 2292 3484
rect 2524 3476 2532 3484
rect 2620 3476 2628 3484
rect 2700 3476 2708 3484
rect 2796 3476 2804 3484
rect 2844 3476 2852 3484
rect 2988 3476 2996 3484
rect 3084 3476 3092 3484
rect 3324 3476 3332 3484
rect 3516 3476 3524 3484
rect 3580 3476 3588 3484
rect 3596 3476 3604 3484
rect 3660 3476 3668 3484
rect 3676 3476 3684 3484
rect 1932 3456 1940 3464
rect 2012 3456 2020 3464
rect 2092 3456 2100 3464
rect 2108 3456 2116 3464
rect 2220 3456 2228 3464
rect 2268 3456 2276 3464
rect 2460 3456 2468 3464
rect 3404 3456 3412 3464
rect 3740 3456 3748 3464
rect 3756 3456 3764 3464
rect 3820 3456 3828 3464
rect 3884 3476 3892 3484
rect 4540 3476 4548 3484
rect 4668 3476 4676 3484
rect 4876 3476 4884 3484
rect 4956 3476 4964 3484
rect 5116 3476 5124 3484
rect 5324 3476 5332 3484
rect 5404 3476 5412 3484
rect 5452 3476 5460 3484
rect 5628 3476 5636 3484
rect 5676 3476 5684 3484
rect 5708 3476 5716 3484
rect 4428 3456 4436 3464
rect 5036 3456 5044 3464
rect 5244 3456 5252 3464
rect 5356 3456 5364 3464
rect 5756 3456 5764 3464
rect 5804 3476 5812 3484
rect 5900 3476 5908 3484
rect 6348 3476 6356 3484
rect 6412 3476 6420 3484
rect 6428 3476 6436 3484
rect 6476 3476 6484 3484
rect 6524 3476 6532 3484
rect 6572 3476 6580 3484
rect 6700 3476 6708 3484
rect 6748 3476 6756 3484
rect 6876 3496 6884 3504
rect 6924 3496 6932 3504
rect 7052 3496 7060 3504
rect 7084 3496 7092 3504
rect 7132 3496 7140 3504
rect 7036 3476 7044 3484
rect 7068 3476 7076 3484
rect 7276 3496 7284 3504
rect 7356 3496 7364 3504
rect 6492 3456 6500 3464
rect 6796 3456 6804 3464
rect 7004 3456 7012 3464
rect 7212 3456 7220 3464
rect 7260 3476 7268 3484
rect 7308 3476 7316 3484
rect 7388 3456 7396 3464
rect 124 3436 132 3444
rect 380 3436 388 3444
rect 460 3436 468 3444
rect 604 3436 612 3444
rect 988 3436 996 3444
rect 1116 3436 1124 3444
rect 1244 3436 1252 3444
rect 1500 3436 1508 3444
rect 1564 3436 1572 3444
rect 1708 3436 1716 3444
rect 1820 3436 1828 3444
rect 1996 3436 2004 3444
rect 2076 3436 2084 3444
rect 2236 3436 2244 3444
rect 2412 3436 2420 3444
rect 2556 3436 2564 3444
rect 2828 3436 2836 3444
rect 3292 3436 3300 3444
rect 3532 3436 3540 3444
rect 3612 3436 3620 3444
rect 4764 3436 4772 3444
rect 4892 3436 4900 3444
rect 5308 3436 5316 3444
rect 5788 3436 5796 3444
rect 6140 3436 6148 3444
rect 6188 3436 6196 3444
rect 6284 3436 6292 3444
rect 6812 3436 6820 3444
rect 7116 3436 7124 3444
rect 7244 3436 7252 3444
rect 556 3416 564 3424
rect 764 3416 772 3424
rect 924 3416 932 3424
rect 940 3416 948 3424
rect 1372 3416 1380 3424
rect 2108 3416 2116 3424
rect 2460 3416 2468 3424
rect 2915 3406 2923 3414
rect 2925 3406 2933 3414
rect 2935 3406 2943 3414
rect 2945 3406 2953 3414
rect 2955 3406 2963 3414
rect 2965 3406 2973 3414
rect 5923 3406 5931 3414
rect 5933 3406 5941 3414
rect 5943 3406 5951 3414
rect 5953 3406 5961 3414
rect 5963 3406 5971 3414
rect 5973 3406 5981 3414
rect 588 3396 596 3404
rect 844 3396 852 3404
rect 1164 3396 1172 3404
rect 1228 3396 1236 3404
rect 108 3376 116 3384
rect 908 3376 916 3384
rect 1212 3376 1220 3384
rect 1436 3376 1444 3384
rect 1676 3376 1684 3384
rect 2732 3376 2740 3384
rect 12 3356 20 3364
rect 76 3356 84 3364
rect 204 3356 212 3364
rect 252 3356 260 3364
rect 444 3356 452 3364
rect 588 3356 596 3364
rect 700 3356 708 3364
rect 844 3356 852 3364
rect 940 3356 948 3364
rect 972 3356 980 3364
rect 1020 3356 1028 3364
rect 1164 3356 1172 3364
rect 1180 3356 1188 3364
rect 1228 3356 1236 3364
rect 1548 3356 1556 3364
rect 1580 3356 1588 3364
rect 1868 3356 1876 3364
rect 140 3336 148 3344
rect 268 3336 276 3344
rect 300 3336 308 3344
rect 444 3336 452 3344
rect 476 3332 484 3340
rect 652 3336 660 3344
rect 684 3336 692 3344
rect 748 3336 756 3344
rect 860 3336 868 3344
rect 1068 3336 1076 3344
rect 1404 3332 1412 3340
rect 1420 3336 1428 3344
rect 1532 3336 1540 3344
rect 1692 3336 1700 3344
rect 2076 3356 2084 3364
rect 2252 3356 2260 3364
rect 2556 3356 2564 3364
rect 3148 3376 3156 3384
rect 3692 3376 3700 3384
rect 4556 3376 4564 3384
rect 5036 3376 5044 3384
rect 5196 3376 5204 3384
rect 5580 3376 5588 3384
rect 5660 3376 5668 3384
rect 6316 3376 6324 3384
rect 6364 3376 6372 3384
rect 6396 3376 6404 3384
rect 6796 3376 6804 3384
rect 6988 3376 6996 3384
rect 7180 3376 7188 3384
rect 3084 3356 3092 3364
rect 3676 3356 3684 3364
rect 4428 3356 4436 3364
rect 4588 3356 4596 3364
rect 4652 3356 4660 3364
rect 4860 3356 4868 3364
rect 5228 3356 5236 3364
rect 6172 3356 6180 3364
rect 6300 3356 6308 3364
rect 6380 3356 6388 3364
rect 1964 3332 1972 3340
rect 1980 3336 1988 3344
rect 1996 3336 2004 3344
rect 2140 3336 2148 3344
rect 2220 3336 2228 3344
rect 2284 3336 2292 3344
rect 2396 3336 2404 3344
rect 2412 3336 2420 3344
rect 2508 3336 2516 3344
rect 2572 3336 2580 3344
rect 2588 3332 2596 3340
rect 3164 3336 3172 3344
rect 3212 3336 3220 3344
rect 3596 3336 3604 3344
rect 3852 3336 3860 3344
rect 4268 3336 4276 3344
rect 4300 3336 4308 3344
rect 4380 3336 4388 3344
rect 4508 3336 4516 3344
rect 4572 3336 4580 3344
rect 4636 3336 4644 3344
rect 4700 3336 4708 3344
rect 4748 3336 4756 3344
rect 4828 3336 4836 3344
rect 4908 3336 4916 3344
rect 4988 3336 4996 3344
rect 5084 3336 5092 3344
rect 5324 3336 5332 3344
rect 5436 3336 5444 3344
rect 5516 3336 5524 3344
rect 5628 3336 5636 3344
rect 5644 3336 5652 3344
rect 5708 3336 5716 3344
rect 5964 3336 5972 3344
rect 5980 3336 5988 3344
rect 6044 3336 6052 3344
rect 6156 3336 6164 3344
rect 6284 3336 6292 3344
rect 6556 3336 6564 3344
rect 6716 3336 6724 3344
rect 6780 3336 6788 3344
rect 156 3316 164 3324
rect 124 3296 132 3304
rect 316 3316 324 3324
rect 412 3316 420 3324
rect 540 3316 548 3324
rect 636 3316 644 3324
rect 668 3316 676 3324
rect 748 3316 756 3324
rect 764 3316 772 3324
rect 796 3316 804 3324
rect 860 3316 868 3324
rect 908 3316 916 3324
rect 1004 3316 1012 3324
rect 1020 3316 1028 3324
rect 1068 3316 1076 3324
rect 1084 3316 1092 3324
rect 1116 3316 1124 3324
rect 1276 3316 1284 3324
rect 1340 3316 1348 3324
rect 1612 3316 1620 3324
rect 204 3296 212 3304
rect 524 3296 532 3304
rect 764 3296 772 3304
rect 1084 3296 1092 3304
rect 1292 3296 1300 3304
rect 1356 3296 1364 3304
rect 1644 3296 1652 3304
rect 1724 3316 1732 3324
rect 1804 3316 1812 3324
rect 1836 3316 1844 3324
rect 2028 3316 2036 3324
rect 2044 3316 2052 3324
rect 2076 3316 2084 3324
rect 2124 3316 2132 3324
rect 2284 3316 2292 3324
rect 2380 3316 2388 3324
rect 2460 3316 2468 3324
rect 2524 3316 2532 3324
rect 2636 3316 2644 3324
rect 2684 3316 2692 3324
rect 2764 3316 2772 3324
rect 2780 3316 2788 3324
rect 2908 3316 2916 3324
rect 2940 3316 2948 3324
rect 3116 3316 3124 3324
rect 3180 3316 3188 3324
rect 3276 3316 3284 3324
rect 3292 3316 3300 3324
rect 3404 3316 3412 3324
rect 3452 3316 3460 3324
rect 3484 3316 3492 3324
rect 3500 3316 3508 3324
rect 3548 3316 3556 3324
rect 3564 3316 3572 3324
rect 3580 3316 3588 3324
rect 3644 3316 3652 3324
rect 3804 3316 3812 3324
rect 3900 3316 3908 3324
rect 3948 3316 3956 3324
rect 3964 3316 3972 3324
rect 3996 3316 4004 3324
rect 4044 3316 4052 3324
rect 4060 3316 4068 3324
rect 4140 3316 4148 3324
rect 4188 3316 4196 3324
rect 4284 3316 4292 3324
rect 1708 3296 1716 3304
rect 1820 3296 1828 3304
rect 4364 3316 4372 3324
rect 4380 3316 4388 3324
rect 4556 3316 4564 3324
rect 4332 3296 4340 3304
rect 4620 3316 4628 3324
rect 4684 3316 4692 3324
rect 4764 3316 4772 3324
rect 4780 3316 4788 3324
rect 4812 3316 4820 3324
rect 4828 3316 4836 3324
rect 4908 3316 4916 3324
rect 4940 3316 4948 3324
rect 4972 3316 4980 3324
rect 5004 3316 5012 3324
rect 5020 3316 5028 3324
rect 5116 3316 5124 3324
rect 5164 3316 5172 3324
rect 5180 3316 5188 3324
rect 5308 3316 5316 3324
rect 5404 3316 5412 3324
rect 5420 3316 5428 3324
rect 5532 3316 5540 3324
rect 5612 3316 5620 3324
rect 5660 3316 5668 3324
rect 5692 3316 5700 3324
rect 5724 3316 5732 3324
rect 5740 3316 5748 3324
rect 5772 3316 5780 3324
rect 5788 3316 5796 3324
rect 5820 3316 5828 3324
rect 5836 3316 5844 3324
rect 5884 3316 5892 3324
rect 5996 3316 6004 3324
rect 6028 3316 6036 3324
rect 6060 3316 6068 3324
rect 6076 3316 6084 3324
rect 6124 3316 6132 3324
rect 6172 3316 6180 3324
rect 6204 3316 6212 3324
rect 6268 3316 6276 3324
rect 6332 3316 6340 3324
rect 6348 3316 6356 3324
rect 6524 3318 6532 3326
rect 6588 3316 6596 3324
rect 6604 3316 6612 3324
rect 6668 3316 6676 3324
rect 6764 3316 6772 3324
rect 6876 3316 6884 3324
rect 6908 3316 6916 3324
rect 7052 3316 7060 3324
rect 7116 3318 7124 3326
rect 7244 3316 7252 3324
rect 7260 3316 7268 3324
rect 4732 3296 4740 3304
rect 4892 3296 4900 3304
rect 5388 3296 5396 3304
rect 5580 3296 5588 3304
rect 6236 3296 6244 3304
rect 6684 3296 6692 3304
rect 6764 3296 6772 3304
rect 524 3276 532 3284
rect 588 3276 596 3284
rect 1260 3276 1268 3284
rect 1324 3276 1332 3284
rect 1356 3276 1364 3284
rect 1740 3276 1748 3284
rect 1788 3276 1796 3284
rect 2044 3276 2052 3284
rect 3628 3276 3636 3284
rect 4012 3276 4020 3284
rect 4252 3276 4260 3284
rect 4828 3276 4836 3284
rect 4972 3276 4980 3284
rect 4716 3256 4724 3264
rect 5500 3256 5508 3264
rect 28 3236 36 3244
rect 60 3236 68 3244
rect 156 3236 164 3244
rect 364 3236 372 3244
rect 508 3236 516 3244
rect 732 3236 740 3244
rect 1004 3236 1012 3244
rect 1196 3236 1204 3244
rect 1244 3236 1252 3244
rect 1340 3236 1348 3244
rect 1756 3236 1764 3244
rect 1804 3236 1812 3244
rect 1916 3236 1924 3244
rect 2156 3236 2164 3244
rect 2524 3236 2532 3244
rect 2620 3236 2628 3244
rect 2668 3236 2676 3244
rect 2716 3236 2724 3244
rect 2812 3236 2820 3244
rect 3372 3236 3380 3244
rect 3436 3236 3444 3244
rect 3516 3236 3524 3244
rect 3916 3236 3924 3244
rect 5564 3236 5572 3244
rect 5996 3236 6004 3244
rect 6092 3236 6100 3244
rect 6620 3236 6628 3244
rect 1411 3206 1419 3214
rect 1421 3206 1429 3214
rect 1431 3206 1439 3214
rect 1441 3206 1449 3214
rect 1451 3206 1459 3214
rect 1461 3206 1469 3214
rect 4419 3206 4427 3214
rect 4429 3206 4437 3214
rect 4439 3206 4447 3214
rect 4449 3206 4457 3214
rect 4459 3206 4467 3214
rect 4469 3206 4477 3214
rect 28 3176 36 3184
rect 3260 3176 3268 3184
rect 4124 3176 4132 3184
rect 4556 3176 4564 3184
rect 4652 3176 4660 3184
rect 5164 3176 5172 3184
rect 5548 3176 5556 3184
rect 5628 3176 5636 3184
rect 5820 3176 5828 3184
rect 6028 3176 6036 3184
rect 6076 3176 6084 3184
rect 6188 3176 6196 3184
rect 6700 3176 6708 3184
rect 6716 3176 6724 3184
rect 6780 3176 6788 3184
rect 620 3156 628 3164
rect 476 3136 484 3144
rect 540 3136 548 3144
rect 668 3136 676 3144
rect 764 3136 772 3144
rect 1084 3136 1092 3144
rect 1148 3156 1156 3164
rect 1932 3156 1940 3164
rect 4716 3156 4724 3164
rect 28 3096 36 3104
rect 76 3116 84 3124
rect 444 3116 452 3124
rect 508 3116 516 3124
rect 636 3116 644 3124
rect 700 3116 708 3124
rect 732 3116 740 3124
rect 796 3116 804 3124
rect 812 3116 820 3124
rect 892 3116 900 3124
rect 1052 3116 1060 3124
rect 1164 3136 1172 3144
rect 1212 3136 1220 3144
rect 1900 3136 1908 3144
rect 2044 3136 2052 3144
rect 3292 3136 3300 3144
rect 4044 3136 4052 3144
rect 4060 3136 4068 3144
rect 4444 3136 4452 3144
rect 5052 3136 5060 3144
rect 5516 3136 5524 3144
rect 6908 3136 6916 3144
rect 7180 3136 7188 3144
rect 1276 3116 1284 3124
rect 1324 3116 1332 3124
rect 1916 3116 1924 3124
rect 1980 3116 1988 3124
rect 2076 3116 2084 3124
rect 2092 3116 2100 3124
rect 2220 3116 2228 3124
rect 2380 3116 2388 3124
rect 2924 3116 2932 3124
rect 3532 3116 3540 3124
rect 3724 3116 3732 3124
rect 108 3096 116 3104
rect 124 3096 132 3104
rect 316 3096 324 3104
rect 348 3096 356 3104
rect 428 3096 436 3104
rect 460 3096 468 3104
rect 524 3096 532 3104
rect 588 3096 596 3104
rect 652 3096 660 3104
rect 780 3096 788 3104
rect 812 3096 820 3104
rect 940 3096 948 3104
rect 972 3096 980 3104
rect 12 3076 20 3084
rect 124 3076 132 3084
rect 156 3076 164 3084
rect 268 3076 276 3084
rect 332 3076 340 3084
rect 380 3076 388 3084
rect 396 3076 404 3084
rect 572 3076 580 3084
rect 700 3076 708 3084
rect 844 3076 852 3084
rect 860 3076 868 3084
rect 956 3076 964 3084
rect 1100 3096 1108 3104
rect 1148 3096 1156 3104
rect 1196 3096 1204 3104
rect 1260 3096 1268 3104
rect 1388 3096 1396 3104
rect 1516 3096 1524 3104
rect 1548 3096 1556 3104
rect 1772 3096 1780 3104
rect 1820 3096 1828 3104
rect 1852 3096 1860 3104
rect 1932 3096 1940 3104
rect 2060 3096 2068 3104
rect 2092 3096 2100 3104
rect 2140 3096 2148 3104
rect 2204 3096 2212 3104
rect 1212 3076 1220 3084
rect 1260 3076 1268 3084
rect 1276 3076 1284 3084
rect 1308 3076 1316 3084
rect 1356 3076 1364 3084
rect 1372 3076 1380 3084
rect 1500 3076 1508 3084
rect 1612 3076 1620 3084
rect 1708 3076 1716 3084
rect 1836 3076 1844 3084
rect 2012 3076 2020 3084
rect 2124 3076 2132 3084
rect 2156 3076 2164 3084
rect 2188 3076 2196 3084
rect 2300 3096 2308 3104
rect 2348 3096 2356 3104
rect 2380 3096 2388 3104
rect 2444 3096 2452 3104
rect 2604 3096 2612 3104
rect 2668 3096 2676 3104
rect 2700 3096 2708 3104
rect 2732 3096 2740 3104
rect 2764 3096 2772 3104
rect 2828 3096 2836 3104
rect 2892 3096 2900 3104
rect 2988 3096 2996 3104
rect 3132 3096 3140 3104
rect 3212 3096 3220 3104
rect 3324 3096 3332 3104
rect 3388 3094 3396 3102
rect 3468 3096 3476 3104
rect 3516 3096 3524 3104
rect 3564 3096 3572 3104
rect 3612 3096 3620 3104
rect 3660 3096 3668 3104
rect 3676 3096 3684 3104
rect 3772 3096 3780 3104
rect 3836 3096 3844 3104
rect 3852 3096 3860 3104
rect 3900 3096 3908 3104
rect 3948 3096 3956 3104
rect 3996 3096 4004 3104
rect 4012 3096 4020 3104
rect 4092 3096 4100 3104
rect 4172 3096 4180 3104
rect 4220 3116 4228 3124
rect 4316 3094 4324 3102
rect 4588 3096 4596 3104
rect 4604 3096 4612 3104
rect 4636 3096 4644 3104
rect 4684 3096 4692 3104
rect 4700 3096 4708 3104
rect 4748 3096 4756 3104
rect 4796 3096 4804 3104
rect 4972 3096 4980 3104
rect 5020 3116 5028 3124
rect 6252 3116 6260 3124
rect 5100 3096 5108 3104
rect 5148 3096 5156 3104
rect 5260 3096 5268 3104
rect 5356 3096 5364 3104
rect 5404 3096 5412 3104
rect 5452 3096 5460 3104
rect 5468 3096 5476 3104
rect 5612 3096 5620 3104
rect 5724 3096 5732 3104
rect 5852 3096 5860 3104
rect 5868 3096 5876 3104
rect 5980 3096 5988 3104
rect 5996 3096 6004 3104
rect 6028 3096 6036 3104
rect 6108 3096 6116 3104
rect 6156 3096 6164 3104
rect 6572 3116 6580 3124
rect 6620 3116 6628 3124
rect 6844 3116 6852 3124
rect 7164 3116 7172 3124
rect 6284 3096 6292 3104
rect 6300 3096 6308 3104
rect 6444 3096 6452 3104
rect 6524 3096 6532 3104
rect 6636 3096 6644 3104
rect 6668 3096 6676 3104
rect 6748 3096 6756 3104
rect 6812 3096 6820 3104
rect 6940 3096 6948 3104
rect 7036 3096 7044 3104
rect 2316 3076 2324 3084
rect 2332 3076 2340 3084
rect 2492 3076 2500 3084
rect 2588 3076 2596 3084
rect 2620 3076 2628 3084
rect 156 3056 164 3064
rect 780 3056 788 3064
rect 908 3056 916 3064
rect 1196 3056 1204 3064
rect 1596 3056 1604 3064
rect 1724 3056 1732 3064
rect 1756 3056 1764 3064
rect 1772 3056 1780 3064
rect 1980 3056 1988 3064
rect 2204 3056 2212 3064
rect 236 3036 244 3044
rect 284 3036 292 3044
rect 460 3036 468 3044
rect 524 3036 532 3044
rect 732 3036 740 3044
rect 844 3036 852 3044
rect 876 3036 884 3044
rect 924 3036 932 3044
rect 1052 3036 1060 3044
rect 1260 3036 1268 3044
rect 1340 3036 1348 3044
rect 1484 3036 1492 3044
rect 1548 3036 1556 3044
rect 1660 3036 1668 3044
rect 2012 3036 2020 3044
rect 2060 3036 2068 3044
rect 2124 3036 2132 3044
rect 2172 3036 2180 3044
rect 2220 3036 2228 3044
rect 2476 3056 2484 3064
rect 2652 3076 2660 3084
rect 2716 3076 2724 3084
rect 2892 3076 2900 3084
rect 2924 3076 2932 3084
rect 3068 3076 3076 3084
rect 3180 3076 3188 3084
rect 3452 3076 3460 3084
rect 3484 3076 3492 3084
rect 3580 3076 3588 3084
rect 3692 3076 3700 3084
rect 3740 3076 3748 3084
rect 3788 3076 3796 3084
rect 2796 3056 2804 3064
rect 2828 3056 2836 3064
rect 2972 3056 2980 3064
rect 3196 3056 3204 3064
rect 3804 3056 3812 3064
rect 3884 3056 3892 3064
rect 3932 3076 3940 3084
rect 3948 3076 3956 3084
rect 4140 3076 4148 3084
rect 4156 3076 4164 3084
rect 4220 3076 4228 3084
rect 4252 3076 4260 3084
rect 4348 3076 4356 3084
rect 4940 3076 4948 3084
rect 4956 3076 4964 3084
rect 5052 3076 5060 3084
rect 5324 3076 5332 3084
rect 5372 3076 5380 3084
rect 5468 3076 5476 3084
rect 5564 3076 5572 3084
rect 5596 3076 5604 3084
rect 5788 3076 5796 3084
rect 6060 3076 6068 3084
rect 6172 3076 6180 3084
rect 6220 3076 6228 3084
rect 6316 3076 6324 3084
rect 6588 3076 6596 3084
rect 6604 3076 6612 3084
rect 6652 3076 6660 3084
rect 6764 3076 6772 3084
rect 6828 3076 6836 3084
rect 6876 3076 6884 3084
rect 7116 3096 7124 3104
rect 7244 3096 7252 3104
rect 7292 3096 7300 3104
rect 7132 3076 7140 3084
rect 7292 3076 7300 3084
rect 5420 3056 5428 3064
rect 5516 3056 5524 3064
rect 5580 3056 5588 3064
rect 5980 3056 5988 3064
rect 6012 3056 6020 3064
rect 6060 3056 6068 3064
rect 6460 3056 6468 3064
rect 6892 3056 6900 3064
rect 6940 3056 6948 3064
rect 6988 3056 6996 3064
rect 7052 3056 7060 3064
rect 7068 3056 7076 3064
rect 7100 3056 7108 3064
rect 7164 3056 7172 3064
rect 2460 3036 2468 3044
rect 2556 3036 2564 3044
rect 2732 3036 2740 3044
rect 3116 3036 3124 3044
rect 3244 3036 3252 3044
rect 3628 3036 3636 3044
rect 3820 3036 3828 3044
rect 4764 3036 4772 3044
rect 4828 3036 4836 3044
rect 5004 3036 5012 3044
rect 5116 3036 5124 3044
rect 6124 3036 6132 3044
rect 6332 3036 6340 3044
rect 6556 3036 6564 3044
rect 6700 3036 6708 3044
rect 6716 3036 6724 3044
rect 6780 3036 6788 3044
rect 6844 3036 6852 3044
rect 6956 3036 6964 3044
rect 1596 3016 1604 3024
rect 2915 3006 2923 3014
rect 2925 3006 2933 3014
rect 2935 3006 2943 3014
rect 2945 3006 2953 3014
rect 2955 3006 2963 3014
rect 2965 3006 2973 3014
rect 5923 3006 5931 3014
rect 5933 3006 5941 3014
rect 5943 3006 5951 3014
rect 5953 3006 5961 3014
rect 5963 3006 5971 3014
rect 5973 3006 5981 3014
rect 2556 2996 2564 3004
rect 1036 2976 1044 2984
rect 1292 2976 1300 2984
rect 1564 2976 1572 2984
rect 1676 2976 1684 2984
rect 1692 2976 1700 2984
rect 2044 2976 2052 2984
rect 2060 2976 2068 2984
rect 2444 2976 2452 2984
rect 2572 2976 2580 2984
rect 3260 2976 3268 2984
rect 3500 2976 3508 2984
rect 3788 2976 3796 2984
rect 5244 2976 5252 2984
rect 5436 2976 5444 2984
rect 6156 2976 6164 2984
rect 6668 2976 6676 2984
rect 6860 2976 6868 2984
rect 6908 2976 6916 2984
rect 7100 2976 7108 2984
rect 7164 2976 7172 2984
rect 7180 2976 7188 2984
rect 12 2956 20 2964
rect 44 2956 52 2964
rect 76 2956 84 2964
rect 172 2956 180 2964
rect 220 2956 228 2964
rect 124 2936 132 2944
rect 972 2956 980 2964
rect 1180 2956 1188 2964
rect 1228 2956 1236 2964
rect 1500 2956 1508 2964
rect 1516 2956 1524 2964
rect 2204 2956 2212 2964
rect 2380 2956 2388 2964
rect 2556 2956 2564 2964
rect 2860 2956 2868 2964
rect 3612 2956 3620 2964
rect 3676 2956 3684 2964
rect 5148 2956 5156 2964
rect 5772 2956 5780 2964
rect 6348 2956 6356 2964
rect 6972 2956 6980 2964
rect 7036 2956 7044 2964
rect 7116 2956 7124 2964
rect 7276 2956 7284 2964
rect 412 2936 420 2944
rect 428 2932 436 2940
rect 28 2916 36 2924
rect 92 2916 100 2924
rect 140 2916 148 2924
rect 172 2916 180 2924
rect 268 2916 276 2924
rect 300 2916 308 2924
rect 364 2916 372 2924
rect 508 2916 516 2924
rect 540 2916 548 2924
rect 604 2916 612 2924
rect 684 2916 692 2924
rect 732 2916 740 2924
rect 812 2916 820 2924
rect 988 2936 996 2944
rect 1036 2936 1044 2944
rect 860 2916 868 2924
rect 924 2916 932 2924
rect 972 2916 980 2924
rect 1036 2916 1044 2924
rect 1084 2916 1092 2924
rect 1244 2936 1252 2944
rect 1292 2936 1300 2944
rect 1132 2916 1140 2924
rect 1212 2916 1220 2924
rect 1228 2916 1236 2924
rect 1292 2916 1300 2924
rect 1340 2916 1348 2924
rect 1516 2936 1524 2944
rect 1564 2936 1572 2944
rect 1580 2936 1588 2944
rect 1692 2936 1700 2944
rect 1996 2936 2004 2944
rect 2060 2936 2068 2944
rect 2108 2936 2116 2944
rect 1388 2916 1396 2924
rect 1500 2916 1508 2924
rect 1564 2916 1572 2924
rect 1596 2916 1604 2924
rect 1644 2916 1652 2924
rect 1724 2916 1732 2924
rect 1772 2916 1780 2924
rect 1836 2916 1844 2924
rect 1884 2916 1892 2924
rect 1948 2916 1956 2924
rect 2012 2916 2020 2924
rect 2060 2916 2068 2924
rect 2396 2936 2404 2944
rect 2444 2936 2452 2944
rect 2460 2936 2468 2944
rect 2156 2916 2164 2924
rect 2204 2916 2212 2924
rect 2236 2916 2244 2924
rect 2284 2916 2292 2924
rect 2332 2916 2340 2924
rect 2380 2916 2388 2924
rect 2444 2916 2452 2924
rect 2460 2916 2468 2924
rect 2508 2916 2516 2924
rect 2652 2932 2660 2940
rect 2684 2936 2692 2944
rect 2780 2936 2788 2944
rect 2892 2936 2900 2944
rect 3212 2936 3220 2944
rect 3276 2936 3284 2944
rect 3292 2936 3300 2944
rect 3388 2936 3396 2944
rect 3420 2936 3428 2944
rect 3516 2936 3524 2944
rect 3564 2936 3572 2944
rect 3596 2936 3604 2944
rect 3644 2936 3652 2944
rect 3756 2936 3764 2944
rect 4220 2936 4228 2944
rect 4252 2936 4260 2944
rect 4636 2936 4644 2944
rect 4668 2936 4676 2944
rect 4700 2936 4708 2944
rect 4828 2936 4836 2944
rect 4924 2936 4932 2944
rect 4956 2936 4964 2944
rect 4988 2936 4996 2944
rect 5052 2936 5060 2944
rect 5164 2936 5172 2944
rect 5228 2936 5236 2944
rect 5452 2936 5460 2944
rect 5596 2936 5604 2944
rect 5628 2936 5636 2944
rect 5660 2936 5668 2944
rect 5724 2936 5732 2944
rect 5836 2936 5844 2944
rect 5980 2936 5988 2944
rect 6316 2936 6324 2944
rect 6380 2936 6388 2944
rect 6428 2936 6436 2944
rect 6492 2936 6500 2944
rect 6588 2936 6596 2944
rect 6652 2936 6660 2944
rect 6828 2936 6836 2944
rect 6892 2936 6900 2944
rect 7084 2936 7092 2944
rect 7228 2936 7236 2944
rect 7276 2936 7284 2944
rect 2780 2916 2788 2924
rect 2812 2916 2820 2924
rect 3180 2918 3188 2926
rect 3276 2916 3284 2924
rect 3340 2916 3348 2924
rect 3404 2916 3412 2924
rect 3436 2916 3444 2924
rect 3532 2916 3540 2924
rect 3580 2916 3588 2924
rect 3660 2916 3668 2924
rect 3708 2916 3716 2924
rect 3772 2916 3780 2924
rect 3900 2916 3908 2924
rect 4044 2916 4052 2924
rect 4092 2916 4100 2924
rect 4204 2916 4212 2924
rect 4268 2916 4276 2924
rect 4300 2916 4308 2924
rect 4348 2916 4356 2924
rect 4364 2916 4372 2924
rect 4508 2916 4516 2924
rect 4556 2916 4564 2924
rect 4652 2916 4660 2924
rect 4716 2916 4724 2924
rect 4844 2916 4852 2924
rect 348 2896 356 2904
rect 524 2896 532 2904
rect 540 2896 548 2904
rect 572 2896 580 2904
rect 716 2896 724 2904
rect 316 2876 324 2884
rect 380 2876 388 2884
rect 460 2876 468 2884
rect 492 2876 500 2884
rect 588 2876 596 2884
rect 700 2876 708 2884
rect 748 2876 756 2884
rect 796 2876 804 2884
rect 908 2896 916 2904
rect 988 2896 996 2904
rect 684 2856 692 2864
rect 876 2876 884 2884
rect 940 2876 948 2884
rect 1068 2876 1076 2884
rect 1148 2876 1156 2884
rect 1244 2876 1252 2884
rect 1324 2876 1332 2884
rect 1724 2896 1732 2904
rect 1740 2896 1748 2904
rect 1852 2896 1860 2904
rect 1868 2896 1876 2904
rect 1932 2896 1940 2904
rect 1996 2896 2004 2904
rect 2140 2896 2148 2904
rect 2300 2896 2308 2904
rect 2316 2896 2324 2904
rect 2476 2896 2484 2904
rect 2572 2896 2580 2904
rect 2796 2896 2804 2904
rect 3244 2896 3252 2904
rect 3340 2896 3348 2904
rect 3468 2896 3476 2904
rect 3548 2896 3556 2904
rect 3612 2896 3620 2904
rect 4684 2896 4692 2904
rect 4716 2896 4724 2904
rect 4988 2896 4996 2904
rect 5036 2916 5044 2924
rect 5100 2916 5108 2924
rect 5116 2916 5124 2924
rect 5212 2916 5220 2924
rect 5324 2916 5332 2924
rect 5356 2916 5364 2924
rect 5564 2918 5572 2926
rect 5660 2896 5668 2904
rect 5708 2916 5716 2924
rect 5740 2916 5748 2924
rect 5820 2916 5828 2924
rect 5852 2916 5860 2924
rect 6092 2916 6100 2924
rect 6108 2916 6116 2924
rect 6284 2918 6292 2926
rect 6396 2916 6404 2924
rect 6428 2896 6436 2904
rect 6476 2916 6484 2924
rect 6508 2916 6516 2924
rect 6636 2916 6644 2924
rect 6748 2916 6756 2924
rect 6940 2916 6948 2924
rect 6972 2916 6980 2924
rect 7116 2916 7124 2924
rect 7212 2916 7220 2924
rect 7244 2916 7252 2924
rect 7308 2916 7316 2924
rect 7324 2916 7332 2924
rect 7340 2916 7348 2924
rect 6556 2896 6564 2904
rect 6636 2896 6644 2904
rect 6860 2896 6868 2904
rect 7052 2896 7060 2904
rect 1404 2876 1412 2884
rect 1772 2876 1780 2884
rect 1820 2876 1828 2884
rect 1836 2876 1844 2884
rect 1964 2876 1972 2884
rect 2108 2876 2116 2884
rect 2172 2876 2180 2884
rect 2268 2876 2276 2884
rect 2348 2876 2356 2884
rect 2828 2876 2836 2884
rect 3820 2876 3828 2884
rect 4332 2876 4340 2884
rect 4748 2876 4756 2884
rect 4956 2876 4964 2884
rect 5180 2876 5188 2884
rect 5788 2876 5796 2884
rect 5996 2876 6004 2884
rect 7084 2876 7092 2884
rect 7228 2876 7236 2884
rect 7404 2876 7412 2884
rect 2236 2856 2244 2864
rect 2396 2856 2404 2864
rect 300 2836 308 2844
rect 364 2836 372 2844
rect 508 2836 516 2844
rect 604 2836 612 2844
rect 732 2836 740 2844
rect 860 2836 868 2844
rect 924 2836 932 2844
rect 1052 2836 1060 2844
rect 1388 2836 1396 2844
rect 1628 2836 1636 2844
rect 1788 2836 1796 2844
rect 1836 2836 1844 2844
rect 1916 2836 1924 2844
rect 2284 2836 2292 2844
rect 2332 2836 2340 2844
rect 2956 2836 2964 2844
rect 3036 2836 3044 2844
rect 3724 2836 3732 2844
rect 4156 2836 4164 2844
rect 4620 2836 4628 2844
rect 5068 2836 5076 2844
rect 5820 2836 5828 2844
rect 6060 2836 6068 2844
rect 6124 2836 6132 2844
rect 6380 2836 6388 2844
rect 6540 2836 6548 2844
rect 7164 2836 7172 2844
rect 1411 2806 1419 2814
rect 1421 2806 1429 2814
rect 1431 2806 1439 2814
rect 1441 2806 1449 2814
rect 1451 2806 1459 2814
rect 1461 2806 1469 2814
rect 4419 2806 4427 2814
rect 4429 2806 4437 2814
rect 4439 2806 4447 2814
rect 4449 2806 4457 2814
rect 4459 2806 4467 2814
rect 4469 2806 4477 2814
rect 156 2776 164 2784
rect 428 2776 436 2784
rect 524 2776 532 2784
rect 716 2776 724 2784
rect 908 2776 916 2784
rect 1196 2776 1204 2784
rect 1372 2776 1380 2784
rect 1532 2776 1540 2784
rect 1692 2776 1700 2784
rect 2124 2776 2132 2784
rect 2252 2776 2260 2784
rect 3500 2776 3508 2784
rect 4316 2776 4324 2784
rect 4508 2776 4516 2784
rect 5244 2776 5252 2784
rect 5420 2776 5428 2784
rect 5580 2776 5588 2784
rect 1004 2756 1012 2764
rect 1324 2756 1332 2764
rect 268 2736 276 2744
rect 300 2736 308 2744
rect 396 2736 404 2744
rect 460 2736 468 2744
rect 508 2736 516 2744
rect 572 2736 580 2744
rect 844 2736 852 2744
rect 1036 2736 1044 2744
rect 1148 2736 1156 2744
rect 1276 2736 1284 2744
rect 1372 2736 1380 2744
rect 1548 2736 1556 2744
rect 1612 2736 1620 2744
rect 1676 2736 1684 2744
rect 1820 2736 1828 2744
rect 1900 2736 1908 2744
rect 1932 2736 1940 2744
rect 1996 2736 2004 2744
rect 2076 2736 2084 2744
rect 2108 2736 2116 2744
rect 2172 2736 2180 2744
rect 2236 2736 2244 2744
rect 2508 2736 2516 2744
rect 3116 2736 3124 2744
rect 3996 2736 4004 2744
rect 4140 2736 4148 2744
rect 4252 2736 4260 2744
rect 6796 2736 6804 2744
rect 6828 2736 6836 2744
rect 124 2716 132 2724
rect 220 2716 228 2724
rect 236 2716 244 2724
rect 604 2716 612 2724
rect 620 2716 628 2724
rect 1068 2716 1076 2724
rect 1132 2716 1140 2724
rect 1260 2716 1268 2724
rect 1836 2716 1844 2724
rect 1964 2716 1972 2724
rect 2028 2716 2036 2724
rect 2204 2716 2212 2724
rect 2348 2716 2356 2724
rect 2540 2716 2548 2724
rect 3116 2716 3124 2724
rect 3164 2716 3172 2724
rect 3292 2716 3300 2724
rect 3420 2716 3428 2724
rect 4028 2716 4036 2724
rect 156 2696 164 2704
rect 220 2696 228 2704
rect 252 2696 260 2704
rect 332 2696 340 2704
rect 12 2676 20 2684
rect 108 2676 116 2684
rect 172 2676 180 2684
rect 188 2676 196 2684
rect 348 2676 356 2684
rect 380 2696 388 2704
rect 460 2696 468 2704
rect 380 2676 388 2684
rect 524 2696 532 2704
rect 588 2696 596 2704
rect 620 2696 628 2704
rect 700 2696 708 2704
rect 748 2696 756 2704
rect 796 2696 804 2704
rect 876 2696 884 2704
rect 892 2696 900 2704
rect 956 2696 964 2704
rect 1004 2696 1012 2704
rect 1052 2696 1060 2704
rect 1116 2696 1124 2704
rect 1180 2696 1188 2704
rect 1228 2696 1236 2704
rect 1260 2696 1268 2704
rect 1308 2696 1316 2704
rect 652 2676 660 2684
rect 908 2676 916 2684
rect 956 2676 964 2684
rect 1116 2676 1124 2684
rect 1372 2696 1380 2704
rect 1516 2696 1524 2704
rect 1564 2696 1572 2704
rect 1484 2676 1492 2684
rect 1628 2696 1636 2704
rect 1692 2696 1700 2704
rect 1740 2696 1748 2704
rect 1788 2696 1796 2704
rect 1820 2696 1828 2704
rect 1868 2696 1876 2704
rect 1948 2696 1956 2704
rect 1980 2696 1988 2704
rect 2012 2696 2020 2704
rect 2044 2696 2052 2704
rect 2124 2696 2132 2704
rect 1724 2676 1732 2684
rect 1852 2676 1860 2684
rect 2188 2696 2196 2704
rect 2252 2696 2260 2704
rect 2332 2696 2340 2704
rect 2364 2696 2372 2704
rect 2476 2696 2484 2704
rect 2524 2696 2532 2704
rect 2556 2696 2564 2704
rect 3100 2696 3108 2704
rect 3260 2696 3268 2704
rect 3356 2696 3364 2704
rect 3388 2696 3396 2704
rect 3484 2696 3492 2704
rect 3628 2694 3636 2702
rect 3724 2696 3732 2704
rect 3788 2696 3796 2704
rect 3868 2696 3876 2704
rect 4588 2716 4596 2724
rect 4780 2716 4788 2724
rect 4908 2716 4916 2724
rect 5212 2716 5220 2724
rect 5788 2716 5796 2724
rect 5820 2716 5828 2724
rect 6140 2716 6148 2724
rect 6172 2716 6180 2724
rect 6332 2716 6340 2724
rect 4092 2696 4100 2704
rect 4124 2696 4132 2704
rect 4172 2696 4180 2704
rect 4204 2696 4212 2704
rect 4220 2696 4228 2704
rect 4268 2696 4276 2704
rect 4284 2696 4292 2704
rect 4316 2696 4324 2704
rect 4348 2696 4356 2704
rect 4380 2696 4388 2704
rect 4540 2696 4548 2704
rect 4556 2696 4564 2704
rect 4588 2696 4596 2704
rect 4652 2696 4660 2704
rect 2380 2676 2388 2684
rect 2476 2676 2484 2684
rect 2604 2676 2612 2684
rect 2700 2676 2708 2684
rect 2716 2676 2724 2684
rect 2812 2676 2820 2684
rect 2828 2676 2836 2684
rect 3020 2676 3028 2684
rect 3132 2676 3140 2684
rect 3228 2676 3236 2684
rect 3244 2676 3252 2684
rect 3340 2676 3348 2684
rect 3372 2676 3380 2684
rect 3468 2676 3476 2684
rect 3660 2676 3668 2684
rect 3772 2676 3780 2684
rect 3820 2676 3828 2684
rect 3996 2676 4004 2684
rect 4044 2676 4052 2684
rect 4092 2676 4100 2684
rect 4300 2676 4308 2684
rect 4364 2676 4372 2684
rect 4524 2676 4532 2684
rect 4604 2676 4612 2684
rect 4652 2676 4660 2684
rect 4732 2696 4740 2704
rect 4748 2696 4756 2704
rect 4796 2696 4804 2704
rect 4828 2696 4836 2704
rect 4876 2696 4884 2704
rect 4892 2696 4900 2704
rect 4940 2696 4948 2704
rect 4972 2696 4980 2704
rect 4988 2696 4996 2704
rect 5052 2696 5060 2704
rect 5068 2696 5076 2704
rect 5084 2696 5092 2704
rect 5180 2696 5188 2704
rect 5244 2696 5252 2704
rect 5276 2696 5284 2704
rect 5308 2696 5316 2704
rect 5372 2696 5380 2704
rect 5388 2696 5396 2704
rect 5404 2696 5412 2704
rect 5452 2696 5460 2704
rect 5484 2696 5492 2704
rect 5500 2696 5508 2704
rect 5548 2696 5556 2704
rect 5708 2694 5716 2702
rect 5788 2696 5796 2704
rect 5900 2696 5908 2704
rect 6108 2696 6116 2704
rect 6140 2696 6148 2704
rect 6204 2696 6212 2704
rect 6236 2696 6244 2704
rect 6284 2696 6292 2704
rect 6460 2696 6468 2704
rect 6572 2696 6580 2704
rect 6604 2696 6612 2704
rect 6652 2696 6660 2704
rect 6668 2696 6676 2704
rect 6684 2696 6692 2704
rect 6780 2696 6788 2704
rect 6924 2694 6932 2702
rect 7100 2696 7108 2704
rect 7308 2694 7316 2702
rect 4796 2676 4804 2684
rect 4876 2676 4884 2684
rect 4972 2676 4980 2684
rect 5132 2676 5140 2684
rect 5164 2676 5172 2684
rect 5196 2676 5204 2684
rect 5260 2676 5268 2684
rect 5356 2676 5364 2684
rect 5676 2676 5684 2684
rect 5740 2676 5748 2684
rect 5772 2676 5780 2684
rect 5852 2676 5860 2684
rect 6092 2676 6100 2684
rect 6220 2676 6228 2684
rect 6268 2676 6276 2684
rect 6300 2676 6308 2684
rect 6508 2676 6516 2684
rect 6700 2676 6708 2684
rect 588 2656 596 2664
rect 668 2656 676 2664
rect 700 2656 708 2664
rect 764 2656 772 2664
rect 828 2656 836 2664
rect 892 2656 900 2664
rect 972 2656 980 2664
rect 1340 2656 1348 2664
rect 1628 2656 1636 2664
rect 1948 2656 1956 2664
rect 2284 2656 2292 2664
rect 2316 2656 2324 2664
rect 2556 2656 2564 2664
rect 3052 2656 3060 2664
rect 3692 2656 3700 2664
rect 4380 2656 4388 2664
rect 4412 2656 4420 2664
rect 4620 2656 4628 2664
rect 4764 2656 4772 2664
rect 4924 2656 4932 2664
rect 4972 2656 4980 2664
rect 5116 2656 5124 2664
rect 5276 2656 5284 2664
rect 6268 2656 6276 2664
rect 6332 2656 6340 2664
rect 6716 2656 6724 2664
rect 6956 2676 6964 2684
rect 7116 2676 7124 2684
rect 7292 2676 7300 2684
rect 6748 2656 6756 2664
rect 6780 2656 6788 2664
rect 6860 2656 6868 2664
rect 76 2636 84 2644
rect 188 2636 196 2644
rect 284 2636 292 2644
rect 652 2636 660 2644
rect 780 2636 788 2644
rect 812 2636 820 2644
rect 956 2636 964 2644
rect 1036 2636 1044 2644
rect 1292 2636 1300 2644
rect 1772 2636 1780 2644
rect 2188 2636 2196 2644
rect 2300 2636 2308 2644
rect 2412 2636 2420 2644
rect 2748 2636 2756 2644
rect 2876 2636 2884 2644
rect 3324 2636 3332 2644
rect 3452 2636 3460 2644
rect 3756 2636 3764 2644
rect 4636 2636 4644 2644
rect 4700 2636 4708 2644
rect 4828 2636 4836 2644
rect 5340 2636 5348 2644
rect 5516 2636 5524 2644
rect 6012 2636 6020 2644
rect 6348 2636 6356 2644
rect 6540 2636 6548 2644
rect 6620 2636 6628 2644
rect 6988 2636 6996 2644
rect 7180 2636 7188 2644
rect 828 2616 836 2624
rect 2915 2606 2923 2614
rect 2925 2606 2933 2614
rect 2935 2606 2943 2614
rect 2945 2606 2953 2614
rect 2955 2606 2963 2614
rect 2965 2606 2973 2614
rect 5923 2606 5931 2614
rect 5933 2606 5941 2614
rect 5943 2606 5951 2614
rect 5953 2606 5961 2614
rect 5963 2606 5971 2614
rect 5973 2606 5981 2614
rect 556 2596 564 2604
rect 588 2596 596 2604
rect 876 2596 884 2604
rect 1004 2596 1012 2604
rect 1260 2596 1268 2604
rect 1564 2596 1572 2604
rect 1692 2596 1700 2604
rect 396 2576 404 2584
rect 412 2576 420 2584
rect 508 2576 516 2584
rect 156 2556 164 2564
rect 556 2556 564 2564
rect 588 2556 596 2564
rect 764 2556 772 2564
rect 796 2556 804 2564
rect 876 2556 884 2564
rect 956 2556 964 2564
rect 1004 2556 1012 2564
rect 1020 2556 1028 2564
rect 1388 2576 1396 2584
rect 1484 2576 1492 2584
rect 1740 2576 1748 2584
rect 1900 2576 1908 2584
rect 2332 2576 2340 2584
rect 2492 2576 2500 2584
rect 2604 2576 2612 2584
rect 2684 2576 2692 2584
rect 2988 2576 2996 2584
rect 3100 2576 3108 2584
rect 3788 2576 3796 2584
rect 3980 2576 3988 2584
rect 4508 2576 4516 2584
rect 4524 2576 4532 2584
rect 4908 2576 4916 2584
rect 5244 2576 5252 2584
rect 5500 2576 5508 2584
rect 5548 2576 5556 2584
rect 6252 2576 6260 2584
rect 6796 2576 6804 2584
rect 7052 2576 7060 2584
rect 7100 2576 7108 2584
rect 1244 2556 1252 2564
rect 1260 2556 1268 2564
rect 1500 2556 1508 2564
rect 1564 2556 1572 2564
rect 1612 2556 1620 2564
rect 1692 2556 1700 2564
rect 1820 2556 1828 2564
rect 1884 2556 1892 2564
rect 2412 2556 2420 2564
rect 2668 2556 2676 2564
rect 3004 2556 3012 2564
rect 3580 2556 3588 2564
rect 3660 2556 3668 2564
rect 3996 2556 4004 2564
rect 4060 2556 4068 2564
rect 4108 2556 4116 2564
rect 5276 2556 5284 2564
rect 5676 2556 5684 2564
rect 6316 2556 6324 2564
rect 6508 2556 6516 2564
rect 6556 2556 6564 2564
rect 6988 2556 6996 2564
rect 7068 2556 7076 2564
rect 7084 2556 7092 2564
rect 44 2532 52 2540
rect 60 2536 68 2544
rect 156 2536 164 2544
rect 348 2536 356 2544
rect 604 2536 612 2544
rect 620 2536 628 2544
rect 652 2536 660 2544
rect 684 2536 692 2544
rect 812 2536 820 2544
rect 1052 2536 1060 2544
rect 1132 2536 1140 2544
rect 1212 2536 1220 2544
rect 1356 2536 1364 2544
rect 1388 2536 1396 2544
rect 1516 2536 1524 2544
rect 1900 2536 1908 2544
rect 12 2516 20 2524
rect 76 2516 84 2524
rect 124 2516 132 2524
rect 204 2516 212 2524
rect 236 2516 244 2524
rect 268 2516 276 2524
rect 300 2516 308 2524
rect 364 2516 372 2524
rect 444 2516 452 2524
rect 460 2516 468 2524
rect 556 2516 564 2524
rect 588 2516 596 2524
rect 636 2516 644 2524
rect 668 2516 676 2524
rect 732 2516 740 2524
rect 812 2516 820 2524
rect 828 2516 836 2524
rect 924 2516 932 2524
rect 956 2516 964 2524
rect 1052 2516 1060 2524
rect 1116 2516 1124 2524
rect 1148 2516 1156 2524
rect 1212 2516 1220 2524
rect 1292 2516 1300 2524
rect 92 2496 100 2504
rect 220 2496 228 2504
rect 284 2496 292 2504
rect 748 2496 756 2504
rect 828 2496 836 2504
rect 860 2496 868 2504
rect 1468 2516 1476 2524
rect 1612 2516 1620 2524
rect 1644 2516 1652 2524
rect 1708 2516 1716 2524
rect 1772 2516 1780 2524
rect 1852 2516 1860 2524
rect 1980 2516 1988 2524
rect 2028 2516 2036 2524
rect 2060 2516 2068 2524
rect 2124 2516 2132 2524
rect 2252 2536 2260 2544
rect 2380 2536 2388 2544
rect 2428 2536 2436 2544
rect 2524 2536 2532 2544
rect 2540 2536 2548 2544
rect 2636 2536 2644 2544
rect 2684 2536 2692 2544
rect 2780 2536 2788 2544
rect 2876 2536 2884 2544
rect 2188 2516 2196 2524
rect 2220 2516 2228 2524
rect 2300 2516 2308 2524
rect 2364 2516 2372 2524
rect 2700 2516 2708 2524
rect 2876 2516 2884 2524
rect 3036 2536 3044 2544
rect 3132 2536 3140 2544
rect 3308 2536 3316 2544
rect 3500 2536 3508 2544
rect 3820 2536 3828 2544
rect 4076 2536 4084 2544
rect 4396 2536 4404 2544
rect 4572 2536 4580 2544
rect 4588 2536 4596 2544
rect 4652 2536 4660 2544
rect 4764 2536 4772 2544
rect 4812 2536 4820 2544
rect 4828 2536 4836 2544
rect 4892 2536 4900 2544
rect 4956 2536 4964 2544
rect 5068 2536 5076 2544
rect 5100 2536 5108 2544
rect 5132 2536 5140 2544
rect 5436 2536 5444 2544
rect 5740 2536 5748 2544
rect 5772 2536 5780 2544
rect 5836 2536 5844 2544
rect 5932 2536 5940 2544
rect 6108 2536 6116 2544
rect 6140 2536 6148 2544
rect 6204 2536 6212 2544
rect 6236 2536 6244 2544
rect 6460 2536 6468 2544
rect 6620 2536 6628 2544
rect 6684 2536 6692 2544
rect 6956 2536 6964 2544
rect 7116 2536 7124 2544
rect 3276 2518 3284 2526
rect 3452 2516 3460 2524
rect 3580 2516 3588 2524
rect 3676 2516 3684 2524
rect 3708 2516 3716 2524
rect 3868 2516 3876 2524
rect 4028 2516 4036 2524
rect 4108 2516 4116 2524
rect 4156 2516 4164 2524
rect 4204 2516 4212 2524
rect 4220 2516 4228 2524
rect 4252 2516 4260 2524
rect 4268 2516 4276 2524
rect 4300 2516 4308 2524
rect 4316 2516 4324 2524
rect 4380 2516 4388 2524
rect 4412 2516 4420 2524
rect 4556 2516 4564 2524
rect 4604 2516 4612 2524
rect 4636 2516 4644 2524
rect 4668 2516 4676 2524
rect 4684 2516 4692 2524
rect 4732 2516 4740 2524
rect 4780 2516 4788 2524
rect 1356 2496 1364 2504
rect 1548 2496 1556 2504
rect 1756 2496 1764 2504
rect 1868 2496 1876 2504
rect 1916 2496 1924 2504
rect 2076 2496 2084 2504
rect 2204 2496 2212 2504
rect 2220 2496 2228 2504
rect 2316 2496 2324 2504
rect 2924 2496 2932 2504
rect 4332 2496 4340 2504
rect 4364 2496 4372 2504
rect 4524 2496 4532 2504
rect 4636 2496 4644 2504
rect 4844 2516 4852 2524
rect 4876 2516 4884 2524
rect 4940 2516 4948 2524
rect 4972 2516 4980 2524
rect 4988 2516 4996 2524
rect 5036 2516 5044 2524
rect 5052 2516 5060 2524
rect 5116 2516 5124 2524
rect 5148 2516 5156 2524
rect 5212 2516 5220 2524
rect 5228 2516 5236 2524
rect 5324 2516 5332 2524
rect 5340 2516 5348 2524
rect 5452 2516 5460 2524
rect 5532 2516 5540 2524
rect 5676 2518 5684 2526
rect 7180 2536 7188 2544
rect 7212 2536 7220 2544
rect 7276 2536 7284 2544
rect 7324 2536 7332 2544
rect 4876 2496 4884 2504
rect 4908 2496 4916 2504
rect 5180 2496 5188 2504
rect 5452 2496 5460 2504
rect 5484 2496 5492 2504
rect 5772 2496 5780 2504
rect 5884 2516 5892 2524
rect 5996 2516 6004 2524
rect 6140 2496 6148 2504
rect 6188 2516 6196 2524
rect 6220 2516 6228 2524
rect 6284 2516 6292 2524
rect 6332 2516 6340 2524
rect 6380 2516 6388 2524
rect 6444 2516 6452 2524
rect 6476 2516 6484 2524
rect 6524 2516 6532 2524
rect 6604 2516 6612 2524
rect 6620 2516 6628 2524
rect 6668 2516 6676 2524
rect 6700 2516 6708 2524
rect 6716 2516 6724 2524
rect 6780 2516 6788 2524
rect 6908 2516 6916 2524
rect 7020 2516 7028 2524
rect 7036 2516 7044 2524
rect 7132 2516 7140 2524
rect 7164 2516 7172 2524
rect 7228 2516 7236 2524
rect 7372 2516 7380 2524
rect 6380 2496 6388 2504
rect 6604 2496 6612 2504
rect 6636 2496 6644 2504
rect 6748 2496 6756 2504
rect 7196 2496 7204 2504
rect 7228 2496 7236 2504
rect 7324 2496 7332 2504
rect 7356 2496 7364 2504
rect 252 2476 260 2484
rect 316 2476 324 2484
rect 492 2476 500 2484
rect 716 2476 724 2484
rect 1788 2476 1796 2484
rect 1836 2476 1844 2484
rect 1996 2476 2004 2484
rect 2044 2476 2052 2484
rect 2108 2476 2116 2484
rect 2172 2476 2180 2484
rect 2284 2476 2292 2484
rect 2844 2476 2852 2484
rect 6108 2476 6116 2484
rect 6572 2476 6580 2484
rect 7020 2476 7028 2484
rect 7260 2476 7268 2484
rect 332 2436 340 2444
rect 412 2436 420 2444
rect 508 2436 516 2444
rect 732 2436 740 2444
rect 1532 2436 1540 2444
rect 1804 2436 1812 2444
rect 2012 2436 2020 2444
rect 2124 2436 2132 2444
rect 2188 2436 2196 2444
rect 2300 2436 2308 2444
rect 2396 2436 2404 2444
rect 3020 2436 3028 2444
rect 3148 2436 3156 2444
rect 3340 2436 3348 2444
rect 3532 2436 3540 2444
rect 3596 2436 3604 2444
rect 4124 2436 4132 2444
rect 4188 2436 4196 2444
rect 4700 2436 4708 2444
rect 5004 2436 5012 2444
rect 6412 2436 6420 2444
rect 6476 2436 6484 2444
rect 6524 2436 6532 2444
rect 6796 2436 6804 2444
rect 7292 2436 7300 2444
rect 1411 2406 1419 2414
rect 1421 2406 1429 2414
rect 1431 2406 1439 2414
rect 1441 2406 1449 2414
rect 1451 2406 1459 2414
rect 1461 2406 1469 2414
rect 4419 2406 4427 2414
rect 4429 2406 4437 2414
rect 4439 2406 4447 2414
rect 4449 2406 4457 2414
rect 4459 2406 4467 2414
rect 4469 2406 4477 2414
rect 604 2376 612 2384
rect 1052 2376 1060 2384
rect 1772 2376 1780 2384
rect 1852 2376 1860 2384
rect 1932 2376 1940 2384
rect 2236 2376 2244 2384
rect 2332 2376 2340 2384
rect 2508 2376 2516 2384
rect 2748 2376 2756 2384
rect 2988 2376 2996 2384
rect 3068 2376 3076 2384
rect 3116 2376 3124 2384
rect 3708 2376 3716 2384
rect 4204 2376 4212 2384
rect 4588 2376 4596 2384
rect 4716 2376 4724 2384
rect 5084 2376 5092 2384
rect 5196 2376 5204 2384
rect 6876 2376 6884 2384
rect 7308 2376 7316 2384
rect 4060 2356 4068 2364
rect 4924 2356 4932 2364
rect 5308 2356 5316 2364
rect 6092 2356 6100 2364
rect 364 2336 372 2344
rect 492 2336 500 2344
rect 556 2336 564 2344
rect 620 2336 628 2344
rect 956 2336 964 2344
rect 1180 2336 1188 2344
rect 2252 2336 2260 2344
rect 2316 2336 2324 2344
rect 2604 2336 2612 2344
rect 3132 2336 3140 2344
rect 4604 2336 4612 2344
rect 5164 2336 5172 2344
rect 5260 2336 5268 2344
rect 5612 2336 5620 2344
rect 6684 2336 6692 2344
rect 7068 2336 7076 2344
rect 44 2296 52 2304
rect 332 2316 340 2324
rect 396 2316 404 2324
rect 524 2316 532 2324
rect 844 2316 852 2324
rect 316 2296 324 2304
rect 348 2296 356 2304
rect 412 2296 420 2304
rect 60 2276 68 2284
rect 76 2276 84 2284
rect 92 2276 100 2284
rect 108 2276 116 2284
rect 140 2276 148 2284
rect 188 2276 196 2284
rect 220 2276 228 2284
rect 316 2276 324 2284
rect 396 2276 404 2284
rect 476 2296 484 2304
rect 556 2296 564 2304
rect 476 2276 484 2284
rect 572 2276 580 2284
rect 604 2296 612 2304
rect 652 2296 660 2304
rect 732 2296 740 2304
rect 748 2296 756 2304
rect 780 2296 788 2304
rect 844 2296 852 2304
rect 892 2316 900 2324
rect 988 2316 996 2324
rect 1084 2316 1092 2324
rect 1148 2316 1156 2324
rect 1324 2316 1332 2324
rect 1596 2316 1604 2324
rect 2156 2316 2164 2324
rect 2220 2316 2228 2324
rect 2284 2316 2292 2324
rect 2348 2316 2356 2324
rect 2556 2316 2564 2324
rect 3372 2316 3380 2324
rect 3564 2316 3572 2324
rect 4092 2316 4100 2324
rect 972 2296 980 2304
rect 1052 2296 1060 2304
rect 1100 2296 1108 2304
rect 1180 2296 1188 2304
rect 1292 2296 1300 2304
rect 1308 2296 1316 2304
rect 1388 2296 1396 2304
rect 1420 2296 1428 2304
rect 924 2276 932 2284
rect 972 2276 980 2284
rect 1404 2276 1412 2284
rect 1628 2296 1636 2304
rect 1692 2296 1700 2304
rect 1756 2296 1764 2304
rect 1804 2296 1812 2304
rect 1820 2296 1828 2304
rect 1868 2296 1876 2304
rect 1884 2296 1892 2304
rect 2012 2296 2020 2304
rect 2060 2296 2068 2304
rect 2204 2296 2212 2304
rect 2236 2296 2244 2304
rect 2300 2296 2308 2304
rect 2412 2296 2420 2304
rect 2444 2296 2452 2304
rect 2508 2296 2516 2304
rect 2588 2296 2596 2304
rect 2652 2296 2660 2304
rect 2844 2296 2852 2304
rect 3020 2296 3028 2304
rect 3036 2296 3044 2304
rect 3084 2296 3092 2304
rect 3260 2294 3268 2302
rect 3340 2296 3348 2304
rect 3372 2296 3380 2304
rect 3436 2296 3444 2304
rect 3452 2296 3460 2304
rect 3532 2296 3540 2304
rect 3628 2296 3636 2304
rect 3676 2296 3684 2304
rect 3868 2296 3876 2304
rect 3948 2296 3956 2304
rect 4092 2296 4100 2304
rect 4140 2316 4148 2324
rect 4636 2316 4644 2324
rect 4236 2296 4244 2304
rect 4300 2296 4308 2304
rect 4476 2296 4484 2304
rect 4956 2316 4964 2324
rect 5228 2316 5236 2324
rect 5548 2316 5556 2324
rect 5692 2316 5700 2324
rect 5932 2316 5940 2324
rect 7292 2316 7300 2324
rect 4684 2296 4692 2304
rect 4844 2294 4852 2302
rect 4908 2296 4916 2304
rect 5004 2296 5012 2304
rect 5020 2296 5028 2304
rect 5068 2296 5076 2304
rect 5116 2296 5124 2304
rect 5132 2296 5140 2304
rect 5260 2296 5268 2304
rect 5356 2296 5364 2304
rect 1708 2276 1716 2284
rect 1756 2276 1764 2284
rect 1964 2276 1972 2284
rect 2028 2276 2036 2284
rect 2076 2276 2084 2284
rect 12 2256 20 2264
rect 204 2256 212 2264
rect 748 2256 756 2264
rect 444 2236 452 2244
rect 684 2236 692 2244
rect 700 2236 708 2244
rect 1100 2256 1108 2264
rect 1132 2256 1140 2264
rect 1228 2256 1236 2264
rect 1244 2256 1252 2264
rect 1340 2256 1348 2264
rect 1532 2256 1540 2264
rect 1548 2256 1556 2264
rect 1580 2256 1588 2264
rect 1676 2256 1684 2264
rect 1900 2256 1908 2264
rect 1916 2256 1924 2264
rect 1948 2256 1956 2264
rect 2076 2256 2084 2264
rect 2380 2276 2388 2284
rect 2396 2276 2404 2284
rect 2604 2276 2612 2284
rect 2668 2276 2676 2284
rect 2780 2276 2788 2284
rect 2828 2276 2836 2284
rect 3292 2276 3300 2284
rect 3324 2276 3332 2284
rect 3420 2276 3428 2284
rect 3468 2276 3476 2284
rect 3516 2276 3524 2284
rect 3612 2276 3620 2284
rect 3820 2276 3828 2284
rect 4076 2276 4084 2284
rect 4172 2276 4180 2284
rect 4220 2276 4228 2284
rect 4252 2276 4260 2284
rect 4428 2276 4436 2284
rect 4524 2276 4532 2284
rect 4604 2276 4612 2284
rect 4636 2276 4644 2284
rect 4700 2276 4708 2284
rect 4844 2276 4852 2284
rect 4908 2276 4916 2284
rect 5052 2276 5060 2284
rect 5212 2276 5220 2284
rect 5292 2276 5300 2284
rect 5324 2276 5332 2284
rect 5388 2296 5396 2304
rect 5452 2296 5460 2304
rect 5500 2296 5508 2304
rect 5580 2296 5588 2304
rect 5612 2296 5620 2304
rect 5644 2296 5652 2304
rect 5724 2296 5732 2304
rect 5756 2296 5764 2304
rect 5804 2296 5812 2304
rect 5868 2296 5876 2304
rect 5900 2296 5908 2304
rect 6012 2296 6020 2304
rect 6060 2296 6068 2304
rect 6204 2296 6212 2304
rect 6284 2296 6292 2304
rect 6348 2296 6356 2304
rect 6396 2296 6404 2304
rect 6428 2296 6436 2304
rect 6444 2296 6452 2304
rect 6492 2296 6500 2304
rect 6508 2296 6516 2304
rect 6524 2296 6532 2304
rect 6604 2296 6612 2304
rect 6668 2296 6676 2304
rect 6748 2296 6756 2304
rect 6796 2296 6804 2304
rect 6956 2296 6964 2304
rect 7004 2294 7012 2302
rect 7132 2296 7140 2304
rect 7196 2294 7204 2302
rect 7356 2296 7364 2304
rect 5388 2276 5396 2284
rect 5484 2276 5492 2284
rect 5500 2276 5508 2284
rect 5628 2276 5636 2284
rect 5708 2276 5716 2284
rect 5740 2276 5748 2284
rect 5756 2276 5764 2284
rect 5820 2276 5828 2284
rect 5884 2276 5892 2284
rect 6044 2276 6052 2284
rect 6076 2276 6084 2284
rect 6252 2276 6260 2284
rect 6332 2276 6340 2284
rect 6652 2276 6660 2284
rect 6844 2276 6852 2284
rect 7260 2276 7268 2284
rect 7372 2276 7380 2284
rect 2172 2256 2180 2264
rect 2492 2256 2500 2264
rect 2540 2256 2548 2264
rect 2828 2256 2836 2264
rect 3500 2256 3508 2264
rect 3932 2256 3940 2264
rect 4396 2256 4404 2264
rect 4972 2256 4980 2264
rect 5340 2256 5348 2264
rect 5436 2256 5444 2264
rect 5644 2256 5652 2264
rect 5676 2256 5684 2264
rect 5836 2256 5844 2264
rect 6284 2256 6292 2264
rect 6316 2256 6324 2264
rect 6524 2256 6532 2264
rect 6556 2256 6564 2264
rect 6572 2256 6580 2264
rect 6636 2256 6644 2264
rect 7308 2256 7316 2264
rect 924 2236 932 2244
rect 1724 2236 1732 2244
rect 1852 2236 1860 2244
rect 2156 2236 2164 2244
rect 2188 2236 2196 2244
rect 2348 2236 2356 2244
rect 2412 2236 2420 2244
rect 2860 2236 2868 2244
rect 3484 2236 3492 2244
rect 3596 2236 3604 2244
rect 3836 2236 3844 2244
rect 4268 2236 4276 2244
rect 5084 2236 5092 2244
rect 5420 2236 5428 2244
rect 5804 2236 5812 2244
rect 5852 2236 5860 2244
rect 6460 2236 6468 2244
rect 7292 2236 7300 2244
rect 1228 2216 1236 2224
rect 1244 2216 1252 2224
rect 1340 2216 1348 2224
rect 1532 2216 1540 2224
rect 2915 2206 2923 2214
rect 2925 2206 2933 2214
rect 2935 2206 2943 2214
rect 2945 2206 2953 2214
rect 2955 2206 2963 2214
rect 2965 2206 2973 2214
rect 5923 2206 5931 2214
rect 5933 2206 5941 2214
rect 5943 2206 5951 2214
rect 5953 2206 5961 2214
rect 5963 2206 5971 2214
rect 5973 2206 5981 2214
rect 908 2196 916 2204
rect 1036 2196 1044 2204
rect 1180 2196 1188 2204
rect 1308 2196 1316 2204
rect 44 2176 52 2184
rect 412 2176 420 2184
rect 492 2176 500 2184
rect 1052 2176 1060 2184
rect 1084 2176 1092 2184
rect 1100 2176 1108 2184
rect 1132 2176 1140 2184
rect 1324 2176 1332 2184
rect 1340 2176 1348 2184
rect 1372 2176 1380 2184
rect 1404 2176 1412 2184
rect 1724 2176 1732 2184
rect 1884 2176 1892 2184
rect 1948 2176 1956 2184
rect 2348 2176 2356 2184
rect 2396 2176 2404 2184
rect 2652 2176 2660 2184
rect 2716 2176 2724 2184
rect 2828 2176 2836 2184
rect 3148 2176 3156 2184
rect 3548 2176 3556 2184
rect 3564 2176 3572 2184
rect 3948 2176 3956 2184
rect 4428 2176 4436 2184
rect 4732 2176 4740 2184
rect 4796 2176 4804 2184
rect 4844 2176 4852 2184
rect 4876 2176 4884 2184
rect 5116 2176 5124 2184
rect 5260 2176 5268 2184
rect 5372 2176 5380 2184
rect 5500 2176 5508 2184
rect 5564 2176 5572 2184
rect 5676 2176 5684 2184
rect 6764 2176 6772 2184
rect 6828 2176 6836 2184
rect 6972 2176 6980 2184
rect 7244 2176 7252 2184
rect 60 2156 68 2164
rect 140 2156 148 2164
rect 156 2156 164 2164
rect 316 2156 324 2164
rect 364 2156 372 2164
rect 428 2156 436 2164
rect 908 2156 916 2164
rect 1036 2156 1044 2164
rect 1148 2156 1156 2164
rect 1180 2156 1188 2164
rect 1228 2156 1236 2164
rect 1308 2156 1316 2164
rect 1532 2156 1540 2164
rect 1708 2156 1716 2164
rect 1836 2156 1844 2164
rect 2172 2156 2180 2164
rect 2204 2156 2212 2164
rect 2220 2156 2228 2164
rect 2508 2156 2516 2164
rect 2636 2156 2644 2164
rect 3020 2156 3028 2164
rect 4012 2156 4020 2164
rect 4572 2156 4580 2164
rect 6380 2156 6388 2164
rect 6844 2156 6852 2164
rect 7276 2156 7284 2164
rect 28 2136 36 2144
rect 76 2136 84 2144
rect 172 2136 180 2144
rect 268 2136 276 2144
rect 396 2136 404 2144
rect 428 2136 436 2144
rect 476 2136 484 2144
rect 492 2136 500 2144
rect 12 2116 20 2124
rect 92 2116 100 2124
rect 124 2116 132 2124
rect 268 2116 276 2124
rect 380 2116 388 2124
rect 556 2116 564 2124
rect 620 2116 628 2124
rect 700 2116 708 2124
rect 748 2116 756 2124
rect 828 2116 836 2124
rect 860 2136 868 2144
rect 972 2136 980 2144
rect 1084 2136 1092 2144
rect 1132 2136 1140 2144
rect 1324 2136 1332 2144
rect 1404 2136 1412 2144
rect 1612 2136 1620 2144
rect 1692 2136 1700 2144
rect 1772 2136 1780 2144
rect 1836 2136 1844 2144
rect 1916 2136 1924 2144
rect 892 2116 900 2124
rect 956 2116 964 2124
rect 988 2116 996 2124
rect 1228 2116 1236 2124
rect 1260 2116 1268 2124
rect 1516 2116 1524 2124
rect 1564 2116 1572 2124
rect 1692 2116 1700 2124
rect 1788 2116 1796 2124
rect 1868 2116 1876 2124
rect 1916 2116 1924 2124
rect 2012 2132 2020 2140
rect 2028 2136 2036 2144
rect 2156 2136 2164 2144
rect 2252 2136 2260 2144
rect 1980 2116 1988 2124
rect 2044 2116 2052 2124
rect 2204 2116 2212 2124
rect 2300 2116 2308 2124
rect 2348 2136 2356 2144
rect 2396 2136 2404 2144
rect 2508 2136 2516 2144
rect 2540 2136 2548 2144
rect 2620 2136 2628 2144
rect 2684 2136 2692 2144
rect 2780 2136 2788 2144
rect 2796 2136 2804 2144
rect 2892 2136 2900 2144
rect 3100 2136 3108 2144
rect 3180 2136 3188 2144
rect 3196 2136 3204 2144
rect 3292 2136 3300 2144
rect 3372 2136 3380 2144
rect 3468 2136 3476 2144
rect 3500 2136 3508 2144
rect 3676 2136 3684 2144
rect 3772 2136 3780 2144
rect 3804 2136 3812 2144
rect 3932 2136 3940 2144
rect 3996 2136 4004 2144
rect 4556 2136 4564 2144
rect 4652 2136 4660 2144
rect 4668 2136 4676 2144
rect 4716 2136 4724 2144
rect 4812 2136 4820 2144
rect 4860 2136 4868 2144
rect 5292 2136 5300 2144
rect 5404 2136 5412 2144
rect 5516 2136 5524 2144
rect 5868 2136 5876 2144
rect 5932 2136 5940 2144
rect 6188 2136 6196 2144
rect 6332 2136 6340 2144
rect 6444 2136 6452 2144
rect 6572 2136 6580 2144
rect 6636 2136 6644 2144
rect 6844 2136 6852 2144
rect 6924 2136 6932 2144
rect 6956 2136 6964 2144
rect 7132 2136 7140 2144
rect 7164 2136 7172 2144
rect 7212 2136 7220 2144
rect 7260 2136 7268 2144
rect 7372 2136 7380 2144
rect 2396 2116 2404 2124
rect 2444 2116 2452 2124
rect 2540 2116 2548 2124
rect 2572 2116 2580 2124
rect 2604 2116 2612 2124
rect 2684 2116 2692 2124
rect 3004 2116 3012 2124
rect 3084 2116 3092 2124
rect 3132 2116 3140 2124
rect 3260 2116 3268 2124
rect 3436 2118 3444 2126
rect 3516 2116 3524 2124
rect 3724 2116 3732 2124
rect 3980 2116 3988 2124
rect 4044 2116 4052 2124
rect 4124 2116 4132 2124
rect 4188 2118 4196 2126
rect 4300 2118 4308 2126
rect 4540 2116 4548 2124
rect 4636 2116 4644 2124
rect 4764 2116 4772 2124
rect 4860 2116 4868 2124
rect 4940 2116 4948 2124
rect 5004 2118 5012 2126
rect 5084 2116 5092 2124
rect 5148 2116 5156 2124
rect 5228 2116 5236 2124
rect 5324 2116 5332 2124
rect 5452 2116 5460 2124
rect 5532 2116 5540 2124
rect 5580 2116 5588 2124
rect 5596 2116 5604 2124
rect 5644 2116 5652 2124
rect 5740 2116 5748 2124
rect 5788 2116 5796 2124
rect 5884 2116 5892 2124
rect 5916 2116 5924 2124
rect 6012 2116 6020 2124
rect 6028 2116 6036 2124
rect 6076 2116 6084 2124
rect 6092 2116 6100 2124
rect 6124 2116 6132 2124
rect 6172 2116 6180 2124
rect 6220 2116 6228 2124
rect 6284 2116 6292 2124
rect 6316 2116 6324 2124
rect 6348 2116 6356 2124
rect 6364 2116 6372 2124
rect 6412 2116 6420 2124
rect 6444 2116 6452 2124
rect 6524 2116 6532 2124
rect 6556 2116 6564 2124
rect 6620 2116 6628 2124
rect 6652 2116 6660 2124
rect 6700 2116 6708 2124
rect 6716 2116 6724 2124
rect 6732 2116 6740 2124
rect 6748 2116 6756 2124
rect 6796 2116 6804 2124
rect 6876 2116 6884 2124
rect 124 2096 132 2104
rect 236 2096 244 2104
rect 364 2096 372 2104
rect 444 2096 452 2104
rect 524 2096 532 2104
rect 604 2096 612 2104
rect 1052 2096 1060 2104
rect 1100 2096 1108 2104
rect 1356 2096 1364 2104
rect 1372 2096 1380 2104
rect 1644 2098 1652 2106
rect 1740 2096 1748 2104
rect 1852 2096 1860 2104
rect 1884 2096 1892 2104
rect 1964 2096 1972 2104
rect 2220 2096 2228 2104
rect 2460 2096 2468 2104
rect 2524 2096 2532 2104
rect 2572 2096 2580 2104
rect 3148 2096 3156 2104
rect 3548 2096 3556 2104
rect 3948 2096 3956 2104
rect 4460 2096 4468 2104
rect 4604 2096 4612 2104
rect 4716 2096 4724 2104
rect 4828 2096 4836 2104
rect 5068 2096 5076 2104
rect 5132 2096 5140 2104
rect 5244 2096 5252 2104
rect 5260 2096 5268 2104
rect 5308 2096 5316 2104
rect 5468 2096 5476 2104
rect 5484 2096 5492 2104
rect 6252 2096 6260 2104
rect 6284 2096 6292 2104
rect 6492 2096 6500 2104
rect 6524 2096 6532 2104
rect 7068 2116 7076 2124
rect 7324 2116 7332 2124
rect 6924 2096 6932 2104
rect 7196 2096 7204 2104
rect 7340 2096 7348 2104
rect 556 2076 564 2084
rect 604 2076 612 2084
rect 636 2076 644 2084
rect 684 2076 692 2084
rect 812 2076 820 2084
rect 1180 2076 1188 2084
rect 2316 2076 2324 2084
rect 2428 2076 2436 2084
rect 4060 2076 4068 2084
rect 4540 2076 4548 2084
rect 5100 2076 5108 2084
rect 5164 2076 5172 2084
rect 5212 2076 5220 2084
rect 2108 2056 2116 2064
rect 5148 2056 5156 2064
rect 5244 2076 5252 2084
rect 5340 2076 5348 2084
rect 5436 2076 5444 2084
rect 5420 2056 5428 2064
rect 556 2036 564 2044
rect 652 2036 660 2044
rect 700 2036 708 2044
rect 780 2036 788 2044
rect 828 2036 836 2044
rect 1420 2036 1428 2044
rect 1548 2036 1556 2044
rect 2076 2036 2084 2044
rect 2188 2036 2196 2044
rect 2300 2036 2308 2044
rect 2444 2036 2452 2044
rect 2908 2036 2916 2044
rect 3036 2036 3044 2044
rect 3052 2036 3060 2044
rect 3308 2036 3316 2044
rect 3612 2036 3620 2044
rect 3916 2036 3924 2044
rect 4044 2036 4052 2044
rect 4588 2036 4596 2044
rect 4636 2036 4644 2044
rect 5612 2036 5620 2044
rect 5916 2036 5924 2044
rect 6044 2036 6052 2044
rect 6140 2036 6148 2044
rect 1411 2006 1419 2014
rect 1421 2006 1429 2014
rect 1431 2006 1439 2014
rect 1441 2006 1449 2014
rect 1451 2006 1459 2014
rect 1461 2006 1469 2014
rect 4419 2006 4427 2014
rect 4429 2006 4437 2014
rect 4439 2006 4447 2014
rect 4449 2006 4457 2014
rect 4459 2006 4467 2014
rect 4469 2006 4477 2014
rect 140 1976 148 1984
rect 428 1976 436 1984
rect 956 1976 964 1984
rect 1596 1976 1604 1984
rect 1724 1976 1732 1984
rect 2028 1976 2036 1984
rect 2108 1976 2116 1984
rect 2444 1976 2452 1984
rect 2828 1976 2836 1984
rect 3020 1976 3028 1984
rect 3212 1976 3220 1984
rect 3356 1976 3364 1984
rect 4268 1976 4276 1984
rect 4364 1976 4372 1984
rect 4716 1976 4724 1984
rect 4892 1976 4900 1984
rect 4972 1976 4980 1984
rect 5052 1976 5060 1984
rect 5324 1976 5332 1984
rect 6204 1976 6212 1984
rect 6412 1976 6420 1984
rect 364 1936 372 1944
rect 524 1936 532 1944
rect 604 1936 612 1944
rect 668 1936 676 1944
rect 1100 1936 1108 1944
rect 1164 1956 1172 1964
rect 1548 1956 1556 1964
rect 3692 1956 3700 1964
rect 6060 1956 6068 1964
rect 7004 1956 7012 1964
rect 12 1896 20 1904
rect 44 1896 52 1904
rect 76 1896 84 1904
rect 172 1916 180 1924
rect 188 1916 196 1924
rect 572 1916 580 1924
rect 636 1916 644 1924
rect 940 1916 948 1924
rect 1180 1936 1188 1944
rect 1388 1936 1396 1944
rect 1404 1936 1412 1944
rect 1644 1936 1652 1944
rect 1964 1936 1972 1944
rect 1996 1936 2004 1944
rect 2124 1936 2132 1944
rect 2460 1936 2468 1944
rect 3900 1936 3908 1944
rect 4252 1936 4260 1944
rect 4700 1936 4708 1944
rect 4812 1936 4820 1944
rect 5340 1936 5348 1944
rect 5532 1936 5540 1944
rect 5900 1936 5908 1944
rect 6796 1936 6804 1944
rect 7196 1936 7204 1944
rect 1212 1916 1220 1924
rect 1340 1916 1348 1924
rect 1484 1916 1492 1924
rect 1580 1916 1588 1924
rect 1692 1916 1700 1924
rect 1788 1916 1796 1924
rect 2012 1916 2020 1924
rect 2156 1916 2164 1924
rect 2668 1916 2676 1924
rect 2764 1916 2772 1924
rect 3116 1916 3124 1924
rect 3164 1916 3172 1924
rect 3468 1916 3476 1924
rect 3580 1916 3588 1924
rect 3756 1916 3764 1924
rect 3820 1916 3828 1924
rect 4092 1916 4100 1924
rect 4284 1916 4292 1924
rect 4348 1916 4356 1924
rect 4492 1916 4500 1924
rect 4556 1916 4564 1924
rect 4620 1916 4628 1924
rect 4732 1916 4740 1924
rect 4796 1916 4804 1924
rect 5308 1916 5316 1924
rect 5372 1916 5380 1924
rect 5980 1916 5988 1924
rect 6092 1916 6100 1924
rect 140 1896 148 1904
rect 236 1896 244 1904
rect 460 1896 468 1904
rect 588 1896 596 1904
rect 652 1896 660 1904
rect 684 1896 692 1904
rect 796 1896 804 1904
rect 860 1896 868 1904
rect 892 1896 900 1904
rect 988 1896 996 1904
rect 1068 1896 1076 1904
rect 1116 1896 1124 1904
rect 44 1876 52 1884
rect 108 1876 116 1884
rect 124 1876 132 1884
rect 204 1876 212 1884
rect 236 1876 244 1884
rect 396 1876 404 1884
rect 444 1876 452 1884
rect 556 1876 564 1884
rect 620 1876 628 1884
rect 700 1876 708 1884
rect 716 1880 724 1888
rect 812 1876 820 1884
rect 876 1876 884 1884
rect 940 1876 948 1884
rect 972 1876 980 1884
rect 1036 1876 1044 1884
rect 1164 1896 1172 1904
rect 1212 1896 1220 1904
rect 1260 1896 1268 1904
rect 1324 1896 1332 1904
rect 1548 1896 1556 1904
rect 1628 1896 1636 1904
rect 1708 1896 1716 1904
rect 1804 1896 1812 1904
rect 1836 1896 1844 1904
rect 1868 1896 1876 1904
rect 1244 1876 1252 1884
rect 1276 1876 1284 1884
rect 1324 1876 1332 1884
rect 1372 1876 1380 1884
rect 1388 1876 1396 1884
rect 1644 1876 1652 1884
rect 1660 1876 1668 1884
rect 1756 1876 1764 1884
rect 1788 1876 1796 1884
rect 1916 1876 1924 1884
rect 12 1856 20 1864
rect 284 1856 292 1864
rect 412 1856 420 1864
rect 1036 1856 1044 1864
rect 1260 1856 1268 1864
rect 1276 1856 1284 1864
rect 1500 1856 1508 1864
rect 1740 1856 1748 1864
rect 1772 1856 1780 1864
rect 1836 1856 1844 1864
rect 1868 1856 1876 1864
rect 2092 1896 2100 1904
rect 2140 1896 2148 1904
rect 1996 1876 2004 1884
rect 2044 1876 2052 1884
rect 2348 1896 2356 1904
rect 2396 1896 2404 1904
rect 2476 1896 2484 1904
rect 2524 1896 2532 1904
rect 2556 1896 2564 1904
rect 2636 1896 2644 1904
rect 2748 1896 2756 1904
rect 2796 1896 2804 1904
rect 3276 1896 3284 1904
rect 3324 1896 3332 1904
rect 3356 1896 3364 1904
rect 3388 1896 3396 1904
rect 3452 1896 3460 1904
rect 3500 1896 3508 1904
rect 3548 1896 3556 1904
rect 3644 1896 3652 1904
rect 3660 1896 3668 1904
rect 3724 1896 3732 1904
rect 3788 1896 3796 1904
rect 3884 1896 3892 1904
rect 3964 1896 3972 1904
rect 4012 1896 4020 1904
rect 4140 1896 4148 1904
rect 4268 1896 4276 1904
rect 4316 1896 4324 1904
rect 4476 1896 4484 1904
rect 4524 1896 4532 1904
rect 4588 1896 4596 1904
rect 4652 1896 4660 1904
rect 4716 1896 4724 1904
rect 4764 1896 4772 1904
rect 4860 1896 4868 1904
rect 5148 1896 5156 1904
rect 5212 1894 5220 1902
rect 5356 1896 5364 1904
rect 5404 1896 5412 1904
rect 5596 1896 5604 1904
rect 5660 1894 5668 1902
rect 5788 1896 5796 1904
rect 6012 1896 6020 1904
rect 6076 1896 6084 1904
rect 6140 1916 6148 1924
rect 6284 1896 6292 1904
rect 6300 1896 6308 1904
rect 6348 1896 6356 1904
rect 6364 1896 6372 1904
rect 6396 1896 6404 1904
rect 6444 1896 6452 1904
rect 6460 1896 6468 1904
rect 6476 1896 6484 1904
rect 6572 1896 6580 1904
rect 6620 1896 6628 1904
rect 6684 1896 6692 1904
rect 6716 1896 6724 1904
rect 6764 1916 6772 1924
rect 7068 1916 7076 1924
rect 7116 1916 7124 1924
rect 6908 1896 6916 1904
rect 7068 1896 7076 1904
rect 7180 1896 7188 1904
rect 7260 1896 7268 1904
rect 7308 1896 7316 1904
rect 2284 1876 2292 1884
rect 2300 1876 2308 1884
rect 2332 1876 2340 1884
rect 2412 1876 2420 1884
rect 2540 1876 2548 1884
rect 2652 1876 2660 1884
rect 2700 1876 2708 1884
rect 2812 1876 2820 1884
rect 2908 1876 2916 1884
rect 2988 1876 2996 1884
rect 3084 1876 3092 1884
rect 3132 1876 3140 1884
rect 3180 1876 3188 1884
rect 3292 1876 3300 1884
rect 3340 1876 3348 1884
rect 3516 1876 3524 1884
rect 3532 1876 3540 1884
rect 3628 1876 3636 1884
rect 3772 1876 3780 1884
rect 3884 1876 3892 1884
rect 4124 1876 4132 1884
rect 4300 1876 4308 1884
rect 4396 1876 4404 1884
rect 4540 1876 4548 1884
rect 4604 1876 4612 1884
rect 4668 1876 4676 1884
rect 4748 1876 4756 1884
rect 4844 1876 4852 1884
rect 4876 1876 4884 1884
rect 4956 1876 4964 1884
rect 5276 1876 5284 1884
rect 5516 1876 5524 1884
rect 5740 1876 5748 1884
rect 5916 1876 5924 1884
rect 6012 1876 6020 1884
rect 6076 1876 6084 1884
rect 6172 1876 6180 1884
rect 6188 1876 6196 1884
rect 6236 1876 6244 1884
rect 2060 1856 2068 1864
rect 2348 1856 2356 1864
rect 2380 1856 2388 1864
rect 2444 1856 2452 1864
rect 2476 1856 2484 1864
rect 2588 1856 2596 1864
rect 2716 1856 2724 1864
rect 2732 1856 2740 1864
rect 2924 1856 2932 1864
rect 3100 1856 3108 1864
rect 3164 1856 3172 1864
rect 3324 1856 3332 1864
rect 3420 1856 3428 1864
rect 4092 1856 4100 1864
rect 4156 1856 4164 1864
rect 4204 1856 4212 1864
rect 4220 1856 4228 1864
rect 6508 1856 6516 1864
rect 6556 1876 6564 1884
rect 6668 1876 6676 1884
rect 6764 1876 6772 1884
rect 6796 1876 6804 1884
rect 6924 1876 6932 1884
rect 6972 1876 6980 1884
rect 7036 1876 7044 1884
rect 7084 1876 7092 1884
rect 7148 1876 7156 1884
rect 6588 1856 6596 1864
rect 7020 1856 7028 1864
rect 7180 1856 7188 1864
rect 748 1836 756 1844
rect 764 1836 772 1844
rect 828 1836 836 1844
rect 1052 1836 1060 1844
rect 1324 1836 1332 1844
rect 1388 1836 1396 1844
rect 1676 1836 1684 1844
rect 1788 1836 1796 1844
rect 2012 1836 2020 1844
rect 2204 1836 2212 1844
rect 2316 1836 2324 1844
rect 2572 1836 2580 1844
rect 2604 1836 2612 1844
rect 2668 1836 2676 1844
rect 3612 1836 3620 1844
rect 3756 1836 3764 1844
rect 3852 1836 3860 1844
rect 4492 1836 4500 1844
rect 4556 1836 4564 1844
rect 4620 1836 4628 1844
rect 5084 1836 5092 1844
rect 5308 1836 5316 1844
rect 6316 1836 6324 1844
rect 6540 1836 6548 1844
rect 6652 1836 6660 1844
rect 1500 1816 1508 1824
rect 2915 1806 2923 1814
rect 2925 1806 2933 1814
rect 2935 1806 2943 1814
rect 2945 1806 2953 1814
rect 2955 1806 2963 1814
rect 2965 1806 2973 1814
rect 5923 1806 5931 1814
rect 5933 1806 5941 1814
rect 5943 1806 5951 1814
rect 5953 1806 5961 1814
rect 5963 1806 5971 1814
rect 5973 1806 5981 1814
rect 12 1776 20 1784
rect 124 1776 132 1784
rect 204 1776 212 1784
rect 236 1776 244 1784
rect 300 1776 308 1784
rect 524 1776 532 1784
rect 700 1776 708 1784
rect 716 1776 724 1784
rect 924 1776 932 1784
rect 1164 1776 1172 1784
rect 1244 1776 1252 1784
rect 1436 1776 1444 1784
rect 1644 1776 1652 1784
rect 2444 1776 2452 1784
rect 2476 1776 2484 1784
rect 2716 1776 2724 1784
rect 3084 1776 3092 1784
rect 3244 1776 3252 1784
rect 3388 1776 3396 1784
rect 3676 1776 3684 1784
rect 3724 1776 3732 1784
rect 3772 1776 3780 1784
rect 4012 1776 4020 1784
rect 4348 1776 4356 1784
rect 4364 1776 4372 1784
rect 4588 1776 4596 1784
rect 4780 1776 4788 1784
rect 4956 1776 4964 1784
rect 5228 1776 5236 1784
rect 5276 1776 5284 1784
rect 5532 1776 5540 1784
rect 5548 1776 5556 1784
rect 5612 1776 5620 1784
rect 5660 1776 5668 1784
rect 5708 1776 5716 1784
rect 5804 1776 5812 1784
rect 6236 1776 6244 1784
rect 6300 1776 6308 1784
rect 6780 1776 6788 1784
rect 6796 1776 6804 1784
rect 7228 1776 7236 1784
rect 60 1756 68 1764
rect 108 1756 116 1764
rect 220 1756 228 1764
rect 332 1756 340 1764
rect 140 1736 148 1744
rect 172 1736 180 1744
rect 284 1736 292 1744
rect 380 1756 388 1764
rect 604 1756 612 1764
rect 1228 1756 1236 1764
rect 1660 1756 1668 1764
rect 2284 1756 2292 1764
rect 2380 1756 2388 1764
rect 2492 1756 2500 1764
rect 2508 1756 2516 1764
rect 2732 1756 2740 1764
rect 2780 1756 2788 1764
rect 460 1732 468 1740
rect 476 1736 484 1744
rect 492 1736 500 1744
rect 588 1736 596 1744
rect 652 1736 660 1744
rect 716 1736 724 1744
rect 924 1736 932 1744
rect 92 1716 100 1724
rect 172 1716 180 1724
rect 252 1716 260 1724
rect 268 1716 276 1724
rect 332 1716 340 1724
rect 348 1716 356 1724
rect 412 1716 420 1724
rect 428 1716 436 1724
rect 636 1716 644 1724
rect 668 1716 676 1724
rect 748 1716 756 1724
rect 780 1716 788 1724
rect 860 1716 868 1724
rect 892 1716 900 1724
rect 972 1716 980 1724
rect 1004 1716 1012 1724
rect 1164 1736 1172 1744
rect 1212 1736 1220 1744
rect 1292 1736 1300 1744
rect 1068 1716 1076 1724
rect 1148 1716 1156 1724
rect 1164 1716 1172 1724
rect 1196 1716 1204 1724
rect 1228 1716 1236 1724
rect 1276 1716 1284 1724
rect 1340 1716 1348 1724
rect 1388 1736 1396 1744
rect 1436 1736 1444 1744
rect 1548 1736 1556 1744
rect 1596 1732 1604 1740
rect 1612 1736 1620 1744
rect 1484 1716 1492 1724
rect 1516 1716 1524 1724
rect 1628 1716 1636 1724
rect 1708 1716 1716 1724
rect 1772 1716 1780 1724
rect 1836 1716 1844 1724
rect 2108 1736 2116 1744
rect 2204 1736 2212 1744
rect 1868 1716 1876 1724
rect 1948 1716 1956 1724
rect 2012 1716 2020 1724
rect 2076 1716 2084 1724
rect 2108 1716 2116 1724
rect 2396 1736 2404 1744
rect 2444 1736 2452 1744
rect 2540 1736 2548 1744
rect 2556 1736 2564 1744
rect 2668 1736 2676 1744
rect 2732 1736 2740 1744
rect 2876 1736 2884 1744
rect 2988 1756 2996 1764
rect 3212 1756 3220 1764
rect 3004 1736 3012 1744
rect 3052 1736 3060 1744
rect 3068 1736 3076 1744
rect 3100 1736 3108 1744
rect 3164 1736 3172 1744
rect 3228 1736 3236 1744
rect 3260 1736 3268 1744
rect 3372 1736 3380 1744
rect 3436 1736 3444 1744
rect 3468 1736 3476 1744
rect 3516 1756 3524 1764
rect 3564 1756 3572 1764
rect 3916 1756 3924 1764
rect 4092 1756 4100 1764
rect 4236 1756 4244 1764
rect 4300 1756 4308 1764
rect 5260 1756 5268 1764
rect 5772 1756 5780 1764
rect 5788 1756 5796 1764
rect 5852 1756 5860 1764
rect 6284 1756 6292 1764
rect 6492 1756 6500 1764
rect 6924 1756 6932 1764
rect 7324 1756 7332 1764
rect 7340 1756 7348 1764
rect 3628 1736 3636 1744
rect 4028 1736 4036 1744
rect 4108 1736 4116 1744
rect 4204 1736 4212 1744
rect 4620 1736 4628 1744
rect 4652 1736 4660 1744
rect 4684 1736 4692 1744
rect 4796 1736 4804 1744
rect 4812 1736 4820 1744
rect 4988 1736 4996 1744
rect 5132 1736 5140 1744
rect 5148 1736 5156 1744
rect 5212 1736 5220 1744
rect 5292 1736 5300 1744
rect 5452 1736 5460 1744
rect 5500 1736 5508 1744
rect 5580 1736 5588 1744
rect 5644 1736 5652 1744
rect 5692 1736 5700 1744
rect 5820 1736 5828 1744
rect 5884 1736 5892 1744
rect 2236 1716 2244 1724
rect 2332 1716 2340 1724
rect 2380 1716 2388 1724
rect 2444 1716 2452 1724
rect 2460 1716 2468 1724
rect 2684 1716 2692 1724
rect 2764 1716 2772 1724
rect 2812 1716 2820 1724
rect 2828 1716 2836 1724
rect 3052 1716 3060 1724
rect 3180 1716 3188 1724
rect 3420 1716 3428 1724
rect 3452 1716 3460 1724
rect 3484 1716 3492 1724
rect 3596 1716 3604 1724
rect 3644 1716 3652 1724
rect 3692 1716 3700 1724
rect 3740 1716 3748 1724
rect 3868 1716 3876 1724
rect 3980 1716 3988 1724
rect 4060 1716 4068 1724
rect 4124 1716 4132 1724
rect 4220 1716 4228 1724
rect 4316 1716 4324 1724
rect 4396 1716 4404 1724
rect 4556 1716 4564 1724
rect 4668 1716 4676 1724
rect 4716 1716 4724 1724
rect 4908 1716 4916 1724
rect 5308 1716 5316 1724
rect 5356 1716 5364 1724
rect 5420 1716 5428 1724
rect 5484 1716 5492 1724
rect 5740 1716 5748 1724
rect 5836 1716 5844 1724
rect 6012 1736 6020 1744
rect 6044 1736 6052 1744
rect 6092 1736 6100 1744
rect 6252 1736 6260 1744
rect 6524 1736 6532 1744
rect 6588 1736 6596 1744
rect 6620 1736 6628 1744
rect 6668 1736 6676 1744
rect 7004 1736 7012 1744
rect 7212 1736 7220 1744
rect 7260 1736 7268 1744
rect 7292 1736 7300 1744
rect 7308 1736 7316 1744
rect 6076 1718 6084 1726
rect 6364 1716 6372 1724
rect 6428 1718 6436 1726
rect 6492 1716 6500 1724
rect 6652 1718 6660 1726
rect 6860 1716 6868 1724
rect 6908 1716 6916 1724
rect 7052 1716 7060 1724
rect 7276 1716 7284 1724
rect 7372 1716 7380 1724
rect 12 1696 20 1704
rect 204 1696 212 1704
rect 748 1696 756 1704
rect 764 1696 772 1704
rect 876 1696 884 1704
rect 892 1696 900 1704
rect 988 1696 996 1704
rect 1004 1696 1012 1704
rect 1964 1696 1972 1704
rect 2028 1696 2036 1704
rect 2092 1696 2100 1704
rect 2316 1696 2324 1704
rect 2508 1696 2516 1704
rect 2716 1696 2724 1704
rect 2844 1696 2852 1704
rect 3132 1696 3140 1704
rect 3260 1696 3268 1704
rect 4156 1696 4164 1704
rect 4572 1696 4580 1704
rect 4588 1696 4596 1704
rect 4636 1696 4644 1704
rect 4748 1696 4756 1704
rect 4764 1696 4772 1704
rect 4892 1696 4900 1704
rect 5180 1696 5188 1704
rect 5372 1696 5380 1704
rect 5436 1696 5444 1704
rect 5532 1696 5540 1704
rect 5980 1696 5988 1704
rect 6220 1696 6228 1704
rect 6252 1696 6260 1704
rect 6556 1696 6564 1704
rect 7180 1696 7188 1704
rect 7228 1696 7236 1704
rect 796 1676 804 1684
rect 844 1676 852 1684
rect 956 1676 964 1684
rect 1084 1676 1092 1684
rect 1116 1676 1124 1684
rect 1324 1676 1332 1684
rect 1692 1676 1700 1684
rect 1756 1676 1764 1684
rect 1820 1676 1828 1684
rect 1900 1676 1908 1684
rect 1932 1676 1940 1684
rect 1996 1676 2004 1684
rect 2060 1676 2068 1684
rect 2220 1676 2228 1684
rect 2316 1676 2324 1684
rect 2348 1676 2356 1684
rect 2588 1676 2596 1684
rect 2780 1676 2788 1684
rect 3788 1676 3796 1684
rect 3820 1676 3828 1684
rect 4092 1676 4100 1684
rect 4540 1676 4548 1684
rect 4700 1676 4708 1684
rect 4716 1676 4724 1684
rect 4924 1676 4932 1684
rect 5340 1676 5348 1684
rect 5404 1676 5412 1684
rect 5548 1676 5556 1684
rect 5644 1676 5652 1684
rect 5692 1676 5700 1684
rect 5724 1676 5732 1684
rect 5852 1676 5860 1684
rect 7132 1676 7140 1684
rect 7196 1676 7204 1684
rect 2332 1656 2340 1664
rect 2396 1656 2404 1664
rect 4556 1656 4564 1664
rect 5356 1656 5364 1664
rect 6204 1656 6212 1664
rect 636 1636 644 1644
rect 780 1636 788 1644
rect 860 1636 868 1644
rect 972 1636 980 1644
rect 1068 1636 1076 1644
rect 1340 1636 1348 1644
rect 1388 1636 1396 1644
rect 1564 1636 1572 1644
rect 1708 1636 1716 1644
rect 1772 1636 1780 1644
rect 1836 1636 1844 1644
rect 1916 1636 1924 1644
rect 1980 1636 1988 1644
rect 2076 1636 2084 1644
rect 2236 1636 2244 1644
rect 2892 1636 2900 1644
rect 3308 1636 3316 1644
rect 3676 1636 3684 1644
rect 3724 1636 3732 1644
rect 4172 1636 4180 1644
rect 4252 1636 4260 1644
rect 4348 1636 4356 1644
rect 4364 1636 4372 1644
rect 4508 1636 4516 1644
rect 4860 1636 4868 1644
rect 5020 1636 5028 1644
rect 5388 1636 5396 1644
rect 7164 1636 7172 1644
rect 7388 1636 7396 1644
rect 1411 1606 1419 1614
rect 1421 1606 1429 1614
rect 1431 1606 1439 1614
rect 1441 1606 1449 1614
rect 1451 1606 1459 1614
rect 1461 1606 1469 1614
rect 4419 1606 4427 1614
rect 4429 1606 4437 1614
rect 4439 1606 4447 1614
rect 4449 1606 4457 1614
rect 4459 1606 4467 1614
rect 4469 1606 4477 1614
rect 108 1576 116 1584
rect 172 1576 180 1584
rect 444 1576 452 1584
rect 748 1576 756 1584
rect 812 1576 820 1584
rect 876 1576 884 1584
rect 892 1576 900 1584
rect 1756 1576 1764 1584
rect 2156 1576 2164 1584
rect 3004 1576 3012 1584
rect 3164 1576 3172 1584
rect 3212 1576 3220 1584
rect 3388 1576 3396 1584
rect 3868 1576 3876 1584
rect 4636 1576 4644 1584
rect 4668 1576 4676 1584
rect 5132 1576 5140 1584
rect 5276 1576 5284 1584
rect 5340 1576 5348 1584
rect 5404 1576 5412 1584
rect 5452 1576 5460 1584
rect 5548 1576 5556 1584
rect 6108 1576 6116 1584
rect 6204 1576 6212 1584
rect 620 1556 628 1564
rect 1308 1556 1316 1564
rect 700 1536 708 1544
rect 732 1536 740 1544
rect 796 1536 804 1544
rect 860 1536 868 1544
rect 956 1536 964 1544
rect 1068 1536 1076 1544
rect 1196 1536 1204 1544
rect 1324 1536 1332 1544
rect 1388 1536 1396 1544
rect 2108 1536 2116 1544
rect 2172 1536 2180 1544
rect 2252 1536 2260 1544
rect 2364 1536 2372 1544
rect 2428 1556 2436 1564
rect 4764 1556 4772 1564
rect 6268 1556 6276 1564
rect 7196 1556 7204 1564
rect 668 1516 676 1524
rect 764 1516 772 1524
rect 828 1516 836 1524
rect 988 1516 996 1524
rect 1228 1516 1236 1524
rect 1356 1516 1364 1524
rect 1596 1516 1604 1524
rect 2172 1516 2180 1524
rect 2284 1516 2292 1524
rect 2444 1536 2452 1544
rect 4604 1536 4612 1544
rect 5116 1536 5124 1544
rect 5324 1536 5332 1544
rect 5388 1536 5396 1544
rect 5660 1536 5668 1544
rect 5804 1536 5812 1544
rect 5884 1536 5892 1544
rect 2492 1516 2500 1524
rect 12 1496 20 1504
rect 44 1496 52 1504
rect 60 1496 68 1504
rect 140 1496 148 1504
rect 268 1496 276 1504
rect 284 1496 292 1504
rect 316 1496 324 1504
rect 332 1496 340 1504
rect 524 1496 532 1504
rect 684 1496 692 1504
rect 716 1496 724 1504
rect 780 1496 788 1504
rect 844 1496 852 1504
rect 924 1496 932 1504
rect 972 1496 980 1504
rect 1036 1496 1044 1504
rect 1052 1496 1060 1504
rect 1132 1496 1140 1504
rect 1212 1496 1220 1504
rect 1276 1496 1284 1504
rect 156 1476 164 1484
rect 204 1476 212 1484
rect 220 1476 228 1484
rect 476 1476 484 1484
rect 540 1476 548 1484
rect 556 1480 564 1488
rect 972 1476 980 1484
rect 1068 1476 1076 1484
rect 1116 1476 1124 1484
rect 1308 1496 1316 1504
rect 1372 1496 1380 1504
rect 1404 1496 1412 1504
rect 1532 1496 1540 1504
rect 1564 1496 1572 1504
rect 1724 1496 1732 1504
rect 1756 1496 1764 1504
rect 1852 1496 1860 1504
rect 1900 1496 1908 1504
rect 2076 1496 2084 1504
rect 2156 1496 2164 1504
rect 2188 1496 2196 1504
rect 2236 1496 2244 1504
rect 2268 1496 2276 1504
rect 2332 1496 2340 1504
rect 2380 1496 2388 1504
rect 1580 1476 1588 1484
rect 1628 1476 1636 1484
rect 1644 1476 1652 1484
rect 1868 1476 1876 1484
rect 1884 1476 1892 1484
rect 1948 1476 1956 1484
rect 2044 1476 2052 1484
rect 2060 1476 2068 1484
rect 2428 1496 2436 1504
rect 2476 1496 2484 1504
rect 2540 1496 2548 1504
rect 2588 1496 2596 1504
rect 2620 1496 2628 1504
rect 2636 1496 2644 1504
rect 2668 1496 2676 1504
rect 2700 1496 2708 1504
rect 2764 1496 2772 1504
rect 2796 1496 2804 1504
rect 2908 1516 2916 1524
rect 3404 1516 3412 1524
rect 3660 1516 3668 1524
rect 3788 1516 3796 1524
rect 3916 1516 3924 1524
rect 4412 1516 4420 1524
rect 4748 1516 4756 1524
rect 5180 1516 5188 1524
rect 5292 1516 5300 1524
rect 5372 1516 5380 1524
rect 5628 1516 5636 1524
rect 5740 1516 5748 1524
rect 5900 1516 5908 1524
rect 5932 1516 5940 1524
rect 6252 1516 6260 1524
rect 6364 1516 6372 1524
rect 2892 1496 2900 1504
rect 3100 1496 3108 1504
rect 3148 1496 3156 1504
rect 3196 1496 3204 1504
rect 3244 1496 3252 1504
rect 2492 1476 2500 1484
rect 2556 1476 2564 1484
rect 2604 1476 2612 1484
rect 2684 1476 2692 1484
rect 12 1456 20 1464
rect 44 1456 52 1464
rect 92 1456 100 1464
rect 220 1456 228 1464
rect 236 1456 244 1464
rect 364 1456 372 1464
rect 492 1456 500 1464
rect 508 1456 516 1464
rect 636 1456 644 1464
rect 652 1456 660 1464
rect 1004 1456 1012 1464
rect 1052 1456 1060 1464
rect 1132 1456 1140 1464
rect 1244 1456 1252 1464
rect 1484 1456 1492 1464
rect 1532 1456 1540 1464
rect 1596 1456 1604 1464
rect 1660 1456 1668 1464
rect 1676 1456 1684 1464
rect 1804 1456 1812 1464
rect 2124 1456 2132 1464
rect 2220 1456 2228 1464
rect 2300 1456 2308 1464
rect 2476 1456 2484 1464
rect 2620 1456 2628 1464
rect 2668 1456 2676 1464
rect 2844 1476 2852 1484
rect 3036 1476 3044 1484
rect 3116 1476 3124 1484
rect 3260 1476 3268 1484
rect 3356 1476 3364 1484
rect 3548 1494 3556 1502
rect 3628 1496 3636 1504
rect 3724 1496 3732 1504
rect 3756 1496 3764 1504
rect 3852 1496 3860 1504
rect 3900 1496 3908 1504
rect 3948 1496 3956 1504
rect 4108 1494 4116 1502
rect 4236 1496 4244 1504
rect 4284 1496 4292 1504
rect 4364 1496 4372 1504
rect 4540 1496 4548 1504
rect 4604 1496 4612 1504
rect 4716 1496 4724 1504
rect 4812 1496 4820 1504
rect 4892 1496 4900 1504
rect 4940 1496 4948 1504
rect 5020 1496 5028 1504
rect 5068 1496 5076 1504
rect 5132 1496 5140 1504
rect 5244 1496 5252 1504
rect 5308 1496 5316 1504
rect 5372 1496 5380 1504
rect 5420 1496 5428 1504
rect 5468 1496 5476 1504
rect 5516 1496 5524 1504
rect 5852 1496 5860 1504
rect 6044 1496 6052 1504
rect 6076 1496 6084 1504
rect 6172 1496 6180 1504
rect 6396 1496 6404 1504
rect 6444 1516 6452 1524
rect 6524 1516 6532 1524
rect 6572 1516 6580 1524
rect 6988 1516 6996 1524
rect 7004 1516 7012 1524
rect 7180 1516 7188 1524
rect 7276 1516 7284 1524
rect 7324 1516 7332 1524
rect 6572 1496 6580 1504
rect 6636 1494 6644 1502
rect 6860 1496 6868 1504
rect 6908 1494 6916 1502
rect 7020 1496 7028 1504
rect 7036 1496 7044 1504
rect 7084 1496 7092 1504
rect 7244 1496 7252 1504
rect 7276 1496 7284 1504
rect 3612 1476 3620 1484
rect 3708 1476 3716 1484
rect 3724 1476 3732 1484
rect 3804 1476 3812 1484
rect 3836 1476 3844 1484
rect 3964 1476 3972 1484
rect 4076 1476 4084 1484
rect 4140 1476 4148 1484
rect 4332 1476 4340 1484
rect 4364 1476 4372 1484
rect 4524 1476 4532 1484
rect 4684 1476 4692 1484
rect 4700 1476 4708 1484
rect 4796 1476 4804 1484
rect 5052 1476 5060 1484
rect 5180 1476 5188 1484
rect 5212 1476 5220 1484
rect 5228 1476 5236 1484
rect 5596 1476 5604 1484
rect 5660 1476 5668 1484
rect 5708 1480 5716 1488
rect 5724 1476 5732 1484
rect 5772 1476 5780 1484
rect 5868 1476 5876 1484
rect 5916 1476 5924 1484
rect 6060 1476 6068 1484
rect 6156 1476 6164 1484
rect 6220 1476 6228 1484
rect 6300 1480 6308 1488
rect 6332 1476 6340 1484
rect 6380 1476 6388 1484
rect 6476 1476 6484 1484
rect 6540 1476 6548 1484
rect 6668 1476 6676 1484
rect 7052 1476 7060 1484
rect 7068 1476 7076 1484
rect 7164 1476 7172 1484
rect 7212 1476 7220 1484
rect 7356 1476 7364 1484
rect 2988 1456 2996 1464
rect 3052 1456 3060 1464
rect 3548 1456 3556 1464
rect 4508 1456 4516 1464
rect 4556 1456 4564 1464
rect 5020 1456 5028 1464
rect 5084 1456 5092 1464
rect 5564 1456 5572 1464
rect 5788 1456 5796 1464
rect 5820 1456 5828 1464
rect 5996 1456 6004 1464
rect 6124 1456 6132 1464
rect 6972 1456 6980 1464
rect 7292 1456 7300 1464
rect 7308 1456 7316 1464
rect 892 1436 900 1444
rect 1020 1436 1028 1444
rect 1116 1436 1124 1444
rect 1148 1436 1156 1444
rect 1260 1436 1268 1444
rect 1820 1436 1828 1444
rect 1932 1436 1940 1444
rect 2012 1436 2020 1444
rect 2316 1436 2324 1444
rect 2556 1436 2564 1444
rect 2860 1436 2868 1444
rect 3068 1436 3076 1444
rect 3420 1436 3428 1444
rect 3692 1436 3700 1444
rect 3916 1436 3924 1444
rect 3980 1436 3988 1444
rect 4172 1436 4180 1444
rect 5004 1436 5012 1444
rect 5500 1436 5508 1444
rect 5580 1436 5588 1444
rect 5740 1436 5748 1444
rect 5836 1436 5844 1444
rect 6012 1436 6020 1444
rect 6140 1436 6148 1444
rect 6204 1436 6212 1444
rect 6236 1436 6244 1444
rect 6364 1436 6372 1444
rect 6428 1436 6436 1444
rect 6508 1436 6516 1444
rect 6764 1436 6772 1444
rect 6780 1436 6788 1444
rect 7116 1436 7124 1444
rect 7148 1436 7156 1444
rect 7324 1436 7332 1444
rect 1484 1416 1492 1424
rect 1660 1416 1668 1424
rect 1676 1416 1684 1424
rect 1804 1416 1812 1424
rect 2915 1406 2923 1414
rect 2925 1406 2933 1414
rect 2935 1406 2943 1414
rect 2945 1406 2953 1414
rect 2955 1406 2963 1414
rect 2965 1406 2973 1414
rect 5923 1406 5931 1414
rect 5933 1406 5941 1414
rect 5943 1406 5951 1414
rect 5953 1406 5961 1414
rect 5963 1406 5971 1414
rect 5973 1406 5981 1414
rect 828 1396 836 1404
rect 76 1376 84 1384
rect 156 1376 164 1384
rect 268 1376 276 1384
rect 316 1376 324 1384
rect 332 1376 340 1384
rect 476 1376 484 1384
rect 652 1376 660 1384
rect 812 1376 820 1384
rect 956 1376 964 1384
rect 988 1376 996 1384
rect 1164 1376 1172 1384
rect 1260 1376 1268 1384
rect 1324 1376 1332 1384
rect 1628 1376 1636 1384
rect 1724 1376 1732 1384
rect 1836 1376 1844 1384
rect 2092 1376 2100 1384
rect 2108 1376 2116 1384
rect 2156 1376 2164 1384
rect 2364 1376 2372 1384
rect 2396 1376 2404 1384
rect 2588 1376 2596 1384
rect 2860 1376 2868 1384
rect 3276 1376 3284 1384
rect 3404 1376 3412 1384
rect 3868 1376 3876 1384
rect 3948 1376 3956 1384
rect 4460 1376 4468 1384
rect 4700 1376 4708 1384
rect 4780 1376 4788 1384
rect 4828 1376 4836 1384
rect 4972 1376 4980 1384
rect 5020 1376 5028 1384
rect 5068 1376 5076 1384
rect 5180 1376 5188 1384
rect 5308 1376 5316 1384
rect 5356 1376 5364 1384
rect 5404 1376 5412 1384
rect 5484 1376 5492 1384
rect 5596 1376 5604 1384
rect 5820 1376 5828 1384
rect 5900 1376 5908 1384
rect 6156 1376 6164 1384
rect 6188 1376 6196 1384
rect 6220 1376 6228 1384
rect 6332 1376 6340 1384
rect 6524 1376 6532 1384
rect 6636 1376 6644 1384
rect 6716 1376 6724 1384
rect 6988 1376 6996 1384
rect 7260 1376 7268 1384
rect 7308 1376 7316 1384
rect 412 1356 420 1364
rect 524 1356 532 1364
rect 700 1356 708 1364
rect 828 1356 836 1364
rect 972 1356 980 1364
rect 1068 1356 1076 1364
rect 1340 1356 1348 1364
rect 1692 1356 1700 1364
rect 1708 1356 1716 1364
rect 1932 1356 1940 1364
rect 2300 1356 2308 1364
rect 2348 1356 2356 1364
rect 2444 1356 2452 1364
rect 2572 1356 2580 1364
rect 92 1336 100 1344
rect 140 1336 148 1344
rect 204 1336 212 1344
rect 220 1336 228 1344
rect 588 1336 596 1344
rect 604 1336 612 1344
rect 44 1316 52 1324
rect 108 1316 116 1324
rect 188 1316 196 1324
rect 236 1316 244 1324
rect 284 1316 292 1324
rect 364 1316 372 1324
rect 380 1316 388 1324
rect 428 1316 436 1324
rect 508 1316 516 1324
rect 556 1316 564 1324
rect 620 1316 628 1324
rect 668 1316 676 1324
rect 732 1316 740 1324
rect 924 1336 932 1344
rect 956 1336 964 1344
rect 1004 1336 1012 1344
rect 876 1316 884 1324
rect 60 1296 68 1304
rect 812 1296 820 1304
rect 1020 1316 1028 1324
rect 1036 1316 1044 1324
rect 1068 1316 1076 1324
rect 1100 1316 1108 1324
rect 1244 1336 1252 1344
rect 1308 1336 1316 1344
rect 1372 1336 1380 1344
rect 1404 1336 1412 1344
rect 1500 1336 1508 1344
rect 1564 1336 1572 1344
rect 1612 1336 1620 1344
rect 1676 1336 1684 1344
rect 1724 1336 1732 1344
rect 1836 1336 1844 1344
rect 1964 1336 1972 1344
rect 2108 1336 2116 1344
rect 2124 1336 2132 1344
rect 2220 1336 2228 1344
rect 2332 1336 2340 1344
rect 2412 1336 2420 1344
rect 2492 1332 2500 1340
rect 2508 1336 2516 1344
rect 2524 1336 2532 1344
rect 2556 1336 2564 1344
rect 2636 1336 2644 1344
rect 2764 1356 2772 1364
rect 2924 1356 2932 1364
rect 3052 1356 3060 1364
rect 3084 1356 3092 1364
rect 3996 1356 4004 1364
rect 4140 1356 4148 1364
rect 4332 1356 4340 1364
rect 4892 1356 4900 1364
rect 5228 1356 5236 1364
rect 5292 1356 5300 1364
rect 5932 1356 5940 1364
rect 6060 1356 6068 1364
rect 6284 1356 6292 1364
rect 6348 1356 6356 1364
rect 6444 1356 6452 1364
rect 6620 1356 6628 1364
rect 6780 1356 6788 1364
rect 6796 1356 6804 1364
rect 2700 1336 2708 1344
rect 2732 1336 2740 1344
rect 2780 1336 2788 1344
rect 2812 1336 2820 1344
rect 2908 1336 2916 1344
rect 2924 1336 2932 1344
rect 3068 1336 3076 1344
rect 3148 1336 3156 1344
rect 3164 1336 3172 1344
rect 3260 1336 3268 1344
rect 3308 1336 3316 1344
rect 3356 1336 3364 1344
rect 3372 1336 3380 1344
rect 3468 1336 3476 1344
rect 3548 1336 3556 1344
rect 3644 1336 3652 1344
rect 3836 1336 3844 1344
rect 3916 1336 3924 1344
rect 3932 1336 3940 1344
rect 4556 1336 4564 1344
rect 4588 1336 4596 1344
rect 4620 1336 4628 1344
rect 4732 1336 4740 1344
rect 4956 1336 4964 1344
rect 4988 1336 4996 1344
rect 5036 1336 5044 1344
rect 5084 1336 5092 1344
rect 5212 1336 5220 1344
rect 5340 1336 5348 1344
rect 5388 1336 5396 1344
rect 5436 1336 5444 1344
rect 5452 1336 5460 1344
rect 5484 1336 5492 1344
rect 5596 1336 5604 1344
rect 5628 1336 5636 1344
rect 5868 1336 5876 1344
rect 1228 1316 1236 1324
rect 1292 1316 1300 1324
rect 1420 1316 1428 1324
rect 1516 1316 1524 1324
rect 1548 1316 1556 1324
rect 1580 1316 1588 1324
rect 1660 1316 1668 1324
rect 1756 1316 1764 1324
rect 1788 1316 1796 1324
rect 1868 1316 1876 1324
rect 1900 1316 1908 1324
rect 1980 1316 1988 1324
rect 2044 1316 2052 1324
rect 2252 1316 2260 1324
rect 2444 1316 2452 1324
rect 2620 1316 2628 1324
rect 2652 1316 2660 1324
rect 2716 1316 2724 1324
rect 2796 1316 2804 1324
rect 3036 1316 3044 1324
rect 3084 1316 3092 1324
rect 3148 1316 3156 1324
rect 3324 1316 3332 1324
rect 3612 1318 3620 1326
rect 3804 1318 3812 1326
rect 3900 1316 3908 1324
rect 4092 1316 4100 1324
rect 4284 1316 4292 1324
rect 4428 1316 4436 1324
rect 4604 1316 4612 1324
rect 4652 1316 4660 1324
rect 4780 1316 4788 1324
rect 4844 1316 4852 1324
rect 4908 1316 4916 1324
rect 5532 1316 5540 1324
rect 5692 1318 5700 1326
rect 5756 1316 5764 1324
rect 6108 1336 6116 1344
rect 6172 1336 6180 1344
rect 6428 1336 6436 1344
rect 6476 1336 6484 1344
rect 6540 1336 6548 1344
rect 6588 1336 6596 1344
rect 6652 1336 6660 1344
rect 6668 1336 6676 1344
rect 6732 1336 6740 1344
rect 6876 1336 6884 1344
rect 7292 1336 7300 1344
rect 7356 1336 7364 1344
rect 924 1296 932 1304
rect 1084 1296 1092 1304
rect 1148 1296 1156 1304
rect 1756 1296 1764 1304
rect 1772 1296 1780 1304
rect 1868 1296 1876 1304
rect 1884 1296 1892 1304
rect 1980 1296 1988 1304
rect 2044 1296 2052 1304
rect 2076 1296 2084 1304
rect 2236 1296 2244 1304
rect 2300 1296 2308 1304
rect 2380 1296 2388 1304
rect 2748 1296 2756 1304
rect 2860 1296 2868 1304
rect 3100 1296 3108 1304
rect 3276 1296 3284 1304
rect 3868 1296 3876 1304
rect 4444 1296 4452 1304
rect 12 1276 20 1284
rect 1116 1276 1124 1284
rect 1804 1276 1812 1284
rect 1916 1276 1924 1284
rect 1996 1276 2004 1284
rect 2028 1276 2036 1284
rect 2060 1276 2068 1284
rect 2268 1276 2276 1284
rect 2444 1276 2452 1284
rect 2636 1276 2644 1284
rect 3228 1276 3236 1284
rect 4012 1276 4020 1284
rect 4412 1276 4420 1284
rect 4572 1296 4580 1304
rect 4636 1296 4644 1304
rect 4796 1296 4804 1304
rect 4956 1296 4964 1304
rect 5004 1296 5012 1304
rect 5052 1296 5060 1304
rect 5180 1296 5188 1304
rect 5276 1296 5284 1304
rect 5484 1296 5492 1304
rect 5836 1296 5844 1304
rect 5916 1296 5924 1304
rect 6252 1316 6260 1324
rect 6300 1316 6308 1324
rect 6380 1316 6388 1324
rect 6396 1316 6404 1324
rect 6412 1316 6420 1324
rect 6540 1316 6548 1324
rect 6604 1316 6612 1324
rect 6668 1316 6676 1324
rect 6684 1316 6692 1324
rect 6748 1316 6756 1324
rect 6844 1316 6852 1324
rect 6876 1316 6884 1324
rect 6892 1316 6900 1324
rect 6956 1316 6964 1324
rect 7020 1316 7028 1324
rect 7132 1316 7140 1324
rect 7164 1316 7172 1324
rect 7340 1316 7348 1324
rect 6156 1296 6164 1304
rect 6380 1296 6388 1304
rect 6524 1296 6532 1304
rect 6924 1296 6932 1304
rect 7004 1296 7012 1304
rect 7260 1296 7268 1304
rect 7308 1296 7316 1304
rect 2252 1256 2260 1264
rect 4668 1276 4676 1284
rect 4764 1276 4772 1284
rect 4828 1276 4836 1284
rect 5308 1276 5316 1284
rect 5356 1276 5364 1284
rect 5388 1276 5396 1284
rect 5596 1276 5604 1284
rect 6204 1276 6212 1284
rect 6588 1276 6596 1284
rect 6780 1276 6788 1284
rect 7036 1276 7044 1284
rect 5148 1256 5156 1264
rect 7020 1256 7028 1264
rect 460 1236 468 1244
rect 540 1236 548 1244
rect 1132 1236 1140 1244
rect 1372 1236 1380 1244
rect 1516 1236 1524 1244
rect 1820 1236 1828 1244
rect 2012 1236 2020 1244
rect 2876 1236 2884 1244
rect 3484 1236 3492 1244
rect 3676 1236 3684 1244
rect 4204 1236 4212 1244
rect 5116 1236 5124 1244
rect 6028 1236 6036 1244
rect 6268 1236 6276 1244
rect 6812 1236 6820 1244
rect 7068 1236 7076 1244
rect 1411 1206 1419 1214
rect 1421 1206 1429 1214
rect 1431 1206 1439 1214
rect 1441 1206 1449 1214
rect 1451 1206 1459 1214
rect 1461 1206 1469 1214
rect 4419 1206 4427 1214
rect 4429 1206 4437 1214
rect 4439 1206 4447 1214
rect 4449 1206 4457 1214
rect 4459 1206 4467 1214
rect 4469 1206 4477 1214
rect 268 1176 276 1184
rect 764 1176 772 1184
rect 860 1176 868 1184
rect 1756 1176 1764 1184
rect 2364 1176 2372 1184
rect 3132 1176 3140 1184
rect 3500 1176 3508 1184
rect 3532 1176 3540 1184
rect 3548 1176 3556 1184
rect 3596 1176 3604 1184
rect 3772 1176 3780 1184
rect 4012 1176 4020 1184
rect 4140 1176 4148 1184
rect 4220 1176 4228 1184
rect 4396 1176 4404 1184
rect 4556 1176 4564 1184
rect 4844 1176 4852 1184
rect 4876 1176 4884 1184
rect 5196 1176 5204 1184
rect 5308 1176 5316 1184
rect 5852 1176 5860 1184
rect 6204 1176 6212 1184
rect 6476 1176 6484 1184
rect 6604 1176 6612 1184
rect 6860 1176 6868 1184
rect 988 1156 996 1164
rect 1836 1156 1844 1164
rect 2348 1156 2356 1164
rect 4748 1156 4756 1164
rect 6540 1156 6548 1164
rect 972 1136 980 1144
rect 1132 1136 1140 1144
rect 2636 1136 2644 1144
rect 2860 1136 2868 1144
rect 4060 1136 4068 1144
rect 4092 1136 4100 1144
rect 4156 1136 4164 1144
rect 4236 1136 4244 1144
rect 4348 1136 4356 1144
rect 4412 1136 4420 1144
rect 4428 1136 4436 1144
rect 4572 1136 4580 1144
rect 4668 1136 4676 1144
rect 4732 1136 4740 1144
rect 6268 1136 6276 1144
rect 6524 1136 6532 1144
rect 6588 1136 6596 1144
rect 7276 1136 7284 1144
rect 236 1116 244 1124
rect 476 1116 484 1124
rect 540 1116 548 1124
rect 924 1116 932 1124
rect 1004 1116 1012 1124
rect 1340 1116 1348 1124
rect 1372 1116 1380 1124
rect 12 1096 20 1104
rect 108 1096 116 1104
rect 220 1096 228 1104
rect 268 1096 276 1104
rect 300 1096 308 1104
rect 348 1096 356 1104
rect 444 1096 452 1104
rect 476 1096 484 1104
rect 588 1096 596 1104
rect 604 1096 612 1104
rect 636 1096 644 1104
rect 668 1096 676 1104
rect 716 1096 724 1104
rect 844 1096 852 1104
rect 876 1096 884 1104
rect 908 1096 916 1104
rect 940 1096 948 1104
rect 988 1096 996 1104
rect 1084 1096 1092 1104
rect 1164 1096 1172 1104
rect 1292 1096 1300 1104
rect 1692 1116 1700 1124
rect 1724 1116 1732 1124
rect 1900 1116 1908 1124
rect 2236 1114 2244 1122
rect 2476 1116 2484 1124
rect 2668 1116 2676 1124
rect 2812 1116 2820 1124
rect 3308 1116 3316 1124
rect 3420 1116 3428 1124
rect 3708 1116 3716 1124
rect 3996 1116 4004 1124
rect 4028 1116 4036 1124
rect 4380 1116 4388 1124
rect 4492 1116 4500 1124
rect 4652 1116 4660 1124
rect 4764 1116 4772 1124
rect 5084 1116 5092 1124
rect 5100 1116 5108 1124
rect 1532 1096 1540 1104
rect 1676 1096 1684 1104
rect 1756 1096 1764 1104
rect 1788 1096 1796 1104
rect 1852 1096 1860 1104
rect 1932 1096 1940 1104
rect 2044 1096 2052 1104
rect 2092 1096 2100 1104
rect 2156 1096 2164 1104
rect 2204 1096 2212 1104
rect 2316 1096 2324 1104
rect 2396 1096 2404 1104
rect 2412 1096 2420 1104
rect 2476 1096 2484 1104
rect 2492 1096 2500 1104
rect 2524 1096 2532 1104
rect 2668 1096 2676 1104
rect 2748 1096 2756 1104
rect 2764 1096 2772 1104
rect 2956 1096 2964 1104
rect 3036 1096 3044 1104
rect 3100 1096 3108 1104
rect 3148 1096 3156 1104
rect 3228 1096 3236 1104
rect 284 1076 292 1084
rect 396 1076 404 1084
rect 492 1076 500 1084
rect 508 1076 516 1084
rect 556 1076 564 1084
rect 620 1076 628 1084
rect 716 1076 724 1084
rect 732 1076 740 1084
rect 764 1076 772 1084
rect 892 1076 900 1084
rect 924 1076 932 1084
rect 1052 1076 1060 1084
rect 1228 1076 1236 1084
rect 1340 1076 1348 1084
rect 1484 1076 1492 1084
rect 108 1056 116 1064
rect 396 1056 404 1064
rect 652 1056 660 1064
rect 700 1056 708 1064
rect 796 1056 804 1064
rect 844 1056 852 1064
rect 1068 1056 1076 1064
rect 1132 1056 1140 1064
rect 1260 1056 1268 1064
rect 1388 1056 1396 1064
rect 1532 1056 1540 1064
rect 1564 1056 1572 1064
rect 1596 1076 1604 1084
rect 1612 1076 1620 1084
rect 1772 1076 1780 1084
rect 1804 1076 1812 1084
rect 1836 1076 1844 1084
rect 1868 1076 1876 1084
rect 1900 1076 1908 1084
rect 3452 1096 3460 1104
rect 3468 1096 3476 1104
rect 3580 1096 3588 1104
rect 3628 1096 3636 1104
rect 3756 1096 3764 1104
rect 3900 1094 3908 1102
rect 4044 1096 4052 1104
rect 4140 1096 4148 1104
rect 4220 1096 4228 1104
rect 4316 1096 4324 1104
rect 4332 1096 4340 1104
rect 4364 1096 4372 1104
rect 4428 1096 4436 1104
rect 4588 1096 4596 1104
rect 4668 1096 4676 1104
rect 4700 1096 4708 1104
rect 4748 1096 4756 1104
rect 4780 1096 4788 1104
rect 4908 1096 4916 1104
rect 5004 1096 5012 1104
rect 5132 1096 5140 1104
rect 5164 1096 5172 1104
rect 5372 1096 5380 1104
rect 5436 1096 5444 1104
rect 5484 1116 5492 1124
rect 5532 1116 5540 1124
rect 5612 1116 5620 1124
rect 5628 1116 5636 1124
rect 5724 1116 5732 1124
rect 5772 1116 5780 1124
rect 5868 1116 5876 1124
rect 6300 1116 6308 1124
rect 6428 1116 6436 1124
rect 6444 1116 6452 1124
rect 6556 1116 6564 1124
rect 6620 1116 6628 1124
rect 6636 1116 6644 1124
rect 6828 1116 6836 1124
rect 6892 1116 6900 1124
rect 7356 1116 7364 1124
rect 5580 1096 5588 1104
rect 5852 1096 5860 1104
rect 6108 1094 6116 1102
rect 6172 1096 6180 1104
rect 6220 1096 6228 1104
rect 6300 1096 6308 1104
rect 6476 1096 6484 1104
rect 6540 1096 6548 1104
rect 6604 1096 6612 1104
rect 6700 1096 6708 1104
rect 6764 1096 6772 1104
rect 6972 1096 6980 1104
rect 7004 1096 7012 1104
rect 7164 1096 7172 1104
rect 7340 1096 7348 1104
rect 1948 1076 1956 1084
rect 1996 1076 2004 1084
rect 2028 1076 2036 1084
rect 2092 1076 2100 1084
rect 2188 1076 2196 1084
rect 2428 1076 2436 1084
rect 1644 1056 1652 1064
rect 1708 1056 1716 1064
rect 1932 1056 1940 1064
rect 1948 1056 1956 1064
rect 1996 1056 2004 1064
rect 2060 1056 2068 1064
rect 2108 1056 2116 1064
rect 2204 1056 2212 1064
rect 2252 1056 2260 1064
rect 2300 1056 2308 1064
rect 2460 1056 2468 1064
rect 2588 1076 2596 1084
rect 2636 1076 2644 1084
rect 2732 1076 2740 1084
rect 2748 1076 2756 1084
rect 2844 1076 2852 1084
rect 2972 1076 2980 1084
rect 3084 1076 3092 1084
rect 2572 1056 2580 1064
rect 2796 1056 2804 1064
rect 3036 1056 3044 1064
rect 3196 1056 3204 1064
rect 3244 1056 3252 1064
rect 3276 1076 3284 1084
rect 3324 1076 3332 1084
rect 3372 1076 3380 1084
rect 3388 1076 3396 1084
rect 3660 1076 3668 1084
rect 3692 1076 3700 1084
rect 3724 1076 3732 1084
rect 3756 1076 3764 1084
rect 4892 1076 4900 1084
rect 4972 1076 4980 1084
rect 5052 1076 5060 1084
rect 5132 1076 5140 1084
rect 5148 1076 5156 1084
rect 5292 1076 5300 1084
rect 5356 1076 5364 1084
rect 5420 1076 5428 1084
rect 5516 1076 5524 1084
rect 5564 1076 5572 1084
rect 5676 1076 5684 1084
rect 5772 1076 5780 1084
rect 5804 1076 5812 1084
rect 5900 1076 5908 1084
rect 6092 1076 6100 1084
rect 6236 1076 6244 1084
rect 6284 1076 6292 1084
rect 6348 1076 6356 1084
rect 6396 1076 6404 1084
rect 6492 1076 6500 1084
rect 6636 1076 6644 1084
rect 6684 1076 6692 1084
rect 6780 1076 6788 1084
rect 6876 1076 6884 1084
rect 6940 1076 6948 1084
rect 6988 1076 6996 1084
rect 7020 1076 7028 1084
rect 7100 1076 7108 1084
rect 7132 1076 7140 1084
rect 7308 1076 7316 1084
rect 3324 1056 3332 1064
rect 3436 1056 3444 1064
rect 3516 1056 3524 1064
rect 3644 1056 3652 1064
rect 3836 1056 3844 1064
rect 3900 1056 3908 1064
rect 3964 1056 3972 1064
rect 3996 1056 4004 1064
rect 4092 1056 4100 1064
rect 4268 1056 4276 1064
rect 4540 1056 4548 1064
rect 4636 1056 4644 1064
rect 4828 1056 4836 1064
rect 5212 1056 5220 1064
rect 5276 1056 5284 1064
rect 5340 1056 5348 1064
rect 5468 1056 5476 1064
rect 5708 1056 5716 1064
rect 5820 1056 5828 1064
rect 5852 1056 5860 1064
rect 6380 1056 6388 1064
rect 6812 1056 6820 1064
rect 7004 1056 7012 1064
rect 7228 1056 7236 1064
rect 7276 1056 7284 1064
rect 44 1036 52 1044
rect 60 1036 68 1044
rect 124 1036 132 1044
rect 156 1036 164 1044
rect 188 1036 196 1044
rect 332 1036 340 1044
rect 540 1036 548 1044
rect 1020 1036 1028 1044
rect 1196 1036 1204 1044
rect 1324 1036 1332 1044
rect 1372 1036 1380 1044
rect 1468 1036 1476 1044
rect 1900 1036 1908 1044
rect 2076 1036 2084 1044
rect 2700 1036 2708 1044
rect 2828 1036 2836 1044
rect 3004 1036 3012 1044
rect 3340 1036 3348 1044
rect 3420 1036 3428 1044
rect 4284 1036 4292 1044
rect 4812 1036 4820 1044
rect 4940 1036 4948 1044
rect 5084 1036 5092 1044
rect 5260 1036 5268 1044
rect 5612 1036 5620 1044
rect 5628 1036 5636 1044
rect 5740 1036 5748 1044
rect 5788 1036 5796 1044
rect 5868 1036 5876 1044
rect 5980 1036 5988 1044
rect 6300 1036 6308 1044
rect 6428 1036 6436 1044
rect 6780 1036 6788 1044
rect 2915 1006 2923 1014
rect 2925 1006 2933 1014
rect 2935 1006 2943 1014
rect 2945 1006 2953 1014
rect 2955 1006 2963 1014
rect 2965 1006 2973 1014
rect 5923 1006 5931 1014
rect 5933 1006 5941 1014
rect 5943 1006 5951 1014
rect 5953 1006 5961 1014
rect 5963 1006 5971 1014
rect 5973 1006 5981 1014
rect 2364 996 2372 1004
rect 2524 996 2532 1004
rect 172 976 180 984
rect 380 976 388 984
rect 476 976 484 984
rect 556 976 564 984
rect 668 976 676 984
rect 956 976 964 984
rect 1036 976 1044 984
rect 1564 976 1572 984
rect 60 956 68 964
rect 124 956 132 964
rect 156 936 164 944
rect 204 956 212 964
rect 332 956 340 964
rect 460 956 468 964
rect 492 956 500 964
rect 508 956 516 964
rect 636 956 644 964
rect 652 956 660 964
rect 684 956 692 964
rect 764 956 772 964
rect 876 956 884 964
rect 908 956 916 964
rect 940 956 948 964
rect 972 956 980 964
rect 1004 956 1012 964
rect 1020 956 1028 964
rect 1100 956 1108 964
rect 1196 956 1204 964
rect 1212 956 1220 964
rect 1276 956 1284 964
rect 268 936 276 944
rect 300 936 308 944
rect 44 916 52 924
rect 92 916 100 924
rect 236 916 244 924
rect 412 936 420 944
rect 556 936 564 944
rect 588 936 596 944
rect 716 936 724 944
rect 812 936 820 944
rect 844 936 852 944
rect 860 936 868 944
rect 1052 936 1060 944
rect 1244 936 1252 944
rect 1292 936 1300 944
rect 1388 956 1396 964
rect 1596 956 1604 964
rect 1788 956 1796 964
rect 1804 956 1812 964
rect 1900 956 1908 964
rect 2172 976 2180 984
rect 2220 976 2228 984
rect 2316 976 2324 984
rect 2476 976 2484 984
rect 2556 976 2564 984
rect 2812 976 2820 984
rect 2924 976 2932 984
rect 3276 976 3284 984
rect 3340 976 3348 984
rect 3404 976 3412 984
rect 3660 976 3668 984
rect 3932 976 3940 984
rect 4108 976 4116 984
rect 4156 976 4164 984
rect 4492 976 4500 984
rect 4812 976 4820 984
rect 4908 976 4916 984
rect 5068 976 5076 984
rect 5132 976 5140 984
rect 5372 976 5380 984
rect 5484 976 5492 984
rect 5756 976 5764 984
rect 6124 976 6132 984
rect 6396 976 6404 984
rect 6972 976 6980 984
rect 7148 976 7156 984
rect 7196 976 7204 984
rect 2044 956 2052 964
rect 2156 956 2164 964
rect 2364 956 2372 964
rect 2492 956 2500 964
rect 2524 956 2532 964
rect 2620 956 2628 964
rect 2764 956 2772 964
rect 2796 956 2804 964
rect 1484 936 1492 944
rect 1500 936 1508 944
rect 1580 936 1588 944
rect 1628 936 1636 944
rect 1708 936 1716 944
rect 1740 936 1748 944
rect 1916 936 1924 944
rect 2060 936 2068 944
rect 2188 936 2196 944
rect 2252 932 2260 940
rect 2268 936 2276 944
rect 2444 936 2452 944
rect 364 916 372 924
rect 428 916 436 924
rect 684 916 692 924
rect 780 916 788 924
rect 796 916 804 924
rect 860 916 868 924
rect 1148 916 1156 924
rect 1308 916 1316 924
rect 1356 916 1364 924
rect 1532 916 1540 924
rect 1564 916 1572 924
rect 1628 916 1636 924
rect 1676 916 1684 924
rect 1724 916 1732 924
rect 1756 916 1764 924
rect 1852 916 1860 924
rect 1868 916 1876 924
rect 1932 916 1940 924
rect 1964 916 1972 924
rect 2076 916 2084 924
rect 2204 916 2212 924
rect 2316 916 2324 924
rect 2396 916 2404 924
rect 2428 916 2436 924
rect 2444 916 2452 924
rect 2556 916 2564 924
rect 2588 916 2596 924
rect 2716 936 2724 944
rect 2860 936 2868 944
rect 3036 936 3044 944
rect 3068 936 3076 944
rect 3116 956 3124 964
rect 3228 956 3236 964
rect 3372 956 3380 964
rect 3532 956 3540 964
rect 3644 956 3652 964
rect 4092 956 4100 964
rect 4140 956 4148 964
rect 4572 956 4580 964
rect 5228 956 5236 964
rect 5276 956 5284 964
rect 3148 936 3156 944
rect 3196 936 3204 944
rect 3356 936 3364 944
rect 3436 936 3444 944
rect 3500 936 3508 944
rect 3548 936 3556 944
rect 3740 936 3748 944
rect 3772 936 3780 944
rect 3836 936 3844 944
rect 3900 936 3908 944
rect 3980 936 3988 944
rect 4028 936 4036 944
rect 4076 936 4084 944
rect 4172 936 4180 944
rect 4204 936 4212 944
rect 4300 936 4308 944
rect 4380 936 4388 944
rect 4604 936 4612 944
rect 4668 936 4676 944
rect 4844 936 4852 944
rect 4940 936 4948 944
rect 5036 936 5044 944
rect 5100 936 5108 944
rect 5196 936 5204 944
rect 5548 956 5556 964
rect 5644 956 5652 964
rect 5692 956 5700 964
rect 5852 956 5860 964
rect 6140 956 6148 964
rect 6284 956 6292 964
rect 6380 956 6388 964
rect 6588 956 6596 964
rect 6652 956 6660 964
rect 6956 956 6964 964
rect 7036 956 7044 964
rect 7132 956 7140 964
rect 7324 956 7332 964
rect 7356 956 7364 964
rect 5356 936 5364 944
rect 5420 936 5428 944
rect 5436 936 5444 944
rect 5580 936 5588 944
rect 5644 936 5652 944
rect 5692 936 5700 944
rect 5772 936 5780 944
rect 5820 936 5828 944
rect 5884 936 5892 944
rect 5916 936 5924 944
rect 5932 936 5940 944
rect 6076 936 6084 944
rect 6108 936 6116 944
rect 6156 936 6164 944
rect 6204 936 6212 944
rect 6252 936 6260 944
rect 6348 936 6356 944
rect 6620 936 6628 944
rect 6732 936 6740 944
rect 6876 936 6884 944
rect 6924 936 6932 944
rect 6988 936 6996 944
rect 7036 936 7044 944
rect 7068 936 7076 944
rect 7164 936 7172 944
rect 7244 936 7252 944
rect 7260 936 7268 944
rect 7276 932 7284 940
rect 2620 916 2628 924
rect 2652 916 2660 924
rect 2716 916 2724 924
rect 2796 916 2804 924
rect 2844 916 2852 924
rect 2908 916 2916 924
rect 3020 916 3028 924
rect 3052 916 3060 924
rect 3084 916 3092 924
rect 3148 916 3156 924
rect 300 896 308 904
rect 380 896 388 904
rect 1468 896 1476 904
rect 1692 896 1700 904
rect 1772 896 1780 904
rect 2332 896 2340 904
rect 2428 896 2436 904
rect 2620 896 2628 904
rect 2684 896 2692 904
rect 2940 896 2948 904
rect 3196 916 3204 924
rect 3244 916 3252 924
rect 3308 916 3316 924
rect 3340 916 3348 924
rect 3500 916 3508 924
rect 3708 916 3716 924
rect 3756 916 3764 924
rect 3820 916 3828 924
rect 3884 916 3892 924
rect 3932 916 3940 924
rect 4092 916 4100 924
rect 4124 916 4132 924
rect 4284 916 4292 924
rect 4396 916 4404 924
rect 4524 916 4532 924
rect 4716 916 4724 924
rect 4764 916 4772 924
rect 4892 916 4900 924
rect 4956 916 4964 924
rect 5164 916 5172 924
rect 5244 916 5252 924
rect 5404 916 5412 924
rect 5452 916 5460 924
rect 5532 916 5540 924
rect 5660 916 5668 924
rect 5724 916 5732 924
rect 5772 916 5780 924
rect 5820 916 5828 924
rect 5868 916 5876 924
rect 5932 916 5940 924
rect 6012 916 6020 924
rect 6076 916 6084 924
rect 6092 916 6100 924
rect 6188 916 6196 924
rect 6204 916 6212 924
rect 6316 916 6324 924
rect 6460 916 6468 924
rect 6524 918 6532 926
rect 6636 916 6644 924
rect 6700 916 6708 924
rect 6716 916 6724 924
rect 6764 916 6772 924
rect 6828 916 6836 924
rect 6876 916 6884 924
rect 6940 916 6948 924
rect 6988 916 6996 924
rect 7052 916 7060 924
rect 7084 916 7092 924
rect 7196 916 7204 924
rect 7228 916 7236 924
rect 7324 916 7332 924
rect 3372 896 3380 904
rect 3436 896 3444 904
rect 3596 898 3604 906
rect 3724 896 3732 904
rect 3788 896 3796 904
rect 3852 896 3860 904
rect 3916 896 3924 904
rect 3980 896 3988 904
rect 4044 896 4052 904
rect 4236 896 4244 904
rect 4252 896 4260 904
rect 4284 896 4292 904
rect 4636 896 4644 904
rect 4732 896 4740 904
rect 4908 896 4916 904
rect 5004 896 5012 904
rect 5020 896 5028 904
rect 5132 896 5140 904
rect 5148 896 5156 904
rect 5260 896 5268 904
rect 5308 896 5316 904
rect 5324 896 5332 904
rect 5628 896 5636 904
rect 5756 896 5764 904
rect 5820 896 5828 904
rect 6060 896 6068 904
rect 6156 896 6164 904
rect 6268 896 6276 904
rect 6300 896 6308 904
rect 6588 896 6596 904
rect 6764 896 6772 904
rect 6828 896 6836 904
rect 7084 896 7092 904
rect 7116 896 7124 904
rect 7196 896 7204 904
rect 12 876 20 884
rect 764 876 772 884
rect 812 876 820 884
rect 972 876 980 884
rect 1100 876 1108 884
rect 1356 876 1364 884
rect 2332 876 2340 884
rect 3916 876 3924 884
rect 4700 876 4708 884
rect 1932 856 1940 864
rect 3820 856 3828 864
rect 4764 876 4772 884
rect 4780 876 4788 884
rect 5100 876 5108 884
rect 6780 876 6788 884
rect 6844 876 6852 884
rect 6860 876 6868 884
rect 6924 876 6932 884
rect 4860 856 4868 864
rect 6764 856 6772 864
rect 1196 836 1204 844
rect 1644 836 1652 844
rect 1804 836 1812 844
rect 2124 836 2132 844
rect 3484 836 3492 844
rect 3676 836 3684 844
rect 3884 836 3892 844
rect 4988 836 4996 844
rect 5500 836 5508 844
rect 5676 836 5684 844
rect 5916 836 5924 844
rect 7308 836 7316 844
rect 1411 806 1419 814
rect 1421 806 1429 814
rect 1431 806 1439 814
rect 1441 806 1449 814
rect 1451 806 1459 814
rect 1461 806 1469 814
rect 4419 806 4427 814
rect 4429 806 4437 814
rect 4439 806 4447 814
rect 4449 806 4457 814
rect 4459 806 4467 814
rect 4469 806 4477 814
rect 316 776 324 784
rect 684 776 692 784
rect 812 776 820 784
rect 1516 776 1524 784
rect 1756 776 1764 784
rect 1948 776 1956 784
rect 1996 776 2004 784
rect 2348 776 2356 784
rect 2460 776 2468 784
rect 2700 776 2708 784
rect 2812 776 2820 784
rect 2892 776 2900 784
rect 3404 776 3412 784
rect 3548 776 3556 784
rect 3692 776 3700 784
rect 4492 776 4500 784
rect 4636 776 4644 784
rect 4700 776 4708 784
rect 4796 776 4804 784
rect 5244 776 5252 784
rect 5324 776 5332 784
rect 5372 776 5380 784
rect 5788 776 5796 784
rect 6092 776 6100 784
rect 6172 776 6180 784
rect 6812 776 6820 784
rect 6908 776 6916 784
rect 7212 776 7220 784
rect 7356 776 7364 784
rect 2316 756 2324 764
rect 5580 756 5588 764
rect 6364 756 6372 764
rect 652 736 660 744
rect 1132 736 1140 744
rect 1148 736 1156 744
rect 1260 736 1268 744
rect 1500 736 1508 744
rect 2092 736 2100 744
rect 2428 736 2436 744
rect 2636 736 2644 744
rect 2684 736 2692 744
rect 2716 736 2724 744
rect 3484 736 3492 744
rect 4140 736 4148 744
rect 4716 736 4724 744
rect 4812 736 4820 744
rect 5228 736 5236 744
rect 6076 736 6084 744
rect 7228 736 7236 744
rect 7276 736 7284 744
rect 284 716 292 724
rect 460 716 468 724
rect 492 716 500 724
rect 636 716 644 724
rect 1084 716 1092 724
rect 1452 716 1460 724
rect 1532 716 1540 724
rect 1692 716 1700 724
rect 1788 716 1796 724
rect 2124 716 2132 724
rect 44 696 52 704
rect 316 696 324 704
rect 396 696 404 704
rect 412 696 420 704
rect 428 696 436 704
rect 540 696 548 704
rect 620 696 628 704
rect 668 696 676 704
rect 732 696 740 704
rect 748 696 756 704
rect 844 696 852 704
rect 892 696 900 704
rect 924 696 932 704
rect 1004 696 1012 704
rect 1036 696 1044 704
rect 1116 696 1124 704
rect 1164 696 1172 704
rect 1244 696 1252 704
rect 1372 696 1380 704
rect 1468 696 1476 704
rect 1516 696 1524 704
rect 1660 696 1668 704
rect 1708 696 1716 704
rect 1756 696 1764 704
rect 1852 696 1860 704
rect 1884 696 1892 704
rect 1980 696 1988 704
rect 2012 696 2020 704
rect 2060 696 2068 704
rect 2108 696 2116 704
rect 2140 696 2148 704
rect 2172 696 2180 704
rect 2204 696 2212 704
rect 2284 696 2292 704
rect 2316 696 2324 704
rect 2684 716 2692 724
rect 2828 716 2836 724
rect 3020 716 3028 724
rect 3372 716 3380 724
rect 3916 716 3924 724
rect 3996 716 4004 724
rect 4044 716 4052 724
rect 4092 716 4100 724
rect 4172 716 4180 724
rect 4252 716 4260 724
rect 4844 716 4852 724
rect 4876 716 4884 724
rect 5004 716 5012 724
rect 5452 716 5460 724
rect 5484 716 5492 724
rect 5548 716 5556 724
rect 5564 716 5572 724
rect 5644 716 5652 724
rect 5708 716 5716 724
rect 5756 716 5764 724
rect 5772 716 5780 724
rect 5804 716 5812 724
rect 6108 716 6116 724
rect 6124 716 6132 724
rect 6492 716 6500 724
rect 6572 716 6580 724
rect 6956 716 6964 724
rect 7148 714 7156 722
rect 7196 716 7204 724
rect 2396 696 2404 704
rect 2428 696 2436 704
rect 2460 696 2468 704
rect 2572 696 2580 704
rect 2588 696 2596 704
rect 2700 696 2708 704
rect 2796 696 2804 704
rect 2876 696 2884 704
rect 2940 696 2948 704
rect 3100 696 3108 704
rect 3148 696 3156 704
rect 3196 696 3204 704
rect 3212 696 3220 704
rect 3244 696 3252 704
rect 3356 696 3364 704
rect 3404 696 3412 704
rect 3436 696 3444 704
rect 3516 696 3524 704
rect 3644 696 3652 704
rect 3820 694 3828 702
rect 3916 696 3924 704
rect 4172 696 4180 704
rect 4236 696 4244 704
rect 4348 694 4356 702
rect 4412 696 4420 704
rect 4604 696 4612 704
rect 4700 696 4708 704
rect 4796 696 4804 704
rect 4844 696 4852 704
rect 4956 696 4964 704
rect 5100 694 5108 702
rect 5292 696 5300 704
rect 5436 696 5444 704
rect 5516 696 5524 704
rect 5676 696 5684 704
rect 5852 696 5860 704
rect 5916 696 5924 704
rect 6012 696 6020 704
rect 6044 696 6052 704
rect 6092 696 6100 704
rect 6236 696 6244 704
rect 6284 696 6292 704
rect 6380 696 6388 704
rect 6444 696 6452 704
rect 6508 696 6516 704
rect 6524 696 6532 704
rect 6700 696 6708 704
rect 6812 696 6820 704
rect 6860 696 6868 704
rect 6924 696 6932 704
rect 6988 696 6996 704
rect 7068 696 7076 704
rect 7116 696 7124 704
rect 7212 696 7220 704
rect 7276 696 7284 704
rect 12 676 20 684
rect 108 676 116 684
rect 332 676 340 684
rect 380 676 388 684
rect 444 676 452 684
rect 556 676 564 684
rect 620 676 628 684
rect 956 676 964 684
rect 1292 676 1300 684
rect 2188 676 2196 684
rect 2204 676 2212 684
rect 2380 676 2388 684
rect 2444 676 2452 684
rect 2540 676 2548 684
rect 2604 676 2612 684
rect 2796 676 2804 684
rect 3052 676 3060 684
rect 3228 676 3236 684
rect 3260 676 3268 684
rect 3308 676 3316 684
rect 3420 676 3428 684
rect 3452 676 3460 684
rect 3852 676 3860 684
rect 3884 676 3892 684
rect 3964 676 3972 684
rect 4028 676 4036 684
rect 4044 676 4052 684
rect 4076 676 4084 684
rect 4124 676 4132 684
rect 4140 676 4148 684
rect 4284 676 4292 684
rect 4380 676 4388 684
rect 4588 676 4596 684
rect 4876 676 4884 684
rect 4924 676 4932 684
rect 4972 676 4980 684
rect 5036 676 5044 684
rect 5068 676 5076 684
rect 5276 676 5284 684
rect 5500 676 5508 684
rect 5596 676 5604 684
rect 5612 676 5620 684
rect 5660 676 5668 684
rect 5724 676 5732 684
rect 5804 676 5812 684
rect 5868 676 5876 684
rect 5884 676 5892 684
rect 6028 676 6036 684
rect 6156 676 6164 684
rect 6460 676 6468 684
rect 6492 676 6500 684
rect 6540 676 6548 684
rect 6716 676 6724 684
rect 6972 676 6980 684
rect 7036 676 7044 684
rect 7100 676 7108 684
rect 7260 676 7268 684
rect 7324 676 7332 684
rect 124 656 132 664
rect 188 656 196 664
rect 204 656 212 664
rect 268 656 276 664
rect 364 656 372 664
rect 556 656 564 664
rect 796 656 804 664
rect 76 636 84 644
rect 140 636 148 644
rect 252 636 260 644
rect 508 636 516 644
rect 700 636 708 644
rect 780 636 788 644
rect 892 656 900 664
rect 956 656 964 664
rect 1340 656 1348 664
rect 1548 656 1556 664
rect 1580 656 1588 664
rect 1612 656 1620 664
rect 1708 656 1716 664
rect 1804 656 1812 664
rect 1884 656 1892 664
rect 1932 656 1940 664
rect 1036 636 1044 644
rect 1196 636 1204 644
rect 1564 636 1572 644
rect 1596 636 1604 644
rect 2012 656 2020 664
rect 2028 656 2036 664
rect 2236 656 2244 664
rect 2252 656 2260 664
rect 2284 656 2292 664
rect 2492 656 2500 664
rect 2508 656 2516 664
rect 2620 656 2628 664
rect 2668 656 2676 664
rect 2844 656 2852 664
rect 3308 656 3316 664
rect 3468 656 3476 664
rect 3532 656 3540 664
rect 3564 656 3572 664
rect 3596 656 3604 664
rect 3628 656 3636 664
rect 3932 656 3940 664
rect 4188 656 4196 664
rect 4556 656 4564 664
rect 4620 656 4628 664
rect 4652 656 4660 664
rect 4748 656 4756 664
rect 4940 656 4948 664
rect 5260 656 5268 664
rect 5340 656 5348 664
rect 5404 656 5412 664
rect 5420 656 5428 664
rect 5548 656 5556 664
rect 5996 656 6004 664
rect 6300 656 6308 664
rect 6380 656 6388 664
rect 6572 656 6580 664
rect 6780 656 6788 664
rect 6828 656 6836 664
rect 6844 656 6852 664
rect 6876 656 6884 664
rect 6924 656 6932 664
rect 6972 656 6980 664
rect 7084 656 7092 664
rect 7340 656 7348 664
rect 7372 656 7380 664
rect 2092 636 2100 644
rect 2748 636 2756 644
rect 3116 636 3124 644
rect 3164 636 3172 644
rect 3676 636 3684 644
rect 3916 636 3924 644
rect 4204 636 4212 644
rect 4508 636 4516 644
rect 4572 636 4580 644
rect 4892 636 4900 644
rect 5628 636 5636 644
rect 5708 636 5716 644
rect 5740 636 5748 644
rect 5820 636 5828 644
rect 6124 636 6132 644
rect 6428 636 6436 644
rect 6588 636 6596 644
rect 7036 636 7044 644
rect 956 616 964 624
rect 1612 616 1620 624
rect 1708 616 1716 624
rect 1804 616 1812 624
rect 1932 616 1940 624
rect 2915 606 2923 614
rect 2925 606 2933 614
rect 2935 606 2943 614
rect 2945 606 2953 614
rect 2955 606 2963 614
rect 2965 606 2973 614
rect 5923 606 5931 614
rect 5933 606 5941 614
rect 5943 606 5951 614
rect 5953 606 5961 614
rect 5963 606 5971 614
rect 5973 606 5981 614
rect 876 596 884 604
rect 1164 596 1172 604
rect 1900 596 1908 604
rect 2012 596 2020 604
rect 2236 596 2244 604
rect 2252 596 2260 604
rect 364 576 372 584
rect 652 576 660 584
rect 716 576 724 584
rect 124 556 132 564
rect 300 556 308 564
rect 348 556 356 564
rect 524 556 532 564
rect 572 556 580 564
rect 604 556 612 564
rect 732 556 740 564
rect 748 556 756 564
rect 876 556 884 564
rect 940 556 948 564
rect 1020 576 1028 584
rect 1068 576 1076 584
rect 1260 576 1268 584
rect 1420 576 1428 584
rect 1548 576 1556 584
rect 1708 576 1716 584
rect 1740 576 1748 584
rect 1756 576 1764 584
rect 1788 576 1796 584
rect 2060 576 2068 584
rect 2108 576 2116 584
rect 2300 576 2308 584
rect 2636 576 2644 584
rect 2716 576 2724 584
rect 3036 576 3044 584
rect 3100 576 3108 584
rect 3292 576 3300 584
rect 3340 576 3348 584
rect 3420 576 3428 584
rect 3868 576 3876 584
rect 4252 576 4260 584
rect 4348 576 4356 584
rect 4604 576 4612 584
rect 4620 576 4628 584
rect 4700 576 4708 584
rect 5004 576 5012 584
rect 5068 576 5076 584
rect 5500 576 5508 584
rect 5612 576 5620 584
rect 5820 576 5828 584
rect 6028 576 6036 584
rect 6076 576 6084 584
rect 7036 576 7044 584
rect 1036 556 1044 564
rect 1052 556 1060 564
rect 1148 556 1156 564
rect 1164 556 1172 564
rect 1308 556 1316 564
rect 1612 556 1620 564
rect 1804 556 1812 564
rect 1900 556 1908 564
rect 2012 556 2020 564
rect 2044 556 2052 564
rect 2092 556 2100 564
rect 2236 556 2244 564
rect 2252 556 2260 564
rect 2364 556 2372 564
rect 2444 556 2452 564
rect 2508 556 2516 564
rect 2684 556 2692 564
rect 2732 556 2740 564
rect 2876 556 2884 564
rect 2892 556 2900 564
rect 3004 556 3012 564
rect 3116 556 3124 564
rect 3132 556 3140 564
rect 3212 556 3220 564
rect 3276 556 3284 564
rect 3372 556 3380 564
rect 3404 556 3412 564
rect 3484 556 3492 564
rect 3676 556 3684 564
rect 3708 556 3716 564
rect 3756 556 3764 564
rect 4812 556 4820 564
rect 5020 556 5028 564
rect 12 536 20 544
rect 108 536 116 544
rect 156 536 164 544
rect 380 536 388 544
rect 412 536 420 544
rect 508 536 516 544
rect 684 536 692 544
rect 764 536 772 544
rect 780 536 788 544
rect 812 536 820 544
rect 892 536 900 544
rect 1132 536 1140 544
rect 1260 536 1268 544
rect 1340 536 1348 544
rect 1372 536 1380 544
rect 1516 536 1524 544
rect 1628 536 1636 544
rect 1740 536 1748 544
rect 1756 536 1764 544
rect 1964 536 1972 544
rect 2140 536 2148 544
rect 2348 536 2356 544
rect 2428 536 2436 544
rect 2444 536 2452 544
rect 2604 536 2612 544
rect 2748 536 2756 544
rect 2812 536 2820 544
rect 2844 536 2852 544
rect 3004 536 3012 544
rect 3020 536 3028 544
rect 3084 536 3092 544
rect 3180 536 3188 544
rect 3196 536 3204 544
rect 3212 536 3220 544
rect 3324 536 3332 544
rect 3436 536 3444 544
rect 3484 536 3492 544
rect 3548 536 3556 544
rect 3580 536 3588 544
rect 3788 536 3796 544
rect 3804 536 3812 544
rect 140 516 148 524
rect 172 516 180 524
rect 220 516 228 524
rect 332 516 340 524
rect 396 516 404 524
rect 556 516 564 524
rect 604 516 612 524
rect 636 516 644 524
rect 780 516 788 524
rect 828 516 836 524
rect 908 516 916 524
rect 940 516 948 524
rect 1004 516 1012 524
rect 1084 516 1092 524
rect 1212 516 1220 524
rect 1228 516 1236 524
rect 1340 516 1348 524
rect 1468 516 1476 524
rect 1500 516 1508 524
rect 1564 516 1572 524
rect 1836 516 1844 524
rect 1900 516 1908 524
rect 1948 516 1956 524
rect 1980 516 1988 524
rect 2076 516 2084 524
rect 2124 516 2132 524
rect 2156 516 2164 524
rect 2172 516 2180 524
rect 2188 516 2196 524
rect 2300 516 2308 524
rect 2332 516 2340 524
rect 2492 516 2500 524
rect 2524 516 2532 524
rect 2540 516 2548 524
rect 2588 516 2596 524
rect 2652 516 2660 524
rect 2780 516 2788 524
rect 2796 516 2804 524
rect 2828 516 2836 524
rect 2860 516 2868 524
rect 3068 516 3076 524
rect 3180 516 3188 524
rect 3276 516 3284 524
rect 3308 516 3316 524
rect 3404 516 3412 524
rect 3516 516 3524 524
rect 3532 516 3540 524
rect 3596 516 3604 524
rect 3628 516 3636 524
rect 3740 516 3748 524
rect 3804 516 3812 524
rect 1292 496 1300 504
rect 1372 496 1380 504
rect 1468 496 1476 504
rect 1708 496 1716 504
rect 1788 496 1796 504
rect 1884 496 1892 504
rect 3052 496 3060 504
rect 3132 496 3140 504
rect 3356 496 3364 504
rect 3468 496 3476 504
rect 3612 496 3620 504
rect 3836 536 3844 544
rect 3852 536 3860 544
rect 3964 536 3972 544
rect 4076 536 4084 544
rect 4300 536 4308 544
rect 4412 536 4420 544
rect 4668 536 4676 544
rect 4716 536 4724 544
rect 5228 556 5236 564
rect 5356 556 5364 564
rect 5404 556 5412 564
rect 5468 556 5476 564
rect 5772 556 5780 564
rect 5804 556 5812 564
rect 5900 556 5908 564
rect 6188 556 6196 564
rect 6268 556 6276 564
rect 6284 556 6292 564
rect 6588 556 6596 564
rect 6684 556 6692 564
rect 7052 556 7060 564
rect 5100 536 5108 544
rect 5196 536 5204 544
rect 5228 536 5236 544
rect 5292 536 5300 544
rect 5308 532 5316 540
rect 5420 536 5428 544
rect 5564 536 5572 544
rect 5692 536 5700 544
rect 5740 536 5748 544
rect 5948 536 5956 544
rect 6092 536 6100 544
rect 6108 536 6116 544
rect 6204 536 6212 544
rect 6236 536 6244 544
rect 6268 536 6276 544
rect 6540 536 6548 544
rect 6620 536 6628 544
rect 6652 536 6660 544
rect 6700 536 6708 544
rect 6716 536 6724 544
rect 6908 536 6916 544
rect 6956 536 6964 544
rect 7004 536 7012 544
rect 7020 536 7028 544
rect 7100 536 7108 544
rect 3996 518 4004 526
rect 4124 516 4132 524
rect 4284 516 4292 524
rect 4316 516 4324 524
rect 4492 516 4500 524
rect 4540 516 4548 524
rect 4764 516 4772 524
rect 4876 518 4884 526
rect 4940 516 4948 524
rect 4620 496 4628 504
rect 4700 496 4708 504
rect 4748 496 4756 504
rect 4812 496 4820 504
rect 5132 496 5140 504
rect 5164 516 5172 524
rect 5276 516 5284 524
rect 5356 516 5364 524
rect 5372 516 5380 524
rect 5468 516 5476 524
rect 5500 516 5508 524
rect 5532 516 5540 524
rect 5580 516 5588 524
rect 5660 516 5668 524
rect 5692 516 5700 524
rect 5756 516 5764 524
rect 5868 516 5876 524
rect 6028 516 6036 524
rect 6060 516 6068 524
rect 6124 516 6132 524
rect 6220 516 6228 524
rect 6332 516 6340 524
rect 6476 516 6484 524
rect 6604 516 6612 524
rect 6668 516 6676 524
rect 6732 516 6740 524
rect 6860 516 6868 524
rect 6940 516 6948 524
rect 7004 516 7012 524
rect 7052 516 7060 524
rect 7100 516 7108 524
rect 7132 516 7140 524
rect 7244 516 7252 524
rect 7292 516 7300 524
rect 5452 496 5460 504
rect 5500 496 5508 504
rect 5612 496 5620 504
rect 5676 496 5684 504
rect 5804 496 5812 504
rect 6044 496 6052 504
rect 6060 496 6068 504
rect 6156 496 6164 504
rect 6172 496 6180 504
rect 6316 496 6324 504
rect 6652 496 6660 504
rect 6988 496 6996 504
rect 7116 496 7124 504
rect 7148 496 7156 504
rect 3644 476 3652 484
rect 3820 476 3828 484
rect 4572 476 4580 484
rect 5644 476 5652 484
rect 5868 476 5876 484
rect 5932 476 5940 484
rect 5980 476 5988 484
rect 6012 476 6020 484
rect 6380 476 6388 484
rect 7116 476 7124 484
rect 7132 456 7140 464
rect 44 436 52 444
rect 444 436 452 444
rect 1100 436 1108 444
rect 1692 436 1700 444
rect 3420 436 3428 444
rect 3580 436 3588 444
rect 3660 436 3668 444
rect 3692 436 3700 444
rect 3724 436 3732 444
rect 3756 436 3764 444
rect 4236 436 4244 444
rect 5388 436 5396 444
rect 5660 436 5668 444
rect 5740 436 5748 444
rect 6124 436 6132 444
rect 6364 436 6372 444
rect 6572 436 6580 444
rect 6748 436 6756 444
rect 7180 436 7188 444
rect 1411 406 1419 414
rect 1421 406 1429 414
rect 1431 406 1439 414
rect 1441 406 1449 414
rect 1451 406 1459 414
rect 1461 406 1469 414
rect 4419 406 4427 414
rect 4429 406 4437 414
rect 4439 406 4447 414
rect 4449 406 4457 414
rect 4459 406 4467 414
rect 4469 406 4477 414
rect 124 376 132 384
rect 188 376 196 384
rect 1196 376 1204 384
rect 1356 376 1364 384
rect 2092 376 2100 384
rect 2428 376 2436 384
rect 2636 376 2644 384
rect 3036 376 3044 384
rect 3116 376 3124 384
rect 3356 376 3364 384
rect 3516 376 3524 384
rect 3804 376 3812 384
rect 3932 376 3940 384
rect 4252 376 4260 384
rect 4300 376 4308 384
rect 4348 376 4356 384
rect 5100 376 5108 384
rect 6140 376 6148 384
rect 6188 376 6196 384
rect 6508 376 6516 384
rect 6780 376 6788 384
rect 7020 376 7028 384
rect 7340 376 7348 384
rect 988 356 996 364
rect 3660 356 3668 364
rect 4764 356 4772 364
rect 5612 356 5620 364
rect 1084 336 1092 344
rect 1180 336 1188 344
rect 44 316 52 324
rect 156 316 164 324
rect 348 316 356 324
rect 380 316 388 324
rect 428 316 436 324
rect 444 316 452 324
rect 492 316 500 324
rect 92 296 100 304
rect 124 296 132 304
rect 172 296 180 304
rect 348 296 356 304
rect 524 296 532 304
rect 604 296 612 304
rect 652 316 660 324
rect 1148 316 1156 324
rect 1244 316 1252 324
rect 1324 336 1332 344
rect 1884 336 1892 344
rect 2076 336 2084 344
rect 3500 336 3508 344
rect 3964 336 3972 344
rect 5468 336 5476 344
rect 5740 336 5748 344
rect 6156 336 6164 344
rect 6220 336 6228 344
rect 6524 336 6532 344
rect 6780 336 6788 344
rect 6796 336 6804 344
rect 6860 336 6868 344
rect 6988 336 6996 344
rect 7036 336 7044 344
rect 1548 316 1556 324
rect 684 296 692 304
rect 860 296 868 304
rect 908 296 916 304
rect 988 296 996 304
rect 1004 296 1012 304
rect 1052 296 1060 304
rect 1164 296 1172 304
rect 1292 296 1300 304
rect 1324 296 1332 304
rect 1388 296 1396 304
rect 1420 296 1428 304
rect 1596 316 1604 324
rect 1740 316 1748 324
rect 1612 296 1620 304
rect 1644 296 1652 304
rect 1788 316 1796 324
rect 1852 316 1860 324
rect 2108 316 2116 324
rect 2284 316 2292 324
rect 2780 316 2788 324
rect 2876 316 2884 324
rect 3292 316 3300 324
rect 3436 316 3444 324
rect 3468 316 3476 324
rect 3580 316 3588 324
rect 3692 316 3700 324
rect 1804 296 1812 304
rect 1884 296 1892 304
rect 1948 296 1956 304
rect 1996 296 2004 304
rect 2028 296 2036 304
rect 2092 296 2100 304
rect 2124 296 2132 304
rect 2156 296 2164 304
rect 2172 296 2180 304
rect 2220 296 2228 304
rect 2444 296 2452 304
rect 2844 296 2852 304
rect 3084 296 3092 304
rect 3164 296 3172 304
rect 3180 296 3188 304
rect 3452 296 3460 304
rect 3628 296 3636 304
rect 3644 296 3652 304
rect 3900 316 3908 324
rect 4332 316 4340 324
rect 4428 316 4436 324
rect 4588 316 4596 324
rect 4668 316 4676 324
rect 4748 316 4756 324
rect 4828 316 4836 324
rect 4908 316 4916 324
rect 5116 316 5124 324
rect 5196 316 5204 324
rect 3836 296 3844 304
rect 3948 296 3956 304
rect 12 276 20 284
rect 60 276 68 284
rect 108 276 116 284
rect 332 276 340 284
rect 396 276 404 284
rect 444 276 452 284
rect 476 276 484 284
rect 508 276 516 284
rect 4092 294 4100 302
rect 4156 296 4164 304
rect 4300 296 4308 304
rect 4396 296 4404 304
rect 4508 296 4516 304
rect 4604 296 4612 304
rect 4972 294 4980 302
rect 5036 296 5044 304
rect 5308 316 5316 324
rect 5436 316 5444 324
rect 5484 316 5492 324
rect 5532 316 5540 324
rect 5548 316 5556 324
rect 5772 316 5780 324
rect 6124 316 6132 324
rect 6348 316 6356 324
rect 6476 316 6484 324
rect 6492 316 6500 324
rect 6684 316 6692 324
rect 6700 316 6708 324
rect 6764 316 6772 324
rect 6828 316 6836 324
rect 7052 316 7060 324
rect 7164 316 7172 324
rect 5244 296 5252 304
rect 5356 296 5364 304
rect 5580 296 5588 304
rect 5644 296 5652 304
rect 5660 296 5668 304
rect 5692 296 5700 304
rect 5756 296 5764 304
rect 5804 296 5812 304
rect 5836 296 5844 304
rect 5900 296 5908 304
rect 5980 296 5988 304
rect 6044 296 6052 304
rect 6108 296 6116 304
rect 6140 296 6148 304
rect 6252 296 6260 304
rect 6316 296 6324 304
rect 6412 296 6420 304
rect 6508 296 6516 304
rect 6572 296 6580 304
rect 6716 296 6724 304
rect 6780 296 6788 304
rect 6876 296 6884 304
rect 7068 296 7076 304
rect 7116 296 7124 304
rect 7292 296 7300 304
rect 700 276 708 284
rect 796 276 804 284
rect 876 276 884 284
rect 1004 276 1012 284
rect 1036 276 1044 284
rect 1068 276 1076 284
rect 1212 276 1220 284
rect 1372 276 1380 284
rect 1436 276 1444 284
rect 1516 276 1524 284
rect 1708 276 1716 284
rect 1884 276 1892 284
rect 2012 276 2020 284
rect 2044 276 2052 284
rect 2172 276 2180 284
rect 2204 276 2212 284
rect 2316 276 2324 284
rect 2412 276 2420 284
rect 2460 276 2468 284
rect 2556 276 2564 284
rect 2604 276 2612 284
rect 2668 276 2676 284
rect 2812 276 2820 284
rect 2828 276 2836 284
rect 2892 276 2900 284
rect 3036 276 3044 284
rect 3260 276 3268 284
rect 3308 276 3316 284
rect 3404 276 3412 284
rect 3436 276 3444 284
rect 3500 276 3508 284
rect 3548 276 3556 284
rect 3708 276 3716 284
rect 3820 276 3828 284
rect 3852 276 3860 284
rect 3948 276 3956 284
rect 4076 276 4084 284
rect 4172 276 4180 284
rect 4268 276 4276 284
rect 4284 276 4292 284
rect 4364 276 4372 284
rect 4412 276 4420 284
rect 4556 276 4564 284
rect 4700 276 4708 284
rect 4716 276 4724 284
rect 4764 276 4772 284
rect 4796 276 4804 284
rect 4860 276 4868 284
rect 4876 276 4884 284
rect 4940 276 4948 284
rect 5164 276 5172 284
rect 5260 276 5268 284
rect 5276 276 5284 284
rect 5340 276 5348 284
rect 5388 276 5396 284
rect 5436 276 5444 284
rect 5484 276 5492 284
rect 5708 276 5716 284
rect 5740 276 5748 284
rect 5820 276 5828 284
rect 5852 276 5860 284
rect 5884 276 5892 284
rect 5996 276 6004 284
rect 6028 276 6036 284
rect 6092 276 6100 284
rect 6204 276 6212 284
rect 6380 276 6388 284
rect 6396 276 6404 284
rect 6556 276 6564 284
rect 6588 276 6596 284
rect 6636 276 6644 284
rect 6652 276 6660 284
rect 6876 276 6884 284
rect 60 256 68 264
rect 204 256 212 264
rect 220 256 228 264
rect 300 256 308 264
rect 444 256 452 264
rect 572 256 580 264
rect 812 256 820 264
rect 940 256 948 264
rect 956 256 964 264
rect 1100 256 1108 264
rect 1116 256 1124 264
rect 1260 256 1268 264
rect 1388 256 1396 264
rect 76 236 84 244
rect 268 236 276 244
rect 636 236 644 244
rect 1212 236 1220 244
rect 1228 236 1236 244
rect 1516 236 1524 244
rect 1676 256 1684 264
rect 1692 256 1700 264
rect 1836 256 1844 264
rect 1932 256 1940 264
rect 1948 256 1956 264
rect 2124 256 2132 264
rect 2252 256 2260 264
rect 2300 256 2308 264
rect 2444 256 2452 264
rect 2572 256 2580 264
rect 2620 256 2628 264
rect 2652 256 2660 264
rect 2972 256 2980 264
rect 2988 256 2996 264
rect 3100 256 3108 264
rect 3132 256 3140 264
rect 3180 256 3188 264
rect 3212 256 3220 264
rect 3340 256 3348 264
rect 3372 256 3380 264
rect 3532 256 3540 264
rect 3580 256 3588 264
rect 3596 256 3604 264
rect 3724 256 3732 264
rect 3772 256 3780 264
rect 3884 256 3892 264
rect 4204 256 4212 264
rect 4364 256 4372 264
rect 4652 256 4660 264
rect 4764 256 4772 264
rect 5292 256 5300 264
rect 5676 256 5684 264
rect 6028 256 6036 264
rect 6188 256 6196 264
rect 6284 256 6292 264
rect 6380 256 6388 264
rect 6620 256 6628 264
rect 6924 276 6932 284
rect 7116 276 7124 284
rect 7196 276 7204 284
rect 7276 276 7284 284
rect 7036 256 7044 264
rect 7228 256 7236 264
rect 7260 256 7268 264
rect 1708 236 1716 244
rect 1884 236 1892 244
rect 2348 236 2356 244
rect 2380 236 2388 244
rect 2700 236 2708 244
rect 2796 236 2804 244
rect 3788 236 3796 244
rect 3868 236 3876 244
rect 4636 236 4644 244
rect 4668 236 4676 244
rect 4892 236 4900 244
rect 5116 236 5124 244
rect 5212 236 5220 244
rect 5308 236 5316 244
rect 5436 236 5444 244
rect 5516 236 5524 244
rect 5548 236 5556 244
rect 5772 236 5780 244
rect 5884 236 5892 244
rect 6012 236 6020 244
rect 6076 236 6084 244
rect 6668 236 6676 244
rect 7212 236 7220 244
rect 812 216 820 224
rect 1836 216 1844 224
rect 1948 216 1956 224
rect 2252 216 2260 224
rect 2915 206 2923 214
rect 2925 206 2933 214
rect 2935 206 2943 214
rect 2945 206 2953 214
rect 2955 206 2963 214
rect 2965 206 2973 214
rect 5923 206 5931 214
rect 5933 206 5941 214
rect 5943 206 5951 214
rect 5953 206 5961 214
rect 5963 206 5971 214
rect 5973 206 5981 214
rect 1180 196 1188 204
rect 1324 196 1332 204
rect 1340 196 1348 204
rect 1580 196 1588 204
rect 1708 196 1716 204
rect 1804 196 1812 204
rect 1916 196 1924 204
rect 1932 196 1940 204
rect 2044 196 2052 204
rect 92 176 100 184
rect 204 176 212 184
rect 300 176 308 184
rect 396 176 404 184
rect 780 176 788 184
rect 892 176 900 184
rect 972 176 980 184
rect 1132 176 1140 184
rect 1356 176 1364 184
rect 284 156 292 164
rect 700 156 708 164
rect 1052 156 1060 164
rect 1180 156 1188 164
rect 1196 156 1204 164
rect 1324 156 1332 164
rect 1340 156 1348 164
rect 1548 176 1556 184
rect 1740 176 1748 184
rect 1868 176 1876 184
rect 2012 176 2020 184
rect 2076 176 2084 184
rect 2108 176 2116 184
rect 2204 176 2212 184
rect 2604 176 2612 184
rect 2924 176 2932 184
rect 3004 176 3012 184
rect 3532 176 3540 184
rect 3948 176 3956 184
rect 4204 176 4212 184
rect 4236 176 4244 184
rect 4476 176 4484 184
rect 4732 176 4740 184
rect 5644 176 5652 184
rect 5804 176 5812 184
rect 6172 176 6180 184
rect 6396 176 6404 184
rect 6508 176 6516 184
rect 6988 176 6996 184
rect 7132 176 7140 184
rect 7356 176 7364 184
rect 60 136 68 144
rect 172 136 180 144
rect 268 136 276 144
rect 332 136 340 144
rect 428 136 436 144
rect 508 136 516 144
rect 524 136 532 144
rect 556 136 564 144
rect 572 136 580 144
rect 620 136 628 144
rect 668 136 676 144
rect 716 136 724 144
rect 828 136 836 144
rect 924 136 932 144
rect 940 136 948 144
rect 1036 136 1044 144
rect 1260 136 1268 144
rect 1388 136 1396 144
rect 1564 156 1572 164
rect 1580 156 1588 164
rect 1708 156 1716 164
rect 1724 156 1732 164
rect 1804 156 1812 164
rect 1916 156 1924 164
rect 1932 156 1940 164
rect 2044 156 2052 164
rect 2092 156 2100 164
rect 2332 156 2340 164
rect 2396 156 2404 164
rect 2508 156 2516 164
rect 2588 156 2596 164
rect 2652 156 2660 164
rect 2716 156 2724 164
rect 2940 156 2948 164
rect 3180 156 3188 164
rect 3260 156 3268 164
rect 3356 156 3364 164
rect 3788 156 3796 164
rect 3916 156 3924 164
rect 4076 156 4084 164
rect 4140 156 4148 164
rect 4252 156 4260 164
rect 4284 156 4292 164
rect 5196 156 5204 164
rect 5660 156 5668 164
rect 5676 156 5684 164
rect 5692 156 5700 164
rect 6156 156 6164 164
rect 6428 156 6436 164
rect 6700 156 6708 164
rect 6780 156 6788 164
rect 6796 156 6804 164
rect 7116 156 7124 164
rect 7164 156 7172 164
rect 1644 136 1652 144
rect 1756 136 1764 144
rect 2172 136 2180 144
rect 2284 136 2292 144
rect 2476 136 2484 144
rect 2620 136 2628 144
rect 2636 136 2644 144
rect 2732 136 2740 144
rect 2828 136 2836 144
rect 2908 136 2916 144
rect 3052 136 3060 144
rect 3116 136 3124 144
rect 3132 136 3140 144
rect 3244 136 3252 144
rect 3340 136 3348 144
rect 3692 136 3700 144
rect 3852 136 3860 144
rect 4108 136 4116 144
rect 4380 136 4388 144
rect 4572 136 4580 144
rect 4796 136 4804 144
rect 4940 136 4948 144
rect 5004 136 5012 144
rect 5164 136 5172 144
rect 5260 136 5268 144
rect 5420 136 5428 144
rect 5468 136 5476 144
rect 5532 136 5540 144
rect 5868 136 5876 144
rect 5964 136 5972 144
rect 6188 136 6196 144
rect 6300 136 6308 144
rect 6604 136 6612 144
rect 6732 136 6740 144
rect 6748 136 6756 144
rect 6828 136 6836 144
rect 6972 136 6980 144
rect 7020 132 7028 140
rect 7244 136 7252 144
rect 284 116 292 124
rect 316 116 324 124
rect 444 116 452 124
rect 492 116 500 124
rect 556 116 564 124
rect 620 116 628 124
rect 668 116 676 124
rect 1100 116 1108 124
rect 1132 116 1140 124
rect 1244 116 1252 124
rect 1276 116 1284 124
rect 1484 116 1492 124
rect 1532 116 1540 124
rect 1628 116 1636 124
rect 1660 116 1668 124
rect 1772 116 1780 124
rect 1820 116 1828 124
rect 1868 116 1876 124
rect 1980 116 1988 124
rect 2012 116 2020 124
rect 2140 116 2148 124
rect 2268 116 2276 124
rect 2364 116 2372 124
rect 2428 116 2436 124
rect 2540 116 2548 124
rect 2636 116 2644 124
rect 2716 116 2724 124
rect 2876 116 2884 124
rect 2892 116 2900 124
rect 3068 116 3076 124
rect 3100 116 3108 124
rect 3164 116 3172 124
rect 3212 116 3220 124
rect 3324 116 3332 124
rect 3388 116 3396 124
rect 3436 116 3444 124
rect 3484 116 3492 124
rect 3660 118 3668 126
rect 3852 116 3860 124
rect 3868 116 3876 124
rect 3884 116 3892 124
rect 3932 116 3940 124
rect 4076 118 4084 126
rect 4188 116 4196 124
rect 4252 116 4260 124
rect 4348 118 4356 126
rect 4636 116 4644 124
rect 4748 116 4756 124
rect 4924 116 4932 124
rect 4972 116 4980 124
rect 4988 116 4996 124
rect 5004 116 5012 124
rect 5212 116 5220 124
rect 5276 116 5284 124
rect 5372 116 5380 124
rect 5452 116 5460 124
rect 5500 116 5508 124
rect 5548 116 5556 124
rect 5596 116 5604 124
rect 5740 116 5748 124
rect 5788 116 5796 124
rect 5932 118 5940 126
rect 6092 116 6100 124
rect 6108 116 6116 124
rect 6204 116 6212 124
rect 6268 118 6276 126
rect 6412 116 6420 124
rect 6476 116 6484 124
rect 6636 118 6644 126
rect 6748 116 6756 124
rect 6844 116 6852 124
rect 6876 116 6884 124
rect 6908 116 6916 124
rect 7100 116 7108 124
rect 7148 116 7156 124
rect 7228 118 7236 126
rect 604 96 612 104
rect 652 96 660 104
rect 1372 96 1380 104
rect 2108 96 2116 104
rect 2316 96 2324 104
rect 2444 96 2452 104
rect 2476 96 2484 104
rect 2524 96 2532 104
rect 3020 96 3028 104
rect 3052 96 3060 104
rect 3132 96 3140 104
rect 3308 96 3316 104
rect 3356 96 3364 104
rect 4156 96 4164 104
rect 4812 96 4820 104
rect 4828 96 4836 104
rect 4892 96 4900 104
rect 4956 96 4964 104
rect 5116 96 5124 104
rect 5308 96 5316 104
rect 5420 96 5428 104
rect 5532 96 5540 104
rect 6492 96 6500 104
rect 6700 96 6708 104
rect 6876 96 6884 104
rect 6892 96 6900 104
rect 6956 96 6964 104
rect 7052 96 7060 104
rect 12 76 20 84
rect 668 76 676 84
rect 2556 76 2564 84
rect 6428 76 6436 84
rect 6460 76 6468 84
rect 6924 76 6932 84
rect 2540 56 2548 64
rect 6908 56 6916 64
rect 476 36 484 44
rect 2844 36 2852 44
rect 3420 36 3428 44
rect 3468 36 3476 44
rect 3516 36 3524 44
rect 3724 36 3732 44
rect 3804 36 3812 44
rect 4844 36 4852 44
rect 5052 36 5060 44
rect 5068 36 5076 44
rect 5244 36 5252 44
rect 5356 36 5364 44
rect 5404 36 5412 44
rect 5580 36 5588 44
rect 5628 36 5636 44
rect 5708 36 5716 44
rect 5756 36 5764 44
rect 6060 36 6068 44
rect 6140 36 6148 44
rect 1411 6 1419 14
rect 1421 6 1429 14
rect 1431 6 1439 14
rect 1441 6 1449 14
rect 1451 6 1459 14
rect 1461 6 1469 14
rect 4419 6 4427 14
rect 4429 6 4437 14
rect 4439 6 4447 14
rect 4449 6 4457 14
rect 4459 6 4467 14
rect 4469 6 4477 14
<< metal2 >>
rect 397 5457 419 5463
rect 413 5384 419 5457
rect 557 5457 579 5463
rect 925 5457 947 5463
rect 973 5457 995 5463
rect 1229 5457 1251 5463
rect 3037 5457 3059 5463
rect 557 5384 563 5457
rect 925 5384 931 5457
rect 973 5384 979 5457
rect 1229 5384 1235 5457
rect 2938 5414 2950 5416
rect 2923 5406 2925 5414
rect 2933 5406 2935 5414
rect 2943 5406 2945 5414
rect 2953 5406 2955 5414
rect 2963 5406 2965 5414
rect 2938 5404 2950 5406
rect 2132 5377 2147 5383
rect 29 5317 44 5323
rect 29 5064 35 5317
rect 61 5304 67 5336
rect 141 5324 147 5336
rect 93 5224 99 5316
rect 173 5304 179 5316
rect 125 5264 131 5276
rect 205 5244 211 5336
rect 221 5284 227 5296
rect 269 5244 275 5336
rect 365 5323 371 5356
rect 365 5317 380 5323
rect 317 5284 323 5316
rect 141 5184 147 5236
rect 317 5164 323 5236
rect 381 5144 387 5316
rect 477 5224 483 5336
rect 509 5324 515 5336
rect 221 5124 227 5136
rect 45 5024 51 5076
rect 93 4984 99 5116
rect 109 5104 115 5116
rect 205 5064 211 5096
rect 148 5057 163 5063
rect 157 4984 163 5057
rect 45 4924 51 4936
rect 13 4884 19 4896
rect 13 4564 19 4676
rect 13 4324 19 4436
rect 13 4284 19 4316
rect 29 4304 35 4636
rect 45 4564 51 4916
rect 77 4744 83 4956
rect 205 4944 211 5056
rect 221 4984 227 5076
rect 253 5064 259 5076
rect 244 5037 259 5043
rect 237 4964 243 5016
rect 205 4744 211 4936
rect 77 4664 83 4736
rect 205 4704 211 4736
rect 93 4664 99 4676
rect 157 4664 163 4696
rect 237 4684 243 4956
rect 253 4824 259 5037
rect 285 4984 291 5096
rect 333 5084 339 5096
rect 301 4804 307 5076
rect 333 4964 339 5076
rect 365 5064 371 5096
rect 381 5084 387 5116
rect 461 5104 467 5216
rect 493 5204 499 5316
rect 445 5084 451 5096
rect 461 5064 467 5096
rect 493 5063 499 5116
rect 477 5057 499 5063
rect 349 4964 355 4996
rect 365 4944 371 5056
rect 461 5004 467 5056
rect 477 4984 483 5057
rect 509 4984 515 5056
rect 509 4964 515 4976
rect 381 4944 387 4956
rect 61 4564 67 4636
rect 125 4563 131 4656
rect 189 4564 195 4636
rect 253 4584 259 4696
rect 365 4684 371 4696
rect 381 4684 387 4936
rect 429 4904 435 4916
rect 493 4903 499 4936
rect 509 4923 515 4956
rect 525 4944 531 5336
rect 589 5304 595 5316
rect 605 5304 611 5336
rect 621 5324 627 5376
rect 1101 5357 1116 5363
rect 637 5324 643 5336
rect 701 5324 707 5336
rect 589 5184 595 5276
rect 637 5104 643 5176
rect 548 5097 563 5103
rect 541 4924 547 4956
rect 509 4917 531 4923
rect 493 4897 515 4903
rect 461 4784 467 4896
rect 381 4664 387 4676
rect 125 4557 140 4563
rect 45 4544 51 4556
rect 125 4544 131 4557
rect 317 4563 323 4636
rect 308 4557 323 4563
rect 397 4563 403 4636
rect 388 4557 403 4563
rect 77 4324 83 4516
rect 189 4504 195 4556
rect 301 4524 307 4556
rect 381 4524 387 4556
rect 397 4524 403 4536
rect 429 4523 435 4696
rect 445 4664 451 4676
rect 445 4564 451 4656
rect 477 4564 483 4656
rect 509 4644 515 4897
rect 525 4704 531 4917
rect 557 4904 563 5097
rect 605 5064 611 5096
rect 573 5044 579 5056
rect 653 5044 659 5296
rect 717 5264 723 5296
rect 749 5284 755 5336
rect 765 5324 771 5356
rect 845 5344 851 5356
rect 845 5184 851 5336
rect 957 5324 963 5336
rect 893 5224 899 5236
rect 685 5124 691 5156
rect 669 5084 675 5116
rect 573 4984 579 5036
rect 685 4984 691 5076
rect 749 5064 755 5156
rect 781 5104 787 5116
rect 845 5104 851 5136
rect 877 5104 883 5216
rect 797 5084 803 5096
rect 813 5084 819 5096
rect 765 4984 771 5036
rect 605 4964 611 4976
rect 589 4924 595 4956
rect 637 4944 643 4976
rect 637 4924 643 4936
rect 653 4904 659 4916
rect 557 4704 563 4836
rect 589 4764 595 4896
rect 589 4704 595 4756
rect 621 4723 627 4836
rect 621 4717 636 4723
rect 525 4664 531 4696
rect 493 4524 499 4636
rect 509 4544 515 4636
rect 589 4624 595 4696
rect 669 4684 675 4936
rect 685 4844 691 4896
rect 701 4744 707 4956
rect 733 4904 739 4936
rect 749 4924 755 4976
rect 797 4963 803 5076
rect 813 4984 819 5076
rect 845 5064 851 5096
rect 877 5084 883 5096
rect 893 5084 899 5096
rect 861 5004 867 5076
rect 925 5064 931 5116
rect 877 4984 883 5016
rect 797 4957 819 4963
rect 660 4657 675 4663
rect 653 4544 659 4636
rect 420 4517 435 4523
rect 93 4324 99 4436
rect 189 4323 195 4476
rect 253 4444 259 4516
rect 317 4364 323 4436
rect 189 4317 204 4323
rect 61 4244 67 4256
rect 13 3884 19 4116
rect 61 3924 67 4236
rect 77 4124 83 4296
rect 205 4284 211 4316
rect 349 4284 355 4316
rect 381 4264 387 4436
rect 429 4344 435 4517
rect 509 4484 515 4516
rect 445 4323 451 4356
rect 436 4317 451 4323
rect 189 4184 195 4236
rect 109 4164 115 4176
rect 205 4164 211 4256
rect 461 4244 467 4276
rect 285 4164 291 4236
rect 180 4157 195 4163
rect 109 4144 115 4156
rect 125 4144 131 4156
rect 189 4143 195 4157
rect 189 4137 204 4143
rect 173 4124 179 4136
rect 285 4084 291 4096
rect 333 4084 339 4156
rect 349 4144 355 4236
rect 365 4104 371 4236
rect 477 4124 483 4316
rect 109 3884 115 3916
rect 77 3764 83 3836
rect 125 3764 131 3836
rect 189 3784 195 4036
rect 237 4024 243 4036
rect 317 3877 332 3883
rect 301 3864 307 3876
rect 317 3864 323 3877
rect 349 3864 355 3876
rect 221 3764 227 3856
rect 365 3784 371 4096
rect 493 4063 499 4436
rect 509 4284 515 4476
rect 525 4284 531 4356
rect 621 4284 627 4296
rect 637 4284 643 4356
rect 653 4344 659 4536
rect 669 4504 675 4657
rect 685 4644 691 4656
rect 701 4644 707 4736
rect 717 4624 723 4676
rect 733 4664 739 4896
rect 717 4564 723 4616
rect 733 4584 739 4636
rect 749 4484 755 4636
rect 797 4563 803 4936
rect 813 4904 819 4957
rect 829 4944 835 4956
rect 893 4944 899 5056
rect 861 4904 867 4936
rect 893 4863 899 4936
rect 909 4884 915 5036
rect 925 4984 931 4996
rect 957 4963 963 5236
rect 973 5084 979 5116
rect 989 5064 995 5356
rect 1021 5323 1027 5336
rect 1012 5317 1027 5323
rect 1005 5284 1011 5316
rect 1069 5304 1075 5316
rect 1005 5144 1011 5276
rect 1101 5184 1107 5357
rect 1117 5324 1123 5336
rect 1149 5164 1155 5336
rect 1213 5264 1219 5336
rect 1405 5326 1411 5376
rect 2141 5364 2147 5377
rect 2436 5377 2451 5383
rect 2445 5364 2451 5377
rect 1629 5344 1635 5356
rect 1437 5324 1443 5336
rect 1117 5084 1123 5096
rect 1021 5064 1027 5076
rect 948 4957 963 4963
rect 941 4903 947 4956
rect 941 4897 963 4903
rect 893 4857 915 4863
rect 893 4784 899 4836
rect 909 4744 915 4857
rect 829 4664 835 4676
rect 813 4584 819 4636
rect 829 4584 835 4616
rect 845 4564 851 4656
rect 893 4644 899 4696
rect 797 4557 812 4563
rect 685 4304 691 4436
rect 525 4124 531 4256
rect 589 4164 595 4236
rect 637 4164 643 4276
rect 605 4157 620 4163
rect 541 4124 547 4136
rect 493 4057 515 4063
rect 445 3923 451 4036
rect 477 3984 483 4036
rect 429 3917 451 3923
rect 381 3864 387 3896
rect 397 3864 403 3916
rect 413 3904 419 3916
rect 397 3764 403 3856
rect 429 3763 435 3917
rect 461 3904 467 3916
rect 461 3864 467 3896
rect 429 3757 444 3763
rect 173 3744 179 3756
rect 13 3404 19 3456
rect 29 3404 35 3736
rect 61 3544 67 3636
rect 93 3404 99 3636
rect 157 3524 163 3636
rect 173 3604 179 3736
rect 189 3704 195 3756
rect 221 3744 227 3756
rect 365 3744 371 3756
rect 253 3704 259 3736
rect 381 3724 387 3736
rect 276 3717 284 3723
rect 237 3624 243 3636
rect 285 3584 291 3716
rect 269 3524 275 3536
rect 109 3504 115 3516
rect 157 3484 163 3516
rect 109 3464 115 3476
rect 29 3224 35 3236
rect 45 3203 51 3396
rect 109 3384 115 3456
rect 125 3384 131 3436
rect 77 3344 83 3356
rect 29 3197 51 3203
rect 29 3184 35 3197
rect 36 3097 51 3103
rect 13 3084 19 3096
rect 13 2964 19 3076
rect 45 2964 51 3097
rect 61 2704 67 3236
rect 77 3124 83 3216
rect 77 2964 83 3076
rect 77 2944 83 2956
rect 93 2943 99 3376
rect 237 3324 243 3496
rect 253 3364 259 3376
rect 301 3344 307 3576
rect 317 3504 323 3596
rect 317 3484 323 3496
rect 333 3484 339 3496
rect 349 3484 355 3636
rect 365 3463 371 3696
rect 381 3524 387 3616
rect 413 3584 419 3636
rect 429 3504 435 3716
rect 445 3504 451 3676
rect 429 3464 435 3476
rect 349 3457 371 3463
rect 301 3304 307 3336
rect 317 3324 323 3376
rect 132 3297 147 3303
rect 109 3084 115 3096
rect 141 3083 147 3297
rect 157 3104 163 3236
rect 349 3104 355 3457
rect 461 3463 467 3636
rect 477 3484 483 3936
rect 493 3904 499 4036
rect 509 3944 515 4057
rect 573 3924 579 4156
rect 605 4143 611 4157
rect 596 4137 611 4143
rect 669 4123 675 4196
rect 685 4144 691 4264
rect 701 4124 707 4216
rect 733 4163 739 4296
rect 749 4284 755 4476
rect 749 4204 755 4236
rect 724 4157 739 4163
rect 660 4117 675 4123
rect 541 3904 547 3916
rect 500 3897 515 3903
rect 493 3724 499 3836
rect 509 3764 515 3897
rect 557 3897 572 3903
rect 525 3744 531 3876
rect 557 3864 563 3897
rect 589 3664 595 4076
rect 605 3904 611 3916
rect 621 3884 627 3896
rect 653 3804 659 4036
rect 669 3884 675 4036
rect 765 3964 771 4516
rect 781 4444 787 4516
rect 781 4304 787 4336
rect 829 4324 835 4436
rect 797 4284 803 4316
rect 877 4304 883 4576
rect 925 4544 931 4656
rect 941 4564 947 4676
rect 957 4624 963 4897
rect 973 4864 979 5036
rect 989 5004 995 5056
rect 996 4957 1011 4963
rect 1005 4903 1011 4957
rect 989 4897 1011 4903
rect 989 4844 995 4897
rect 1021 4844 1027 4996
rect 1037 4964 1043 4996
rect 1053 4984 1059 5076
rect 1037 4924 1043 4956
rect 1069 4904 1075 5036
rect 1085 4984 1091 5056
rect 1165 4984 1171 5136
rect 1197 5104 1203 5256
rect 1213 5084 1219 5136
rect 1229 5104 1235 5116
rect 1245 5084 1251 5216
rect 1261 5124 1267 5316
rect 1277 5244 1283 5296
rect 1277 5224 1283 5236
rect 1565 5224 1571 5336
rect 1581 5304 1587 5316
rect 1434 5214 1446 5216
rect 1419 5206 1421 5214
rect 1429 5206 1431 5214
rect 1439 5206 1441 5214
rect 1449 5206 1451 5214
rect 1459 5206 1461 5214
rect 1434 5204 1446 5206
rect 1389 5183 1395 5196
rect 1389 5177 1404 5183
rect 1277 5124 1283 5176
rect 1309 5084 1315 5156
rect 1581 5144 1587 5256
rect 1428 5137 1443 5143
rect 1341 5104 1347 5136
rect 1325 5084 1331 5096
rect 1389 5083 1395 5116
rect 1412 5097 1427 5103
rect 1421 5084 1427 5097
rect 1389 5077 1411 5083
rect 1357 5064 1363 5076
rect 1085 4904 1091 4916
rect 989 4604 995 4696
rect 1005 4684 1011 4836
rect 1037 4784 1043 4896
rect 1165 4884 1171 4896
rect 1197 4884 1203 4916
rect 1213 4864 1219 4936
rect 1069 4704 1075 4756
rect 1069 4604 1075 4696
rect 1085 4644 1091 4656
rect 957 4524 963 4536
rect 973 4524 979 4536
rect 989 4524 995 4556
rect 925 4364 931 4516
rect 989 4384 995 4516
rect 925 4304 931 4356
rect 797 4124 803 4256
rect 813 4164 819 4276
rect 685 3864 691 3916
rect 765 3904 771 3956
rect 669 3784 675 3836
rect 701 3784 707 3836
rect 621 3764 627 3776
rect 733 3764 739 3836
rect 749 3764 755 3836
rect 797 3784 803 4116
rect 813 4004 819 4136
rect 861 4104 867 4236
rect 973 4224 979 4296
rect 1053 4284 1059 4556
rect 1069 4504 1075 4596
rect 1117 4583 1123 4636
rect 1101 4577 1123 4583
rect 1085 4524 1091 4576
rect 1101 4504 1107 4577
rect 1149 4564 1155 4676
rect 1165 4544 1171 4736
rect 1197 4724 1203 4836
rect 1229 4824 1235 4916
rect 1181 4684 1187 4696
rect 1149 4464 1155 4516
rect 1181 4484 1187 4636
rect 1213 4544 1219 4636
rect 1245 4544 1251 4836
rect 1309 4804 1315 4916
rect 1357 4884 1363 4956
rect 1373 4904 1379 4956
rect 1357 4744 1363 4836
rect 1389 4704 1395 5036
rect 1405 4984 1411 5077
rect 1437 5044 1443 5137
rect 1517 5064 1523 5136
rect 1597 5084 1603 5336
rect 1613 5224 1619 5316
rect 1805 5264 1811 5336
rect 1965 5324 1971 5336
rect 2013 5324 2019 5356
rect 1709 5104 1715 5116
rect 1821 5104 1827 5156
rect 1645 5024 1651 5036
rect 1469 4904 1475 4936
rect 1485 4824 1491 4956
rect 1565 4864 1571 4956
rect 1581 4924 1587 4936
rect 1597 4924 1603 4936
rect 1434 4814 1446 4816
rect 1419 4806 1421 4814
rect 1429 4806 1431 4814
rect 1439 4806 1441 4814
rect 1449 4806 1451 4814
rect 1459 4806 1461 4814
rect 1434 4804 1446 4806
rect 1581 4804 1587 4916
rect 1373 4684 1379 4696
rect 1613 4683 1619 5016
rect 1645 4944 1651 4956
rect 1661 4944 1667 5076
rect 1677 4984 1683 5036
rect 1693 5003 1699 5096
rect 1725 5084 1731 5096
rect 1709 5064 1715 5076
rect 1709 5024 1715 5056
rect 1693 4997 1731 5003
rect 1693 4944 1699 4956
rect 1709 4944 1715 4976
rect 1661 4904 1667 4916
rect 1629 4844 1635 4876
rect 1613 4677 1628 4683
rect 1389 4644 1395 4656
rect 1252 4517 1267 4523
rect 1149 4444 1155 4456
rect 1085 4344 1091 4436
rect 1197 4364 1203 4516
rect 1261 4504 1267 4517
rect 1277 4504 1283 4516
rect 1245 4464 1251 4496
rect 1309 4483 1315 4636
rect 1341 4524 1347 4536
rect 1357 4524 1363 4536
rect 1389 4484 1395 4616
rect 1421 4504 1427 4636
rect 1453 4544 1459 4576
rect 1485 4544 1491 4556
rect 1517 4484 1523 4676
rect 1581 4663 1587 4676
rect 1645 4664 1651 4696
rect 1661 4684 1667 4796
rect 1677 4704 1683 4736
rect 1693 4703 1699 4936
rect 1725 4924 1731 4997
rect 1741 4984 1747 5036
rect 1773 4964 1779 5096
rect 1837 5084 1843 5236
rect 1789 4943 1795 5016
rect 1805 4963 1811 5056
rect 1885 5044 1891 5056
rect 1821 4984 1827 5016
rect 1805 4957 1827 4963
rect 1780 4937 1795 4943
rect 1805 4924 1811 4936
rect 1741 4903 1747 4916
rect 1741 4897 1788 4903
rect 1805 4864 1811 4916
rect 1821 4884 1827 4957
rect 1853 4904 1859 5036
rect 1901 4924 1907 5156
rect 1949 5084 1955 5176
rect 2061 5104 2067 5276
rect 2093 5104 2099 5276
rect 2141 5244 2147 5356
rect 2221 5324 2227 5336
rect 2317 5324 2323 5356
rect 2445 5344 2451 5356
rect 2877 5344 2883 5376
rect 2525 5324 2531 5336
rect 2573 5324 2579 5336
rect 2669 5324 2675 5336
rect 2237 5144 2243 5316
rect 1949 5044 1955 5076
rect 1949 4944 1955 4976
rect 1693 4697 1708 4703
rect 1741 4684 1747 4716
rect 1773 4684 1779 4776
rect 1805 4724 1811 4736
rect 1837 4704 1843 4876
rect 1844 4697 1859 4703
rect 1853 4684 1859 4697
rect 1581 4657 1596 4663
rect 1549 4584 1555 4636
rect 1533 4557 1548 4563
rect 1533 4544 1539 4557
rect 1581 4544 1587 4556
rect 1677 4544 1683 4556
rect 1556 4537 1571 4543
rect 1300 4477 1315 4483
rect 1133 4284 1139 4296
rect 909 4164 915 4176
rect 845 3984 851 3996
rect 893 3884 899 4156
rect 925 4104 931 4136
rect 957 4084 963 4196
rect 1005 4164 1011 4256
rect 1053 4104 1059 4196
rect 1101 4184 1107 4236
rect 1133 4164 1139 4276
rect 1213 4204 1219 4296
rect 1229 4284 1235 4316
rect 1277 4304 1283 4436
rect 1373 4384 1379 4456
rect 1261 4264 1267 4296
rect 1309 4264 1315 4336
rect 1325 4244 1331 4296
rect 1389 4264 1395 4476
rect 1533 4464 1539 4516
rect 1565 4484 1571 4537
rect 1581 4504 1587 4536
rect 1597 4524 1603 4536
rect 1434 4414 1446 4416
rect 1419 4406 1421 4414
rect 1429 4406 1431 4414
rect 1439 4406 1441 4414
rect 1449 4406 1451 4414
rect 1459 4406 1461 4414
rect 1434 4404 1446 4406
rect 1325 4224 1331 4236
rect 1117 4124 1123 4156
rect 1341 4144 1347 4156
rect 1149 4124 1155 4136
rect 941 3923 947 4036
rect 1069 3984 1075 4036
rect 973 3924 979 3936
rect 925 3917 947 3923
rect 925 3884 931 3917
rect 836 3857 851 3863
rect 621 3724 627 3756
rect 685 3744 691 3756
rect 669 3724 675 3736
rect 765 3704 771 3716
rect 445 3457 467 3463
rect 365 3164 371 3236
rect 381 3124 387 3436
rect 413 3324 419 3376
rect 429 3104 435 3416
rect 445 3384 451 3457
rect 445 3344 451 3356
rect 445 3304 451 3336
rect 461 3304 467 3436
rect 477 3340 483 3376
rect 461 3104 467 3276
rect 477 3104 483 3136
rect 269 3084 275 3096
rect 141 3077 156 3083
rect 125 3064 131 3076
rect 141 3043 147 3077
rect 317 3064 323 3096
rect 397 3084 403 3096
rect 461 3064 467 3096
rect 125 3037 147 3043
rect 125 2944 131 3037
rect 93 2937 115 2943
rect 109 2723 115 2937
rect 141 2924 147 2936
rect 157 2784 163 3036
rect 173 2964 179 3056
rect 173 2924 179 2956
rect 221 2944 227 2956
rect 237 2904 243 3036
rect 285 2923 291 3036
rect 365 2924 371 3056
rect 493 3044 499 3496
rect 509 3484 515 3536
rect 541 3444 547 3456
rect 557 3424 563 3456
rect 589 3424 595 3636
rect 605 3504 611 3516
rect 605 3404 611 3436
rect 589 3364 595 3396
rect 637 3324 643 3516
rect 653 3484 659 3656
rect 717 3504 723 3516
rect 669 3484 675 3496
rect 685 3463 691 3496
rect 749 3484 755 3636
rect 797 3464 803 3636
rect 845 3584 851 3857
rect 861 3783 867 3836
rect 909 3824 915 3856
rect 941 3784 947 3896
rect 1021 3884 1027 3976
rect 861 3777 883 3783
rect 877 3764 883 3777
rect 861 3704 867 3756
rect 909 3724 915 3736
rect 893 3604 899 3636
rect 829 3517 844 3523
rect 829 3504 835 3517
rect 669 3457 691 3463
rect 653 3344 659 3356
rect 669 3324 675 3457
rect 765 3424 771 3456
rect 685 3344 691 3376
rect 701 3364 707 3396
rect 749 3344 755 3416
rect 781 3323 787 3416
rect 772 3317 787 3323
rect 541 3284 547 3316
rect 749 3303 755 3316
rect 749 3297 764 3303
rect 509 3224 515 3236
rect 509 3124 515 3196
rect 525 3104 531 3276
rect 461 2944 467 3036
rect 525 2943 531 3036
rect 509 2937 531 2943
rect 276 2917 291 2923
rect 301 2884 307 2916
rect 221 2724 227 2856
rect 301 2764 307 2836
rect 317 2804 323 2876
rect 365 2863 371 2916
rect 413 2903 419 2936
rect 509 2924 515 2937
rect 525 2917 540 2923
rect 525 2904 531 2917
rect 413 2897 435 2903
rect 365 2857 387 2863
rect 381 2844 387 2857
rect 109 2717 124 2723
rect 237 2703 243 2716
rect 253 2704 259 2756
rect 228 2697 243 2703
rect 109 2684 115 2696
rect 13 2583 19 2676
rect 76 2664 84 2670
rect 13 2577 35 2583
rect 29 2283 35 2577
rect 61 2544 67 2616
rect 77 2564 83 2636
rect 157 2564 163 2616
rect 157 2524 163 2536
rect 125 2304 131 2516
rect 93 2284 99 2296
rect 29 2277 51 2283
rect 45 2184 51 2277
rect 61 2203 67 2276
rect 93 2264 99 2276
rect 61 2197 83 2203
rect 61 2164 67 2176
rect 77 2144 83 2197
rect 61 2137 76 2143
rect 13 1904 19 2116
rect 13 1864 19 1876
rect 13 1784 19 1856
rect 61 1764 67 2137
rect 93 2124 99 2156
rect 77 2117 92 2123
rect 77 1904 83 2117
rect 109 2103 115 2276
rect 125 2143 131 2176
rect 157 2164 163 2256
rect 173 2184 179 2676
rect 189 2644 195 2676
rect 189 2284 195 2616
rect 205 2424 211 2516
rect 221 2504 227 2556
rect 237 2384 243 2516
rect 253 2464 259 2476
rect 301 2464 307 2516
rect 317 2484 323 2796
rect 365 2704 371 2836
rect 397 2584 403 2716
rect 413 2584 419 2876
rect 429 2784 435 2897
rect 557 2903 563 3156
rect 589 3104 595 3276
rect 733 3144 739 3236
rect 781 3164 787 3317
rect 797 3264 803 3316
rect 765 3144 771 3156
rect 813 3144 819 3456
rect 845 3424 851 3496
rect 845 3364 851 3396
rect 877 3264 883 3496
rect 893 3323 899 3516
rect 925 3424 931 3456
rect 941 3424 947 3456
rect 941 3364 947 3416
rect 893 3317 908 3323
rect 653 2984 659 3096
rect 605 2904 611 2916
rect 557 2897 572 2903
rect 468 2877 492 2883
rect 301 2344 307 2456
rect 349 2444 355 2536
rect 445 2524 451 2816
rect 509 2764 515 2836
rect 525 2784 531 2876
rect 541 2864 547 2896
rect 589 2804 595 2876
rect 605 2743 611 2836
rect 589 2737 611 2743
rect 509 2584 515 2736
rect 525 2704 531 2736
rect 573 2724 579 2736
rect 589 2704 595 2737
rect 621 2724 627 2856
rect 669 2804 675 3136
rect 820 3117 835 3123
rect 733 3104 739 3116
rect 781 3104 787 3116
rect 797 3103 803 3116
rect 797 3097 812 3103
rect 701 3084 707 3096
rect 685 2924 691 2976
rect 733 2924 739 3036
rect 717 2864 723 2896
rect 749 2884 755 2916
rect 797 2884 803 2996
rect 813 2924 819 2976
rect 717 2784 723 2836
rect 605 2703 611 2716
rect 605 2697 620 2703
rect 653 2644 659 2676
rect 669 2664 675 2756
rect 733 2704 739 2836
rect 557 2564 563 2596
rect 589 2564 595 2596
rect 653 2544 659 2556
rect 621 2524 627 2536
rect 461 2464 467 2516
rect 557 2504 563 2516
rect 333 2364 339 2436
rect 413 2384 419 2436
rect 317 2317 332 2323
rect 317 2304 323 2317
rect 349 2304 355 2376
rect 413 2344 419 2376
rect 397 2303 403 2316
rect 397 2297 412 2303
rect 205 2264 211 2296
rect 221 2264 227 2276
rect 317 2164 323 2276
rect 349 2184 355 2296
rect 413 2184 419 2236
rect 157 2144 163 2156
rect 445 2144 451 2236
rect 125 2137 147 2143
rect 109 2097 124 2103
rect 141 1984 147 2137
rect 173 2124 179 2136
rect 269 2124 275 2136
rect 397 2124 403 2136
rect 109 1884 115 1896
rect 141 1884 147 1896
rect 125 1784 131 1876
rect 13 1504 19 1696
rect 61 1464 67 1496
rect 61 1304 67 1456
rect 77 1384 83 1736
rect 93 1724 99 1756
rect 109 1584 115 1756
rect 141 1744 147 1756
rect 189 1724 195 1916
rect 205 1784 211 1856
rect 237 1784 243 1876
rect 269 1864 275 2116
rect 365 2084 371 2096
rect 381 2064 387 2116
rect 429 1984 435 2076
rect 445 2064 451 2096
rect 461 2024 467 2456
rect 509 2363 515 2436
rect 557 2364 563 2496
rect 637 2444 643 2516
rect 701 2483 707 2656
rect 749 2543 755 2696
rect 813 2683 819 2856
rect 829 2724 835 3117
rect 861 3084 867 3216
rect 941 3104 947 3136
rect 957 3084 963 3456
rect 989 3323 995 3436
rect 1005 3344 1011 3836
rect 1037 3783 1043 3836
rect 1021 3777 1043 3783
rect 1021 3744 1027 3777
rect 1069 3764 1075 3776
rect 1053 3744 1059 3756
rect 1101 3744 1107 4016
rect 1133 3923 1139 4036
rect 1165 3924 1171 4136
rect 1197 4124 1203 4136
rect 1245 4124 1251 4136
rect 1405 4124 1411 4376
rect 1565 4284 1571 4476
rect 1581 4304 1587 4356
rect 1661 4304 1667 4396
rect 1677 4304 1683 4516
rect 1693 4504 1699 4676
rect 1885 4664 1891 4856
rect 1917 4844 1923 4916
rect 1981 4904 1987 4956
rect 1997 4904 2003 4976
rect 2013 4924 2019 5016
rect 2061 4904 2067 5056
rect 2093 4944 2099 5056
rect 2116 5037 2131 5043
rect 2109 4944 2115 4956
rect 2125 4924 2131 5037
rect 2173 4984 2179 5116
rect 2317 5104 2323 5216
rect 2349 5124 2355 5296
rect 2237 5084 2243 5094
rect 2221 4984 2227 5016
rect 2301 4984 2307 5076
rect 2349 5024 2355 5116
rect 2493 5104 2499 5116
rect 2397 5084 2403 5096
rect 2173 4964 2179 4976
rect 2317 4964 2323 4976
rect 2109 4917 2124 4923
rect 1949 4784 1955 4896
rect 2029 4884 2035 4896
rect 1933 4684 1939 4696
rect 1741 4644 1747 4656
rect 1725 4637 1740 4643
rect 1725 4524 1731 4637
rect 1741 4524 1747 4536
rect 1789 4524 1795 4636
rect 1821 4543 1827 4636
rect 1869 4564 1875 4576
rect 1885 4564 1891 4656
rect 1837 4544 1843 4556
rect 1901 4544 1907 4636
rect 1805 4537 1827 4543
rect 1741 4344 1747 4516
rect 1805 4504 1811 4537
rect 1773 4484 1779 4496
rect 1821 4464 1827 4516
rect 1917 4504 1923 4516
rect 1757 4404 1763 4436
rect 1677 4264 1683 4276
rect 1469 4124 1475 4176
rect 1533 4123 1539 4236
rect 1645 4204 1651 4236
rect 1693 4184 1699 4336
rect 1725 4304 1731 4316
rect 1773 4284 1779 4456
rect 1805 4284 1811 4336
rect 1821 4304 1827 4316
rect 1853 4284 1859 4336
rect 1869 4284 1875 4436
rect 1933 4384 1939 4676
rect 1965 4604 1971 4836
rect 2013 4824 2019 4836
rect 2013 4784 2019 4796
rect 2109 4764 2115 4917
rect 2221 4884 2227 4936
rect 2237 4924 2243 4956
rect 1997 4644 2003 4656
rect 1981 4564 1987 4596
rect 1949 4524 1955 4556
rect 1981 4524 1987 4536
rect 1949 4344 1955 4376
rect 1997 4344 2003 4636
rect 2013 4543 2019 4756
rect 2093 4724 2099 4736
rect 2125 4684 2131 4876
rect 2189 4704 2195 4716
rect 2237 4704 2243 4916
rect 2253 4744 2259 4936
rect 2349 4904 2355 4936
rect 2365 4924 2371 4936
rect 2397 4924 2403 5076
rect 2413 5064 2419 5096
rect 2429 5004 2435 5036
rect 2429 4944 2435 4956
rect 2333 4784 2339 4856
rect 2365 4764 2371 4836
rect 2221 4697 2236 4703
rect 2221 4684 2227 4697
rect 2180 4677 2195 4683
rect 2029 4564 2035 4676
rect 2061 4604 2067 4670
rect 2141 4564 2147 4636
rect 2189 4584 2195 4677
rect 2221 4584 2227 4676
rect 2093 4544 2099 4556
rect 2157 4544 2163 4576
rect 2253 4544 2259 4736
rect 2285 4724 2291 4756
rect 2413 4744 2419 4936
rect 2461 4924 2467 5036
rect 2525 4944 2531 5316
rect 2541 5224 2547 5316
rect 2557 5184 2563 5316
rect 2525 4784 2531 4916
rect 2317 4664 2323 4736
rect 2381 4724 2387 4736
rect 2372 4697 2387 4703
rect 2269 4584 2275 4636
rect 2285 4564 2291 4636
rect 2317 4584 2323 4616
rect 2013 4537 2035 4543
rect 2029 4524 2035 4537
rect 1549 4164 1555 4176
rect 1741 4164 1747 4236
rect 1677 4124 1683 4156
rect 1741 4144 1747 4156
rect 1524 4117 1539 4123
rect 1117 3917 1139 3923
rect 1117 3884 1123 3917
rect 1165 3884 1171 3916
rect 1181 3904 1187 4016
rect 1277 3923 1283 4036
rect 1357 3984 1363 4036
rect 1434 4014 1446 4016
rect 1419 4006 1421 4014
rect 1429 4006 1431 4014
rect 1439 4006 1441 4014
rect 1449 4006 1451 4014
rect 1459 4006 1461 4014
rect 1434 4004 1446 4006
rect 1261 3917 1283 3923
rect 1197 3864 1203 3876
rect 1197 3764 1203 3856
rect 1021 3724 1027 3736
rect 1213 3704 1219 3896
rect 1229 3864 1235 3876
rect 1245 3744 1251 3796
rect 1261 3744 1267 3917
rect 1277 3884 1283 3896
rect 1309 3864 1315 3916
rect 1341 3884 1347 3896
rect 1389 3864 1395 3876
rect 1309 3804 1315 3836
rect 1437 3764 1443 3836
rect 1357 3744 1363 3756
rect 1021 3424 1027 3496
rect 1037 3484 1043 3596
rect 1069 3484 1075 3576
rect 1085 3504 1091 3636
rect 1165 3523 1171 3636
rect 1261 3524 1267 3736
rect 1437 3724 1443 3756
rect 1165 3517 1187 3523
rect 1149 3484 1155 3496
rect 1165 3484 1171 3496
rect 1108 3457 1132 3463
rect 1021 3364 1027 3376
rect 1085 3324 1091 3416
rect 1117 3344 1123 3436
rect 1165 3364 1171 3396
rect 1181 3364 1187 3517
rect 1213 3384 1219 3476
rect 1261 3464 1267 3496
rect 1277 3484 1283 3596
rect 1373 3564 1379 3716
rect 1434 3614 1446 3616
rect 1419 3606 1421 3614
rect 1429 3606 1431 3614
rect 1439 3606 1441 3614
rect 1449 3606 1451 3614
rect 1459 3606 1461 3614
rect 1434 3604 1446 3606
rect 1389 3584 1395 3596
rect 1229 3364 1235 3396
rect 989 3317 1004 3323
rect 845 3044 851 3076
rect 877 2923 883 3036
rect 925 2943 931 3036
rect 925 2937 947 2943
rect 868 2917 883 2923
rect 861 2704 867 2836
rect 909 2784 915 2876
rect 925 2864 931 2916
rect 941 2884 947 2937
rect 877 2704 883 2776
rect 797 2677 819 2683
rect 749 2537 771 2543
rect 701 2477 716 2483
rect 733 2463 739 2516
rect 749 2484 755 2496
rect 733 2457 755 2463
rect 605 2384 611 2436
rect 733 2384 739 2436
rect 493 2357 515 2363
rect 493 2344 499 2357
rect 493 2144 499 2176
rect 477 2124 483 2136
rect 477 1964 483 2116
rect 509 2084 515 2136
rect 541 2123 547 2356
rect 557 2244 563 2296
rect 541 2117 556 2123
rect 525 1984 531 2096
rect 573 2044 579 2276
rect 557 2004 563 2036
rect 525 1924 531 1936
rect 573 1924 579 1936
rect 173 1704 179 1716
rect 173 1584 179 1696
rect 109 1504 115 1576
rect 141 1464 147 1496
rect 221 1484 227 1756
rect 285 1744 291 1856
rect 301 1784 307 1916
rect 589 1904 595 2156
rect 605 2124 611 2296
rect 621 2124 627 2156
rect 637 2084 643 2376
rect 653 2304 659 2356
rect 685 2244 691 2336
rect 749 2304 755 2457
rect 765 2304 771 2537
rect 781 2344 787 2636
rect 797 2564 803 2677
rect 813 2544 819 2636
rect 829 2624 835 2656
rect 877 2644 883 2696
rect 893 2664 899 2696
rect 909 2684 915 2756
rect 925 2644 931 2836
rect 877 2564 883 2596
rect 836 2517 851 2523
rect 813 2503 819 2516
rect 813 2497 828 2503
rect 845 2483 851 2517
rect 829 2477 851 2483
rect 781 2304 787 2316
rect 829 2303 835 2477
rect 829 2297 844 2303
rect 685 2084 691 2236
rect 701 2164 707 2236
rect 749 2204 755 2256
rect 845 2244 851 2296
rect 605 1944 611 2076
rect 653 1924 659 2036
rect 333 1744 339 1756
rect 333 1724 339 1736
rect 93 1424 99 1456
rect 157 1424 163 1476
rect 205 1464 211 1476
rect 93 1344 99 1416
rect 205 1344 211 1436
rect 221 1424 227 1456
rect 237 1444 243 1456
rect 221 1344 227 1396
rect 141 1324 147 1336
rect 221 1324 227 1336
rect 237 1324 243 1436
rect 253 1384 259 1716
rect 381 1704 387 1756
rect 397 1724 403 1876
rect 445 1864 451 1876
rect 429 1724 435 1736
rect 269 1404 275 1496
rect 285 1383 291 1496
rect 317 1384 323 1476
rect 333 1444 339 1496
rect 381 1484 387 1696
rect 445 1584 451 1856
rect 461 1844 467 1896
rect 557 1884 563 1896
rect 701 1884 707 2036
rect 781 1884 787 2036
rect 829 1884 835 2036
rect 525 1784 531 1836
rect 701 1764 707 1776
rect 605 1744 611 1756
rect 717 1744 723 1776
rect 477 1704 483 1736
rect 493 1604 499 1736
rect 589 1704 595 1736
rect 637 1704 643 1716
rect 653 1644 659 1736
rect 669 1664 675 1716
rect 333 1384 339 1436
rect 365 1404 371 1456
rect 477 1444 483 1476
rect 493 1423 499 1456
rect 525 1444 531 1496
rect 541 1484 547 1596
rect 477 1417 499 1423
rect 477 1384 483 1417
rect 276 1377 291 1383
rect 541 1363 547 1476
rect 637 1464 643 1636
rect 733 1564 739 1816
rect 749 1764 755 1836
rect 765 1744 771 1836
rect 756 1717 771 1723
rect 765 1704 771 1717
rect 781 1684 787 1716
rect 797 1684 803 1756
rect 749 1584 755 1676
rect 781 1604 787 1636
rect 813 1584 819 1716
rect 829 1684 835 1836
rect 845 1764 851 2236
rect 861 2224 867 2496
rect 893 2284 899 2316
rect 909 2223 915 2636
rect 925 2324 931 2516
rect 941 2364 947 2816
rect 957 2764 963 2936
rect 973 2924 979 2956
rect 989 2904 995 2916
rect 1005 2783 1011 3236
rect 1021 2804 1027 3316
rect 1069 3303 1075 3316
rect 1069 3297 1084 3303
rect 1117 3264 1123 3316
rect 1245 3263 1251 3436
rect 1293 3424 1299 3496
rect 1309 3464 1315 3476
rect 1325 3443 1331 3496
rect 1309 3437 1331 3443
rect 1261 3284 1267 3296
rect 1277 3284 1283 3316
rect 1293 3304 1299 3336
rect 1309 3264 1315 3437
rect 1373 3424 1379 3456
rect 1405 3340 1411 3376
rect 1421 3364 1427 3516
rect 1437 3384 1443 3456
rect 1421 3344 1427 3356
rect 1325 3284 1331 3296
rect 1341 3284 1347 3316
rect 1357 3304 1363 3316
rect 1229 3257 1251 3263
rect 1197 3184 1203 3236
rect 1149 3144 1155 3156
rect 1037 2944 1043 2976
rect 1053 2964 1059 3036
rect 1085 3004 1091 3136
rect 1101 2984 1107 3096
rect 1149 3084 1155 3096
rect 1197 3064 1203 3096
rect 1101 2964 1107 2976
rect 1085 2924 1091 2956
rect 1133 2924 1139 2956
rect 1149 2884 1155 2996
rect 1213 2944 1219 3076
rect 1229 2984 1235 3257
rect 1245 3004 1251 3236
rect 1309 3084 1315 3156
rect 1325 3144 1331 3276
rect 1261 3044 1267 3076
rect 1229 2924 1235 2956
rect 989 2777 1011 2783
rect 957 2704 963 2716
rect 957 2644 963 2676
rect 957 2444 963 2516
rect 989 2324 995 2777
rect 1037 2744 1043 2756
rect 1053 2723 1059 2836
rect 1069 2724 1075 2796
rect 1037 2717 1059 2723
rect 1037 2704 1043 2717
rect 1117 2704 1123 2736
rect 1133 2724 1139 2856
rect 1149 2804 1155 2876
rect 1213 2824 1219 2916
rect 1197 2784 1203 2796
rect 1261 2724 1267 2976
rect 1293 2944 1299 2976
rect 1293 2884 1299 2916
rect 1325 2904 1331 3116
rect 1341 3104 1347 3236
rect 1357 3084 1363 3276
rect 1434 3214 1446 3216
rect 1419 3206 1421 3214
rect 1429 3206 1431 3214
rect 1439 3206 1441 3214
rect 1449 3206 1451 3214
rect 1459 3206 1461 3214
rect 1434 3204 1446 3206
rect 1341 2964 1347 3036
rect 1277 2744 1283 2756
rect 1309 2704 1315 2816
rect 1325 2804 1331 2876
rect 1373 2784 1379 3076
rect 1485 3064 1491 3776
rect 1533 3764 1539 3836
rect 1533 3724 1539 3736
rect 1533 3484 1539 3716
rect 1549 3704 1555 3716
rect 1565 3604 1571 4116
rect 1581 3844 1587 3896
rect 1613 3844 1619 3916
rect 1629 3864 1635 3976
rect 1597 3744 1603 3756
rect 1629 3723 1635 3856
rect 1645 3724 1651 3836
rect 1661 3764 1667 3836
rect 1677 3764 1683 4116
rect 1757 4104 1763 4116
rect 1789 4104 1795 4276
rect 1901 4263 1907 4296
rect 1965 4284 1971 4296
rect 1997 4264 2003 4316
rect 2029 4283 2035 4516
rect 2052 4497 2067 4503
rect 2013 4277 2035 4283
rect 1844 4257 1907 4263
rect 1917 4224 1923 4256
rect 1901 4144 1907 4156
rect 1917 4144 1923 4216
rect 1997 4163 2003 4196
rect 1988 4157 2003 4163
rect 1869 4084 1875 4136
rect 1965 4104 1971 4116
rect 1901 4004 1907 4036
rect 1693 3904 1699 3976
rect 1668 3757 1676 3763
rect 1620 3717 1635 3723
rect 1597 3524 1603 3716
rect 1629 3484 1635 3556
rect 1645 3504 1651 3636
rect 1517 3244 1523 3476
rect 1645 3444 1651 3456
rect 1533 3344 1539 3376
rect 1565 3324 1571 3436
rect 1501 3084 1507 3176
rect 1517 3104 1523 3236
rect 1549 3104 1555 3196
rect 1565 3044 1571 3276
rect 1581 3084 1587 3356
rect 1613 3324 1619 3396
rect 1613 3084 1619 3316
rect 1645 3304 1651 3336
rect 1661 3284 1667 3736
rect 1677 3504 1683 3556
rect 1677 3384 1683 3476
rect 1693 3424 1699 3896
rect 1709 3864 1715 3896
rect 1773 3884 1779 3896
rect 1837 3884 1843 3916
rect 1853 3904 1859 3916
rect 1821 3844 1827 3876
rect 1709 3404 1715 3436
rect 1725 3343 1731 3636
rect 1757 3563 1763 3836
rect 1805 3744 1811 3796
rect 1821 3724 1827 3836
rect 1853 3764 1859 3796
rect 1933 3784 1939 3836
rect 1869 3724 1875 3756
rect 1997 3744 2003 4157
rect 2013 3904 2019 4277
rect 2045 4264 2051 4296
rect 2045 4224 2051 4256
rect 2061 4184 2067 4497
rect 2205 4384 2211 4516
rect 2301 4504 2307 4516
rect 2349 4504 2355 4516
rect 2381 4464 2387 4697
rect 2541 4684 2547 5076
rect 2557 5064 2563 5094
rect 2589 5084 2595 5236
rect 2701 5164 2707 5236
rect 2557 4984 2563 4996
rect 2573 4963 2579 5016
rect 2557 4957 2579 4963
rect 2557 4904 2563 4957
rect 2621 4923 2627 5036
rect 2685 4924 2691 5096
rect 2749 4984 2755 5316
rect 2781 5304 2787 5316
rect 2893 5224 2899 5336
rect 2909 5224 2915 5316
rect 2989 5284 2995 5316
rect 3037 5304 3043 5316
rect 2877 5104 2883 5116
rect 3005 5084 3011 5136
rect 2989 5024 2995 5076
rect 2938 5014 2950 5016
rect 2923 5006 2925 5014
rect 2933 5006 2935 5014
rect 2943 5006 2945 5014
rect 2953 5006 2955 5014
rect 2963 5006 2965 5014
rect 2938 5004 2950 5006
rect 2813 4964 2819 4996
rect 3021 4984 3027 5096
rect 2884 4937 2899 4943
rect 2612 4917 2627 4923
rect 2845 4904 2851 4936
rect 2557 4764 2563 4896
rect 2573 4884 2579 4896
rect 2605 4704 2611 4776
rect 2621 4704 2627 4796
rect 2669 4704 2675 4776
rect 2733 4724 2739 4756
rect 2749 4704 2755 4896
rect 2861 4804 2867 4916
rect 2893 4884 2899 4937
rect 3037 4924 3043 4936
rect 2925 4784 2931 4896
rect 2765 4697 2780 4703
rect 2605 4684 2611 4696
rect 2477 4544 2483 4676
rect 2580 4657 2595 4663
rect 2365 4364 2371 4436
rect 2093 4284 2099 4336
rect 2189 4304 2195 4336
rect 2221 4304 2227 4336
rect 2141 4264 2147 4276
rect 2093 4204 2099 4256
rect 2141 4203 2147 4256
rect 2141 4197 2156 4203
rect 2045 4144 2051 4176
rect 2157 4164 2163 4196
rect 2173 4184 2179 4216
rect 2173 4164 2179 4176
rect 2093 4124 2099 4156
rect 2221 4144 2227 4296
rect 2237 4184 2243 4296
rect 2301 4224 2307 4276
rect 2253 4144 2259 4216
rect 2285 4144 2291 4156
rect 2045 3943 2051 4076
rect 2045 3937 2067 3943
rect 2061 3924 2067 3937
rect 2093 3904 2099 3976
rect 2029 3884 2035 3896
rect 2109 3784 2115 3856
rect 2141 3824 2147 3936
rect 2189 3884 2195 3916
rect 2285 3884 2291 4136
rect 2301 4044 2307 4116
rect 2317 4104 2323 4256
rect 2381 4124 2387 4456
rect 2477 4304 2483 4536
rect 2493 4526 2499 4556
rect 2557 4544 2563 4576
rect 2589 4544 2595 4657
rect 2653 4584 2659 4676
rect 2669 4664 2675 4696
rect 2749 4684 2755 4696
rect 2733 4544 2739 4556
rect 2557 4384 2563 4496
rect 2397 4204 2403 4276
rect 2436 4257 2451 4263
rect 2445 4224 2451 4257
rect 2397 4184 2403 4196
rect 2445 4184 2451 4216
rect 2333 3944 2339 4036
rect 2349 3904 2355 4036
rect 2413 3884 2419 3896
rect 2221 3844 2227 3876
rect 2253 3844 2259 3856
rect 2173 3764 2179 3836
rect 2205 3764 2211 3776
rect 1901 3604 1907 3636
rect 1757 3557 1779 3563
rect 1741 3523 1747 3536
rect 1741 3517 1763 3523
rect 1757 3504 1763 3517
rect 1741 3484 1747 3496
rect 1709 3337 1731 3343
rect 1709 3304 1715 3337
rect 1725 3184 1731 3316
rect 1741 3224 1747 3276
rect 1757 3083 1763 3236
rect 1773 3124 1779 3557
rect 1789 3444 1795 3516
rect 1805 3484 1811 3516
rect 1789 3364 1795 3436
rect 1821 3324 1827 3436
rect 1837 3324 1843 3376
rect 1853 3284 1859 3596
rect 1901 3464 1907 3516
rect 1933 3464 1939 3516
rect 1949 3484 1955 3556
rect 1965 3464 1971 3480
rect 1933 3344 1939 3456
rect 1965 3344 1971 3376
rect 1981 3364 1987 3596
rect 1997 3484 2003 3636
rect 2013 3564 2019 3636
rect 2045 3544 2051 3736
rect 2061 3544 2067 3756
rect 2285 3743 2291 3876
rect 2301 3804 2307 3836
rect 2301 3764 2307 3796
rect 2285 3737 2300 3743
rect 2173 3544 2179 3736
rect 2013 3524 2019 3536
rect 2061 3504 2067 3536
rect 2093 3464 2099 3476
rect 2141 3464 2147 3476
rect 1981 3344 1987 3356
rect 1997 3344 2003 3396
rect 2029 3324 2035 3416
rect 2077 3364 2083 3436
rect 2109 3424 2115 3456
rect 2141 3344 2147 3456
rect 1789 3224 1795 3276
rect 1805 3144 1811 3236
rect 1853 3104 1859 3256
rect 1780 3097 1795 3103
rect 1741 3077 1763 3083
rect 1389 2924 1395 2956
rect 1405 2884 1411 2956
rect 1485 2864 1491 3036
rect 1549 3024 1555 3036
rect 1597 3024 1603 3056
rect 1725 3044 1731 3056
rect 1501 2924 1507 2956
rect 1565 2944 1571 2976
rect 1517 2924 1523 2936
rect 1389 2824 1395 2836
rect 1434 2814 1446 2816
rect 1419 2806 1421 2814
rect 1429 2806 1431 2814
rect 1439 2806 1441 2814
rect 1449 2806 1451 2814
rect 1459 2806 1461 2814
rect 1434 2804 1446 2806
rect 1037 2604 1043 2636
rect 1005 2564 1011 2596
rect 1053 2544 1059 2696
rect 1133 2544 1139 2556
rect 1053 2384 1059 2516
rect 1117 2444 1123 2516
rect 1181 2504 1187 2696
rect 1213 2544 1219 2696
rect 925 2244 931 2276
rect 893 2217 915 2223
rect 861 2124 867 2136
rect 893 2124 899 2217
rect 909 2164 915 2196
rect 941 2104 947 2276
rect 957 2144 963 2316
rect 980 2297 995 2303
rect 989 2264 995 2297
rect 973 2144 979 2196
rect 957 2124 963 2136
rect 861 1904 867 1916
rect 893 1904 899 2016
rect 845 1684 851 1736
rect 877 1717 892 1723
rect 861 1683 867 1716
rect 877 1704 883 1717
rect 861 1677 883 1683
rect 861 1584 867 1636
rect 877 1584 883 1677
rect 893 1624 899 1636
rect 893 1584 899 1616
rect 701 1544 707 1556
rect 733 1544 739 1556
rect 797 1544 803 1556
rect 861 1544 867 1556
rect 749 1537 787 1543
rect 749 1523 755 1537
rect 781 1524 787 1537
rect 701 1517 755 1523
rect 701 1504 707 1517
rect 685 1444 691 1496
rect 532 1357 547 1363
rect 13 1284 19 1296
rect 109 1244 115 1316
rect 109 1104 115 1236
rect 269 1184 275 1356
rect 589 1344 595 1436
rect 653 1384 659 1436
rect 813 1384 819 1476
rect 829 1364 835 1396
rect 605 1344 611 1356
rect 509 1324 515 1336
rect 589 1324 595 1336
rect 669 1324 675 1336
rect 516 1317 531 1323
rect 285 1124 291 1316
rect 365 1284 371 1316
rect 349 1124 355 1176
rect 221 1104 227 1116
rect 237 1084 243 1116
rect 349 1104 355 1116
rect 45 1044 51 1056
rect 45 924 51 1036
rect 61 964 67 1036
rect 125 1004 131 1036
rect 13 884 19 896
rect 45 704 51 916
rect 61 724 67 956
rect 109 684 115 936
rect 125 744 131 956
rect 157 944 163 1036
rect 173 984 179 1076
rect 269 1064 275 1096
rect 189 963 195 1036
rect 189 957 204 963
rect 205 944 211 956
rect 237 924 243 996
rect 301 924 307 936
rect 13 544 19 676
rect 109 664 115 676
rect 125 664 131 696
rect 205 664 211 736
rect 269 724 275 876
rect 317 784 323 1076
rect 365 924 371 1276
rect 381 1164 387 1316
rect 429 1244 435 1316
rect 381 1104 387 1156
rect 461 1103 467 1236
rect 452 1097 467 1103
rect 461 1064 467 1097
rect 381 1004 387 1056
rect 381 984 387 996
rect 397 964 403 1056
rect 477 984 483 1096
rect 493 1044 499 1076
rect 509 983 515 1076
rect 493 977 515 983
rect 413 944 419 976
rect 493 964 499 977
rect 372 917 380 923
rect 525 864 531 1317
rect 564 1317 579 1323
rect 541 1124 547 1236
rect 557 884 563 936
rect 269 664 275 716
rect 285 704 291 716
rect 397 704 403 716
rect 317 664 323 696
rect 77 584 83 636
rect 109 544 115 656
rect 141 563 147 636
rect 253 584 259 636
rect 132 557 147 563
rect 157 544 163 576
rect 301 564 307 576
rect 317 564 323 656
rect 333 624 339 676
rect 381 664 387 676
rect 429 644 435 696
rect 365 584 371 636
rect 45 444 51 516
rect 45 324 51 436
rect 125 384 131 476
rect 141 323 147 516
rect 189 384 195 496
rect 141 317 156 323
rect 125 304 131 316
rect 173 284 179 296
rect 13 224 19 276
rect 221 264 227 276
rect 61 184 67 256
rect 285 243 291 516
rect 317 263 323 556
rect 349 484 355 556
rect 413 544 419 556
rect 445 550 451 656
rect 509 544 515 636
rect 525 584 531 856
rect 573 744 579 1317
rect 733 1264 739 1316
rect 669 1104 675 1116
rect 612 1097 636 1103
rect 685 1083 691 1216
rect 765 1184 771 1336
rect 669 1077 691 1083
rect 589 944 595 1016
rect 621 964 627 1076
rect 637 984 643 1076
rect 637 964 643 976
rect 653 964 659 996
rect 669 984 675 1077
rect 701 1064 707 1096
rect 765 1084 771 1136
rect 845 1123 851 1396
rect 877 1324 883 1516
rect 893 1324 899 1436
rect 909 1303 915 2096
rect 957 1984 963 2076
rect 941 1884 947 1916
rect 973 1884 979 1976
rect 1005 1903 1011 2356
rect 1053 2304 1059 2316
rect 1053 2244 1059 2296
rect 1085 2243 1091 2316
rect 1101 2304 1107 2336
rect 1085 2237 1107 2243
rect 1037 2164 1043 2196
rect 1053 2184 1059 2216
rect 1101 2184 1107 2237
rect 1085 2144 1091 2176
rect 1117 2164 1123 2376
rect 1149 2204 1155 2316
rect 1165 2224 1171 2496
rect 1229 2484 1235 2696
rect 1341 2664 1347 2716
rect 1485 2684 1491 2696
rect 1501 2663 1507 2816
rect 1533 2784 1539 2836
rect 1517 2704 1523 2776
rect 1549 2763 1555 2936
rect 1565 2884 1571 2916
rect 1565 2784 1571 2876
rect 1581 2844 1587 2936
rect 1597 2924 1603 2996
rect 1533 2757 1555 2763
rect 1517 2664 1523 2696
rect 1485 2657 1507 2663
rect 1261 2564 1267 2596
rect 1293 2584 1299 2636
rect 1485 2584 1491 2657
rect 1389 2544 1395 2576
rect 1533 2543 1539 2757
rect 1565 2723 1571 2776
rect 1613 2764 1619 3036
rect 1524 2537 1539 2543
rect 1549 2717 1571 2723
rect 1357 2524 1363 2536
rect 1549 2524 1555 2717
rect 1565 2564 1571 2596
rect 1181 2304 1187 2316
rect 1197 2304 1203 2336
rect 1213 2304 1219 2436
rect 1293 2324 1299 2516
rect 1293 2304 1299 2316
rect 1309 2304 1315 2516
rect 1133 2144 1139 2176
rect 1181 2164 1187 2196
rect 1213 2124 1219 2296
rect 1229 2224 1235 2256
rect 1245 2224 1251 2256
rect 1261 2144 1267 2156
rect 1261 2124 1267 2136
rect 1220 2117 1228 2123
rect 996 1897 1011 1903
rect 941 1824 947 1876
rect 1021 1863 1027 1996
rect 1101 1944 1107 2036
rect 1165 1944 1171 1956
rect 1037 1904 1043 1936
rect 1069 1904 1075 1936
rect 1037 1884 1043 1896
rect 1021 1857 1036 1863
rect 925 1744 931 1776
rect 925 1544 931 1576
rect 925 1504 931 1536
rect 941 1524 947 1756
rect 989 1717 1004 1723
rect 989 1704 995 1717
rect 1021 1703 1027 1756
rect 1012 1697 1027 1703
rect 957 1604 963 1636
rect 973 1544 979 1636
rect 957 1524 963 1536
rect 989 1524 995 1596
rect 1005 1464 1011 1536
rect 1053 1524 1059 1836
rect 1069 1744 1075 1876
rect 1069 1724 1075 1736
rect 1101 1683 1107 1936
rect 1181 1864 1187 1936
rect 1213 1784 1219 1876
rect 1245 1784 1251 1876
rect 1261 1864 1267 1896
rect 1277 1884 1283 2236
rect 1293 2144 1299 2296
rect 1325 2203 1331 2316
rect 1341 2224 1347 2256
rect 1325 2197 1347 2203
rect 1309 2164 1315 2196
rect 1341 2184 1347 2197
rect 1325 2144 1331 2176
rect 1357 2104 1363 2496
rect 1434 2414 1446 2416
rect 1419 2406 1421 2414
rect 1429 2406 1431 2414
rect 1439 2406 1441 2414
rect 1449 2406 1451 2414
rect 1459 2406 1461 2414
rect 1434 2404 1446 2406
rect 1421 2284 1427 2296
rect 1373 2184 1379 2196
rect 1389 2184 1395 2276
rect 1405 2264 1411 2276
rect 1405 2144 1411 2176
rect 1421 2164 1427 2276
rect 1341 1924 1347 2036
rect 1325 1844 1331 1876
rect 1165 1744 1171 1776
rect 1213 1744 1219 1776
rect 1341 1763 1347 1916
rect 1373 1884 1379 1976
rect 1389 1944 1395 2116
rect 1469 2084 1475 2316
rect 1434 2014 1446 2016
rect 1419 2006 1421 2014
rect 1429 2006 1431 2014
rect 1439 2006 1441 2014
rect 1449 2006 1451 2014
rect 1459 2006 1461 2014
rect 1434 2004 1446 2006
rect 1485 1924 1491 2096
rect 1501 2084 1507 2516
rect 1517 2164 1523 2476
rect 1533 2384 1539 2436
rect 1581 2404 1587 2656
rect 1645 2643 1651 2916
rect 1661 2884 1667 3036
rect 1677 2984 1683 2996
rect 1693 2944 1699 2976
rect 1741 2944 1747 3077
rect 1789 3064 1795 3097
rect 1837 3064 1843 3076
rect 1732 2917 1747 2923
rect 1741 2904 1747 2917
rect 1725 2884 1731 2896
rect 1693 2784 1699 2796
rect 1629 2637 1651 2643
rect 1565 2264 1571 2336
rect 1597 2324 1603 2376
rect 1613 2304 1619 2516
rect 1629 2364 1635 2637
rect 1533 2224 1539 2256
rect 1533 2164 1539 2176
rect 1517 2124 1523 2156
rect 1485 1883 1491 1896
rect 1501 1883 1507 2076
rect 1549 2063 1555 2176
rect 1565 2124 1571 2256
rect 1581 2204 1587 2256
rect 1533 2057 1555 2063
rect 1485 1877 1507 1883
rect 1389 1844 1395 1876
rect 1325 1757 1347 1763
rect 1117 1684 1123 1696
rect 1092 1677 1107 1683
rect 1117 1664 1123 1676
rect 1069 1604 1075 1636
rect 1085 1524 1091 1636
rect 1133 1504 1139 1716
rect 1149 1644 1155 1716
rect 1197 1544 1203 1716
rect 1213 1564 1219 1736
rect 1229 1724 1235 1756
rect 1277 1624 1283 1716
rect 1293 1704 1299 1736
rect 1325 1684 1331 1757
rect 1389 1744 1395 1776
rect 1437 1744 1443 1776
rect 1341 1724 1347 1736
rect 1485 1724 1491 1877
rect 1501 1824 1507 1856
rect 1517 1724 1523 1916
rect 1229 1524 1235 1556
rect 1037 1484 1043 1496
rect 1053 1464 1059 1496
rect 1117 1444 1123 1476
rect 1021 1424 1027 1436
rect 989 1384 995 1416
rect 957 1344 963 1376
rect 973 1364 979 1376
rect 925 1324 931 1336
rect 909 1297 924 1303
rect 925 1204 931 1296
rect 1005 1224 1011 1336
rect 1021 1324 1027 1396
rect 1069 1364 1075 1416
rect 1069 1297 1084 1303
rect 861 1184 867 1196
rect 989 1144 995 1156
rect 829 1117 851 1123
rect 861 1137 915 1143
rect 685 964 691 1056
rect 733 1044 739 1076
rect 765 964 771 1016
rect 797 964 803 1056
rect 717 944 723 956
rect 797 924 803 936
rect 685 784 691 916
rect 541 704 547 736
rect 621 644 627 676
rect 605 637 620 643
rect 381 504 387 536
rect 397 504 403 516
rect 333 284 339 356
rect 445 324 451 436
rect 509 364 515 536
rect 557 524 563 576
rect 605 564 611 637
rect 573 544 579 556
rect 429 304 435 316
rect 477 284 483 296
rect 493 284 499 316
rect 509 284 515 316
rect 525 284 531 296
rect 308 257 323 263
rect 285 237 307 243
rect 205 184 211 216
rect 269 184 275 236
rect 285 164 291 196
rect 301 184 307 237
rect 317 224 323 257
rect 493 244 499 276
rect 397 184 403 196
rect 173 144 179 156
rect 285 124 291 136
rect 317 124 323 156
rect 364 150 372 156
rect 445 124 451 216
rect 477 164 483 236
rect 493 124 499 176
rect 509 144 515 276
rect 557 224 563 496
rect 605 284 611 296
rect 621 264 627 636
rect 637 564 643 656
rect 653 584 659 736
rect 637 524 643 556
rect 685 544 691 756
rect 749 744 755 836
rect 749 704 755 736
rect 717 584 723 616
rect 733 564 739 576
rect 765 563 771 876
rect 813 784 819 816
rect 829 744 835 1117
rect 861 1103 867 1137
rect 877 1104 883 1116
rect 909 1104 915 1137
rect 932 1117 956 1123
rect 852 1097 867 1103
rect 893 1084 899 1096
rect 925 1084 931 1096
rect 900 1077 915 1083
rect 845 1064 851 1076
rect 845 1044 851 1056
rect 845 944 851 976
rect 877 964 883 1056
rect 909 964 915 1077
rect 989 1064 995 1096
rect 1069 1083 1075 1297
rect 1133 1283 1139 1436
rect 1149 1324 1155 1436
rect 1165 1384 1171 1496
rect 1245 1464 1251 1516
rect 1293 1503 1299 1656
rect 1325 1544 1331 1676
rect 1341 1664 1347 1716
rect 1341 1523 1347 1636
rect 1389 1544 1395 1636
rect 1434 1614 1446 1616
rect 1419 1606 1421 1614
rect 1429 1606 1431 1614
rect 1439 1606 1441 1614
rect 1449 1606 1451 1614
rect 1459 1606 1461 1614
rect 1434 1604 1446 1606
rect 1341 1517 1356 1523
rect 1293 1497 1308 1503
rect 1373 1484 1379 1496
rect 1181 1424 1187 1456
rect 1309 1344 1315 1436
rect 1485 1424 1491 1456
rect 1373 1344 1379 1416
rect 1124 1277 1139 1283
rect 1085 1104 1091 1276
rect 1133 1204 1139 1236
rect 1069 1077 1091 1083
rect 1053 1064 1059 1076
rect 957 984 963 996
rect 973 964 979 996
rect 1021 983 1027 1036
rect 1037 984 1043 1056
rect 1069 1024 1075 1056
rect 1005 977 1027 983
rect 1005 964 1011 977
rect 909 764 915 956
rect 845 664 851 696
rect 804 657 819 663
rect 781 584 787 636
rect 756 557 771 563
rect 653 244 659 316
rect 701 284 707 556
rect 813 544 819 657
rect 877 564 883 596
rect 788 537 803 543
rect 797 524 803 537
rect 909 524 915 736
rect 925 704 931 736
rect 973 683 979 876
rect 1005 704 1011 796
rect 964 677 979 683
rect 957 624 963 656
rect 1021 584 1027 696
rect 1037 684 1043 696
rect 1037 583 1043 636
rect 1053 604 1059 936
rect 1085 824 1091 1077
rect 1101 984 1107 1196
rect 1117 1157 1155 1163
rect 1117 1144 1123 1157
rect 1149 1143 1155 1157
rect 1149 1137 1171 1143
rect 1165 1124 1171 1137
rect 1085 704 1091 716
rect 1069 584 1075 656
rect 1037 577 1059 583
rect 1053 564 1059 577
rect 1101 564 1107 876
rect 1117 723 1123 1116
rect 1133 1044 1139 1056
rect 1149 924 1155 1116
rect 1165 964 1171 1096
rect 1181 764 1187 1316
rect 1197 1244 1203 1296
rect 1229 1143 1235 1316
rect 1220 1137 1235 1143
rect 1213 964 1219 1136
rect 1229 1084 1235 1096
rect 1245 1084 1251 1336
rect 1229 924 1235 1076
rect 1245 944 1251 1076
rect 1261 1064 1267 1236
rect 1293 1224 1299 1316
rect 1341 1124 1347 1156
rect 1373 1124 1379 1236
rect 1389 1204 1395 1416
rect 1405 1244 1411 1336
rect 1421 1324 1427 1356
rect 1501 1344 1507 1376
rect 1517 1324 1523 1596
rect 1533 1524 1539 2057
rect 1549 2024 1555 2036
rect 1597 1984 1603 2216
rect 1613 2184 1619 2296
rect 1629 2244 1635 2296
rect 1645 2284 1651 2516
rect 1661 2384 1667 2756
rect 1693 2564 1699 2596
rect 1709 2464 1715 2516
rect 1725 2464 1731 2576
rect 1693 2304 1699 2436
rect 1645 2183 1651 2276
rect 1677 2244 1683 2256
rect 1709 2223 1715 2276
rect 1741 2244 1747 2516
rect 1757 2504 1763 3056
rect 1773 2924 1779 2956
rect 1821 2903 1827 2996
rect 1837 2924 1843 2936
rect 1853 2904 1859 3056
rect 1869 2904 1875 3316
rect 2045 3284 2051 3296
rect 1901 3144 1907 3216
rect 1885 2924 1891 2936
rect 1821 2897 1843 2903
rect 1837 2884 1843 2897
rect 1773 2844 1779 2876
rect 1821 2864 1827 2876
rect 1837 2864 1843 2876
rect 1789 2724 1795 2836
rect 1805 2644 1811 2776
rect 1837 2744 1843 2836
rect 1821 2724 1827 2736
rect 1773 2544 1779 2636
rect 1821 2564 1827 2656
rect 1837 2644 1843 2716
rect 1885 2704 1891 2916
rect 1901 2844 1907 3136
rect 1917 3124 1923 3236
rect 2125 3184 2131 3316
rect 2189 3244 2195 3496
rect 2205 3484 2211 3676
rect 2237 3484 2243 3636
rect 2253 3584 2259 3636
rect 2301 3604 2307 3716
rect 2413 3664 2419 3876
rect 2429 3723 2435 3796
rect 2445 3783 2451 4036
rect 2461 3904 2467 4216
rect 2541 4144 2547 4276
rect 2557 4224 2563 4236
rect 2573 4144 2579 4516
rect 2621 4444 2627 4516
rect 2676 4497 2691 4503
rect 2557 4124 2563 4136
rect 2605 4124 2611 4216
rect 2477 4083 2483 4116
rect 2477 4077 2499 4083
rect 2461 3804 2467 3896
rect 2477 3884 2483 4056
rect 2493 3984 2499 4077
rect 2621 3984 2627 4436
rect 2653 4344 2659 4436
rect 2669 4184 2675 4296
rect 2653 4164 2659 4176
rect 2653 4124 2659 4136
rect 2685 4104 2691 4497
rect 2717 4484 2723 4536
rect 2765 4524 2771 4697
rect 2797 4684 2803 4736
rect 2925 4724 2931 4776
rect 2941 4704 2947 4916
rect 3053 4864 3059 5457
rect 5946 5414 5958 5416
rect 5931 5406 5933 5414
rect 5941 5406 5943 5414
rect 5951 5406 5953 5414
rect 5961 5406 5963 5414
rect 5971 5406 5973 5414
rect 5946 5404 5958 5406
rect 3677 5364 3683 5376
rect 3997 5364 4003 5376
rect 3197 5283 3203 5316
rect 3213 5304 3219 5336
rect 3197 5277 3219 5283
rect 3101 5124 3107 5216
rect 3101 5104 3107 5116
rect 3117 5084 3123 5116
rect 3165 5084 3171 5136
rect 3181 5124 3187 5176
rect 3197 5104 3203 5236
rect 3213 5184 3219 5277
rect 3293 5144 3299 5236
rect 3149 4984 3155 5056
rect 3085 4977 3139 4983
rect 3085 4944 3091 4977
rect 3133 4964 3139 4977
rect 3165 4964 3171 5076
rect 3181 4984 3187 5096
rect 3245 5084 3251 5096
rect 3325 5083 3331 5336
rect 3373 5284 3379 5316
rect 3693 5304 3699 5316
rect 3405 5184 3411 5196
rect 3485 5164 3491 5236
rect 3709 5224 3715 5336
rect 3789 5224 3795 5316
rect 3885 5204 3891 5356
rect 3997 5344 4003 5356
rect 4285 5344 4291 5376
rect 5101 5344 5107 5376
rect 5213 5344 5219 5356
rect 3933 5326 3939 5336
rect 3965 5324 3971 5336
rect 4077 5304 4083 5316
rect 4109 5284 4115 5316
rect 3357 5104 3363 5116
rect 3309 5077 3331 5083
rect 3117 4944 3123 4956
rect 3076 4917 3091 4923
rect 3085 4884 3091 4917
rect 3021 4704 3027 4856
rect 2813 4604 2819 4696
rect 2909 4684 2915 4696
rect 2941 4684 2947 4696
rect 2861 4644 2867 4656
rect 2781 4544 2787 4596
rect 2877 4524 2883 4636
rect 2938 4614 2950 4616
rect 2923 4606 2925 4614
rect 2933 4606 2935 4614
rect 2943 4606 2945 4614
rect 2953 4606 2955 4614
rect 2963 4606 2965 4614
rect 2938 4604 2950 4606
rect 2765 4223 2771 4516
rect 2781 4344 2787 4516
rect 2749 4217 2771 4223
rect 2749 4124 2755 4217
rect 2845 4184 2851 4296
rect 2861 4284 2867 4516
rect 3021 4303 3027 4696
rect 3021 4297 3036 4303
rect 2938 4214 2950 4216
rect 2923 4206 2925 4214
rect 2933 4206 2935 4214
rect 2943 4206 2945 4214
rect 2953 4206 2955 4214
rect 2963 4206 2965 4214
rect 2938 4204 2950 4206
rect 2765 4124 2771 4136
rect 2781 4124 2787 4136
rect 2877 4124 2883 4176
rect 2893 4144 2899 4156
rect 2909 4124 2915 4136
rect 2589 3904 2595 3956
rect 2637 3924 2643 4096
rect 2701 4044 2707 4116
rect 2445 3777 2460 3783
rect 2429 3717 2444 3723
rect 2541 3704 2547 3836
rect 2653 3784 2659 3956
rect 2685 3884 2691 3936
rect 2749 3924 2755 4116
rect 2989 4104 2995 4236
rect 3037 4184 3043 4256
rect 3101 4184 3107 4294
rect 3133 4284 3139 4676
rect 3149 4284 3155 4936
rect 3213 4883 3219 4936
rect 3197 4877 3219 4883
rect 3197 4684 3203 4877
rect 3245 4683 3251 4936
rect 3245 4677 3260 4683
rect 3245 4584 3251 4677
rect 3277 4624 3283 4696
rect 3309 4684 3315 5077
rect 3357 4944 3363 5096
rect 3485 5064 3491 5096
rect 3501 5064 3507 5076
rect 3437 5003 3443 5056
rect 3437 4997 3507 5003
rect 3380 4977 3459 4983
rect 3453 4964 3459 4977
rect 3501 4963 3507 4997
rect 3501 4957 3523 4963
rect 3437 4944 3443 4956
rect 3485 4944 3491 4956
rect 3444 4937 3459 4943
rect 3405 4903 3411 4916
rect 3396 4897 3411 4903
rect 3373 4824 3379 4896
rect 3421 4844 3427 4916
rect 3437 4744 3443 4836
rect 3357 4704 3363 4716
rect 3309 4544 3315 4676
rect 3405 4583 3411 4676
rect 3453 4604 3459 4937
rect 3501 4884 3507 4936
rect 3517 4924 3523 4957
rect 3533 4924 3539 5076
rect 3549 5064 3555 5156
rect 3549 4864 3555 4916
rect 3581 4884 3587 4896
rect 3549 4704 3555 4836
rect 3597 4784 3603 5096
rect 3629 5064 3635 5136
rect 3661 5104 3667 5116
rect 3693 5064 3699 5096
rect 3709 5084 3715 5116
rect 3805 5104 3811 5116
rect 3741 5064 3747 5096
rect 3789 5064 3795 5096
rect 3821 5084 3827 5116
rect 3885 5084 3891 5196
rect 3645 5057 3683 5063
rect 3645 5044 3651 5057
rect 3677 5043 3683 5057
rect 3677 5037 3724 5043
rect 3869 5024 3875 5076
rect 3629 4944 3635 4956
rect 3613 4924 3619 4936
rect 3645 4904 3651 4956
rect 3661 4924 3667 4976
rect 3853 4963 3859 5016
rect 3901 4984 3907 5096
rect 3853 4957 3875 4963
rect 3725 4943 3731 4956
rect 3725 4937 3740 4943
rect 3613 4724 3619 4736
rect 3485 4664 3491 4696
rect 3405 4577 3427 4583
rect 3325 4544 3331 4576
rect 3421 4544 3427 4577
rect 3565 4564 3571 4696
rect 3629 4684 3635 4716
rect 3661 4704 3667 4736
rect 3677 4684 3683 4716
rect 3693 4684 3699 4896
rect 3709 4784 3715 4816
rect 3581 4644 3587 4676
rect 3661 4584 3667 4656
rect 3677 4604 3683 4676
rect 3149 4144 3155 4276
rect 3165 4264 3171 4516
rect 3373 4503 3379 4516
rect 3364 4497 3379 4503
rect 3229 4224 3235 4236
rect 3181 4164 3187 4216
rect 3149 4124 3155 4136
rect 3069 4104 3075 4116
rect 2813 3924 2819 4096
rect 3117 3924 3123 3976
rect 2733 3884 2739 3896
rect 2253 3564 2259 3576
rect 2221 3464 2227 3476
rect 2253 3444 2259 3496
rect 2285 3484 2291 3536
rect 2333 3524 2339 3636
rect 2349 3497 2364 3503
rect 2221 3324 2227 3336
rect 2157 3164 2163 3236
rect 1933 3124 1939 3156
rect 1933 3004 1939 3096
rect 2013 3044 2019 3076
rect 1933 2904 1939 2956
rect 1949 2924 1955 2936
rect 1965 2884 1971 2996
rect 2045 2984 2051 3136
rect 2061 3104 2067 3136
rect 2077 3103 2083 3116
rect 2077 3097 2092 3103
rect 2061 3024 2067 3036
rect 2061 2944 2067 2976
rect 1981 2937 1996 2943
rect 1965 2864 1971 2876
rect 1869 2684 1875 2696
rect 1917 2684 1923 2836
rect 1981 2804 1987 2937
rect 1997 2917 2012 2923
rect 1997 2904 2003 2917
rect 1997 2744 2003 2836
rect 1901 2544 1907 2576
rect 1853 2484 1859 2516
rect 1764 2337 1779 2343
rect 1757 2304 1763 2336
rect 1709 2217 1731 2223
rect 1725 2184 1731 2217
rect 1629 2177 1651 2183
rect 1581 1924 1587 1936
rect 1597 1924 1603 1976
rect 1613 1904 1619 2136
rect 1629 2063 1635 2177
rect 1677 2137 1692 2143
rect 1645 2084 1651 2098
rect 1629 2057 1651 2063
rect 1645 1944 1651 2057
rect 1661 1944 1667 2016
rect 1677 1924 1683 2137
rect 1709 2024 1715 2156
rect 1693 1924 1699 1976
rect 1741 1963 1747 2096
rect 1757 2024 1763 2276
rect 1773 2144 1779 2337
rect 1789 2144 1795 2396
rect 1805 2383 1811 2436
rect 1869 2424 1875 2496
rect 1917 2424 1923 2496
rect 1853 2384 1859 2396
rect 1933 2384 1939 2676
rect 1965 2564 1971 2716
rect 1997 2584 2003 2736
rect 2029 2724 2035 2936
rect 2077 2923 2083 3056
rect 2125 3044 2131 3076
rect 2141 3064 2147 3096
rect 2157 3084 2163 3136
rect 2189 3044 2195 3076
rect 2205 3064 2211 3096
rect 2109 2944 2115 3036
rect 2093 2937 2108 2943
rect 2093 2924 2099 2937
rect 2157 2924 2163 2956
rect 2068 2917 2083 2923
rect 2061 2764 2067 2916
rect 2045 2684 2051 2696
rect 1997 2484 2003 2536
rect 2045 2484 2051 2576
rect 1949 2424 1955 2476
rect 1805 2377 1827 2383
rect 1805 2304 1811 2356
rect 1821 2344 1827 2377
rect 2013 2344 2019 2436
rect 1821 2264 1827 2296
rect 1869 2264 1875 2296
rect 1789 2124 1795 2136
rect 1725 1957 1747 1963
rect 1629 1904 1635 1916
rect 1709 1904 1715 1956
rect 1597 1897 1612 1903
rect 1549 1864 1555 1896
rect 1597 1804 1603 1897
rect 1565 1644 1571 1756
rect 1597 1740 1603 1796
rect 1629 1724 1635 1896
rect 1661 1884 1667 1896
rect 1645 1803 1651 1876
rect 1645 1797 1667 1803
rect 1661 1764 1667 1797
rect 1629 1644 1635 1696
rect 1565 1564 1571 1636
rect 1597 1524 1603 1536
rect 1533 1504 1539 1516
rect 1677 1504 1683 1836
rect 1725 1824 1731 1957
rect 1757 1884 1763 1936
rect 1789 1884 1795 1916
rect 1821 1883 1827 2236
rect 1837 2164 1843 2196
rect 1837 1944 1843 2136
rect 1853 2124 1859 2236
rect 1869 2143 1875 2256
rect 1901 2244 1907 2256
rect 1885 2184 1891 2196
rect 1917 2164 1923 2236
rect 1917 2144 1923 2156
rect 1869 2137 1891 2143
rect 1805 1877 1827 1883
rect 1693 1684 1699 1736
rect 1709 1724 1715 1736
rect 1741 1663 1747 1856
rect 1757 1744 1763 1876
rect 1757 1723 1763 1736
rect 1757 1717 1772 1723
rect 1741 1657 1763 1663
rect 1709 1484 1715 1636
rect 1725 1504 1731 1516
rect 1629 1384 1635 1476
rect 1549 1324 1555 1356
rect 1434 1214 1446 1216
rect 1419 1206 1421 1214
rect 1429 1206 1431 1214
rect 1439 1206 1441 1214
rect 1449 1206 1451 1214
rect 1459 1206 1461 1214
rect 1434 1204 1446 1206
rect 1485 1204 1491 1296
rect 1565 1244 1571 1336
rect 1613 1324 1619 1336
rect 1517 1183 1523 1236
rect 1581 1184 1587 1316
rect 1501 1177 1523 1183
rect 1501 1164 1507 1177
rect 1517 1124 1523 1156
rect 1533 1104 1539 1116
rect 1613 1104 1619 1316
rect 1629 1224 1635 1336
rect 1645 1163 1651 1456
rect 1661 1424 1667 1456
rect 1677 1424 1683 1456
rect 1725 1344 1731 1376
rect 1645 1157 1667 1163
rect 1261 1004 1267 1056
rect 1341 1044 1347 1076
rect 1389 1064 1395 1096
rect 1485 1084 1491 1096
rect 1565 1064 1571 1096
rect 1613 1064 1619 1076
rect 1645 1064 1651 1136
rect 1293 944 1299 1016
rect 1325 1004 1331 1036
rect 1373 984 1379 1036
rect 1389 964 1395 1056
rect 1469 924 1475 1036
rect 1549 964 1555 996
rect 1565 984 1571 996
rect 1501 944 1507 956
rect 1581 944 1587 956
rect 1597 944 1603 956
rect 1565 924 1571 936
rect 1613 923 1619 976
rect 1613 917 1628 923
rect 1133 744 1139 756
rect 1117 717 1139 723
rect 1117 664 1123 696
rect 1133 664 1139 717
rect 1165 704 1171 716
rect 1197 704 1203 836
rect 1213 724 1219 796
rect 781 384 787 516
rect 829 284 835 516
rect 909 444 915 516
rect 909 304 915 376
rect 861 284 867 296
rect 797 264 803 276
rect 877 264 883 276
rect 557 144 563 216
rect 573 144 579 176
rect 557 104 563 116
rect 605 104 611 236
rect 637 164 643 236
rect 813 224 819 256
rect 781 184 787 196
rect 701 164 707 176
rect 621 144 627 156
rect 829 144 835 256
rect 925 144 931 556
rect 941 544 947 556
rect 1005 524 1011 536
rect 941 304 947 516
rect 1037 484 1043 556
rect 1133 544 1139 596
rect 1149 564 1155 696
rect 1293 684 1299 916
rect 1533 904 1539 916
rect 1357 884 1363 896
rect 1469 884 1475 896
rect 1434 814 1446 816
rect 1419 806 1421 814
rect 1429 806 1431 814
rect 1439 806 1441 814
rect 1449 806 1451 814
rect 1459 806 1461 814
rect 1434 804 1446 806
rect 1485 783 1491 816
rect 1517 784 1523 876
rect 1469 777 1491 783
rect 1165 564 1171 596
rect 1005 324 1011 436
rect 1005 304 1011 316
rect 989 264 995 296
rect 1021 283 1027 336
rect 1012 277 1027 283
rect 1037 264 1043 276
rect 1069 264 1075 276
rect 1101 264 1107 436
rect 941 224 947 256
rect 973 184 979 216
rect 941 144 947 176
rect 989 156 995 236
rect 1037 144 1043 196
rect 1133 184 1139 476
rect 1149 324 1155 356
rect 1181 344 1187 656
rect 1197 544 1203 636
rect 1261 544 1267 576
rect 1293 564 1299 676
rect 1309 564 1315 696
rect 1341 644 1347 656
rect 1213 484 1219 516
rect 1197 384 1203 436
rect 1245 324 1251 496
rect 1165 244 1171 296
rect 1261 283 1267 376
rect 1325 344 1331 616
rect 1341 544 1347 596
rect 1357 384 1363 656
rect 1373 564 1379 696
rect 1421 584 1427 696
rect 1437 544 1443 636
rect 1373 524 1379 536
rect 1373 504 1379 516
rect 1453 503 1459 716
rect 1469 704 1475 777
rect 1533 643 1539 716
rect 1533 637 1555 643
rect 1469 524 1475 596
rect 1549 584 1555 637
rect 1565 624 1571 636
rect 1453 497 1468 503
rect 1485 424 1491 476
rect 1434 414 1446 416
rect 1419 406 1421 414
rect 1429 406 1431 414
rect 1439 406 1441 414
rect 1449 406 1451 414
rect 1459 406 1461 414
rect 1434 404 1446 406
rect 1421 304 1427 316
rect 1293 284 1299 296
rect 1245 277 1267 283
rect 1213 244 1219 276
rect 1181 164 1187 196
rect 1197 164 1203 176
rect 1229 164 1235 236
rect 1053 144 1059 156
rect 1245 144 1251 277
rect 1325 264 1331 296
rect 1437 284 1443 336
rect 1357 277 1372 283
rect 1261 144 1267 256
rect 1325 164 1331 196
rect 1341 164 1347 196
rect 1357 184 1363 277
rect 1389 264 1395 276
rect 676 137 691 143
rect 685 104 691 137
rect 717 124 723 136
rect 1101 124 1107 136
rect 1245 124 1251 136
rect 1373 104 1379 156
rect 1485 124 1491 416
rect 1549 324 1555 496
rect 1581 444 1587 656
rect 1597 604 1603 636
rect 1613 624 1619 656
rect 1645 564 1651 836
rect 1661 704 1667 1157
rect 1709 1104 1715 1336
rect 1741 1224 1747 1616
rect 1757 1584 1763 1657
rect 1773 1564 1779 1636
rect 1789 1464 1795 1836
rect 1805 1624 1811 1877
rect 1837 1724 1843 1736
rect 1837 1504 1843 1636
rect 1853 1544 1859 1936
rect 1869 1904 1875 2116
rect 1885 2104 1891 2137
rect 1917 1884 1923 2076
rect 1869 1864 1875 1876
rect 1917 1864 1923 1876
rect 1869 1724 1875 1776
rect 1917 1724 1923 1856
rect 1933 1764 1939 2336
rect 2045 2324 2051 2436
rect 2061 2384 2067 2516
rect 2077 2364 2083 2496
rect 1965 2284 1971 2296
rect 1949 2244 1955 2256
rect 1965 2184 1971 2276
rect 2013 2140 2019 2256
rect 2029 2144 2035 2156
rect 1981 2124 1987 2136
rect 1965 1944 1971 2096
rect 1997 1944 2003 2116
rect 2013 2024 2019 2132
rect 2045 2124 2051 2176
rect 2061 2164 2067 2296
rect 2077 2284 2083 2296
rect 2093 2284 2099 2916
rect 2125 2897 2140 2903
rect 2125 2784 2131 2897
rect 2173 2903 2179 3036
rect 2205 2964 2211 3016
rect 2221 2964 2227 3036
rect 2237 3004 2243 3436
rect 2253 3364 2259 3376
rect 2269 3337 2284 3343
rect 2269 2944 2275 3337
rect 2301 3203 2307 3476
rect 2285 3197 2307 3203
rect 2285 2944 2291 3197
rect 2301 3104 2307 3176
rect 2317 3084 2323 3456
rect 2333 3084 2339 3156
rect 2349 3104 2355 3497
rect 2381 3324 2387 3656
rect 2413 3523 2419 3636
rect 2397 3517 2419 3523
rect 2397 3384 2403 3517
rect 2509 3484 2515 3496
rect 2525 3484 2531 3656
rect 2637 3584 2643 3636
rect 2461 3424 2467 3456
rect 2397 3344 2403 3376
rect 2509 3344 2515 3456
rect 2557 3364 2563 3436
rect 2589 3340 2595 3396
rect 2621 3384 2627 3476
rect 2349 3084 2355 3096
rect 2212 2917 2236 2923
rect 2157 2897 2179 2903
rect 2109 2484 2115 2736
rect 2125 2524 2131 2696
rect 2157 2483 2163 2897
rect 2253 2784 2259 2896
rect 2269 2864 2275 2876
rect 2285 2864 2291 2916
rect 2301 2904 2307 2996
rect 2333 2924 2339 2976
rect 2365 2904 2371 3236
rect 2413 3184 2419 3336
rect 2509 3143 2515 3336
rect 2493 3137 2515 3143
rect 2445 3104 2451 3116
rect 2381 3024 2387 3096
rect 2493 3084 2499 3137
rect 2525 3104 2531 3236
rect 2573 3204 2579 3336
rect 2589 3084 2595 3176
rect 2605 3104 2611 3356
rect 2621 3264 2627 3376
rect 2637 3324 2643 3516
rect 2669 3504 2675 3576
rect 2669 3323 2675 3476
rect 2685 3344 2691 3876
rect 2701 3844 2707 3856
rect 2717 3724 2723 3836
rect 2749 3664 2755 3896
rect 2765 3864 2771 3876
rect 2813 3764 2819 3836
rect 2877 3744 2883 3896
rect 3117 3884 3123 3896
rect 3133 3884 3139 4116
rect 3197 4084 3203 4116
rect 3165 3904 3171 3976
rect 3172 3877 3180 3883
rect 2893 3744 2899 3876
rect 3021 3864 3027 3876
rect 3021 3844 3027 3856
rect 2938 3814 2950 3816
rect 2923 3806 2925 3814
rect 2933 3806 2935 3814
rect 2943 3806 2945 3814
rect 2953 3806 2955 3814
rect 2963 3806 2965 3814
rect 2938 3804 2950 3806
rect 3165 3744 3171 3876
rect 2701 3484 2707 3556
rect 2797 3484 2803 3576
rect 2845 3484 2851 3696
rect 2877 3444 2883 3736
rect 2893 3584 2899 3676
rect 2733 3384 2739 3436
rect 2765 3324 2771 3376
rect 2781 3324 2787 3416
rect 2829 3383 2835 3436
rect 2829 3377 2851 3383
rect 2669 3317 2684 3323
rect 2621 3144 2627 3236
rect 2669 3124 2675 3236
rect 2381 2924 2387 2956
rect 2397 2944 2403 3036
rect 2445 2944 2451 2976
rect 2461 2964 2467 3036
rect 2349 2864 2355 2876
rect 2285 2804 2291 2836
rect 2333 2704 2339 2836
rect 2445 2764 2451 2916
rect 2461 2904 2467 2916
rect 2477 2904 2483 3056
rect 2557 2964 2563 2996
rect 2573 2884 2579 2896
rect 2589 2764 2595 3076
rect 2653 3064 2659 3076
rect 2685 2944 2691 3256
rect 2717 3184 2723 3236
rect 2765 3184 2771 3316
rect 2765 3104 2771 3136
rect 2701 3083 2707 3096
rect 2733 3084 2739 3096
rect 2701 3077 2716 3083
rect 2733 2984 2739 3036
rect 2781 2944 2787 3136
rect 2797 3084 2803 3196
rect 2813 3103 2819 3236
rect 2829 3104 2835 3116
rect 2813 3097 2828 3103
rect 2797 3064 2803 3076
rect 2813 2924 2819 3036
rect 2781 2903 2787 2916
rect 2781 2897 2796 2903
rect 2829 2903 2835 2976
rect 2845 2963 2851 3377
rect 2845 2957 2860 2963
rect 2877 2924 2883 3436
rect 2893 3104 2899 3576
rect 2938 3414 2950 3416
rect 2923 3406 2925 3414
rect 2933 3406 2935 3414
rect 2943 3406 2945 3414
rect 2953 3406 2955 3414
rect 2963 3406 2965 3414
rect 2938 3404 2950 3406
rect 2909 3324 2915 3376
rect 2989 3344 2995 3476
rect 2941 3324 2947 3336
rect 3021 3304 3027 3716
rect 3037 3704 3043 3716
rect 3053 3224 3059 3494
rect 3085 3484 3091 3716
rect 3165 3443 3171 3736
rect 3213 3504 3219 3876
rect 3261 3744 3267 3776
rect 3277 3744 3283 4216
rect 3325 4164 3331 4276
rect 3357 4184 3363 4496
rect 3389 4404 3395 4536
rect 3517 4443 3523 4536
rect 3517 4437 3539 4443
rect 3373 4302 3379 4316
rect 3469 4304 3475 4316
rect 3405 4264 3411 4276
rect 3437 4164 3443 4296
rect 3501 4244 3507 4256
rect 3325 4126 3331 4136
rect 3389 4124 3395 4136
rect 3437 4104 3443 4136
rect 3469 4124 3475 4176
rect 3485 4144 3491 4156
rect 3501 4143 3507 4236
rect 3501 4137 3523 4143
rect 3373 3904 3379 3936
rect 3300 3897 3315 3903
rect 3309 3784 3315 3897
rect 3373 3764 3379 3896
rect 3229 3704 3235 3716
rect 3165 3437 3180 3443
rect 3165 3324 3171 3336
rect 3181 3324 3187 3436
rect 3213 3344 3219 3496
rect 3229 3404 3235 3696
rect 3277 3604 3283 3716
rect 3165 3184 3171 3316
rect 3261 3184 3267 3596
rect 3293 3584 3299 3736
rect 3405 3724 3411 3776
rect 3421 3724 3427 4096
rect 3437 3984 3443 4076
rect 3485 4064 3491 4136
rect 3517 4124 3523 4137
rect 3501 4024 3507 4116
rect 3533 3984 3539 4437
rect 3549 4304 3555 4456
rect 3565 4124 3571 4296
rect 3597 4284 3603 4436
rect 3629 4304 3635 4356
rect 3645 4324 3651 4536
rect 3661 4504 3667 4516
rect 3613 4244 3619 4296
rect 3645 4284 3651 4316
rect 3597 4124 3603 4136
rect 3613 4024 3619 4116
rect 3645 4104 3651 4276
rect 3661 4124 3667 4236
rect 3677 4124 3683 4556
rect 3693 4244 3699 4676
rect 3709 4564 3715 4696
rect 3725 4564 3731 4636
rect 3757 4524 3763 4916
rect 3773 4824 3779 4916
rect 3821 4904 3827 4916
rect 3805 4704 3811 4776
rect 3821 4684 3827 4716
rect 3837 4704 3843 4916
rect 3853 4884 3859 4936
rect 3869 4924 3875 4957
rect 3780 4677 3804 4683
rect 3837 4664 3843 4696
rect 3773 4644 3779 4656
rect 3837 4584 3843 4616
rect 3853 4604 3859 4696
rect 3885 4624 3891 4656
rect 3901 4604 3907 4976
rect 3917 4704 3923 5216
rect 3933 5104 3939 5116
rect 3933 5084 3939 5096
rect 3965 5084 3971 5096
rect 3981 5064 3987 5076
rect 3997 5044 4003 5096
rect 4013 5084 4019 5096
rect 3940 4937 3964 4943
rect 3981 4884 3987 4896
rect 3933 4624 3939 4836
rect 3965 4704 3971 4856
rect 3981 4724 3987 4836
rect 3981 4704 3987 4716
rect 3965 4684 3971 4696
rect 3981 4663 3987 4696
rect 3997 4684 4003 4956
rect 4029 4944 4035 5016
rect 4045 4944 4051 5196
rect 4093 5184 4099 5276
rect 4237 5264 4243 5336
rect 4397 5304 4403 5316
rect 4237 5244 4243 5256
rect 4237 5204 4243 5236
rect 4141 5144 4147 5156
rect 4157 5124 4163 5156
rect 4093 5084 4099 5096
rect 4061 4924 4067 4936
rect 4077 4844 4083 5076
rect 4189 5064 4195 5076
rect 4109 4964 4115 5056
rect 4221 4983 4227 5136
rect 4253 5064 4259 5076
rect 4285 5064 4291 5156
rect 4301 5084 4307 5096
rect 4237 4984 4243 5016
rect 4205 4977 4227 4983
rect 4093 4884 4099 4896
rect 4061 4824 4067 4836
rect 4045 4764 4051 4816
rect 4109 4784 4115 4956
rect 4132 4917 4140 4923
rect 4125 4844 4131 4916
rect 4141 4884 4147 4896
rect 4157 4884 4163 4936
rect 4205 4924 4211 4977
rect 4228 4937 4243 4943
rect 4221 4904 4227 4916
rect 4173 4764 4179 4836
rect 4237 4824 4243 4937
rect 4253 4924 4259 5056
rect 4317 4964 4323 5076
rect 4333 4984 4339 5096
rect 4349 4984 4355 5096
rect 4013 4704 4019 4716
rect 4013 4663 4019 4696
rect 4061 4684 4067 4696
rect 4093 4684 4099 4736
rect 3965 4657 3987 4663
rect 3997 4657 4019 4663
rect 3933 4544 3939 4616
rect 3805 4524 3811 4536
rect 3949 4524 3955 4636
rect 3757 4384 3763 4516
rect 3757 4304 3763 4356
rect 3773 4324 3779 4496
rect 3789 4304 3795 4376
rect 3805 4364 3811 4516
rect 3869 4317 3884 4323
rect 3709 4284 3715 4296
rect 3773 4284 3779 4296
rect 3741 4144 3747 4236
rect 3821 4204 3827 4256
rect 3821 4164 3827 4196
rect 3565 3904 3571 4016
rect 3677 4004 3683 4116
rect 3725 4084 3731 4116
rect 3453 3884 3459 3896
rect 3453 3724 3459 3736
rect 3469 3724 3475 3896
rect 3549 3884 3555 3896
rect 3549 3784 3555 3876
rect 3501 3724 3507 3776
rect 3549 3724 3555 3736
rect 3565 3724 3571 3896
rect 3581 3864 3587 3876
rect 3629 3864 3635 3916
rect 3581 3744 3587 3856
rect 3341 3584 3347 3716
rect 3565 3684 3571 3716
rect 3309 3444 3315 3496
rect 3325 3484 3331 3576
rect 3373 3504 3379 3576
rect 3437 3524 3443 3636
rect 3501 3504 3507 3676
rect 3533 3504 3539 3516
rect 3405 3464 3411 3496
rect 3293 3424 3299 3436
rect 3405 3424 3411 3456
rect 3405 3324 3411 3416
rect 3453 3364 3459 3496
rect 3549 3483 3555 3556
rect 3565 3504 3571 3616
rect 3581 3504 3587 3716
rect 3597 3564 3603 3636
rect 3613 3624 3619 3796
rect 3629 3744 3635 3836
rect 3645 3744 3651 3856
rect 3661 3804 3667 3836
rect 3597 3484 3603 3516
rect 3613 3504 3619 3536
rect 3549 3477 3580 3483
rect 3629 3483 3635 3696
rect 3645 3524 3651 3736
rect 3661 3724 3667 3756
rect 3613 3477 3635 3483
rect 3453 3324 3459 3356
rect 3485 3324 3491 3476
rect 3517 3464 3523 3476
rect 3613 3464 3619 3477
rect 3645 3463 3651 3496
rect 3661 3484 3667 3536
rect 3677 3504 3683 3996
rect 3725 3904 3731 3916
rect 3757 3904 3763 4036
rect 3773 3984 3779 4036
rect 3693 3864 3699 3876
rect 3709 3763 3715 3836
rect 3693 3757 3715 3763
rect 3693 3724 3699 3757
rect 3725 3744 3731 3776
rect 3709 3564 3715 3676
rect 3709 3503 3715 3556
rect 3700 3497 3715 3503
rect 3677 3464 3683 3476
rect 3741 3464 3747 3776
rect 3773 3683 3779 3896
rect 3757 3677 3779 3683
rect 3757 3483 3763 3677
rect 3789 3664 3795 4076
rect 3837 4064 3843 4276
rect 3853 4163 3859 4296
rect 3869 4184 3875 4317
rect 3917 4304 3923 4336
rect 3901 4244 3907 4296
rect 3853 4157 3875 4163
rect 3805 3824 3811 3896
rect 3821 3783 3827 3956
rect 3837 3884 3843 3936
rect 3853 3924 3859 4116
rect 3869 4104 3875 4157
rect 3901 4144 3907 4236
rect 3965 4124 3971 4657
rect 3981 4184 3987 4196
rect 3876 4097 3891 4103
rect 3885 3984 3891 4097
rect 3805 3777 3827 3783
rect 3805 3724 3811 3777
rect 3821 3744 3827 3756
rect 3805 3704 3811 3716
rect 3821 3704 3827 3736
rect 3773 3504 3779 3536
rect 3757 3477 3779 3483
rect 3645 3457 3667 3463
rect 3501 3324 3507 3356
rect 2925 3084 2931 3116
rect 3261 3104 3267 3176
rect 3277 3124 3283 3316
rect 3293 3144 3299 3316
rect 3373 3104 3379 3236
rect 3437 3204 3443 3236
rect 2989 3084 2995 3096
rect 2973 3064 2979 3076
rect 3133 3044 3139 3096
rect 3245 3044 3251 3076
rect 2938 3014 2950 3016
rect 2923 3006 2925 3014
rect 2933 3006 2935 3014
rect 2943 3006 2945 3014
rect 2953 3006 2955 3014
rect 2963 3006 2965 3014
rect 2938 3004 2950 3006
rect 2829 2897 2851 2903
rect 2829 2824 2835 2876
rect 2189 2543 2195 2636
rect 2253 2544 2259 2556
rect 2189 2537 2211 2543
rect 2205 2504 2211 2537
rect 2301 2543 2307 2636
rect 2285 2537 2307 2543
rect 2317 2543 2323 2656
rect 2333 2564 2339 2576
rect 2317 2537 2339 2543
rect 2221 2484 2227 2496
rect 2157 2477 2172 2483
rect 2109 2184 2115 2456
rect 2125 2404 2131 2436
rect 2141 2104 2147 2296
rect 2173 2264 2179 2336
rect 2189 2303 2195 2436
rect 2221 2324 2227 2396
rect 2237 2384 2243 2416
rect 2189 2297 2204 2303
rect 2157 2144 2163 2236
rect 2029 1984 2035 2096
rect 2189 2064 2195 2236
rect 2205 2164 2211 2256
rect 2237 2244 2243 2296
rect 2253 2184 2259 2336
rect 2269 2324 2275 2496
rect 2285 2484 2291 2537
rect 2301 2464 2307 2516
rect 2301 2424 2307 2436
rect 2333 2384 2339 2537
rect 2349 2504 2355 2576
rect 2381 2544 2387 2676
rect 2477 2584 2483 2676
rect 2493 2584 2499 2656
rect 2509 2604 2515 2736
rect 2605 2684 2611 2696
rect 2813 2684 2819 2736
rect 2701 2664 2707 2676
rect 2701 2624 2707 2656
rect 2685 2584 2691 2596
rect 2717 2584 2723 2676
rect 2429 2544 2435 2576
rect 2669 2564 2675 2576
rect 2749 2544 2755 2636
rect 2845 2584 2851 2897
rect 2781 2544 2787 2576
rect 2877 2564 2883 2636
rect 2381 2504 2387 2536
rect 2429 2524 2435 2536
rect 2525 2504 2531 2536
rect 2205 2124 2211 2136
rect 2221 2084 2227 2096
rect 1965 1924 1971 1936
rect 2077 1904 2083 2036
rect 2093 1904 2099 2056
rect 2109 1984 2115 2036
rect 2189 1944 2195 2036
rect 2253 2023 2259 2136
rect 2285 2104 2291 2316
rect 2301 2304 2307 2316
rect 2317 2224 2323 2336
rect 2349 2324 2355 2476
rect 2333 2143 2339 2276
rect 2349 2264 2355 2316
rect 2333 2137 2348 2143
rect 2301 2124 2307 2136
rect 2253 2017 2275 2023
rect 2045 1884 2051 1896
rect 1997 1864 2003 1876
rect 1949 1724 1955 1796
rect 1965 1704 1971 1816
rect 2013 1724 2019 1796
rect 2061 1744 2067 1856
rect 2077 1724 2083 1796
rect 2125 1784 2131 1936
rect 2141 1844 2147 1896
rect 2269 1884 2275 2017
rect 2301 1944 2307 2036
rect 2301 1884 2307 1916
rect 2317 1904 2323 2076
rect 2349 1943 2355 2136
rect 2365 2104 2371 2356
rect 2381 2284 2387 2336
rect 2397 2284 2403 2436
rect 2509 2304 2515 2316
rect 2525 2284 2531 2496
rect 2541 2304 2547 2536
rect 2589 2324 2595 2516
rect 2589 2304 2595 2316
rect 2653 2304 2659 2536
rect 2701 2364 2707 2516
rect 2749 2384 2755 2516
rect 2893 2304 2899 2936
rect 2957 2684 2963 2836
rect 2938 2614 2950 2616
rect 2923 2606 2925 2614
rect 2933 2606 2935 2614
rect 2943 2606 2945 2614
rect 2953 2606 2955 2614
rect 2963 2606 2965 2614
rect 2938 2604 2950 2606
rect 2989 2584 2995 2676
rect 3037 2663 3043 2836
rect 3117 2744 3123 3036
rect 3181 2926 3187 2936
rect 3213 2904 3219 2936
rect 3245 2904 3251 3036
rect 3261 2984 3267 3036
rect 3277 2944 3283 3056
rect 3293 2884 3299 2936
rect 3325 2903 3331 3096
rect 3389 3044 3395 3094
rect 3453 3084 3459 3276
rect 3485 3204 3491 3316
rect 3517 3284 3523 3456
rect 3661 3443 3667 3457
rect 3693 3443 3699 3456
rect 3661 3437 3699 3443
rect 3469 3104 3475 3196
rect 3421 2944 3427 3056
rect 3453 2984 3459 3076
rect 3485 3064 3491 3076
rect 3501 2984 3507 3216
rect 3517 3164 3523 3236
rect 3533 3164 3539 3436
rect 3549 3324 3555 3376
rect 3613 3364 3619 3436
rect 3693 3384 3699 3416
rect 3741 3403 3747 3456
rect 3741 3397 3763 3403
rect 3677 3377 3692 3383
rect 3677 3364 3683 3377
rect 3645 3324 3651 3336
rect 3565 3224 3571 3316
rect 3645 3204 3651 3316
rect 3517 3024 3523 3096
rect 3533 2984 3539 3116
rect 3565 3104 3571 3196
rect 3661 3104 3667 3156
rect 3677 3104 3683 3156
rect 3693 3104 3699 3336
rect 3725 3124 3731 3396
rect 3725 3104 3731 3116
rect 3581 3044 3587 3076
rect 3565 2944 3571 2956
rect 3581 2944 3587 3036
rect 3597 2944 3603 3076
rect 3613 3064 3619 3096
rect 3693 3084 3699 3096
rect 3741 3084 3747 3116
rect 3757 3064 3763 3397
rect 3773 3224 3779 3477
rect 3789 3464 3795 3496
rect 3821 3464 3827 3616
rect 3869 3503 3875 3596
rect 3917 3564 3923 4116
rect 3949 3904 3955 3936
rect 3965 3864 3971 4096
rect 3997 3964 4003 4657
rect 4173 4624 4179 4696
rect 4061 4464 4067 4556
rect 4077 4544 4083 4596
rect 4205 4584 4211 4696
rect 4317 4684 4323 4916
rect 4365 4904 4371 4918
rect 4397 4744 4403 5296
rect 4445 5284 4451 5336
rect 4637 5284 4643 5336
rect 4442 5214 4454 5216
rect 4427 5206 4429 5214
rect 4437 5206 4439 5214
rect 4447 5206 4449 5214
rect 4457 5206 4459 5214
rect 4467 5206 4469 5214
rect 4442 5204 4454 5206
rect 4637 5144 4643 5176
rect 4413 5084 4419 5136
rect 4509 5104 4515 5136
rect 4541 4963 4547 5016
rect 4557 4984 4563 5096
rect 4541 4957 4563 4963
rect 4493 4944 4499 4956
rect 4557 4944 4563 4957
rect 4573 4944 4579 5096
rect 4573 4923 4579 4936
rect 4589 4924 4595 5076
rect 4557 4917 4579 4923
rect 4493 4883 4499 4916
rect 4493 4877 4515 4883
rect 4442 4814 4454 4816
rect 4427 4806 4429 4814
rect 4437 4806 4439 4814
rect 4447 4806 4449 4814
rect 4457 4806 4459 4814
rect 4467 4806 4469 4814
rect 4442 4804 4454 4806
rect 4189 4544 4195 4556
rect 4077 4524 4083 4536
rect 4013 4284 4019 4296
rect 4061 4264 4067 4276
rect 4061 4124 4067 4256
rect 4109 4244 4115 4516
rect 4125 4464 4131 4536
rect 4157 4524 4163 4536
rect 4237 4524 4243 4556
rect 4173 4404 4179 4516
rect 4237 4504 4243 4516
rect 4173 4364 4179 4396
rect 4125 4244 4131 4296
rect 4141 4204 4147 4316
rect 4157 4183 4163 4236
rect 4141 4177 4163 4183
rect 4109 4126 4115 4136
rect 4013 3943 4019 4076
rect 3997 3937 4019 3943
rect 3997 3884 4003 3937
rect 3933 3584 3939 3696
rect 3949 3684 3955 3716
rect 3965 3604 3971 3836
rect 4029 3764 4035 3876
rect 4029 3584 4035 3716
rect 4045 3704 4051 3716
rect 3997 3504 4003 3556
rect 3869 3497 3884 3503
rect 3869 3444 3875 3497
rect 3901 3484 3907 3496
rect 3885 3464 3891 3476
rect 3853 3344 3859 3376
rect 3789 3084 3795 3316
rect 3805 3284 3811 3316
rect 3885 3283 3891 3456
rect 3917 3424 3923 3496
rect 3949 3464 3955 3496
rect 3901 3324 3907 3356
rect 3949 3324 3955 3396
rect 3965 3344 3971 3496
rect 3981 3364 3987 3496
rect 4013 3424 4019 3496
rect 4029 3424 4035 3536
rect 4061 3523 4067 3936
rect 4093 3884 4099 3916
rect 4109 3884 4115 4016
rect 4141 3904 4147 4177
rect 4173 4104 4179 4316
rect 4189 4304 4195 4476
rect 4253 4304 4259 4596
rect 4301 4524 4307 4556
rect 4189 4244 4195 4296
rect 4237 4244 4243 4296
rect 4285 4264 4291 4336
rect 4157 3904 4163 4036
rect 4221 3984 4227 4076
rect 4237 4064 4243 4136
rect 4260 4117 4275 4123
rect 4237 4024 4243 4056
rect 4253 3924 4259 4096
rect 4269 4064 4275 4117
rect 4285 4084 4291 4236
rect 4333 4164 4339 4336
rect 4349 4304 4355 4536
rect 4365 4524 4371 4576
rect 4381 4424 4387 4616
rect 4413 4584 4419 4676
rect 4477 4564 4483 4636
rect 4445 4524 4451 4556
rect 4461 4464 4467 4516
rect 4493 4444 4499 4736
rect 4397 4437 4412 4443
rect 4365 4284 4371 4316
rect 4381 4304 4387 4416
rect 4397 4323 4403 4437
rect 4442 4414 4454 4416
rect 4427 4406 4429 4414
rect 4437 4406 4439 4414
rect 4447 4406 4449 4414
rect 4457 4406 4459 4414
rect 4467 4406 4469 4414
rect 4442 4404 4454 4406
rect 4493 4364 4499 4396
rect 4397 4317 4419 4323
rect 4397 4244 4403 4296
rect 4397 4144 4403 4156
rect 4301 4124 4307 4136
rect 4333 4004 4339 4116
rect 4141 3864 4147 3876
rect 4077 3724 4083 3776
rect 4093 3744 4099 3796
rect 4109 3744 4115 3856
rect 4173 3744 4179 3756
rect 4189 3744 4195 3836
rect 4205 3723 4211 3916
rect 4253 3904 4259 3916
rect 4196 3717 4211 3723
rect 4221 3877 4236 3883
rect 4173 3703 4179 3716
rect 4221 3703 4227 3877
rect 4253 3804 4259 3836
rect 4269 3824 4275 3896
rect 4285 3803 4291 3896
rect 4301 3824 4307 3876
rect 4285 3797 4307 3803
rect 4237 3724 4243 3756
rect 4269 3724 4275 3776
rect 4285 3704 4291 3736
rect 4173 3697 4195 3703
rect 4221 3697 4243 3703
rect 4189 3684 4195 3697
rect 4045 3517 4067 3523
rect 4045 3364 4051 3517
rect 4061 3344 4067 3496
rect 4077 3383 4083 3656
rect 4141 3584 4147 3616
rect 4125 3504 4131 3516
rect 4077 3377 4099 3383
rect 3869 3277 3891 3283
rect 3853 3124 3859 3196
rect 3869 3184 3875 3277
rect 3965 3264 3971 3316
rect 3997 3304 4003 3316
rect 4029 3284 4035 3316
rect 3853 3104 3859 3116
rect 3837 3044 3843 3096
rect 3341 2924 3347 2936
rect 3389 2924 3395 2936
rect 3405 2924 3411 2936
rect 3316 2897 3331 2903
rect 3021 2657 3043 2663
rect 3005 2564 3011 2636
rect 2925 2484 2931 2496
rect 2653 2284 2659 2296
rect 2669 2284 2675 2296
rect 2397 2144 2403 2176
rect 2413 2164 2419 2236
rect 2493 2204 2499 2256
rect 2541 2244 2547 2256
rect 2445 2124 2451 2196
rect 2653 2184 2659 2236
rect 2717 2184 2723 2196
rect 2829 2184 2835 2256
rect 2973 2244 2979 2536
rect 2989 2384 2995 2536
rect 3021 2463 3027 2657
rect 3053 2644 3059 2656
rect 3101 2584 3107 2696
rect 3133 2684 3139 2696
rect 3229 2684 3235 2876
rect 3261 2684 3267 2696
rect 3133 2564 3139 2676
rect 3164 2664 3172 2670
rect 3037 2504 3043 2536
rect 3037 2484 3043 2496
rect 3021 2457 3043 2463
rect 3021 2404 3027 2436
rect 2989 2324 2995 2376
rect 3021 2304 3027 2316
rect 3037 2304 3043 2457
rect 3053 2344 3059 2416
rect 3069 2384 3075 2516
rect 3085 2304 3091 2416
rect 3117 2384 3123 2476
rect 3133 2384 3139 2536
rect 3229 2524 3235 2676
rect 3245 2484 3251 2676
rect 3277 2526 3283 2576
rect 3309 2544 3315 2896
rect 3341 2724 3347 2896
rect 3357 2704 3363 2736
rect 3469 2724 3475 2896
rect 3501 2784 3507 2936
rect 3517 2924 3523 2936
rect 3325 2584 3331 2636
rect 3373 2564 3379 2676
rect 3149 2424 3155 2436
rect 3133 2324 3139 2336
rect 3005 2297 3020 2303
rect 2861 2224 2867 2236
rect 2938 2214 2950 2216
rect 2923 2206 2925 2214
rect 2933 2206 2935 2214
rect 2943 2206 2945 2214
rect 2953 2206 2955 2214
rect 2963 2206 2965 2214
rect 2938 2204 2950 2206
rect 2637 2144 2643 2156
rect 2797 2144 2803 2176
rect 2516 2137 2540 2143
rect 2605 2124 2611 2136
rect 2397 2104 2403 2116
rect 2541 2104 2547 2116
rect 2621 2104 2627 2136
rect 2685 2124 2691 2136
rect 2685 2083 2691 2116
rect 2685 2077 2707 2083
rect 2429 2064 2435 2076
rect 2445 2024 2451 2036
rect 2445 1984 2451 1996
rect 2349 1937 2371 1943
rect 2349 1904 2355 1916
rect 2285 1844 2291 1876
rect 2349 1864 2355 1896
rect 2205 1824 2211 1836
rect 2317 1804 2323 1836
rect 2109 1744 2115 1776
rect 2205 1744 2211 1796
rect 2029 1704 2035 1716
rect 2100 1697 2108 1703
rect 1853 1504 1859 1516
rect 1869 1484 1875 1556
rect 1917 1503 1923 1636
rect 1981 1524 1987 1636
rect 1997 1504 2003 1676
rect 2077 1504 2083 1636
rect 2157 1584 2163 1716
rect 2221 1684 2227 1716
rect 2237 1684 2243 1716
rect 2116 1537 2172 1543
rect 1908 1497 1923 1503
rect 1885 1484 1891 1496
rect 1805 1424 1811 1456
rect 1789 1324 1795 1336
rect 1764 1317 1779 1323
rect 1773 1304 1779 1317
rect 1821 1283 1827 1436
rect 1933 1383 1939 1436
rect 1917 1377 1939 1383
rect 1837 1344 1843 1376
rect 1876 1317 1891 1323
rect 1885 1304 1891 1317
rect 1917 1284 1923 1377
rect 1812 1277 1827 1283
rect 1725 1124 1731 1216
rect 1757 1184 1763 1256
rect 1677 1084 1683 1096
rect 1709 1064 1715 1096
rect 1757 1064 1763 1096
rect 1773 1084 1779 1156
rect 1789 1063 1795 1096
rect 1805 1084 1811 1096
rect 1821 1064 1827 1236
rect 1844 1157 1875 1163
rect 1853 1104 1859 1136
rect 1869 1084 1875 1157
rect 1789 1057 1811 1063
rect 1677 864 1683 916
rect 1693 904 1699 1056
rect 1805 1043 1811 1057
rect 1805 1037 1827 1043
rect 1709 977 1811 983
rect 1709 944 1715 977
rect 1805 964 1811 977
rect 1725 924 1731 956
rect 1741 824 1747 936
rect 1757 784 1763 916
rect 1789 904 1795 956
rect 1821 924 1827 1037
rect 1853 863 1859 896
rect 1869 884 1875 916
rect 1885 904 1891 1216
rect 1908 1117 1939 1123
rect 1933 1104 1939 1117
rect 1949 1104 1955 1476
rect 1981 1344 1987 1436
rect 2045 1384 2051 1476
rect 2061 1344 2067 1376
rect 2077 1324 2083 1456
rect 2093 1384 2099 1516
rect 2125 1444 2131 1456
rect 2157 1384 2163 1496
rect 2205 1444 2211 1556
rect 2221 1524 2227 1676
rect 2237 1523 2243 1636
rect 2253 1544 2259 1736
rect 2333 1724 2339 1756
rect 2365 1744 2371 1937
rect 2397 1904 2403 1936
rect 2381 1864 2387 1896
rect 2413 1884 2419 1916
rect 2637 1904 2643 2036
rect 2653 1904 2659 2016
rect 2669 1924 2675 1976
rect 2477 1884 2483 1896
rect 2445 1864 2451 1876
rect 2381 1724 2387 1756
rect 2445 1744 2451 1776
rect 2461 1724 2467 1876
rect 2493 1864 2499 1896
rect 2637 1884 2643 1896
rect 2653 1884 2659 1896
rect 2701 1884 2707 2077
rect 2781 1984 2787 2136
rect 2797 2044 2803 2136
rect 2893 2124 2899 2136
rect 3005 2124 3011 2297
rect 3037 2264 3043 2296
rect 2829 1984 2835 2096
rect 2893 2024 2899 2116
rect 3005 2104 3011 2116
rect 2781 1924 2787 1956
rect 2797 1904 2803 1956
rect 2589 1864 2595 1876
rect 2477 1824 2483 1856
rect 2573 1824 2579 1836
rect 2493 1764 2499 1816
rect 2605 1784 2611 1836
rect 2541 1744 2547 1776
rect 2669 1744 2675 1836
rect 2701 1824 2707 1876
rect 2717 1864 2723 1876
rect 2717 1784 2723 1836
rect 2781 1824 2787 1856
rect 2877 1844 2883 1996
rect 2909 1944 2915 2036
rect 3021 1984 3027 2136
rect 3085 2124 3091 2296
rect 3149 2184 3155 2296
rect 3037 2024 3043 2036
rect 2909 1884 2915 1936
rect 2925 1904 2931 1976
rect 2909 1864 2915 1876
rect 2925 1864 2931 1896
rect 2989 1884 2995 1956
rect 3037 1924 3043 1976
rect 3053 1904 3059 2036
rect 3085 1924 3091 2116
rect 3133 2044 3139 2116
rect 3165 2104 3171 2436
rect 3261 2284 3267 2294
rect 3325 2284 3331 2376
rect 3421 2324 3427 2716
rect 3485 2704 3491 2736
rect 3469 2684 3475 2696
rect 3453 2524 3459 2636
rect 3437 2304 3443 2356
rect 3469 2304 3475 2676
rect 3533 2624 3539 2916
rect 3565 2563 3571 2796
rect 3581 2704 3587 2916
rect 3565 2557 3580 2563
rect 3533 2324 3539 2436
rect 3373 2284 3379 2296
rect 3293 2264 3299 2276
rect 3389 2264 3395 2296
rect 3469 2264 3475 2276
rect 3293 2184 3299 2196
rect 3293 2144 3299 2176
rect 3373 2144 3379 2256
rect 3485 2184 3491 2236
rect 3501 2184 3507 2256
rect 3517 2204 3523 2276
rect 3533 2264 3539 2296
rect 3533 2183 3539 2256
rect 3565 2184 3571 2196
rect 3517 2177 3539 2183
rect 3181 2124 3187 2136
rect 3437 2126 3443 2176
rect 3469 2144 3475 2156
rect 3517 2124 3523 2177
rect 3149 2064 3155 2096
rect 3213 1984 3219 2056
rect 3357 1984 3363 1996
rect 3101 1864 3107 1896
rect 3133 1884 3139 1936
rect 2781 1764 2787 1816
rect 2938 1814 2950 1816
rect 2923 1806 2925 1814
rect 2933 1806 2935 1814
rect 2943 1806 2945 1814
rect 2953 1806 2955 1814
rect 2963 1806 2965 1814
rect 2938 1804 2950 1806
rect 3085 1784 3091 1856
rect 3181 1843 3187 1876
rect 3181 1837 3203 1843
rect 2685 1724 2691 1756
rect 2877 1744 2883 1756
rect 2669 1717 2684 1723
rect 2269 1544 2275 1716
rect 2237 1517 2259 1523
rect 2253 1383 2259 1517
rect 2269 1504 2275 1536
rect 2285 1504 2291 1516
rect 2237 1377 2259 1383
rect 2109 1344 2115 1376
rect 1965 1203 1971 1316
rect 1981 1224 1987 1296
rect 2004 1277 2028 1283
rect 2045 1263 2051 1296
rect 2061 1284 2067 1316
rect 2045 1257 2067 1263
rect 1997 1237 2012 1243
rect 1997 1203 2003 1237
rect 1965 1197 2003 1203
rect 1956 1077 1971 1083
rect 1933 1064 1939 1076
rect 1965 1064 1971 1077
rect 1901 964 1907 1036
rect 1917 1023 1923 1056
rect 1917 1017 1939 1023
rect 1917 963 1923 996
rect 1908 957 1923 963
rect 1933 943 1939 1017
rect 1933 937 1980 943
rect 1917 924 1923 936
rect 1933 904 1939 916
rect 1853 857 1932 863
rect 1805 784 1811 836
rect 1949 784 1955 916
rect 1965 744 1971 916
rect 1997 784 2003 896
rect 1693 603 1699 716
rect 1709 704 1715 716
rect 1709 624 1715 656
rect 1693 597 1715 603
rect 1709 584 1715 597
rect 1789 584 1795 716
rect 1853 704 1859 736
rect 1805 624 1811 656
rect 1741 544 1747 576
rect 1757 544 1763 576
rect 1805 564 1811 616
rect 1837 524 1843 696
rect 1933 624 1939 656
rect 1901 564 1907 596
rect 1949 524 1955 696
rect 1965 583 1971 736
rect 1981 704 1987 716
rect 2013 704 2019 1216
rect 2029 1084 2035 1156
rect 2045 1104 2051 1116
rect 2061 1083 2067 1257
rect 2045 1077 2067 1083
rect 2045 1064 2051 1077
rect 2077 1063 2083 1216
rect 2093 1104 2099 1296
rect 2125 1084 2131 1336
rect 2157 1104 2163 1216
rect 2068 1057 2083 1063
rect 2045 964 2051 996
rect 2077 984 2083 1036
rect 2061 884 2067 936
rect 2077 784 2083 916
rect 2093 744 2099 1076
rect 2109 944 2115 1056
rect 2173 984 2179 1316
rect 2221 1283 2227 1316
rect 2237 1304 2243 1377
rect 2253 1324 2259 1356
rect 2269 1324 2275 1476
rect 2317 1464 2323 1676
rect 2349 1664 2355 1676
rect 2333 1504 2339 1556
rect 2365 1524 2371 1536
rect 2381 1504 2387 1536
rect 2221 1277 2243 1283
rect 2237 1122 2243 1277
rect 2253 1264 2259 1296
rect 2269 1284 2275 1296
rect 2189 1084 2195 1116
rect 2212 1097 2275 1103
rect 2269 1064 2275 1097
rect 2212 1057 2252 1063
rect 2285 984 2291 1436
rect 2301 1384 2307 1436
rect 2317 1203 2323 1436
rect 2349 1364 2355 1416
rect 2365 1384 2371 1416
rect 2397 1404 2403 1536
rect 2445 1524 2451 1536
rect 2461 1517 2492 1523
rect 2429 1384 2435 1496
rect 2461 1484 2467 1517
rect 2541 1504 2547 1716
rect 2589 1504 2595 1516
rect 2477 1464 2483 1496
rect 2557 1444 2563 1476
rect 2621 1464 2627 1496
rect 2637 1444 2643 1496
rect 2653 1464 2659 1656
rect 2669 1504 2675 1717
rect 2829 1704 2835 1716
rect 2989 1704 2995 1756
rect 3005 1744 3011 1756
rect 3069 1744 3075 1776
rect 2333 1344 2339 1356
rect 2445 1344 2451 1356
rect 2317 1197 2339 1203
rect 2317 1104 2323 1176
rect 2333 1003 2339 1197
rect 2365 1184 2371 1236
rect 2397 1123 2403 1336
rect 2413 1324 2419 1336
rect 2381 1117 2403 1123
rect 2333 997 2355 1003
rect 2317 984 2323 996
rect 2189 944 2195 956
rect 2253 940 2259 956
rect 2269 944 2275 956
rect 2093 697 2108 703
rect 2029 664 2035 676
rect 2093 664 2099 697
rect 2125 683 2131 716
rect 2109 677 2131 683
rect 1965 577 1987 583
rect 1965 544 1971 556
rect 1981 524 1987 577
rect 2013 564 2019 596
rect 2061 584 2067 656
rect 2109 584 2115 677
rect 2093 564 2099 576
rect 2141 544 2147 556
rect 2157 524 2163 936
rect 2189 924 2195 936
rect 2205 844 2211 916
rect 2173 704 2179 716
rect 2205 704 2211 716
rect 2189 664 2195 676
rect 2221 524 2227 916
rect 2317 903 2323 916
rect 2333 904 2339 976
rect 2308 897 2323 903
rect 2349 883 2355 997
rect 2365 964 2371 996
rect 2381 924 2387 1117
rect 2397 1044 2403 1096
rect 2413 1064 2419 1096
rect 2429 1084 2435 1196
rect 2413 924 2419 1056
rect 2445 944 2451 1276
rect 2461 1204 2467 1436
rect 2477 1124 2483 1376
rect 2493 1340 2499 1416
rect 2509 1344 2515 1436
rect 2541 1344 2547 1376
rect 2557 1344 2563 1416
rect 2573 1364 2579 1436
rect 2669 1424 2675 1456
rect 2685 1444 2691 1476
rect 2701 1464 2707 1496
rect 2781 1403 2787 1676
rect 2797 1464 2803 1496
rect 2660 1397 2675 1403
rect 2781 1397 2803 1403
rect 2589 1364 2595 1376
rect 2589 1283 2595 1336
rect 2605 1324 2611 1356
rect 2653 1324 2659 1376
rect 2669 1324 2675 1397
rect 2701 1344 2707 1376
rect 2733 1344 2739 1356
rect 2589 1277 2636 1283
rect 2493 1104 2499 1116
rect 2477 1083 2483 1096
rect 2509 1083 2515 1116
rect 2525 1104 2531 1116
rect 2477 1077 2515 1083
rect 2573 1064 2579 1116
rect 2589 1084 2595 1196
rect 2644 1137 2659 1143
rect 2637 1084 2643 1116
rect 2653 1103 2659 1137
rect 2669 1124 2675 1196
rect 2653 1097 2668 1103
rect 2461 964 2467 1056
rect 2493 964 2499 976
rect 2525 964 2531 996
rect 2429 924 2435 936
rect 2388 917 2396 923
rect 2445 903 2451 916
rect 2436 897 2451 903
rect 2340 877 2355 883
rect 2349 784 2355 836
rect 2253 664 2259 716
rect 2429 684 2435 696
rect 2445 684 2451 796
rect 2461 784 2467 916
rect 2461 704 2467 736
rect 2477 704 2483 736
rect 2381 664 2387 676
rect 2493 664 2499 696
rect 2541 684 2547 716
rect 2237 564 2243 596
rect 2253 564 2259 596
rect 2285 544 2291 656
rect 1597 283 1603 316
rect 1613 304 1619 416
rect 1693 344 1699 436
rect 1629 297 1644 303
rect 1629 283 1635 297
rect 1725 303 1731 456
rect 1741 324 1747 496
rect 1837 424 1843 516
rect 1725 297 1747 303
rect 1597 277 1635 283
rect 1517 244 1523 276
rect 1549 184 1555 236
rect 1581 164 1587 196
rect 1693 184 1699 256
rect 1709 244 1715 276
rect 1709 164 1715 196
rect 1741 184 1747 297
rect 1789 283 1795 316
rect 1805 304 1811 416
rect 1853 324 1859 496
rect 1885 344 1891 496
rect 1853 297 1884 303
rect 1853 283 1859 297
rect 1789 277 1859 283
rect 1805 164 1811 196
rect 1645 144 1651 156
rect 1533 124 1539 136
rect 1629 124 1635 136
rect 1725 104 1731 156
rect 1757 144 1763 156
rect 1821 144 1827 256
rect 1837 224 1843 256
rect 1885 244 1891 276
rect 1917 264 1923 356
rect 1949 344 1955 516
rect 1981 364 1987 516
rect 2093 384 2099 416
rect 2157 324 2163 516
rect 1949 317 2051 323
rect 1949 304 1955 317
rect 2045 303 2051 317
rect 2116 317 2131 323
rect 2125 304 2131 317
rect 2173 304 2179 316
rect 2045 297 2092 303
rect 1997 284 2003 296
rect 2029 284 2035 296
rect 2157 284 2163 296
rect 2189 283 2195 316
rect 2221 304 2227 516
rect 2301 504 2307 516
rect 2301 464 2307 496
rect 2317 284 2323 536
rect 2333 524 2339 576
rect 2445 564 2451 656
rect 2525 564 2531 676
rect 2413 557 2428 563
rect 2349 524 2355 536
rect 2333 384 2339 516
rect 2413 284 2419 557
rect 2429 544 2435 556
rect 2509 544 2515 556
rect 2429 384 2435 516
rect 2493 444 2499 516
rect 2541 444 2547 516
rect 2557 504 2563 916
rect 2573 904 2579 976
rect 2685 964 2691 1336
rect 2717 1324 2723 1336
rect 2749 1304 2755 1316
rect 2765 1204 2771 1356
rect 2797 1324 2803 1397
rect 2829 1364 2835 1516
rect 2845 1484 2851 1696
rect 2893 1504 2899 1636
rect 2989 1464 2995 1696
rect 3005 1584 3011 1716
rect 3133 1704 3139 1756
rect 3165 1704 3171 1736
rect 3181 1724 3187 1736
rect 3053 1524 3059 1636
rect 3165 1584 3171 1696
rect 2861 1423 2867 1436
rect 2845 1417 2867 1423
rect 2845 1324 2851 1417
rect 2861 1384 2867 1396
rect 2877 1384 2883 1436
rect 2893 1364 2899 1456
rect 2938 1414 2950 1416
rect 2923 1406 2925 1414
rect 2933 1406 2935 1414
rect 2943 1406 2945 1414
rect 2953 1406 2955 1414
rect 2963 1406 2965 1414
rect 2938 1404 2950 1406
rect 2861 1324 2867 1356
rect 2909 1344 2915 1376
rect 2845 1303 2851 1316
rect 2845 1297 2860 1303
rect 2797 1217 2835 1223
rect 2797 1143 2803 1217
rect 2829 1204 2835 1217
rect 2877 1204 2883 1236
rect 2765 1137 2803 1143
rect 2765 1123 2771 1137
rect 2813 1124 2819 1196
rect 2861 1124 2867 1136
rect 2749 1117 2771 1123
rect 2749 1104 2755 1117
rect 2628 917 2643 923
rect 2605 723 2611 916
rect 2637 904 2643 917
rect 2621 844 2627 896
rect 2653 883 2659 916
rect 2637 877 2659 883
rect 2637 764 2643 877
rect 2589 717 2611 723
rect 2621 723 2627 736
rect 2653 723 2659 836
rect 2685 804 2691 896
rect 2701 803 2707 1036
rect 2733 984 2739 1076
rect 2749 1064 2755 1076
rect 2765 1064 2771 1096
rect 2845 1064 2851 1076
rect 2797 964 2803 1056
rect 2813 984 2819 1056
rect 2829 984 2835 1036
rect 2893 1024 2899 1196
rect 2941 1084 2947 1356
rect 3005 1143 3011 1516
rect 3021 1477 3036 1483
rect 3021 1244 3027 1477
rect 3053 1464 3059 1516
rect 3037 1324 3043 1416
rect 3085 1364 3091 1536
rect 3101 1504 3107 1576
rect 3181 1504 3187 1716
rect 3197 1704 3203 1837
rect 3229 1744 3235 1796
rect 3261 1744 3267 1756
rect 3213 1737 3228 1743
rect 3213 1584 3219 1737
rect 3277 1724 3283 1896
rect 3293 1884 3299 1956
rect 3389 1904 3395 1916
rect 3517 1904 3523 2116
rect 3581 2103 3587 2516
rect 3597 2484 3603 2936
rect 3629 2804 3635 3036
rect 3677 2964 3683 3036
rect 3821 3024 3827 3036
rect 3869 3024 3875 3176
rect 3885 3004 3891 3056
rect 3789 2984 3795 2996
rect 3645 2924 3651 2936
rect 3661 2904 3667 2916
rect 3709 2864 3715 2916
rect 3757 2864 3763 2936
rect 3901 2924 3907 3096
rect 3725 2724 3731 2836
rect 3629 2702 3635 2716
rect 3725 2684 3731 2696
rect 3661 2564 3667 2676
rect 3693 2584 3699 2656
rect 3789 2644 3795 2696
rect 3821 2684 3827 2876
rect 3917 2744 3923 3236
rect 3933 3084 3939 3116
rect 3949 3104 3955 3176
rect 3965 3164 3971 3256
rect 4061 3224 4067 3316
rect 4061 3144 4067 3156
rect 4045 3124 4051 3136
rect 4061 3104 4067 3136
rect 3949 3024 3955 3076
rect 3869 2704 3875 2716
rect 3949 2684 3955 3016
rect 3997 2924 4003 3096
rect 4045 2924 4051 2996
rect 3997 2704 4003 2736
rect 4029 2724 4035 2776
rect 3997 2684 4003 2696
rect 4045 2684 4051 2716
rect 3661 2544 3667 2556
rect 3597 2384 3603 2436
rect 3629 2304 3635 2316
rect 3677 2304 3683 2496
rect 3597 2124 3603 2236
rect 3581 2097 3603 2103
rect 3549 2064 3555 2096
rect 3581 1924 3587 2056
rect 3325 1804 3331 1856
rect 3373 1744 3379 1816
rect 3389 1784 3395 1876
rect 3421 1824 3427 1856
rect 3437 1744 3443 1796
rect 3261 1704 3267 1716
rect 3197 1504 3203 1576
rect 3213 1524 3219 1576
rect 3309 1544 3315 1636
rect 3389 1584 3395 1736
rect 3453 1724 3459 1856
rect 3501 1783 3507 1896
rect 3517 1824 3523 1876
rect 3533 1804 3539 1876
rect 3581 1864 3587 1916
rect 3501 1777 3516 1783
rect 3517 1764 3523 1776
rect 3565 1764 3571 1816
rect 3597 1744 3603 2097
rect 3645 1904 3651 2256
rect 3677 2144 3683 2156
rect 3693 2123 3699 2556
rect 3757 2524 3763 2636
rect 3821 2544 3827 2676
rect 3988 2577 4003 2583
rect 3997 2564 4003 2577
rect 3869 2524 3875 2556
rect 3997 2544 4003 2556
rect 4077 2544 4083 3116
rect 4093 3104 4099 3377
rect 4125 3184 4131 3436
rect 4141 3324 4147 3336
rect 4157 3324 4163 3636
rect 4205 3423 4211 3496
rect 4189 3417 4211 3423
rect 4189 3384 4195 3417
rect 4189 3324 4195 3376
rect 4157 3084 4163 3176
rect 4141 3024 4147 3076
rect 4189 2944 4195 3316
rect 4221 3084 4227 3096
rect 4093 2924 4099 2936
rect 4205 2924 4211 2956
rect 4221 2944 4227 2996
rect 4237 2884 4243 3697
rect 4285 3684 4291 3696
rect 4253 3464 4259 3496
rect 4301 3484 4307 3797
rect 4333 3744 4339 3816
rect 4349 3804 4355 3896
rect 4365 3784 4371 4116
rect 4381 4104 4387 4136
rect 4413 4123 4419 4317
rect 4445 4224 4451 4296
rect 4429 4124 4435 4156
rect 4404 4117 4419 4123
rect 4317 3724 4323 3736
rect 4381 3644 4387 4076
rect 4461 4044 4467 4236
rect 4442 4014 4454 4016
rect 4427 4006 4429 4014
rect 4437 4006 4439 4014
rect 4447 4006 4449 4014
rect 4457 4006 4459 4014
rect 4467 4006 4469 4014
rect 4442 4004 4454 4006
rect 4509 3984 4515 4877
rect 4541 4544 4547 4916
rect 4557 4784 4563 4917
rect 4589 4804 4595 4896
rect 4589 4704 4595 4716
rect 4589 4544 4595 4696
rect 4541 4384 4547 4536
rect 4605 4524 4611 5096
rect 4637 5044 4643 5136
rect 4685 5124 4691 5316
rect 4797 5164 4803 5236
rect 4685 5084 4691 5096
rect 4621 4924 4627 5016
rect 4685 4963 4691 5036
rect 4701 5004 4707 5076
rect 4733 5024 4739 5076
rect 4685 4957 4700 4963
rect 4749 4924 4755 4936
rect 4765 4924 4771 4956
rect 4637 4644 4643 4836
rect 4669 4824 4675 4916
rect 4669 4623 4675 4796
rect 4685 4664 4691 4916
rect 4733 4844 4739 4916
rect 4749 4884 4755 4896
rect 4733 4763 4739 4836
rect 4749 4784 4755 4876
rect 4765 4824 4771 4836
rect 4733 4757 4755 4763
rect 4749 4644 4755 4757
rect 4669 4617 4691 4623
rect 4637 4524 4643 4536
rect 4557 4364 4563 4456
rect 4557 4124 4563 4356
rect 4589 4344 4595 4476
rect 4637 4363 4643 4516
rect 4653 4404 4659 4536
rect 4621 4357 4643 4363
rect 4573 4164 4579 4296
rect 4589 4184 4595 4276
rect 4621 4124 4627 4357
rect 4685 4344 4691 4617
rect 4765 4604 4771 4796
rect 4781 4763 4787 5076
rect 4813 4964 4819 5336
rect 4877 5324 4883 5336
rect 4829 5264 4835 5316
rect 4877 5264 4883 5296
rect 4941 5284 4947 5336
rect 4925 4964 4931 5176
rect 5069 5084 5075 5276
rect 5101 5224 5107 5336
rect 5181 5324 5187 5336
rect 5181 5204 5187 5316
rect 5069 5064 5075 5076
rect 5101 5064 5107 5136
rect 5133 5104 5139 5176
rect 5181 5084 5187 5176
rect 5197 5044 5203 5096
rect 5229 5064 5235 5076
rect 5069 4977 5139 4983
rect 5069 4963 5075 4977
rect 5021 4957 5075 4963
rect 5085 4957 5116 4963
rect 5021 4943 5027 4957
rect 4989 4937 5027 4943
rect 4797 4844 4803 4916
rect 4813 4904 4819 4936
rect 4861 4924 4867 4936
rect 4797 4784 4803 4816
rect 4877 4804 4883 4916
rect 4893 4884 4899 4936
rect 4989 4924 4995 4937
rect 5085 4943 5091 4957
rect 5069 4937 5091 4943
rect 5037 4924 5043 4936
rect 5069 4924 5075 4937
rect 5101 4923 5107 4936
rect 5101 4917 5116 4923
rect 5021 4903 5027 4916
rect 5053 4904 5059 4916
rect 5005 4897 5027 4903
rect 4893 4824 4899 4876
rect 4909 4784 4915 4816
rect 4973 4764 4979 4836
rect 4781 4757 4803 4763
rect 4781 4684 4787 4696
rect 4637 4324 4643 4336
rect 4701 4324 4707 4376
rect 4733 4304 4739 4336
rect 4429 3824 4435 3836
rect 4413 3684 4419 3716
rect 4365 3584 4371 3636
rect 4442 3614 4454 3616
rect 4427 3606 4429 3614
rect 4437 3606 4439 3614
rect 4447 3606 4449 3614
rect 4457 3606 4459 3614
rect 4467 3606 4469 3614
rect 4442 3604 4454 3606
rect 4493 3604 4499 3856
rect 4509 3744 4515 3876
rect 4557 3804 4563 3894
rect 4589 3884 4595 3996
rect 4605 3944 4611 4056
rect 4621 4004 4627 4076
rect 4541 3726 4547 3756
rect 4637 3724 4643 4016
rect 4653 3984 4659 4296
rect 4749 4284 4755 4396
rect 4765 4384 4771 4596
rect 4669 4144 4675 4236
rect 4653 3904 4659 3976
rect 4669 3904 4675 4136
rect 4701 4124 4707 4236
rect 4717 4164 4723 4256
rect 4685 3783 4691 4116
rect 4717 3904 4723 4116
rect 4749 4084 4755 4276
rect 4781 4083 4787 4636
rect 4797 4584 4803 4757
rect 4925 4702 4931 4736
rect 4989 4684 4995 4876
rect 4797 4564 4803 4576
rect 4877 4544 4883 4576
rect 4925 4564 4931 4656
rect 5005 4624 5011 4897
rect 5085 4844 5091 4916
rect 5117 4904 5123 4916
rect 5133 4904 5139 4977
rect 5197 4964 5203 5036
rect 5149 4937 5164 4943
rect 5149 4884 5155 4937
rect 5172 4917 5187 4923
rect 5021 4704 5027 4716
rect 5021 4624 5027 4696
rect 5085 4684 5091 4776
rect 5085 4664 5091 4676
rect 4893 4304 4899 4316
rect 4925 4304 4931 4556
rect 4941 4524 4947 4536
rect 5005 4384 5011 4616
rect 5021 4344 5027 4616
rect 5053 4524 5059 4656
rect 5117 4604 5123 4696
rect 5149 4643 5155 4856
rect 5165 4704 5171 4716
rect 5181 4704 5187 4917
rect 5229 4784 5235 4836
rect 5277 4724 5283 5356
rect 5405 5344 5411 5376
rect 6013 5364 6019 5396
rect 5876 5357 5891 5363
rect 5293 5024 5299 5096
rect 5309 5084 5315 5336
rect 5405 5284 5411 5336
rect 5453 5244 5459 5356
rect 5501 5324 5507 5336
rect 5581 5326 5587 5336
rect 5629 5317 5644 5323
rect 5405 5144 5411 5196
rect 5501 5184 5507 5316
rect 5517 5163 5523 5316
rect 5501 5157 5523 5163
rect 5437 5137 5484 5143
rect 5309 4964 5315 5076
rect 5373 4964 5379 4976
rect 5405 4964 5411 5136
rect 5437 5084 5443 5137
rect 5453 5084 5459 5116
rect 5485 5104 5491 5116
rect 5501 5004 5507 5157
rect 5533 5137 5548 5143
rect 5533 5124 5539 5137
rect 5549 5104 5555 5116
rect 5517 5043 5523 5096
rect 5556 5077 5571 5083
rect 5517 5037 5539 5043
rect 5405 4924 5411 4956
rect 5453 4944 5459 4956
rect 5309 4884 5315 4918
rect 5277 4704 5283 4716
rect 5149 4637 5164 4643
rect 5117 4584 5123 4596
rect 5117 4564 5123 4576
rect 4829 4264 4835 4276
rect 4861 4124 4867 4236
rect 4877 4184 4883 4296
rect 5005 4284 5011 4336
rect 5037 4324 5043 4516
rect 5021 4303 5027 4316
rect 5021 4297 5043 4303
rect 5037 4284 5043 4297
rect 4925 4184 4931 4216
rect 4877 4143 4883 4156
rect 4877 4137 4892 4143
rect 4820 4117 4844 4123
rect 4765 4077 4787 4083
rect 4749 3984 4755 3996
rect 4765 3984 4771 4077
rect 4717 3884 4723 3896
rect 4749 3824 4755 3856
rect 4685 3777 4707 3783
rect 4605 3704 4611 3716
rect 4637 3703 4643 3716
rect 4621 3697 4643 3703
rect 4397 3504 4403 3536
rect 4349 3404 4355 3496
rect 4253 3284 4259 3316
rect 4269 3204 4275 3336
rect 4285 3324 4291 3396
rect 4365 3324 4371 3456
rect 4381 3344 4387 3356
rect 4333 3304 4339 3316
rect 4365 3184 4371 3256
rect 4253 3084 4259 3116
rect 4253 2944 4259 2956
rect 4093 2704 4099 2776
rect 4093 2644 4099 2676
rect 4109 2564 4115 2796
rect 4157 2724 4163 2836
rect 4125 2704 4131 2716
rect 4173 2684 4179 2696
rect 4173 2604 4179 2676
rect 4189 2604 4195 2876
rect 4269 2824 4275 2916
rect 4285 2903 4291 2976
rect 4349 2944 4355 3076
rect 4365 2924 4371 3176
rect 4381 3044 4387 3316
rect 4413 3264 4419 3496
rect 4429 3364 4435 3456
rect 4493 3364 4499 3596
rect 4525 3444 4531 3496
rect 4541 3484 4547 3676
rect 4621 3624 4627 3697
rect 4653 3604 4659 3736
rect 4701 3724 4707 3777
rect 4717 3744 4723 3756
rect 4733 3744 4739 3816
rect 4765 3803 4771 3936
rect 4781 3924 4787 4036
rect 4797 3944 4803 3976
rect 4813 3904 4819 4116
rect 4877 4004 4883 4137
rect 4893 4124 4899 4136
rect 4893 4004 4899 4096
rect 4893 3984 4899 3996
rect 4909 3964 4915 4136
rect 4925 4104 4931 4116
rect 4957 3963 4963 4256
rect 4973 4157 4988 4163
rect 4973 4124 4979 4157
rect 4996 4137 5020 4143
rect 4941 3957 4963 3963
rect 4893 3904 4899 3936
rect 4909 3904 4915 3916
rect 4797 3864 4803 3896
rect 4845 3824 4851 3876
rect 4749 3797 4771 3803
rect 4669 3684 4675 3696
rect 4749 3684 4755 3797
rect 4781 3784 4787 3796
rect 4829 3744 4835 3756
rect 4813 3704 4819 3716
rect 4708 3637 4723 3643
rect 4621 3524 4627 3536
rect 4589 3504 4595 3516
rect 4653 3504 4659 3516
rect 4557 3484 4563 3496
rect 4669 3484 4675 3616
rect 4685 3584 4691 3596
rect 4557 3384 4563 3396
rect 4429 3344 4435 3356
rect 4445 3304 4451 3336
rect 4397 3257 4412 3263
rect 4397 3224 4403 3257
rect 4493 3223 4499 3356
rect 4509 3344 4515 3356
rect 4493 3217 4515 3223
rect 4442 3214 4454 3216
rect 4427 3206 4429 3214
rect 4437 3206 4439 3214
rect 4447 3206 4449 3214
rect 4457 3206 4459 3214
rect 4467 3206 4469 3214
rect 4442 3204 4454 3206
rect 4445 3124 4451 3136
rect 4493 3084 4499 3196
rect 4308 2917 4323 2923
rect 4285 2897 4307 2903
rect 4221 2704 4227 2716
rect 4205 2683 4211 2696
rect 4205 2677 4227 2683
rect 4077 2524 4083 2536
rect 4205 2524 4211 2536
rect 4221 2524 4227 2677
rect 4237 2644 4243 2816
rect 4253 2724 4259 2736
rect 4269 2684 4275 2696
rect 4164 2517 4172 2523
rect 3709 2384 3715 2516
rect 4109 2484 4115 2516
rect 3949 2304 3955 2316
rect 3805 2277 3820 2283
rect 3805 2144 3811 2277
rect 3677 2117 3699 2123
rect 3661 1904 3667 1916
rect 3629 1884 3635 1896
rect 3469 1724 3475 1736
rect 3117 1484 3123 1496
rect 3053 1304 3059 1356
rect 3037 1244 3043 1296
rect 2957 1137 3011 1143
rect 2957 1104 2963 1137
rect 3005 1123 3011 1137
rect 3005 1117 3027 1123
rect 2973 1084 2979 1116
rect 3021 1103 3027 1117
rect 3021 1097 3036 1103
rect 2938 1014 2950 1016
rect 2923 1006 2925 1014
rect 2933 1006 2935 1014
rect 2943 1006 2945 1014
rect 2953 1006 2955 1014
rect 2963 1006 2965 1014
rect 2938 1004 2950 1006
rect 2845 963 2851 996
rect 2893 964 2899 996
rect 2813 957 2851 963
rect 2717 944 2723 956
rect 2813 903 2819 957
rect 2861 944 2867 956
rect 2797 897 2819 903
rect 2797 844 2803 897
rect 2701 797 2723 803
rect 2685 744 2691 796
rect 2621 717 2659 723
rect 2589 704 2595 717
rect 2605 684 2611 696
rect 2612 657 2620 663
rect 2605 544 2611 656
rect 2637 584 2643 676
rect 2669 664 2675 696
rect 2685 684 2691 716
rect 2701 704 2707 756
rect 2717 744 2723 797
rect 2797 704 2803 796
rect 2813 784 2819 836
rect 2829 724 2835 756
rect 2845 704 2851 916
rect 2861 844 2867 916
rect 2893 904 2899 936
rect 2877 784 2883 896
rect 2893 784 2899 836
rect 2909 804 2915 916
rect 2941 844 2947 896
rect 2877 704 2883 736
rect 2669 604 2675 656
rect 2717 584 2723 676
rect 2797 664 2803 676
rect 2733 564 2739 596
rect 2749 564 2755 636
rect 2180 277 2195 283
rect 2013 264 2019 276
rect 1933 244 1939 256
rect 1949 224 1955 256
rect 1917 164 1923 196
rect 1933 164 1939 196
rect 1821 124 1827 136
rect 1981 124 1987 256
rect 2013 184 2019 236
rect 2045 164 2051 196
rect 2077 184 2083 276
rect 2253 224 2259 256
rect 2109 184 2115 196
rect 2093 164 2099 176
rect 660 97 675 103
rect 13 84 19 96
rect 669 84 675 97
rect 1773 84 1779 116
rect 2109 104 2115 156
rect 2173 144 2179 196
rect 2317 163 2323 276
rect 2317 157 2332 163
rect 2333 144 2339 156
rect 2285 124 2291 136
rect 2349 104 2355 236
rect 2413 184 2419 276
rect 2445 264 2451 296
rect 2605 284 2611 456
rect 2461 244 2467 276
rect 2509 164 2515 176
rect 2429 124 2435 156
rect 2541 124 2547 236
rect 2557 184 2563 276
rect 2605 224 2611 276
rect 2621 264 2627 556
rect 2813 544 2819 556
rect 2845 544 2851 656
rect 2877 584 2883 616
rect 2893 604 2899 676
rect 2941 664 2947 696
rect 2938 614 2950 616
rect 2923 606 2925 614
rect 2933 606 2935 614
rect 2943 606 2945 614
rect 2953 606 2955 614
rect 2963 606 2965 614
rect 2938 604 2950 606
rect 2637 384 2643 516
rect 2653 464 2659 516
rect 2797 464 2803 516
rect 2829 504 2835 516
rect 2861 484 2867 516
rect 2893 344 2899 556
rect 2989 483 2995 1076
rect 3005 944 3011 1036
rect 3037 1003 3043 1056
rect 3053 1024 3059 1296
rect 3085 1283 3091 1316
rect 3101 1304 3107 1336
rect 3117 1283 3123 1396
rect 3085 1277 3123 1283
rect 3101 1104 3107 1196
rect 3133 1184 3139 1456
rect 3149 1344 3155 1416
rect 3197 1384 3203 1496
rect 3261 1464 3267 1476
rect 3357 1403 3363 1476
rect 3341 1397 3363 1403
rect 3277 1384 3283 1396
rect 3149 1304 3155 1316
rect 3133 1104 3139 1176
rect 3149 1104 3155 1196
rect 3165 1124 3171 1336
rect 3229 1284 3235 1296
rect 3117 1024 3123 1056
rect 3037 997 3059 1003
rect 3021 964 3027 996
rect 3053 964 3059 997
rect 3117 964 3123 1016
rect 3037 924 3043 936
rect 3053 924 3059 936
rect 3181 884 3187 1196
rect 3229 1104 3235 1116
rect 3197 944 3203 1016
rect 3229 984 3235 1056
rect 3229 964 3235 976
rect 3261 964 3267 1336
rect 3277 1024 3283 1076
rect 3277 984 3283 1016
rect 3005 804 3011 836
rect 3021 724 3027 736
rect 3005 624 3011 696
rect 3005 564 3011 616
rect 3037 584 3043 796
rect 3053 684 3059 716
rect 3101 704 3107 716
rect 3197 704 3203 796
rect 3213 704 3219 736
rect 3245 704 3251 756
rect 3277 744 3283 796
rect 3293 724 3299 1376
rect 3309 1344 3315 1396
rect 3341 1164 3347 1397
rect 3389 1384 3395 1476
rect 3405 1384 3411 1516
rect 3421 1484 3427 1716
rect 3485 1424 3491 1716
rect 3613 1504 3619 1836
rect 3629 1744 3635 1776
rect 3645 1564 3651 1716
rect 3661 1684 3667 1896
rect 3677 1784 3683 2117
rect 3693 1724 3699 1736
rect 3677 1644 3683 1656
rect 3661 1524 3667 1636
rect 3677 1604 3683 1636
rect 3709 1504 3715 1876
rect 3757 1864 3763 1916
rect 3725 1784 3731 1856
rect 3757 1804 3763 1836
rect 3773 1784 3779 1876
rect 3741 1724 3747 1756
rect 3789 1684 3795 1716
rect 3725 1604 3731 1636
rect 3725 1504 3731 1536
rect 3709 1484 3715 1496
rect 3613 1464 3619 1476
rect 3404 1350 3412 1356
rect 3373 1204 3379 1336
rect 3405 1117 3420 1123
rect 3309 924 3315 1116
rect 3405 1104 3411 1117
rect 3469 1104 3475 1276
rect 3485 1124 3491 1236
rect 3501 1204 3507 1416
rect 3549 1344 3555 1456
rect 3725 1444 3731 1476
rect 3597 1344 3603 1436
rect 3693 1364 3699 1436
rect 3773 1364 3779 1616
rect 3789 1524 3795 1596
rect 3805 1544 3811 1956
rect 3821 1864 3827 1916
rect 3837 1904 3843 2236
rect 3869 1944 3875 2296
rect 4077 2284 4083 2476
rect 4125 2324 4131 2436
rect 4173 2364 4179 2516
rect 4221 2504 4227 2516
rect 4205 2384 4211 2496
rect 4141 2304 4147 2316
rect 3933 2144 3939 2256
rect 3949 2184 3955 2196
rect 3885 1904 3891 1996
rect 3901 1924 3907 1936
rect 3917 1904 3923 2036
rect 3853 1723 3859 1836
rect 3917 1764 3923 1896
rect 3981 1784 3987 2116
rect 3997 2104 4003 2136
rect 3853 1717 3868 1723
rect 3821 1484 3827 1676
rect 3869 1584 3875 1696
rect 3949 1504 3955 1776
rect 3981 1724 3987 1756
rect 3837 1484 3843 1496
rect 3549 1284 3555 1316
rect 3501 1184 3507 1196
rect 3533 1184 3539 1196
rect 3549 1184 3555 1276
rect 3565 1204 3571 1316
rect 3581 1104 3587 1196
rect 3597 1184 3603 1336
rect 3613 1326 3619 1356
rect 3373 1084 3379 1096
rect 3332 1077 3347 1083
rect 3341 1064 3347 1077
rect 3389 1064 3395 1076
rect 3341 1024 3347 1036
rect 3405 984 3411 1096
rect 3437 1043 3443 1056
rect 3437 1037 3459 1043
rect 3357 977 3395 983
rect 3357 963 3363 977
rect 3341 957 3363 963
rect 3341 943 3347 957
rect 3325 937 3347 943
rect 3325 904 3331 937
rect 3341 904 3347 916
rect 3389 904 3395 977
rect 3421 964 3427 1036
rect 3437 884 3443 896
rect 3405 784 3411 876
rect 3453 764 3459 1037
rect 3501 944 3507 1016
rect 3517 1004 3523 1056
rect 3581 1044 3587 1096
rect 3549 944 3555 976
rect 3485 824 3491 836
rect 3485 724 3491 736
rect 3357 704 3363 716
rect 3213 677 3228 683
rect 3085 584 3091 676
rect 3101 584 3107 676
rect 3117 624 3123 636
rect 3085 544 3091 556
rect 3117 544 3123 556
rect 3028 537 3043 543
rect 2973 477 2995 483
rect 2861 317 2876 323
rect 2781 284 2787 316
rect 2813 284 2819 296
rect 2669 264 2675 276
rect 2621 164 2627 256
rect 2653 244 2659 256
rect 2861 244 2867 317
rect 2717 164 2723 216
rect 2797 204 2803 236
rect 2589 144 2595 156
rect 2829 144 2835 156
rect 2621 124 2627 136
rect 2877 124 2883 296
rect 2973 264 2979 477
rect 2989 264 2995 456
rect 3037 384 3043 537
rect 3069 524 3075 536
rect 3117 497 3132 503
rect 3117 484 3123 497
rect 3117 384 3123 476
rect 3165 464 3171 636
rect 3213 564 3219 677
rect 3261 624 3267 676
rect 3181 544 3187 556
rect 3181 504 3187 516
rect 3037 284 3043 336
rect 3165 304 3171 436
rect 3213 324 3219 536
rect 3261 344 3267 616
rect 3277 564 3283 676
rect 3293 584 3299 696
rect 3341 584 3347 676
rect 3325 544 3331 556
rect 3357 544 3363 696
rect 3373 684 3379 716
rect 3389 624 3395 716
rect 3405 684 3411 696
rect 3421 684 3427 696
rect 3437 663 3443 696
rect 3421 657 3443 663
rect 3389 563 3395 616
rect 3421 584 3427 657
rect 3389 557 3404 563
rect 3437 544 3443 556
rect 3277 524 3283 536
rect 3357 504 3363 516
rect 3357 384 3363 496
rect 3213 284 3219 316
rect 3261 304 3267 336
rect 3293 284 3299 316
rect 3309 284 3315 296
rect 3181 264 3187 276
rect 3213 264 3219 276
rect 3261 264 3267 276
rect 2938 214 2950 216
rect 2923 206 2925 214
rect 2933 206 2935 214
rect 2943 206 2945 214
rect 2953 206 2955 214
rect 2963 206 2965 214
rect 2938 204 2950 206
rect 2893 124 2899 196
rect 3005 184 3011 256
rect 2909 124 2915 136
rect 2365 104 2371 116
rect 2525 104 2531 116
rect 2637 104 2643 116
rect 3021 104 3027 116
rect 3053 104 3059 136
rect 3101 124 3107 236
rect 3181 164 3187 176
rect 3245 144 3251 156
rect 3309 144 3315 276
rect 3341 264 3347 296
rect 3405 284 3411 316
rect 3421 283 3427 436
rect 3453 304 3459 656
rect 3485 564 3491 636
rect 3501 344 3507 916
rect 3613 864 3619 1116
rect 3629 1104 3635 1236
rect 3645 1064 3651 1216
rect 3773 1184 3779 1356
rect 3805 1326 3811 1476
rect 3821 1403 3827 1476
rect 3901 1464 3907 1496
rect 3821 1397 3843 1403
rect 3837 1344 3843 1397
rect 3869 1384 3875 1396
rect 3949 1384 3955 1496
rect 3965 1484 3971 1636
rect 3981 1584 3987 1716
rect 3997 1644 4003 2096
rect 4013 2044 4019 2156
rect 4045 2124 4051 2156
rect 4125 2124 4131 2136
rect 4141 2044 4147 2296
rect 4173 2284 4179 2356
rect 4237 2304 4243 2636
rect 4285 2564 4291 2696
rect 4301 2684 4307 2897
rect 4317 2784 4323 2917
rect 4349 2904 4355 2916
rect 4333 2884 4339 2896
rect 4365 2864 4371 2916
rect 4317 2704 4323 2736
rect 4381 2704 4387 3036
rect 4509 2964 4515 3217
rect 4493 2824 4499 2916
rect 4442 2814 4454 2816
rect 4427 2806 4429 2814
rect 4437 2806 4439 2814
rect 4447 2806 4449 2814
rect 4457 2806 4459 2814
rect 4467 2806 4469 2814
rect 4442 2804 4454 2806
rect 4509 2784 4515 2796
rect 4525 2724 4531 3256
rect 4541 2884 4547 3376
rect 4557 3184 4563 3316
rect 4573 3104 4579 3336
rect 4621 3324 4627 3456
rect 4637 3344 4643 3476
rect 4685 3463 4691 3476
rect 4669 3457 4691 3463
rect 4637 3264 4643 3336
rect 4653 3184 4659 3296
rect 4669 3184 4675 3457
rect 4701 3443 4707 3596
rect 4717 3504 4723 3637
rect 4749 3604 4755 3676
rect 4685 3437 4707 3443
rect 4685 3324 4691 3437
rect 4717 3403 4723 3496
rect 4733 3484 4739 3496
rect 4749 3404 4755 3496
rect 4701 3397 4723 3403
rect 4701 3384 4707 3397
rect 4765 3383 4771 3436
rect 4717 3377 4771 3383
rect 4781 3383 4787 3596
rect 4797 3404 4803 3496
rect 4813 3484 4819 3696
rect 4845 3624 4851 3636
rect 4829 3524 4835 3596
rect 4861 3584 4867 3616
rect 4877 3544 4883 3876
rect 4909 3524 4915 3856
rect 4925 3843 4931 3896
rect 4941 3864 4947 3957
rect 4957 3884 4963 3936
rect 4989 3924 4995 4116
rect 5021 3964 5027 4076
rect 5005 3904 5011 3956
rect 5037 3944 5043 4096
rect 5053 3984 5059 4516
rect 5069 4504 5075 4536
rect 5149 4524 5155 4536
rect 5149 4504 5155 4516
rect 5165 4483 5171 4636
rect 5181 4523 5187 4696
rect 5213 4604 5219 4696
rect 5261 4677 5276 4683
rect 5197 4564 5203 4576
rect 5261 4544 5267 4677
rect 5309 4624 5315 4696
rect 5405 4684 5411 4694
rect 5373 4544 5379 4676
rect 5261 4524 5267 4536
rect 5181 4517 5203 4523
rect 5149 4477 5171 4483
rect 5149 4384 5155 4477
rect 5085 4304 5091 4316
rect 5085 4224 5091 4296
rect 5101 4244 5107 4276
rect 5117 4184 5123 4296
rect 5076 4117 5091 4123
rect 5037 3924 5043 3936
rect 4973 3884 4979 3896
rect 4925 3837 4972 3843
rect 5037 3764 5043 3856
rect 5069 3803 5075 3996
rect 5085 3944 5091 4117
rect 5101 4103 5107 4136
rect 5133 4123 5139 4356
rect 5165 4264 5171 4296
rect 5181 4184 5187 4436
rect 5197 4384 5203 4517
rect 5261 4483 5267 4516
rect 5261 4477 5283 4483
rect 5245 4384 5251 4416
rect 5261 4384 5267 4436
rect 5197 4324 5203 4376
rect 5213 4244 5219 4296
rect 5277 4264 5283 4477
rect 5357 4464 5363 4496
rect 5293 4304 5299 4396
rect 5325 4244 5331 4296
rect 5229 4157 5244 4163
rect 5229 4144 5235 4157
rect 5261 4143 5267 4236
rect 5341 4204 5347 4236
rect 5252 4137 5267 4143
rect 5181 4124 5187 4136
rect 5261 4124 5267 4137
rect 5124 4117 5139 4123
rect 5149 4104 5155 4116
rect 5101 4097 5123 4103
rect 5117 4044 5123 4097
rect 5085 3904 5091 3936
rect 5101 3844 5107 3856
rect 5069 3797 5091 3803
rect 4925 3624 4931 3716
rect 4941 3544 4947 3756
rect 5069 3724 5075 3756
rect 5085 3744 5091 3797
rect 5101 3784 5107 3796
rect 5117 3784 5123 3876
rect 5133 3724 5139 3736
rect 5165 3704 5171 3876
rect 5165 3684 5171 3696
rect 4925 3504 4931 3536
rect 4941 3504 4947 3536
rect 4861 3484 4867 3496
rect 4781 3377 4803 3383
rect 4701 3264 4707 3336
rect 4717 3284 4723 3377
rect 4733 3304 4739 3356
rect 4765 3304 4771 3316
rect 4797 3284 4803 3377
rect 4813 3364 4819 3476
rect 4877 3463 4883 3476
rect 4973 3463 4979 3676
rect 4989 3584 4995 3616
rect 5117 3504 5123 3616
rect 5005 3484 5011 3496
rect 4845 3457 4883 3463
rect 4957 3457 4979 3463
rect 4829 3344 4835 3436
rect 4813 3303 4819 3316
rect 4813 3297 4835 3303
rect 4829 3284 4835 3297
rect 4605 3104 4611 3156
rect 4637 3104 4643 3116
rect 4589 3064 4595 3096
rect 4685 3064 4691 3096
rect 4717 3064 4723 3116
rect 4749 3104 4755 3116
rect 4797 3084 4803 3096
rect 4733 2964 4739 3076
rect 4765 2984 4771 3036
rect 4621 2957 4675 2963
rect 4557 2924 4563 2936
rect 4621 2924 4627 2957
rect 4669 2944 4675 2957
rect 4701 2944 4707 2956
rect 4829 2944 4835 3036
rect 4845 2964 4851 3457
rect 4861 3184 4867 3356
rect 4877 2984 4883 3376
rect 4893 3324 4899 3436
rect 4909 3344 4915 3376
rect 4925 3344 4931 3436
rect 4941 3384 4947 3436
rect 4893 3024 4899 3276
rect 4909 3044 4915 3316
rect 4925 2963 4931 3316
rect 4941 3304 4947 3316
rect 4957 3284 4963 3457
rect 4973 3324 4979 3376
rect 4989 3224 4995 3336
rect 5005 3324 5011 3456
rect 5037 3444 5043 3456
rect 5021 3363 5027 3436
rect 5021 3357 5043 3363
rect 5037 3304 5043 3357
rect 5069 3324 5075 3436
rect 5101 3404 5107 3436
rect 5117 3384 5123 3476
rect 5085 3344 5091 3356
rect 5117 3324 5123 3336
rect 5165 3324 5171 3596
rect 5197 3403 5203 4056
rect 5213 3984 5219 4116
rect 5245 4004 5251 4116
rect 5261 3904 5267 4116
rect 5277 4084 5283 4136
rect 5357 4124 5363 4396
rect 5373 4304 5379 4476
rect 5389 4384 5395 4616
rect 5389 4304 5395 4376
rect 5373 4124 5379 4276
rect 5389 4223 5395 4296
rect 5421 4284 5427 4756
rect 5437 4304 5443 4936
rect 5469 4924 5475 4976
rect 5485 4924 5491 4996
rect 5517 4984 5523 5016
rect 5533 4984 5539 5037
rect 5501 4884 5507 4936
rect 5549 4884 5555 4916
rect 5501 4644 5507 4876
rect 5565 4844 5571 5077
rect 5581 4964 5587 5036
rect 5517 4637 5532 4643
rect 5517 4544 5523 4637
rect 5549 4643 5555 4716
rect 5581 4644 5587 4676
rect 5549 4637 5571 4643
rect 5469 4504 5475 4516
rect 5469 4444 5475 4496
rect 5485 4323 5491 4536
rect 5533 4524 5539 4536
rect 5501 4324 5507 4416
rect 5517 4364 5523 4516
rect 5549 4404 5555 4436
rect 5565 4384 5571 4637
rect 5581 4604 5587 4636
rect 5597 4584 5603 4636
rect 5613 4544 5619 4916
rect 5629 4644 5635 5317
rect 5853 5264 5859 5336
rect 5869 5204 5875 5236
rect 5757 5137 5804 5143
rect 5661 5064 5667 5096
rect 5725 5084 5731 5094
rect 5757 5084 5763 5137
rect 5853 5117 5868 5123
rect 5812 5097 5827 5103
rect 5645 4904 5651 4916
rect 5661 4704 5667 5056
rect 5677 4924 5683 4956
rect 5709 4924 5715 5016
rect 5773 4964 5779 5036
rect 5789 5004 5795 5076
rect 5725 4904 5731 4936
rect 5741 4904 5747 4916
rect 5741 4784 5747 4896
rect 5581 4537 5596 4543
rect 5581 4444 5587 4537
rect 5629 4543 5635 4636
rect 5629 4537 5651 4543
rect 5597 4444 5603 4516
rect 5476 4317 5491 4323
rect 5469 4304 5475 4316
rect 5517 4304 5523 4336
rect 5405 4264 5411 4276
rect 5389 4217 5411 4223
rect 5389 4144 5395 4196
rect 5309 4084 5315 4116
rect 5405 3944 5411 4217
rect 5421 4104 5427 4136
rect 5229 3884 5235 3894
rect 5373 3884 5379 3896
rect 5373 3864 5379 3876
rect 5213 3744 5219 3856
rect 5389 3844 5395 3896
rect 5229 3724 5235 3796
rect 5405 3784 5411 3836
rect 5309 3724 5315 3736
rect 5341 3724 5347 3776
rect 5421 3723 5427 3736
rect 5412 3717 5427 3723
rect 5213 3464 5219 3716
rect 5229 3624 5235 3716
rect 5245 3604 5251 3716
rect 5229 3584 5235 3596
rect 5229 3457 5244 3463
rect 5197 3397 5219 3403
rect 5181 3324 5187 3396
rect 5197 3344 5203 3376
rect 5213 3284 5219 3397
rect 5229 3364 5235 3457
rect 4957 3084 4963 3196
rect 5021 3124 5027 3136
rect 4909 2957 4931 2963
rect 4637 2884 4643 2936
rect 4692 2897 4716 2903
rect 4541 2704 4547 2736
rect 4557 2704 4563 2796
rect 4596 2717 4611 2723
rect 4605 2704 4611 2717
rect 4301 2664 4307 2676
rect 4349 2664 4355 2696
rect 4301 2524 4307 2536
rect 4317 2524 4323 2556
rect 4333 2504 4339 2656
rect 4365 2504 4371 2676
rect 4413 2664 4419 2696
rect 4509 2677 4524 2683
rect 4509 2584 4515 2677
rect 4589 2677 4604 2683
rect 4381 2504 4387 2516
rect 4253 2284 4259 2296
rect 4189 2084 4195 2118
rect 4045 1984 4051 2036
rect 4013 1904 4019 1916
rect 4029 1904 4035 1976
rect 4013 1784 4019 1816
rect 4029 1744 4035 1876
rect 4061 1864 4067 1936
rect 4141 1904 4147 1936
rect 4221 1904 4227 2276
rect 4269 2164 4275 2236
rect 4269 1984 4275 2136
rect 4301 2126 4307 2156
rect 4317 1964 4323 2356
rect 4093 1864 4099 1876
rect 4029 1724 4035 1736
rect 4061 1724 4067 1856
rect 4093 1764 4099 1836
rect 4109 1704 4115 1736
rect 4125 1724 4131 1876
rect 4157 1864 4163 1876
rect 4237 1864 4243 1936
rect 3885 1303 3891 1376
rect 3965 1344 3971 1476
rect 3981 1444 3987 1456
rect 3876 1297 3891 1303
rect 3901 1163 3907 1316
rect 3933 1264 3939 1336
rect 3885 1157 3907 1163
rect 3661 1084 3667 1136
rect 3709 1104 3715 1116
rect 3885 1104 3891 1157
rect 3764 1077 3779 1083
rect 3725 1064 3731 1076
rect 3645 1044 3651 1056
rect 3661 984 3667 996
rect 3517 704 3523 856
rect 3549 784 3555 836
rect 3565 664 3571 716
rect 3629 664 3635 956
rect 3645 804 3651 956
rect 3645 704 3651 736
rect 3677 664 3683 836
rect 3693 784 3699 1036
rect 3741 944 3747 1036
rect 3773 944 3779 1077
rect 3709 924 3715 936
rect 3773 897 3788 903
rect 3725 844 3731 896
rect 3693 764 3699 776
rect 3693 724 3699 756
rect 3533 624 3539 656
rect 3565 644 3571 656
rect 3549 524 3555 536
rect 3517 504 3523 516
rect 3517 384 3523 496
rect 3533 484 3539 516
rect 3517 324 3523 376
rect 3421 277 3436 283
rect 3380 257 3395 263
rect 3357 164 3363 176
rect 3341 144 3347 156
rect 3117 123 3123 136
rect 3389 124 3395 257
rect 3453 224 3459 296
rect 3533 264 3539 436
rect 3565 283 3571 636
rect 3597 524 3603 656
rect 3629 524 3635 656
rect 3757 564 3763 676
rect 3773 584 3779 897
rect 3613 504 3619 516
rect 3677 484 3683 556
rect 3805 544 3811 976
rect 3837 964 3843 1056
rect 3885 924 3891 1096
rect 3901 1024 3907 1056
rect 3933 984 3939 1236
rect 3965 1084 3971 1336
rect 3981 1124 3987 1436
rect 4013 1284 4019 1296
rect 4013 1184 4019 1196
rect 4045 1123 4051 1676
rect 4157 1604 4163 1696
rect 4077 1264 4083 1356
rect 4093 1324 4099 1556
rect 4173 1524 4179 1636
rect 4109 1502 4115 1516
rect 4141 1364 4147 1476
rect 4189 1423 4195 1836
rect 4205 1784 4211 1856
rect 4221 1844 4227 1856
rect 4253 1844 4259 1936
rect 4269 1884 4275 1896
rect 4205 1724 4211 1736
rect 4221 1724 4227 1756
rect 4237 1624 4243 1756
rect 4253 1584 4259 1636
rect 4237 1484 4243 1496
rect 4237 1423 4243 1436
rect 4173 1417 4195 1423
rect 4221 1417 4243 1423
rect 4045 1117 4067 1123
rect 3965 984 3971 1056
rect 3981 923 3987 936
rect 3940 917 3987 923
rect 3901 877 3916 883
rect 3885 824 3891 836
rect 3885 684 3891 796
rect 3853 664 3859 676
rect 3821 503 3827 636
rect 3853 544 3859 576
rect 3869 564 3875 576
rect 3805 497 3827 503
rect 3581 364 3587 436
rect 3661 384 3667 436
rect 3693 404 3699 436
rect 3588 317 3603 323
rect 3556 277 3571 283
rect 3597 264 3603 317
rect 3645 304 3651 356
rect 3629 284 3635 296
rect 3725 284 3731 436
rect 3725 264 3731 276
rect 3533 184 3539 256
rect 3437 124 3443 136
rect 3485 124 3491 156
rect 3693 144 3699 156
rect 3757 124 3763 436
rect 3805 384 3811 497
rect 3821 343 3827 476
rect 3853 404 3859 536
rect 3885 444 3891 676
rect 3805 337 3827 343
rect 3789 164 3795 236
rect 3117 117 3164 123
rect 3069 104 3075 116
rect 3213 104 3219 116
rect 2557 84 2563 96
rect 2541 64 2547 76
rect 3805 64 3811 337
rect 3821 284 3827 316
rect 3837 304 3843 396
rect 3901 364 3907 877
rect 3933 664 3939 676
rect 3933 644 3939 656
rect 3917 604 3923 636
rect 3949 583 3955 896
rect 3933 577 3955 583
rect 3837 124 3843 296
rect 3901 284 3907 316
rect 3853 264 3859 276
rect 3869 184 3875 236
rect 3885 144 3891 256
rect 3917 164 3923 396
rect 3933 384 3939 577
rect 3965 544 3971 656
rect 3949 337 3964 343
rect 3949 324 3955 337
rect 3949 304 3955 316
rect 3981 284 3987 896
rect 3997 884 4003 1056
rect 4029 944 4035 956
rect 3997 724 4003 836
rect 4045 763 4051 896
rect 4061 764 4067 1117
rect 4077 944 4083 1256
rect 4093 1144 4099 1256
rect 4141 1184 4147 1296
rect 4173 1204 4179 1417
rect 4205 1184 4211 1236
rect 4221 1184 4227 1417
rect 4253 1403 4259 1576
rect 4237 1397 4259 1403
rect 4237 1144 4243 1397
rect 4269 1244 4275 1876
rect 4285 1504 4291 1836
rect 4301 1824 4307 1876
rect 4317 1824 4323 1896
rect 4333 1804 4339 2416
rect 4349 1964 4355 2376
rect 4365 2104 4371 2316
rect 4381 2264 4387 2316
rect 4397 2264 4403 2536
rect 4413 2524 4419 2556
rect 4557 2524 4563 2556
rect 4589 2544 4595 2677
rect 4621 2664 4627 2836
rect 4653 2744 4659 2796
rect 4653 2704 4659 2736
rect 4749 2723 4755 2876
rect 4909 2804 4915 2957
rect 4909 2743 4915 2796
rect 4893 2737 4915 2743
rect 4749 2717 4771 2723
rect 4637 2683 4643 2696
rect 4637 2677 4652 2683
rect 4525 2464 4531 2496
rect 4442 2414 4454 2416
rect 4427 2406 4429 2414
rect 4437 2406 4439 2414
rect 4447 2406 4449 2414
rect 4457 2406 4459 2414
rect 4467 2406 4469 2414
rect 4442 2404 4454 2406
rect 4397 2184 4403 2256
rect 4461 2104 4467 2376
rect 4493 2364 4499 2456
rect 4573 2443 4579 2536
rect 4589 2464 4595 2536
rect 4637 2524 4643 2636
rect 4653 2544 4659 2576
rect 4669 2524 4675 2696
rect 4701 2624 4707 2636
rect 4733 2624 4739 2696
rect 4765 2664 4771 2717
rect 4733 2524 4739 2596
rect 4685 2503 4691 2516
rect 4781 2504 4787 2516
rect 4644 2497 4691 2503
rect 4573 2437 4595 2443
rect 4589 2384 4595 2437
rect 4701 2384 4707 2436
rect 4477 2284 4483 2296
rect 4493 2264 4499 2296
rect 4365 1984 4371 2076
rect 4397 2024 4403 2076
rect 4442 2014 4454 2016
rect 4427 2006 4429 2014
rect 4437 2006 4439 2014
rect 4447 2006 4449 2014
rect 4457 2006 4459 2014
rect 4467 2006 4469 2014
rect 4442 2004 4454 2006
rect 4493 1983 4499 2176
rect 4525 2164 4531 2276
rect 4573 2164 4579 2336
rect 4605 2284 4611 2336
rect 4477 1977 4499 1983
rect 4349 1883 4355 1916
rect 4477 1904 4483 1977
rect 4493 1924 4499 1956
rect 4509 1904 4515 1956
rect 4525 1904 4531 2116
rect 4557 1924 4563 1936
rect 4349 1877 4371 1883
rect 4349 1784 4355 1816
rect 4365 1784 4371 1877
rect 4397 1824 4403 1876
rect 4573 1864 4579 1996
rect 4589 1924 4595 2036
rect 4605 2024 4611 2096
rect 4621 1984 4627 2336
rect 4637 2304 4643 2316
rect 4733 2184 4739 2456
rect 4637 1924 4643 2036
rect 4285 1324 4291 1456
rect 4301 1364 4307 1756
rect 4317 1724 4323 1776
rect 4333 1504 4339 1776
rect 4397 1724 4403 1736
rect 4493 1724 4499 1836
rect 4557 1764 4563 1836
rect 4589 1784 4595 1796
rect 4621 1744 4627 1816
rect 4637 1723 4643 1776
rect 4653 1763 4659 1896
rect 4669 1884 4675 2136
rect 4733 2083 4739 2096
rect 4717 2077 4739 2083
rect 4717 1984 4723 2077
rect 4749 1984 4755 2436
rect 4781 2404 4787 2496
rect 4797 2464 4803 2676
rect 4829 2664 4835 2696
rect 4829 2604 4835 2636
rect 4845 2604 4851 2716
rect 4861 2683 4867 2736
rect 4877 2704 4883 2716
rect 4893 2704 4899 2737
rect 4861 2677 4876 2683
rect 4925 2664 4931 2936
rect 4941 2704 4947 3036
rect 4957 3004 4963 3076
rect 4957 2884 4963 2936
rect 4973 2903 4979 3096
rect 5005 3004 5011 3036
rect 4989 2924 4995 2936
rect 4973 2897 4988 2903
rect 4973 2784 4979 2897
rect 4957 2677 4972 2683
rect 4868 2657 4915 2663
rect 4909 2643 4915 2657
rect 4957 2643 4963 2677
rect 4909 2637 4963 2643
rect 4813 2503 4819 2536
rect 4845 2524 4851 2576
rect 4861 2503 4867 2536
rect 4877 2524 4883 2596
rect 4909 2584 4915 2596
rect 4989 2584 4995 2696
rect 4941 2524 4947 2556
rect 4813 2497 4867 2503
rect 4893 2503 4899 2516
rect 4884 2497 4899 2503
rect 4957 2503 4963 2536
rect 4989 2524 4995 2536
rect 5005 2503 5011 2956
rect 5037 2924 5043 3136
rect 5069 3123 5075 3176
rect 5053 3117 5075 3123
rect 5053 3084 5059 3117
rect 5037 2904 5043 2916
rect 5021 2684 5027 2736
rect 5037 2724 5043 2796
rect 5053 2704 5059 2816
rect 5069 2744 5075 2836
rect 5085 2744 5091 3276
rect 5149 3104 5155 3136
rect 5101 3024 5107 3096
rect 5229 3064 5235 3216
rect 5261 3144 5267 3516
rect 5277 3504 5283 3556
rect 5117 2924 5123 3036
rect 5133 2824 5139 3036
rect 5149 2804 5155 2956
rect 5229 2944 5235 3056
rect 5245 2984 5251 3036
rect 5261 3004 5267 3096
rect 5165 2924 5171 2936
rect 5213 2884 5219 2916
rect 5085 2704 5091 2716
rect 4957 2497 4979 2503
rect 4909 2464 4915 2496
rect 4797 2184 4803 2356
rect 4845 2184 4851 2236
rect 4877 2184 4883 2436
rect 4909 2304 4915 2396
rect 4973 2384 4979 2497
rect 4989 2497 5011 2503
rect 4941 2303 4947 2316
rect 4941 2297 4963 2303
rect 4868 2137 4883 2143
rect 4813 2024 4819 2136
rect 4676 1877 4691 1883
rect 4653 1757 4675 1763
rect 4669 1724 4675 1757
rect 4685 1744 4691 1877
rect 4701 1784 4707 1936
rect 4717 1904 4723 1916
rect 4733 1904 4739 1916
rect 4733 1877 4748 1883
rect 4637 1717 4659 1723
rect 4541 1684 4547 1696
rect 4589 1664 4595 1696
rect 4637 1684 4643 1696
rect 4653 1663 4659 1717
rect 4637 1657 4659 1663
rect 4349 1543 4355 1636
rect 4365 1604 4371 1636
rect 4442 1614 4454 1616
rect 4427 1606 4429 1614
rect 4437 1606 4439 1614
rect 4447 1606 4449 1614
rect 4457 1606 4459 1614
rect 4467 1606 4469 1614
rect 4442 1604 4454 1606
rect 4365 1563 4371 1596
rect 4365 1557 4387 1563
rect 4349 1537 4371 1543
rect 4365 1504 4371 1537
rect 4381 1524 4387 1557
rect 4093 984 4099 1056
rect 4109 984 4115 996
rect 4157 984 4163 1076
rect 4173 1004 4179 1116
rect 4317 1104 4323 1396
rect 4333 1364 4339 1476
rect 4349 1144 4355 1236
rect 4365 1184 4371 1476
rect 4397 1184 4403 1356
rect 4429 1324 4435 1416
rect 4461 1384 4467 1536
rect 4493 1444 4499 1616
rect 4509 1484 4515 1636
rect 4637 1584 4643 1657
rect 4669 1584 4675 1676
rect 4685 1584 4691 1736
rect 4717 1724 4723 1836
rect 4717 1624 4723 1676
rect 4605 1544 4611 1576
rect 4525 1484 4531 1496
rect 4557 1424 4563 1456
rect 4653 1444 4659 1576
rect 4717 1484 4723 1496
rect 4685 1443 4691 1476
rect 4701 1464 4707 1476
rect 4733 1463 4739 1877
rect 4781 1784 4787 1956
rect 4804 1917 4819 1923
rect 4797 1744 4803 1836
rect 4813 1744 4819 1917
rect 4829 1804 4835 1916
rect 4861 1904 4867 1976
rect 4877 1944 4883 2137
rect 4893 1984 4899 2116
rect 4909 1964 4915 2176
rect 4941 2124 4947 2156
rect 4957 2144 4963 2297
rect 4973 2284 4979 2376
rect 4973 2264 4979 2276
rect 4941 1904 4947 2116
rect 4973 2104 4979 2236
rect 4989 2083 4995 2497
rect 5005 2424 5011 2436
rect 5021 2323 5027 2676
rect 5037 2563 5043 2696
rect 5053 2664 5059 2696
rect 5069 2564 5075 2696
rect 5085 2624 5091 2676
rect 5117 2664 5123 2796
rect 5229 2723 5235 2936
rect 5245 2784 5251 2916
rect 5277 2824 5283 3396
rect 5293 3124 5299 3696
rect 5325 3484 5331 3696
rect 5357 3544 5363 3596
rect 5341 3504 5347 3536
rect 5341 3444 5347 3496
rect 5357 3464 5363 3536
rect 5309 3324 5315 3436
rect 5373 3403 5379 3676
rect 5389 3544 5395 3716
rect 5389 3484 5395 3496
rect 5405 3444 5411 3476
rect 5421 3464 5427 3717
rect 5437 3584 5443 4256
rect 5453 4204 5459 4276
rect 5517 4184 5523 4296
rect 5533 4244 5539 4316
rect 5565 4284 5571 4296
rect 5581 4284 5587 4416
rect 5597 4384 5603 4396
rect 5613 4364 5619 4516
rect 5629 4464 5635 4516
rect 5629 4364 5635 4436
rect 5613 4284 5619 4296
rect 5469 4124 5475 4136
rect 5485 4084 5491 4136
rect 5517 3904 5523 4136
rect 5549 4104 5555 4118
rect 5453 3724 5459 3736
rect 5469 3724 5475 3836
rect 5501 3784 5507 3896
rect 5517 3884 5523 3896
rect 5533 3824 5539 3936
rect 5533 3764 5539 3776
rect 5565 3743 5571 4276
rect 5645 4144 5651 4537
rect 5677 4524 5683 4576
rect 5661 4304 5667 4436
rect 5693 4344 5699 4776
rect 5725 4684 5731 4694
rect 5757 4624 5763 4916
rect 5821 4904 5827 5097
rect 5837 4944 5843 5116
rect 5853 5104 5859 5117
rect 5853 4984 5859 5076
rect 5853 4944 5859 4976
rect 5821 4784 5827 4896
rect 5853 4884 5859 4916
rect 5709 4524 5715 4536
rect 5725 4464 5731 4516
rect 5773 4404 5779 4616
rect 5789 4524 5795 4676
rect 5837 4604 5843 4876
rect 5869 4863 5875 5096
rect 5853 4857 5875 4863
rect 5853 4744 5859 4857
rect 5869 4824 5875 4836
rect 5805 4544 5811 4596
rect 5828 4537 5843 4543
rect 5821 4524 5827 4536
rect 5757 4344 5763 4396
rect 5773 4384 5779 4396
rect 5693 4304 5699 4336
rect 5789 4324 5795 4336
rect 5789 4304 5795 4316
rect 5741 4264 5747 4296
rect 5821 4263 5827 4316
rect 5837 4304 5843 4537
rect 5853 4524 5859 4736
rect 5885 4724 5891 5357
rect 5901 5344 5907 5356
rect 6141 5264 6147 5316
rect 6045 5204 6051 5236
rect 6029 5124 6035 5156
rect 5901 5104 5907 5116
rect 5946 5014 5958 5016
rect 5931 5006 5933 5014
rect 5941 5006 5943 5014
rect 5951 5006 5953 5014
rect 5961 5006 5963 5014
rect 5971 5006 5973 5014
rect 5946 5004 5958 5006
rect 5997 4943 6003 5096
rect 6029 5063 6035 5116
rect 6029 5057 6044 5063
rect 6013 4964 6019 4996
rect 6029 4964 6035 5057
rect 6061 5004 6067 5156
rect 6077 5123 6083 5136
rect 6077 5117 6099 5123
rect 6093 5104 6099 5117
rect 6141 5104 6147 5116
rect 6173 5104 6179 5376
rect 6077 5004 6083 5076
rect 6045 4944 6051 4956
rect 5997 4937 6019 4943
rect 5901 4924 5907 4936
rect 5933 4904 5939 4916
rect 5981 4784 5987 4856
rect 5997 4824 6003 4916
rect 5869 4704 5875 4716
rect 5869 4624 5875 4696
rect 5885 4664 5891 4676
rect 5869 4544 5875 4596
rect 5885 4564 5891 4656
rect 5946 4614 5958 4616
rect 5931 4606 5933 4614
rect 5941 4606 5943 4614
rect 5951 4606 5953 4614
rect 5961 4606 5963 4614
rect 5971 4606 5973 4614
rect 5946 4604 5958 4606
rect 5901 4523 5907 4576
rect 5892 4517 5907 4523
rect 5917 4344 5923 4576
rect 5933 4464 5939 4536
rect 5997 4524 6003 4816
rect 6013 4684 6019 4937
rect 6093 4924 6099 5036
rect 6109 4904 6115 4936
rect 6141 4924 6147 5036
rect 6013 4624 6019 4636
rect 5997 4464 6003 4516
rect 6013 4344 6019 4616
rect 6045 4564 6051 4776
rect 6109 4604 6115 4896
rect 6125 4764 6131 4916
rect 6157 4903 6163 5076
rect 6141 4897 6163 4903
rect 6141 4844 6147 4897
rect 6157 4804 6163 4836
rect 6173 4744 6179 5056
rect 6189 4804 6195 5316
rect 6237 5104 6243 5116
rect 6253 5064 6259 5096
rect 6221 4984 6227 4996
rect 6237 4923 6243 4996
rect 6253 4924 6259 5056
rect 6269 5023 6275 5236
rect 6349 5044 6355 5096
rect 6269 5017 6291 5023
rect 6269 4944 6275 4956
rect 6285 4924 6291 5017
rect 6317 4924 6323 5036
rect 6333 4944 6339 4956
rect 6228 4917 6243 4923
rect 6228 4897 6243 4903
rect 6237 4844 6243 4897
rect 6253 4864 6259 4916
rect 6237 4784 6243 4836
rect 6301 4744 6307 4776
rect 6141 4623 6147 4694
rect 6173 4684 6179 4736
rect 6205 4643 6211 4696
rect 6253 4684 6259 4716
rect 6269 4684 6275 4696
rect 6253 4663 6259 4676
rect 6253 4657 6275 4663
rect 6189 4637 6211 4643
rect 6141 4617 6163 4623
rect 6109 4544 6115 4556
rect 5876 4297 5891 4303
rect 5853 4263 5859 4276
rect 5821 4257 5859 4263
rect 5725 4244 5731 4256
rect 5789 4244 5795 4256
rect 5613 4124 5619 4136
rect 5597 4004 5603 4036
rect 5597 3864 5603 3996
rect 5629 3864 5635 3896
rect 5629 3784 5635 3796
rect 5661 3743 5667 4236
rect 5677 4184 5683 4196
rect 5741 4184 5747 4196
rect 5789 4164 5795 4236
rect 5716 4117 5731 4123
rect 5725 4044 5731 4117
rect 5741 4104 5747 4136
rect 5757 4083 5763 4116
rect 5741 4077 5763 4083
rect 5709 3984 5715 3996
rect 5693 3904 5699 3956
rect 5725 3903 5731 4036
rect 5709 3897 5731 3903
rect 5693 3864 5699 3876
rect 5565 3737 5587 3743
rect 5469 3603 5475 3716
rect 5485 3704 5491 3736
rect 5581 3724 5587 3737
rect 5645 3737 5667 3743
rect 5485 3684 5491 3696
rect 5453 3597 5475 3603
rect 5453 3504 5459 3597
rect 5373 3397 5395 3403
rect 5325 3344 5331 3376
rect 5325 3084 5331 3336
rect 5357 3264 5363 3376
rect 5389 3324 5395 3397
rect 5421 3344 5427 3456
rect 5421 3324 5427 3336
rect 5389 3304 5395 3316
rect 5405 3304 5411 3316
rect 5437 3284 5443 3336
rect 5453 3104 5459 3476
rect 5469 3264 5475 3436
rect 5469 3104 5475 3196
rect 5485 3184 5491 3576
rect 5501 3304 5507 3576
rect 5533 3324 5539 3716
rect 5565 3684 5571 3716
rect 5501 3144 5507 3256
rect 5325 3064 5331 3076
rect 5357 3063 5363 3096
rect 5357 3057 5379 3063
rect 5325 2924 5331 3056
rect 5373 2944 5379 3057
rect 5220 2717 5235 2723
rect 5133 2624 5139 2676
rect 5149 2603 5155 2716
rect 5277 2704 5283 2736
rect 5229 2697 5244 2703
rect 5181 2624 5187 2696
rect 5133 2597 5155 2603
rect 5037 2557 5059 2563
rect 5037 2524 5043 2536
rect 5053 2524 5059 2557
rect 5133 2544 5139 2597
rect 5069 2503 5075 2536
rect 5117 2504 5123 2516
rect 5053 2497 5075 2503
rect 5037 2444 5043 2496
rect 5005 2317 5027 2323
rect 5005 2304 5011 2317
rect 5005 2284 5011 2296
rect 4973 2077 4995 2083
rect 4973 1984 4979 2077
rect 4845 1884 4851 1896
rect 4765 1684 4771 1696
rect 4749 1524 4755 1616
rect 4717 1457 4739 1463
rect 4781 1463 4787 1696
rect 4797 1484 4803 1676
rect 4813 1624 4819 1736
rect 4845 1684 4851 1876
rect 4877 1864 4883 1876
rect 4957 1784 4963 1876
rect 5005 1804 5011 2118
rect 4909 1724 4915 1756
rect 4989 1724 4995 1736
rect 4845 1637 4860 1643
rect 4813 1504 4819 1536
rect 4781 1457 4803 1463
rect 4685 1437 4707 1443
rect 4413 1264 4419 1276
rect 4442 1214 4454 1216
rect 4427 1206 4429 1214
rect 4437 1206 4439 1214
rect 4447 1206 4449 1214
rect 4457 1206 4459 1214
rect 4467 1206 4469 1214
rect 4442 1204 4454 1206
rect 4365 1164 4371 1176
rect 4381 1124 4387 1136
rect 4413 1104 4419 1136
rect 4493 1124 4499 1296
rect 4365 1084 4371 1096
rect 4077 804 4083 936
rect 4093 924 4099 956
rect 4125 943 4131 976
rect 4141 964 4147 976
rect 4109 937 4131 943
rect 4036 757 4051 763
rect 4029 684 4035 756
rect 4109 723 4115 937
rect 4125 904 4131 916
rect 4173 904 4179 936
rect 4141 744 4147 896
rect 4173 724 4179 836
rect 4100 717 4115 723
rect 4077 584 4083 676
rect 3949 184 3955 276
rect 3853 104 3859 116
rect 3885 104 3891 116
rect 477 -17 483 36
rect 1434 14 1446 16
rect 1419 6 1421 14
rect 1429 6 1431 14
rect 1439 6 1441 14
rect 1449 6 1451 14
rect 1459 6 1461 14
rect 1434 4 1446 6
rect 461 -23 483 -17
rect 2845 -17 2851 36
rect 3421 -17 3427 36
rect 3469 -17 3475 36
rect 3517 -17 3523 36
rect 2845 -23 2867 -17
rect 3405 -23 3427 -17
rect 3453 -23 3475 -17
rect 3501 -23 3523 -17
rect 3725 -17 3731 36
rect 3725 -23 3747 -17
rect 3805 -23 3811 36
rect 3837 -23 3843 56
rect 4061 44 4067 396
rect 4077 284 4083 536
rect 4109 404 4115 717
rect 4141 564 4147 676
rect 4189 664 4195 976
rect 4205 944 4211 956
rect 4253 904 4259 1016
rect 4237 844 4243 896
rect 4269 723 4275 1056
rect 4285 984 4291 1036
rect 4429 1024 4435 1096
rect 4365 824 4371 1016
rect 4260 717 4275 723
rect 4189 644 4195 656
rect 4205 524 4211 636
rect 4253 584 4259 676
rect 4125 444 4131 516
rect 4237 444 4243 536
rect 4157 304 4163 376
rect 4077 164 4083 276
rect 4093 244 4099 294
rect 4237 264 4243 436
rect 4253 384 4259 476
rect 4269 364 4275 717
rect 4349 584 4355 694
rect 4381 684 4387 936
rect 4442 814 4454 816
rect 4427 806 4429 814
rect 4437 806 4439 814
rect 4447 806 4449 814
rect 4457 806 4459 814
rect 4467 806 4469 814
rect 4442 804 4454 806
rect 4493 784 4499 816
rect 4509 724 4515 1416
rect 4573 1363 4579 1416
rect 4557 1357 4579 1363
rect 4557 1344 4563 1357
rect 4621 1344 4627 1436
rect 4573 1304 4579 1336
rect 4653 1324 4659 1376
rect 4557 1184 4563 1216
rect 4573 1144 4579 1236
rect 4589 1104 4595 1236
rect 4637 1204 4643 1296
rect 4669 1284 4675 1436
rect 4701 1384 4707 1437
rect 4717 1284 4723 1457
rect 4733 1344 4739 1376
rect 4589 1084 4595 1096
rect 4637 1064 4643 1156
rect 4669 1144 4675 1256
rect 4733 1164 4739 1316
rect 4765 1303 4771 1376
rect 4781 1324 4787 1336
rect 4797 1304 4803 1457
rect 4765 1297 4787 1303
rect 4765 1224 4771 1276
rect 4781 1224 4787 1297
rect 4813 1283 4819 1476
rect 4829 1384 4835 1436
rect 4845 1404 4851 1637
rect 4877 1423 4883 1556
rect 4941 1504 4947 1516
rect 4861 1417 4883 1423
rect 4797 1277 4819 1283
rect 4413 544 4419 696
rect 4317 524 4323 536
rect 4493 524 4499 536
rect 4509 524 4515 636
rect 4541 524 4547 676
rect 4557 664 4563 956
rect 4605 843 4611 936
rect 4589 837 4611 843
rect 4589 684 4595 837
rect 4605 704 4611 716
rect 4621 683 4627 1056
rect 4637 864 4643 896
rect 4653 823 4659 1116
rect 4669 944 4675 976
rect 4637 817 4659 823
rect 4637 784 4643 817
rect 4596 677 4611 683
rect 4621 677 4643 683
rect 4573 544 4579 636
rect 4301 384 4307 456
rect 4349 384 4355 436
rect 4442 414 4454 416
rect 4427 406 4429 414
rect 4437 406 4439 414
rect 4447 406 4449 414
rect 4457 406 4459 414
rect 4467 406 4469 414
rect 4442 404 4454 406
rect 4356 317 4371 323
rect 4301 284 4307 296
rect 4205 184 4211 236
rect 4237 184 4243 236
rect 4253 164 4259 276
rect 4285 264 4291 276
rect 4333 244 4339 316
rect 4365 284 4371 317
rect 4509 304 4515 516
rect 4397 284 4403 296
rect 4413 264 4419 276
rect 4285 164 4291 196
rect 4477 184 4483 276
rect 4141 124 4147 156
rect 4077 104 4083 118
rect 4061 -23 4067 16
rect 4093 -23 4099 36
rect 4253 -23 4259 16
rect 4442 14 4454 16
rect 4427 6 4429 14
rect 4437 6 4439 14
rect 4447 6 4449 14
rect 4457 6 4459 14
rect 4467 6 4469 14
rect 4442 4 4454 6
rect 4541 -23 4547 256
rect 4573 144 4579 476
rect 4589 324 4595 616
rect 4605 603 4611 677
rect 4621 624 4627 656
rect 4605 597 4627 603
rect 4621 584 4627 597
rect 4589 203 4595 316
rect 4605 244 4611 296
rect 4589 197 4611 203
rect 4605 -17 4611 197
rect 4589 -23 4611 -17
rect 4621 -17 4627 496
rect 4637 264 4643 677
rect 4653 504 4659 656
rect 4637 124 4643 236
rect 4685 203 4691 1156
rect 4733 1104 4739 1136
rect 4765 1124 4771 1196
rect 4717 884 4723 916
rect 4733 904 4739 1076
rect 4749 1024 4755 1096
rect 4765 1084 4771 1116
rect 4797 983 4803 1277
rect 4829 1264 4835 1276
rect 4845 1244 4851 1316
rect 4861 1223 4867 1417
rect 4900 1417 4963 1423
rect 4957 1363 4963 1417
rect 4973 1384 4979 1616
rect 5021 1524 5027 1636
rect 5037 1544 5043 2376
rect 5053 2364 5059 2497
rect 5069 2304 5075 2476
rect 5085 2384 5091 2396
rect 5085 2124 5091 2196
rect 5101 2144 5107 2396
rect 5133 2324 5139 2536
rect 5149 2524 5155 2576
rect 5165 2544 5171 2616
rect 5197 2384 5203 2596
rect 5213 2524 5219 2656
rect 5229 2524 5235 2697
rect 5309 2684 5315 2696
rect 5261 2604 5267 2676
rect 5236 2517 5251 2523
rect 5165 2324 5171 2336
rect 5133 2284 5139 2296
rect 5117 2184 5123 2196
rect 5213 2184 5219 2276
rect 5245 2244 5251 2517
rect 5261 2384 5267 2576
rect 5277 2564 5283 2656
rect 5261 2244 5267 2296
rect 5133 2104 5139 2116
rect 5053 1984 5059 2076
rect 5069 1704 5075 2096
rect 5149 2064 5155 2076
rect 5165 2024 5171 2076
rect 5181 1984 5187 2136
rect 5229 2084 5235 2116
rect 5261 2083 5267 2096
rect 5252 2077 5267 2083
rect 5213 1984 5219 2076
rect 5085 1764 5091 1836
rect 5213 1823 5219 1894
rect 5277 1884 5283 2456
rect 5293 2284 5299 2376
rect 5309 2364 5315 2636
rect 5325 2524 5331 2916
rect 5373 2704 5379 2936
rect 5405 2924 5411 3096
rect 5453 3084 5459 3096
rect 5421 3044 5427 3056
rect 5453 3044 5459 3076
rect 5437 2964 5443 2976
rect 5421 2784 5427 2876
rect 5389 2704 5395 2736
rect 5453 2704 5459 2936
rect 5469 2724 5475 3076
rect 5501 2924 5507 3116
rect 5517 3064 5523 3076
rect 5533 2884 5539 3296
rect 5549 3184 5555 3616
rect 5581 3584 5587 3716
rect 5645 3664 5651 3737
rect 5677 3724 5683 3736
rect 5613 3584 5619 3636
rect 5565 3463 5571 3496
rect 5581 3484 5587 3496
rect 5565 3457 5587 3463
rect 5581 3384 5587 3457
rect 5597 3444 5603 3536
rect 5629 3504 5635 3636
rect 5661 3584 5667 3716
rect 5693 3624 5699 3856
rect 5709 3784 5715 3897
rect 5741 3823 5747 4077
rect 5773 3923 5779 4156
rect 5805 4144 5811 4196
rect 5885 4164 5891 4297
rect 5901 4263 5907 4296
rect 5917 4284 5923 4296
rect 5933 4264 5939 4336
rect 5949 4264 5955 4316
rect 5901 4257 5923 4263
rect 5917 4243 5923 4257
rect 5917 4237 5932 4243
rect 5988 4237 6003 4243
rect 5853 4124 5859 4156
rect 5869 4117 5884 4123
rect 5821 3963 5827 4036
rect 5805 3957 5827 3963
rect 5773 3917 5795 3923
rect 5741 3817 5763 3823
rect 5757 3784 5763 3817
rect 5757 3764 5763 3776
rect 5725 3704 5731 3716
rect 5661 3443 5667 3516
rect 5725 3504 5731 3616
rect 5757 3524 5763 3576
rect 5773 3564 5779 3636
rect 5789 3524 5795 3917
rect 5805 3784 5811 3957
rect 5821 3904 5827 3936
rect 5805 3724 5811 3736
rect 5821 3724 5827 3816
rect 5837 3724 5843 3936
rect 5869 3924 5875 4117
rect 5901 3944 5907 4236
rect 5946 4214 5958 4216
rect 5931 4206 5933 4214
rect 5941 4206 5943 4214
rect 5951 4206 5953 4214
rect 5961 4206 5963 4214
rect 5971 4206 5973 4214
rect 5946 4204 5958 4206
rect 5997 4204 6003 4237
rect 6013 4224 6019 4276
rect 6029 4164 6035 4336
rect 6045 4304 6051 4536
rect 6093 4504 6099 4516
rect 6141 4503 6147 4596
rect 6157 4584 6163 4617
rect 6173 4504 6179 4616
rect 6125 4497 6147 4503
rect 6077 4364 6083 4436
rect 6125 4304 6131 4497
rect 6141 4304 6147 4456
rect 6189 4304 6195 4637
rect 6269 4584 6275 4657
rect 6205 4464 6211 4576
rect 6269 4544 6275 4576
rect 6301 4524 6307 4676
rect 6221 4504 6227 4516
rect 6084 4297 6099 4303
rect 6045 4244 6051 4276
rect 6061 4224 6067 4276
rect 6093 4244 6099 4297
rect 6109 4264 6115 4296
rect 6125 4284 6131 4296
rect 6157 4277 6172 4283
rect 6157 4264 6163 4277
rect 6173 4244 6179 4256
rect 5997 3984 6003 4116
rect 6013 4004 6019 4136
rect 6093 4124 6099 4176
rect 6189 4144 6195 4256
rect 6109 4103 6115 4136
rect 6205 4124 6211 4296
rect 6109 4097 6124 4103
rect 6157 4044 6163 4116
rect 6013 3984 6019 3996
rect 5869 3864 5875 3916
rect 5885 3724 5891 3776
rect 5821 3624 5827 3716
rect 5901 3704 5907 3896
rect 5946 3814 5958 3816
rect 5931 3806 5933 3814
rect 5941 3806 5943 3814
rect 5951 3806 5953 3814
rect 5961 3806 5963 3814
rect 5971 3806 5973 3814
rect 5946 3804 5958 3806
rect 5853 3584 5859 3636
rect 5821 3504 5827 3536
rect 5732 3497 5747 3503
rect 5645 3437 5667 3443
rect 5645 3344 5651 3437
rect 5661 3384 5667 3416
rect 5677 3344 5683 3476
rect 5693 3464 5699 3496
rect 5709 3444 5715 3476
rect 5741 3464 5747 3497
rect 5757 3464 5763 3496
rect 5805 3464 5811 3476
rect 5613 3284 5619 3316
rect 5565 3124 5571 3236
rect 5581 3204 5587 3276
rect 5629 3204 5635 3336
rect 5645 3324 5651 3336
rect 5725 3324 5731 3456
rect 5757 3444 5763 3456
rect 5741 3324 5747 3416
rect 5773 3404 5779 3436
rect 5789 3404 5795 3436
rect 5789 3324 5795 3336
rect 5549 3077 5564 3083
rect 5549 2903 5555 3077
rect 5581 3064 5587 3196
rect 5629 3184 5635 3196
rect 5613 3104 5619 3176
rect 5597 2944 5603 3056
rect 5629 2944 5635 2956
rect 5565 2926 5571 2936
rect 5549 2897 5571 2903
rect 5508 2697 5523 2703
rect 5341 2524 5347 2636
rect 5357 2584 5363 2676
rect 5325 2444 5331 2516
rect 5325 2244 5331 2276
rect 5341 2264 5347 2456
rect 5357 2404 5363 2516
rect 5373 2484 5379 2696
rect 5405 2684 5411 2696
rect 5485 2683 5491 2696
rect 5517 2684 5523 2697
rect 5485 2677 5507 2683
rect 5405 2464 5411 2676
rect 5437 2544 5443 2596
rect 5501 2584 5507 2677
rect 5517 2624 5523 2636
rect 5533 2604 5539 2736
rect 5453 2524 5459 2556
rect 5501 2524 5507 2576
rect 5549 2564 5555 2576
rect 5389 2364 5395 2436
rect 5389 2304 5395 2356
rect 5453 2304 5459 2356
rect 5373 2184 5379 2236
rect 5213 1817 5235 1823
rect 5229 1784 5235 1817
rect 5293 1804 5299 2136
rect 5325 2124 5331 2156
rect 5389 2104 5395 2276
rect 5437 2264 5443 2296
rect 5421 2164 5427 2236
rect 5469 2184 5475 2456
rect 5485 2297 5500 2303
rect 5485 2284 5491 2297
rect 5517 2283 5523 2376
rect 5533 2364 5539 2516
rect 5549 2324 5555 2496
rect 5565 2484 5571 2897
rect 5629 2884 5635 2916
rect 5645 2903 5651 3196
rect 5693 3104 5699 3316
rect 5805 3263 5811 3456
rect 5837 3424 5843 3436
rect 5837 3324 5843 3416
rect 5853 3404 5859 3516
rect 5885 3363 5891 3696
rect 5917 3524 5923 3676
rect 5901 3504 5907 3516
rect 5869 3357 5891 3363
rect 5821 3284 5827 3316
rect 5805 3257 5827 3263
rect 5821 3184 5827 3257
rect 5725 3104 5731 3136
rect 5789 3064 5795 3076
rect 5837 3024 5843 3236
rect 5853 3104 5859 3356
rect 5869 3264 5875 3357
rect 5885 3324 5891 3336
rect 5869 3104 5875 3256
rect 5901 3064 5907 3476
rect 5933 3464 5939 3736
rect 6013 3724 6019 3896
rect 6045 3823 6051 3896
rect 6029 3817 6051 3823
rect 5997 3684 6003 3716
rect 6029 3704 6035 3817
rect 6061 3743 6067 4036
rect 6125 3904 6131 3936
rect 6045 3737 6067 3743
rect 6045 3724 6051 3737
rect 6077 3724 6083 3856
rect 6093 3824 6099 3836
rect 6109 3764 6115 3776
rect 6013 3504 6019 3536
rect 5946 3414 5958 3416
rect 5931 3406 5933 3414
rect 5941 3406 5943 3414
rect 5951 3406 5953 3414
rect 5961 3406 5963 3414
rect 5971 3406 5973 3414
rect 5946 3404 5958 3406
rect 5997 3343 6003 3416
rect 6029 3404 6035 3656
rect 6061 3624 6067 3716
rect 6045 3483 6051 3616
rect 6093 3544 6099 3716
rect 6125 3684 6131 3736
rect 6141 3724 6147 3896
rect 6157 3864 6163 4036
rect 6189 4004 6195 4076
rect 6205 3904 6211 4116
rect 6221 4024 6227 4496
rect 6237 4484 6243 4516
rect 6301 4504 6307 4516
rect 6285 4304 6291 4316
rect 6317 4304 6323 4916
rect 6333 4764 6339 4936
rect 6349 4824 6355 4916
rect 6365 4703 6371 5336
rect 6381 5124 6387 5276
rect 6397 5264 6403 5318
rect 6381 5104 6387 5116
rect 6397 5063 6403 5216
rect 6429 5104 6435 5236
rect 6381 5057 6403 5063
rect 6381 4964 6387 5057
rect 6461 5044 6467 5236
rect 6397 5024 6403 5036
rect 6445 4944 6451 4956
rect 6429 4924 6435 4936
rect 6397 4903 6403 4916
rect 6445 4903 6451 4916
rect 6397 4897 6451 4903
rect 6477 4824 6483 5356
rect 6589 5284 6595 5318
rect 6621 5204 6627 5336
rect 6653 5164 6659 5236
rect 6525 5104 6531 5116
rect 6557 5104 6563 5136
rect 6621 5104 6627 5116
rect 6717 5102 6723 5116
rect 6541 5064 6547 5096
rect 6557 5084 6563 5096
rect 6493 4924 6499 4936
rect 6509 4904 6515 4936
rect 6541 4864 6547 5056
rect 6573 4944 6579 5056
rect 6589 5004 6595 5056
rect 6605 4943 6611 5016
rect 6653 4984 6659 5096
rect 6669 4984 6675 5016
rect 6621 4944 6627 4956
rect 6596 4937 6611 4943
rect 6445 4704 6451 4736
rect 6365 4697 6387 4703
rect 6333 4604 6339 4676
rect 6349 4524 6355 4696
rect 6381 4523 6387 4697
rect 6365 4517 6387 4523
rect 6333 4344 6339 4476
rect 6237 4103 6243 4296
rect 6253 4184 6259 4296
rect 6317 4264 6323 4276
rect 6317 4244 6323 4256
rect 6333 4244 6339 4256
rect 6301 4204 6307 4236
rect 6253 4124 6259 4176
rect 6285 4104 6291 4136
rect 6237 4097 6275 4103
rect 6221 4004 6227 4016
rect 6253 3984 6259 4016
rect 6221 3904 6227 3936
rect 6237 3923 6243 3976
rect 6237 3917 6259 3923
rect 6173 3824 6179 3896
rect 6237 3864 6243 3896
rect 6157 3744 6163 3796
rect 6173 3724 6179 3796
rect 6253 3744 6259 3917
rect 6269 3884 6275 4097
rect 6285 4024 6291 4096
rect 6301 4064 6307 4116
rect 6317 4044 6323 4136
rect 6333 4124 6339 4196
rect 6365 4123 6371 4517
rect 6397 4144 6403 4516
rect 6349 4117 6371 4123
rect 6333 3904 6339 3996
rect 6285 3884 6291 3896
rect 6301 3884 6307 3896
rect 6333 3864 6339 3896
rect 6349 3764 6355 4117
rect 6372 4097 6387 4103
rect 6365 3904 6371 3916
rect 6196 3737 6211 3743
rect 6205 3704 6211 3737
rect 6269 3724 6275 3756
rect 6093 3504 6099 3536
rect 6045 3477 6067 3483
rect 6045 3344 6051 3456
rect 5988 3337 6003 3343
rect 6029 3324 6035 3336
rect 5997 3284 6003 3316
rect 6045 3304 6051 3336
rect 6061 3324 6067 3477
rect 6141 3464 6147 3516
rect 6157 3504 6163 3616
rect 6173 3504 6179 3576
rect 6205 3464 6211 3696
rect 6221 3684 6227 3716
rect 6141 3424 6147 3436
rect 6077 3324 6083 3396
rect 6189 3384 6195 3436
rect 6173 3344 6179 3356
rect 6125 3324 6131 3336
rect 5997 3224 6003 3236
rect 6029 3184 6035 3276
rect 5981 3104 5987 3176
rect 6029 3104 6035 3116
rect 6061 3103 6067 3316
rect 6157 3304 6163 3336
rect 6205 3324 6211 3396
rect 6237 3324 6243 3576
rect 6253 3504 6259 3636
rect 6285 3624 6291 3716
rect 6285 3584 6291 3616
rect 6301 3544 6307 3736
rect 6317 3684 6323 3736
rect 6365 3724 6371 3756
rect 6381 3744 6387 4097
rect 6413 4064 6419 4136
rect 6429 4124 6435 4616
rect 6477 4524 6483 4636
rect 6445 4284 6451 4476
rect 6461 4302 6467 4336
rect 6461 4177 6476 4183
rect 6461 4164 6467 4177
rect 6461 4144 6467 4156
rect 6429 4084 6435 4096
rect 6413 3984 6419 3996
rect 6301 3504 6307 3536
rect 6333 3524 6339 3536
rect 6397 3524 6403 3876
rect 6413 3523 6419 3736
rect 6429 3724 6435 3856
rect 6445 3744 6451 3976
rect 6477 3844 6483 4116
rect 6461 3744 6467 3756
rect 6461 3684 6467 3716
rect 6413 3517 6428 3523
rect 6285 3363 6291 3436
rect 6317 3384 6323 3396
rect 6365 3384 6371 3496
rect 6397 3464 6403 3496
rect 6413 3484 6419 3517
rect 6301 3364 6307 3376
rect 6381 3364 6387 3376
rect 6269 3357 6291 3363
rect 6269 3324 6275 3357
rect 6397 3344 6403 3376
rect 6077 3184 6083 3276
rect 6061 3097 6083 3103
rect 5709 2904 5715 2916
rect 5645 2897 5660 2903
rect 5741 2884 5747 2916
rect 5581 2784 5587 2796
rect 5709 2702 5715 2716
rect 5773 2684 5779 2936
rect 5821 2924 5827 2936
rect 5837 2904 5843 2936
rect 5853 2924 5859 3056
rect 5933 3044 5939 3076
rect 5981 3064 5987 3096
rect 6013 3044 6019 3056
rect 5946 3014 5958 3016
rect 5931 3006 5933 3014
rect 5941 3006 5943 3014
rect 5951 3006 5953 3014
rect 5961 3006 5963 3014
rect 5971 3006 5973 3014
rect 5946 3004 5958 3006
rect 5789 2804 5795 2876
rect 5821 2724 5827 2836
rect 5853 2684 5859 2916
rect 5556 2317 5571 2323
rect 5508 2277 5523 2283
rect 5565 2264 5571 2317
rect 5645 2304 5651 2636
rect 5677 2564 5683 2676
rect 5773 2644 5779 2676
rect 5741 2544 5747 2556
rect 5837 2544 5843 2636
rect 5853 2544 5859 2676
rect 5773 2524 5779 2536
rect 5661 2377 5699 2383
rect 5661 2364 5667 2377
rect 5588 2297 5603 2303
rect 5597 2263 5603 2297
rect 5613 2284 5619 2296
rect 5629 2264 5635 2276
rect 5597 2257 5619 2263
rect 5405 2084 5411 2136
rect 5380 2077 5395 2083
rect 5389 2063 5395 2077
rect 5389 2057 5420 2063
rect 5437 2024 5443 2076
rect 5341 1944 5347 2016
rect 5316 1917 5331 1923
rect 5277 1784 5283 1796
rect 5149 1744 5155 1756
rect 5053 1484 5059 1596
rect 5133 1584 5139 1676
rect 5181 1664 5187 1696
rect 5085 1483 5091 1516
rect 5069 1477 5091 1483
rect 5005 1444 5011 1476
rect 5053 1384 5059 1476
rect 5069 1384 5075 1477
rect 5085 1444 5091 1456
rect 4957 1357 4979 1363
rect 4893 1304 4899 1356
rect 4916 1317 4931 1323
rect 4845 1217 4867 1223
rect 4845 1184 4851 1217
rect 4877 1184 4883 1296
rect 4925 1224 4931 1317
rect 4909 1104 4915 1116
rect 4900 1077 4915 1083
rect 4813 1004 4819 1036
rect 4797 977 4812 983
rect 4749 917 4764 923
rect 4749 904 4755 917
rect 4765 884 4771 896
rect 4788 877 4803 883
rect 4701 784 4707 876
rect 4797 784 4803 877
rect 4701 584 4707 656
rect 4701 504 4707 516
rect 4701 424 4707 496
rect 4701 284 4707 396
rect 4717 284 4723 536
rect 4749 524 4755 656
rect 4829 604 4835 1056
rect 4909 984 4915 1077
rect 4845 944 4851 976
rect 4925 824 4931 1216
rect 4941 1144 4947 1356
rect 4973 1324 4979 1357
rect 4957 1304 4963 1316
rect 4941 964 4947 1036
rect 4941 904 4947 936
rect 4957 924 4963 1056
rect 4893 683 4899 796
rect 4925 684 4931 736
rect 4973 684 4979 996
rect 4989 864 4995 1296
rect 5053 1204 5059 1296
rect 5117 1264 5123 1536
rect 5181 1524 5187 1656
rect 5213 1604 5219 1736
rect 5261 1724 5267 1756
rect 5293 1684 5299 1736
rect 5309 1724 5315 1836
rect 5325 1664 5331 1917
rect 5341 1764 5347 1936
rect 5373 1924 5379 1976
rect 5453 1924 5459 2116
rect 5485 2104 5491 2196
rect 5501 2184 5507 2256
rect 5565 2184 5571 2256
rect 5613 2243 5619 2257
rect 5645 2243 5651 2256
rect 5613 2237 5651 2243
rect 5661 2204 5667 2336
rect 5677 2264 5683 2356
rect 5693 2344 5699 2377
rect 5693 2264 5699 2316
rect 5741 2284 5747 2456
rect 5837 2444 5843 2536
rect 5885 2524 5891 2956
rect 5981 2864 5987 2936
rect 5997 2924 6003 3016
rect 5997 2884 6003 2896
rect 6013 2824 6019 2996
rect 6029 2924 6035 3096
rect 6061 3044 6067 3056
rect 6061 2804 6067 2836
rect 5901 2644 5907 2696
rect 6013 2644 6019 2656
rect 5946 2614 5958 2616
rect 5931 2606 5933 2614
rect 5941 2606 5943 2614
rect 5951 2606 5953 2614
rect 5961 2606 5963 2614
rect 5971 2606 5973 2614
rect 5946 2604 5958 2606
rect 5885 2504 5891 2516
rect 5757 2304 5763 2416
rect 5517 2064 5523 2136
rect 5581 2124 5587 2136
rect 5597 2124 5603 2196
rect 5789 2184 5795 2336
rect 5805 2304 5811 2336
rect 5821 2264 5827 2276
rect 5837 2264 5843 2356
rect 5869 2304 5875 2316
rect 5885 2284 5891 2456
rect 5789 2124 5795 2156
rect 5645 2104 5651 2116
rect 5533 1944 5539 1996
rect 5357 1904 5363 1916
rect 5357 1744 5363 1896
rect 5469 1864 5475 1936
rect 5533 1924 5539 1936
rect 5341 1723 5347 1736
rect 5341 1717 5356 1723
rect 5389 1704 5395 1776
rect 5341 1584 5347 1676
rect 5357 1664 5363 1676
rect 5293 1524 5299 1556
rect 5373 1524 5379 1696
rect 5405 1684 5411 1756
rect 5421 1724 5427 1736
rect 5421 1683 5427 1716
rect 5437 1704 5443 1776
rect 5453 1724 5459 1736
rect 5485 1724 5491 1736
rect 5421 1677 5443 1683
rect 5405 1663 5411 1676
rect 5405 1657 5427 1663
rect 5389 1544 5395 1636
rect 5405 1584 5411 1596
rect 5133 1244 5139 1496
rect 5213 1464 5219 1476
rect 5245 1463 5251 1496
rect 5373 1484 5379 1496
rect 5220 1457 5251 1463
rect 5181 1384 5187 1416
rect 5197 1324 5203 1416
rect 5229 1364 5235 1457
rect 5293 1364 5299 1476
rect 5309 1384 5315 1416
rect 5245 1324 5251 1356
rect 5005 1104 5011 1156
rect 5085 1124 5091 1176
rect 5101 1104 5107 1116
rect 5117 1064 5123 1236
rect 5197 1184 5203 1236
rect 5005 904 5011 1016
rect 5037 944 5043 956
rect 5085 924 5091 1036
rect 5133 984 5139 1076
rect 5165 1064 5171 1096
rect 5101 944 5107 956
rect 5197 944 5203 1076
rect 4989 724 4995 836
rect 4996 717 5004 723
rect 5037 684 5043 716
rect 5069 684 5075 916
rect 5149 904 5155 916
rect 5101 824 5107 876
rect 5165 844 5171 916
rect 5213 804 5219 1056
rect 5229 964 5235 1296
rect 5261 1224 5267 1356
rect 5293 1283 5299 1356
rect 5277 1277 5299 1283
rect 5277 1084 5283 1277
rect 5309 1244 5315 1276
rect 5309 1184 5315 1216
rect 5293 1084 5299 1096
rect 5277 1064 5283 1076
rect 5261 1024 5267 1036
rect 5261 964 5267 1016
rect 5277 964 5283 1056
rect 5325 944 5331 1476
rect 5405 1384 5411 1556
rect 5421 1544 5427 1657
rect 5437 1504 5443 1677
rect 5453 1604 5459 1656
rect 5453 1584 5459 1596
rect 5421 1444 5427 1496
rect 5341 1064 5347 1236
rect 5357 1104 5363 1276
rect 5373 1164 5379 1196
rect 5373 1104 5379 1156
rect 5373 1024 5379 1096
rect 5245 784 5251 916
rect 5325 884 5331 896
rect 5325 784 5331 796
rect 5229 724 5235 736
rect 5277 704 5283 736
rect 5277 684 5283 696
rect 5293 684 5299 696
rect 4884 677 4899 683
rect 4669 197 4691 203
rect 4621 -23 4643 -17
rect 4669 -23 4675 197
rect 4733 184 4739 396
rect 4797 384 4803 596
rect 4877 584 4883 676
rect 4973 664 4979 676
rect 5261 664 5267 676
rect 4804 377 4819 383
rect 4749 324 4755 376
rect 4749 124 4755 156
rect 4813 123 4819 377
rect 4845 264 4851 556
rect 4893 524 4899 636
rect 4877 504 4883 518
rect 4861 284 4867 376
rect 4909 324 4915 616
rect 4941 564 4947 656
rect 5069 584 5075 596
rect 5021 524 5027 556
rect 4941 284 4947 516
rect 5021 384 5027 516
rect 4973 302 4979 356
rect 5133 343 5139 496
rect 5165 424 5171 516
rect 5261 404 5267 656
rect 5309 644 5315 776
rect 5277 524 5283 576
rect 5293 524 5299 536
rect 5124 337 5139 343
rect 5117 324 5123 336
rect 5197 304 5203 316
rect 5245 304 5251 336
rect 4797 117 4819 123
rect 4717 -23 4723 76
rect 4749 -23 4755 16
rect 4797 -23 4803 117
rect 4829 104 4835 216
rect 4877 144 4883 276
rect 4893 104 4899 236
rect 4925 124 4931 176
rect 4989 124 4995 276
rect 5037 244 5043 296
rect 5117 104 5123 236
rect 5165 144 5171 276
rect 5261 264 5267 276
rect 5293 264 5299 456
rect 5325 443 5331 736
rect 5341 724 5347 916
rect 5373 784 5379 816
rect 5389 804 5395 1276
rect 5421 1264 5427 1436
rect 5469 1364 5475 1496
rect 5485 1404 5491 1716
rect 5501 1483 5507 1736
rect 5517 1704 5523 1856
rect 5533 1784 5539 1876
rect 5549 1784 5555 1836
rect 5533 1677 5548 1683
rect 5533 1584 5539 1677
rect 5549 1584 5555 1656
rect 5565 1643 5571 2056
rect 5597 1923 5603 2016
rect 5613 1944 5619 2036
rect 5597 1917 5619 1923
rect 5613 1784 5619 1917
rect 5741 1884 5747 2116
rect 5805 2104 5811 2236
rect 5853 2204 5859 2236
rect 5869 2144 5875 2176
rect 5885 2124 5891 2196
rect 5901 2064 5907 2296
rect 5933 2244 5939 2316
rect 5946 2214 5958 2216
rect 5931 2206 5933 2214
rect 5941 2206 5943 2214
rect 5951 2206 5953 2214
rect 5961 2206 5963 2214
rect 5971 2206 5973 2214
rect 5946 2204 5958 2206
rect 5917 2124 5923 2156
rect 5933 2144 5939 2156
rect 5949 2104 5955 2136
rect 5917 2024 5923 2036
rect 5997 1944 6003 2496
rect 6013 2304 6019 2436
rect 6029 2184 6035 2396
rect 6077 2303 6083 3097
rect 6093 3004 6099 3236
rect 6109 3104 6115 3156
rect 6093 2924 6099 2976
rect 6109 2884 6115 2916
rect 6125 2864 6131 3036
rect 6125 2703 6131 2836
rect 6141 2724 6147 3296
rect 6173 3224 6179 3316
rect 6285 3264 6291 3336
rect 6157 3104 6163 3196
rect 6189 3184 6195 3196
rect 6157 3084 6163 3096
rect 6173 2963 6179 3076
rect 6221 3044 6227 3076
rect 6253 3064 6259 3116
rect 6301 3064 6307 3096
rect 6317 3084 6323 3296
rect 6333 3144 6339 3316
rect 6349 3184 6355 3316
rect 6317 3024 6323 3076
rect 6157 2957 6179 2963
rect 6125 2697 6140 2703
rect 6093 2664 6099 2676
rect 6109 2564 6115 2696
rect 6109 2484 6115 2536
rect 6141 2524 6147 2536
rect 6109 2384 6115 2476
rect 6125 2384 6131 2436
rect 6077 2297 6099 2303
rect 6029 2143 6035 2176
rect 6013 2137 6035 2143
rect 6013 2124 6019 2137
rect 6045 2123 6051 2276
rect 6061 2244 6067 2296
rect 6061 2144 6067 2216
rect 6077 2164 6083 2276
rect 6093 2124 6099 2297
rect 6045 2117 6076 2123
rect 6029 2103 6035 2116
rect 6125 2104 6131 2116
rect 6013 2097 6035 2103
rect 6013 2024 6019 2097
rect 6029 1964 6035 2056
rect 5789 1904 5795 1936
rect 5901 1904 5907 1936
rect 5661 1784 5667 1816
rect 5709 1784 5715 1796
rect 5741 1784 5747 1876
rect 5805 1784 5811 1896
rect 5933 1884 5939 1936
rect 5988 1917 6003 1923
rect 5581 1704 5587 1736
rect 5645 1704 5651 1736
rect 5693 1704 5699 1736
rect 5581 1664 5587 1696
rect 5565 1637 5587 1643
rect 5524 1497 5539 1503
rect 5501 1477 5523 1483
rect 5501 1364 5507 1436
rect 5517 1384 5523 1477
rect 5421 944 5427 1076
rect 5453 1004 5459 1336
rect 5469 1124 5475 1316
rect 5485 1304 5491 1336
rect 5533 1324 5539 1497
rect 5581 1463 5587 1637
rect 5597 1524 5603 1676
rect 5597 1484 5603 1516
rect 5581 1457 5603 1463
rect 5581 1324 5587 1436
rect 5597 1384 5603 1457
rect 5533 1124 5539 1276
rect 5597 1184 5603 1276
rect 5613 1124 5619 1636
rect 5629 1604 5635 1656
rect 5629 1524 5635 1596
rect 5645 1563 5651 1676
rect 5693 1604 5699 1676
rect 5709 1624 5715 1756
rect 5741 1724 5747 1736
rect 5725 1564 5731 1676
rect 5645 1557 5667 1563
rect 5661 1544 5667 1557
rect 5661 1504 5667 1536
rect 5661 1384 5667 1476
rect 5709 1384 5715 1480
rect 5725 1464 5731 1476
rect 5533 1104 5539 1116
rect 5629 1103 5635 1116
rect 5588 1097 5635 1103
rect 5469 924 5475 976
rect 5405 904 5411 916
rect 5501 844 5507 936
rect 5533 924 5539 1016
rect 5565 924 5571 956
rect 5341 664 5347 716
rect 5357 564 5363 776
rect 5405 664 5411 696
rect 5421 664 5427 796
rect 5453 724 5459 756
rect 5357 524 5363 556
rect 5421 544 5427 636
rect 5453 563 5459 716
rect 5469 604 5475 816
rect 5501 684 5507 836
rect 5533 804 5539 916
rect 5613 903 5619 1036
rect 5629 1024 5635 1036
rect 5645 984 5651 1176
rect 5645 964 5651 976
rect 5693 964 5699 1176
rect 5709 1064 5715 1236
rect 5725 1124 5731 1136
rect 5741 1064 5747 1436
rect 5757 1324 5763 1776
rect 5789 1724 5795 1756
rect 5821 1684 5827 1736
rect 5837 1724 5843 1876
rect 5853 1724 5859 1756
rect 5901 1744 5907 1816
rect 5946 1814 5958 1816
rect 5931 1806 5933 1814
rect 5941 1806 5943 1814
rect 5951 1806 5953 1814
rect 5961 1806 5963 1814
rect 5971 1806 5973 1814
rect 5946 1804 5958 1806
rect 5997 1783 6003 1917
rect 6013 1904 6019 1916
rect 6029 1883 6035 1956
rect 6020 1877 6035 1883
rect 6045 1804 6051 2036
rect 6077 1964 6083 1996
rect 6141 1984 6147 2036
rect 6077 1904 6083 1936
rect 6141 1924 6147 1936
rect 6157 1903 6163 2957
rect 6269 2904 6275 2996
rect 6349 2964 6355 2976
rect 6317 2944 6323 2956
rect 6381 2944 6387 2976
rect 6397 2924 6403 3176
rect 6461 3083 6467 3656
rect 6477 3504 6483 3716
rect 6493 3664 6499 4656
rect 6525 4264 6531 4276
rect 6509 3884 6515 4076
rect 6509 3704 6515 3836
rect 6541 3784 6547 4816
rect 6589 4663 6595 4916
rect 6605 4884 6611 4916
rect 6637 4904 6643 4916
rect 6653 4844 6659 4936
rect 6669 4844 6675 4896
rect 6605 4684 6611 4756
rect 6653 4704 6659 4716
rect 6669 4684 6675 4696
rect 6685 4684 6691 5076
rect 6717 4964 6723 5056
rect 6717 4944 6723 4956
rect 6749 4924 6755 4996
rect 6765 4944 6771 4956
rect 6701 4864 6707 4916
rect 6589 4657 6611 4663
rect 6605 4584 6611 4657
rect 6685 4584 6691 4616
rect 6573 4284 6579 4336
rect 6589 4283 6595 4476
rect 6605 4384 6611 4436
rect 6605 4304 6611 4316
rect 6621 4284 6627 4536
rect 6701 4524 6707 4856
rect 6781 4704 6787 5318
rect 6845 5164 6851 5236
rect 6909 5204 6915 5316
rect 6845 5004 6851 5036
rect 6845 4924 6851 4996
rect 6829 4864 6835 4916
rect 6861 4844 6867 5096
rect 6893 5064 6899 5096
rect 6797 4704 6803 4736
rect 6717 4544 6723 4696
rect 6653 4504 6659 4516
rect 6717 4484 6723 4516
rect 6749 4484 6755 4596
rect 6701 4477 6716 4483
rect 6637 4324 6643 4336
rect 6653 4324 6659 4476
rect 6685 4304 6691 4376
rect 6701 4304 6707 4477
rect 6589 4277 6611 4283
rect 6589 4124 6595 4196
rect 6605 4043 6611 4277
rect 6637 4144 6643 4156
rect 6669 4124 6675 4296
rect 6717 4204 6723 4436
rect 6765 4364 6771 4516
rect 6749 4304 6755 4356
rect 6781 4343 6787 4656
rect 6829 4564 6835 4836
rect 6797 4404 6803 4516
rect 6765 4337 6787 4343
rect 6685 4144 6691 4196
rect 6669 4084 6675 4096
rect 6605 4037 6627 4043
rect 6605 3884 6611 3896
rect 6589 3784 6595 3796
rect 6525 3724 6531 3756
rect 6573 3724 6579 3756
rect 6477 3264 6483 3476
rect 6493 3344 6499 3456
rect 6509 3244 6515 3696
rect 6557 3624 6563 3716
rect 6525 3504 6531 3516
rect 6525 3326 6531 3476
rect 6541 3464 6547 3516
rect 6557 3464 6563 3616
rect 6605 3544 6611 3876
rect 6621 3724 6627 4037
rect 6637 3904 6643 3916
rect 6653 3844 6659 3896
rect 6701 3884 6707 4116
rect 6717 3964 6723 4136
rect 6653 3784 6659 3816
rect 6621 3684 6627 3716
rect 6685 3664 6691 3836
rect 6701 3824 6707 3856
rect 6573 3484 6579 3536
rect 6669 3504 6675 3516
rect 6589 3484 6595 3496
rect 6589 3324 6595 3456
rect 6621 3444 6627 3496
rect 6605 3437 6620 3443
rect 6605 3324 6611 3437
rect 6669 3324 6675 3496
rect 6685 3484 6691 3496
rect 6701 3304 6707 3476
rect 6717 3464 6723 3776
rect 6749 3624 6755 4196
rect 6765 3864 6771 4337
rect 6797 4304 6803 4316
rect 6781 4244 6787 4276
rect 6797 4124 6803 4296
rect 6813 3964 6819 4536
rect 6861 4524 6867 4576
rect 6845 4384 6851 4516
rect 6877 4463 6883 5036
rect 6909 4984 6915 5096
rect 6925 5084 6931 5176
rect 6909 4904 6915 4936
rect 6925 4924 6931 5076
rect 6957 5023 6963 5056
rect 6973 5044 6979 5056
rect 6941 5017 6963 5023
rect 6941 4984 6947 5017
rect 6957 4924 6963 4956
rect 6964 4917 6979 4923
rect 6925 4683 6931 4916
rect 6973 4884 6979 4917
rect 6909 4677 6931 4683
rect 6909 4624 6915 4677
rect 6989 4644 6995 4696
rect 6925 4584 6931 4636
rect 6957 4524 6963 4576
rect 6909 4484 6915 4516
rect 6877 4457 6899 4463
rect 6877 4424 6883 4436
rect 6845 4284 6851 4296
rect 6877 4284 6883 4336
rect 6877 4264 6883 4276
rect 6829 4144 6835 4156
rect 6797 3904 6803 3956
rect 6829 3903 6835 4136
rect 6813 3897 6835 3903
rect 6781 3884 6787 3896
rect 6781 3844 6787 3876
rect 6765 3724 6771 3836
rect 6813 3744 6819 3897
rect 6836 3877 6851 3883
rect 6845 3724 6851 3877
rect 6877 3864 6883 3936
rect 6733 3564 6739 3596
rect 6717 3344 6723 3376
rect 6509 3143 6515 3236
rect 6621 3224 6627 3236
rect 6669 3164 6675 3176
rect 6509 3137 6531 3143
rect 6525 3104 6531 3137
rect 6605 3084 6611 3136
rect 6669 3104 6675 3156
rect 6653 3084 6659 3096
rect 6445 3077 6467 3083
rect 6285 2904 6291 2918
rect 6429 2923 6435 2936
rect 6413 2917 6435 2923
rect 6173 2124 6179 2716
rect 6237 2704 6243 2816
rect 6205 2624 6211 2696
rect 6205 2544 6211 2556
rect 6237 2544 6243 2696
rect 6269 2644 6275 2656
rect 6253 2584 6259 2636
rect 6189 2504 6195 2516
rect 6205 2304 6211 2476
rect 6269 2464 6275 2636
rect 6285 2564 6291 2696
rect 6301 2684 6307 2816
rect 6333 2664 6339 2676
rect 6317 2564 6323 2656
rect 6285 2524 6291 2536
rect 6381 2524 6387 2836
rect 6397 2783 6403 2916
rect 6413 2904 6419 2917
rect 6397 2777 6419 2783
rect 6413 2544 6419 2777
rect 6445 2644 6451 3077
rect 6461 2964 6467 3056
rect 6557 3044 6563 3056
rect 6493 2964 6499 2996
rect 6461 2784 6467 2956
rect 6493 2924 6499 2936
rect 6509 2924 6515 2976
rect 6557 2924 6563 3036
rect 6477 2904 6483 2916
rect 6557 2904 6563 2916
rect 6461 2704 6467 2716
rect 6285 2304 6291 2436
rect 6333 2344 6339 2516
rect 6461 2504 6467 2536
rect 6477 2524 6483 2876
rect 6509 2684 6515 2776
rect 6541 2664 6547 2836
rect 6573 2704 6579 3016
rect 6589 2944 6595 2976
rect 6589 2684 6595 2936
rect 6605 2704 6611 2716
rect 6621 2683 6627 2936
rect 6605 2677 6627 2683
rect 6509 2564 6515 2596
rect 6525 2524 6531 2536
rect 6509 2517 6524 2523
rect 6397 2304 6403 2396
rect 6221 2284 6227 2296
rect 6253 2284 6259 2296
rect 6189 2103 6195 2136
rect 6221 2124 6227 2276
rect 6333 2264 6339 2276
rect 6349 2264 6355 2296
rect 6253 2144 6259 2256
rect 6253 2104 6259 2136
rect 6285 2124 6291 2256
rect 6317 2244 6323 2256
rect 6173 2097 6195 2103
rect 6173 1984 6179 2097
rect 6301 2103 6307 2176
rect 6317 2124 6323 2176
rect 6381 2144 6387 2156
rect 6413 2124 6419 2436
rect 6429 2304 6435 2336
rect 6445 2304 6451 2336
rect 6333 2117 6348 2123
rect 6333 2103 6339 2117
rect 6429 2123 6435 2296
rect 6445 2264 6451 2296
rect 6461 2264 6467 2496
rect 6477 2464 6483 2516
rect 6477 2424 6483 2436
rect 6493 2304 6499 2396
rect 6509 2324 6515 2517
rect 6525 2384 6531 2436
rect 6516 2317 6531 2323
rect 6525 2304 6531 2317
rect 6509 2284 6515 2296
rect 6461 2204 6467 2236
rect 6493 2164 6499 2256
rect 6452 2137 6467 2143
rect 6429 2117 6444 2123
rect 6301 2097 6339 2103
rect 6445 2064 6451 2116
rect 6205 1984 6211 1996
rect 6173 1904 6179 1976
rect 6301 1904 6307 1936
rect 6365 1904 6371 2056
rect 6413 1984 6419 2036
rect 6461 1984 6467 2137
rect 6477 1943 6483 2136
rect 6493 2104 6499 2156
rect 6509 2144 6515 2276
rect 6525 2124 6531 2256
rect 6509 2103 6515 2116
rect 6509 2097 6524 2103
rect 6541 2084 6547 2636
rect 6557 2604 6563 2676
rect 6557 2564 6563 2596
rect 6589 2584 6595 2656
rect 6557 2264 6563 2416
rect 6573 2364 6579 2476
rect 6573 2264 6579 2336
rect 6589 2303 6595 2576
rect 6605 2544 6611 2677
rect 6621 2624 6627 2636
rect 6637 2543 6643 2796
rect 6653 2764 6659 2936
rect 6685 2924 6691 3296
rect 6701 3184 6707 3236
rect 6733 3183 6739 3556
rect 6749 3464 6755 3476
rect 6749 3244 6755 3456
rect 6781 3363 6787 3656
rect 6861 3604 6867 3856
rect 6877 3764 6883 3776
rect 6877 3504 6883 3736
rect 6797 3443 6803 3456
rect 6797 3437 6812 3443
rect 6797 3424 6803 3437
rect 6765 3357 6787 3363
rect 6765 3324 6771 3357
rect 6781 3324 6787 3336
rect 6724 3177 6739 3183
rect 6797 3183 6803 3356
rect 6877 3344 6883 3496
rect 6893 3484 6899 4457
rect 6925 4164 6931 4176
rect 6957 4124 6963 4136
rect 6957 3924 6963 4116
rect 6925 3903 6931 3916
rect 6916 3897 6931 3903
rect 6909 3784 6915 3816
rect 6925 3744 6931 3897
rect 6925 3724 6931 3736
rect 6941 3704 6947 3716
rect 6925 3504 6931 3536
rect 6973 3424 6979 3796
rect 6989 3564 6995 4616
rect 7005 4544 7011 5316
rect 7037 5204 7043 5236
rect 7037 4964 7043 5196
rect 7101 5104 7107 5316
rect 7053 4924 7059 5036
rect 7069 4884 7075 5096
rect 7101 5084 7107 5096
rect 7085 4944 7091 5076
rect 7172 5037 7187 5043
rect 7005 4484 7011 4516
rect 7005 4264 7011 4476
rect 7021 4284 7027 4636
rect 7053 4623 7059 4694
rect 7085 4684 7091 4936
rect 7149 4683 7155 4876
rect 7165 4744 7171 4956
rect 7181 4864 7187 5037
rect 7245 4984 7251 5316
rect 7357 5224 7363 5336
rect 7213 4924 7219 4976
rect 7197 4884 7203 4916
rect 7149 4677 7171 4683
rect 7053 4617 7075 4623
rect 7069 4584 7075 4617
rect 7101 4564 7107 4576
rect 7053 4544 7059 4556
rect 7037 4504 7043 4516
rect 7117 4504 7123 4676
rect 7133 4544 7139 4556
rect 7133 4524 7139 4536
rect 7085 4284 7091 4356
rect 7021 4124 7027 4236
rect 7053 4144 7059 4236
rect 7101 4184 7107 4396
rect 7117 4324 7123 4336
rect 7117 4304 7123 4316
rect 7053 4044 7059 4136
rect 7005 3584 7011 3636
rect 7005 3464 7011 3476
rect 6989 3384 6995 3396
rect 6877 3324 6883 3336
rect 6909 3304 6915 3316
rect 6788 3177 6803 3183
rect 6749 3104 6755 3136
rect 6765 3064 6771 3076
rect 6829 3064 6835 3076
rect 6685 2704 6691 2756
rect 6701 2704 6707 3036
rect 6717 3024 6723 3036
rect 6749 2904 6755 2916
rect 6765 2904 6771 3056
rect 6877 3044 6883 3076
rect 6941 3064 6947 3096
rect 6781 2924 6787 3036
rect 6861 2964 6867 2976
rect 6893 2944 6899 3036
rect 6941 3004 6947 3056
rect 6909 2984 6915 2996
rect 6957 2984 6963 3036
rect 6973 2964 6979 3116
rect 6989 3024 6995 3056
rect 6653 2644 6659 2696
rect 6669 2684 6675 2696
rect 6628 2537 6643 2543
rect 6605 2524 6611 2536
rect 6669 2524 6675 2656
rect 6685 2564 6691 2696
rect 6701 2684 6707 2696
rect 6701 2564 6707 2676
rect 6685 2544 6691 2556
rect 6621 2484 6627 2516
rect 6685 2503 6691 2536
rect 6717 2524 6723 2636
rect 6749 2604 6755 2656
rect 6669 2497 6691 2503
rect 6701 2503 6707 2516
rect 6701 2497 6723 2503
rect 6605 2304 6611 2316
rect 6589 2297 6604 2303
rect 6653 2284 6659 2316
rect 6669 2304 6675 2497
rect 6676 2297 6691 2303
rect 6557 2244 6563 2256
rect 6573 2144 6579 2156
rect 6637 2124 6643 2136
rect 6621 2104 6627 2116
rect 6461 1937 6483 1943
rect 6397 1904 6403 1936
rect 6461 1904 6467 1937
rect 6541 1924 6547 2076
rect 6477 1904 6483 1916
rect 6141 1897 6163 1903
rect 6077 1824 6083 1876
rect 5981 1777 6003 1783
rect 5885 1644 5891 1736
rect 5981 1704 5987 1777
rect 6013 1763 6019 1796
rect 5997 1757 6019 1763
rect 5997 1744 6003 1757
rect 6045 1744 6051 1776
rect 6013 1703 6019 1736
rect 5997 1697 6019 1703
rect 5981 1664 5987 1696
rect 5892 1537 5923 1543
rect 5917 1523 5923 1537
rect 5997 1524 6003 1697
rect 6077 1684 6083 1718
rect 5917 1517 5932 1523
rect 5773 1464 5779 1476
rect 5789 1464 5795 1496
rect 5853 1484 5859 1496
rect 5869 1464 5875 1476
rect 5837 1304 5843 1436
rect 5901 1384 5907 1496
rect 5997 1464 6003 1516
rect 6045 1504 6051 1536
rect 6061 1464 6067 1476
rect 5946 1414 5958 1416
rect 5931 1406 5933 1414
rect 5941 1406 5943 1414
rect 5951 1406 5953 1414
rect 5961 1406 5963 1414
rect 5971 1406 5973 1414
rect 5946 1404 5958 1406
rect 6013 1384 6019 1436
rect 6061 1424 6067 1456
rect 6077 1444 6083 1496
rect 5933 1364 5939 1376
rect 6061 1364 6067 1416
rect 5837 1184 5843 1296
rect 5853 1184 5859 1276
rect 5757 1064 5763 1096
rect 5613 897 5628 903
rect 5501 664 5507 676
rect 5469 564 5475 596
rect 5501 584 5507 596
rect 5533 584 5539 796
rect 5645 744 5651 936
rect 5565 724 5571 736
rect 5677 704 5683 836
rect 5693 704 5699 936
rect 5741 884 5747 1036
rect 5757 984 5763 996
rect 5773 984 5779 1076
rect 5789 883 5795 1036
rect 5805 984 5811 1076
rect 5821 1064 5827 1076
rect 5853 964 5859 1056
rect 5869 943 5875 1036
rect 5885 963 5891 996
rect 5901 984 5907 1076
rect 5988 1037 6003 1043
rect 5946 1014 5958 1016
rect 5931 1006 5933 1014
rect 5941 1006 5943 1014
rect 5951 1006 5953 1014
rect 5961 1006 5963 1014
rect 5971 1006 5973 1014
rect 5946 1004 5958 1006
rect 5917 963 5923 976
rect 5885 957 5923 963
rect 5933 944 5939 956
rect 5853 937 5875 943
rect 5789 877 5811 883
rect 5789 784 5795 856
rect 5709 724 5715 756
rect 5805 724 5811 877
rect 5821 864 5827 896
rect 5853 864 5859 937
rect 5437 557 5459 563
rect 5316 437 5331 443
rect 5309 324 5315 436
rect 5357 304 5363 396
rect 5389 344 5395 436
rect 5341 257 5347 276
rect 5197 164 5203 196
rect 5213 124 5219 236
rect 5261 144 5267 256
rect 5277 124 5283 136
rect 5309 104 5315 236
rect 5357 164 5363 296
rect 5421 283 5427 536
rect 5437 324 5443 557
rect 5565 544 5571 696
rect 5613 684 5619 696
rect 5805 684 5811 696
rect 5837 683 5843 836
rect 5853 704 5859 756
rect 5885 684 5891 696
rect 5837 677 5859 683
rect 5597 544 5603 676
rect 5613 584 5619 616
rect 5453 504 5459 536
rect 5469 504 5475 516
rect 5581 504 5587 516
rect 5629 503 5635 636
rect 5620 497 5635 503
rect 5645 484 5651 576
rect 5661 524 5667 556
rect 5693 544 5699 596
rect 5677 504 5683 516
rect 5629 477 5644 483
rect 5629 464 5635 477
rect 5485 324 5491 356
rect 5549 324 5555 336
rect 5485 284 5491 316
rect 5421 277 5436 283
rect 5405 164 5411 196
rect 5421 124 5427 136
rect 5437 103 5443 236
rect 5453 124 5459 196
rect 5469 144 5475 256
rect 5501 124 5507 156
rect 5428 97 5443 103
rect 5517 103 5523 236
rect 5549 124 5555 236
rect 5597 224 5603 436
rect 5645 404 5651 456
rect 5645 304 5651 396
rect 5661 364 5667 436
rect 5677 264 5683 496
rect 5693 304 5699 516
rect 5709 504 5715 636
rect 5741 563 5747 636
rect 5821 624 5827 636
rect 5725 557 5747 563
rect 5709 284 5715 416
rect 5725 324 5731 557
rect 5773 504 5779 536
rect 5741 424 5747 436
rect 5757 264 5763 296
rect 5661 164 5667 216
rect 5677 184 5683 236
rect 5693 164 5699 236
rect 5773 204 5779 236
rect 5597 124 5603 136
rect 5741 124 5747 196
rect 5789 124 5795 616
rect 5805 564 5811 576
rect 5805 304 5811 396
rect 5821 384 5827 556
rect 5821 284 5827 376
rect 5837 304 5843 616
rect 5853 284 5859 677
rect 5869 564 5875 676
rect 5901 624 5907 916
rect 5933 824 5939 916
rect 5917 704 5923 796
rect 5933 664 5939 796
rect 5997 784 6003 1037
rect 6013 924 6019 976
rect 6077 944 6083 1236
rect 6093 1084 6099 1736
rect 6109 1584 6115 1676
rect 6125 1464 6131 1576
rect 6141 1504 6147 1897
rect 6173 1884 6179 1896
rect 6189 1824 6195 1876
rect 6237 1784 6243 1876
rect 6349 1864 6355 1896
rect 6445 1864 6451 1896
rect 6541 1883 6547 1916
rect 6621 1904 6627 1916
rect 6573 1884 6579 1896
rect 6669 1884 6675 1916
rect 6685 1904 6691 2297
rect 6717 2124 6723 2497
rect 6765 2204 6771 2856
rect 6829 2784 6835 2936
rect 6941 2884 6947 2916
rect 6973 2804 6979 2916
rect 6829 2744 6835 2776
rect 6797 2724 6803 2736
rect 6781 2524 6787 2656
rect 6797 2584 6803 2596
rect 6813 2544 6819 2596
rect 6861 2544 6867 2656
rect 6797 2404 6803 2436
rect 6877 2384 6883 2696
rect 6909 2524 6915 2656
rect 6925 2624 6931 2694
rect 6957 2544 6963 2676
rect 6989 2544 6995 2556
rect 7005 2544 7011 3416
rect 7021 2664 7027 3776
rect 7037 3684 7043 3756
rect 7053 3684 7059 3956
rect 7117 3924 7123 4296
rect 7069 3724 7075 3816
rect 7085 3764 7091 3876
rect 7085 3744 7091 3756
rect 7037 3484 7043 3496
rect 7069 3484 7075 3696
rect 7085 3504 7091 3656
rect 7117 3643 7123 3896
rect 7133 3784 7139 4376
rect 7149 4284 7155 4516
rect 7165 4344 7171 4677
rect 7181 4584 7187 4736
rect 7181 4343 7187 4536
rect 7197 4383 7203 4836
rect 7213 4604 7219 4856
rect 7261 4744 7267 5096
rect 7325 4964 7331 5156
rect 7357 4964 7363 5196
rect 7277 4884 7283 4916
rect 7325 4884 7331 4916
rect 7245 4684 7251 4696
rect 7213 4564 7219 4596
rect 7245 4584 7251 4676
rect 7277 4624 7283 4836
rect 7245 4524 7251 4556
rect 7197 4377 7219 4383
rect 7181 4337 7203 4343
rect 7156 4277 7171 4283
rect 7165 4243 7171 4277
rect 7181 4243 7187 4276
rect 7165 4237 7187 4243
rect 7149 3984 7155 4036
rect 7165 3904 7171 4237
rect 7197 4223 7203 4337
rect 7181 4217 7203 4223
rect 7181 4084 7187 4217
rect 7149 3897 7164 3903
rect 7149 3724 7155 3897
rect 7165 3744 7171 3836
rect 7181 3784 7187 4016
rect 7197 3863 7203 4176
rect 7213 4164 7219 4377
rect 7213 3984 7219 4076
rect 7229 3904 7235 4136
rect 7229 3884 7235 3896
rect 7197 3857 7212 3863
rect 7245 3724 7251 3836
rect 7149 3704 7155 3716
rect 7101 3637 7123 3643
rect 7069 3303 7075 3476
rect 7101 3364 7107 3637
rect 7117 3524 7123 3616
rect 7133 3504 7139 3676
rect 7117 3326 7123 3436
rect 7133 3404 7139 3496
rect 7053 3297 7075 3303
rect 7053 3204 7059 3297
rect 7069 3144 7075 3256
rect 7069 3064 7075 3136
rect 7117 3084 7123 3096
rect 7053 3044 7059 3056
rect 7133 3044 7139 3076
rect 7101 2984 7107 2996
rect 7037 2944 7043 2956
rect 7053 2904 7059 2976
rect 7117 2964 7123 3036
rect 7149 2984 7155 3656
rect 7165 3584 7171 3716
rect 7245 3484 7251 3716
rect 7261 3504 7267 4516
rect 7277 4304 7283 4576
rect 7293 4484 7299 4496
rect 7309 4384 7315 4516
rect 7309 4304 7315 4316
rect 7277 3584 7283 3636
rect 7261 3464 7267 3476
rect 7213 3444 7219 3456
rect 7197 3184 7203 3396
rect 7213 3384 7219 3436
rect 7245 3343 7251 3436
rect 7245 3337 7267 3343
rect 7261 3324 7267 3337
rect 7165 2984 7171 3036
rect 7197 2983 7203 3176
rect 7188 2977 7203 2983
rect 7053 2584 7059 2856
rect 6797 2264 6803 2296
rect 6829 2184 6835 2216
rect 6845 2164 6851 2256
rect 6733 2124 6739 2136
rect 6701 2104 6707 2116
rect 6541 1877 6556 1883
rect 6301 1784 6307 1856
rect 6173 1524 6179 1656
rect 6173 1504 6179 1516
rect 6157 1424 6163 1476
rect 6157 1384 6163 1396
rect 6189 1384 6195 1736
rect 6221 1624 6227 1696
rect 6285 1664 6291 1756
rect 6317 1724 6323 1836
rect 6365 1724 6371 1776
rect 6205 1584 6211 1596
rect 6301 1488 6307 1616
rect 6461 1564 6467 1836
rect 6493 1764 6499 1836
rect 6509 1804 6515 1856
rect 6525 1644 6531 1736
rect 6541 1724 6547 1836
rect 6621 1744 6627 1776
rect 6653 1764 6659 1836
rect 6701 1804 6707 2096
rect 6717 2064 6723 2116
rect 6749 2104 6755 2116
rect 6765 2024 6771 2096
rect 6765 1924 6771 2016
rect 6717 1904 6723 1916
rect 6765 1884 6771 1896
rect 6797 1884 6803 1936
rect 6845 1884 6851 2136
rect 6877 2124 6883 2196
rect 6909 2144 6915 2476
rect 6957 2304 6963 2536
rect 7021 2524 7027 2576
rect 7069 2564 7075 2636
rect 7085 2604 7091 2876
rect 7101 2704 7107 2736
rect 7101 2584 7107 2616
rect 7037 2524 7043 2556
rect 7085 2504 7091 2556
rect 7117 2544 7123 2576
rect 7021 2484 7027 2496
rect 7133 2484 7139 2516
rect 7149 2344 7155 2956
rect 7213 2943 7219 2996
rect 7197 2937 7219 2943
rect 7165 2824 7171 2836
rect 7181 2584 7187 2636
rect 7197 2523 7203 2937
rect 7229 2924 7235 2936
rect 7245 2924 7251 3016
rect 7213 2884 7219 2916
rect 7220 2877 7228 2883
rect 7213 2544 7219 2796
rect 7229 2524 7235 2596
rect 7245 2524 7251 2916
rect 7197 2517 7219 2523
rect 6957 2284 6963 2296
rect 7005 2244 7011 2294
rect 7133 2284 7139 2296
rect 6957 2177 6972 2183
rect 6957 2144 6963 2177
rect 7133 2144 7139 2276
rect 7165 2144 7171 2156
rect 6957 2124 6963 2136
rect 7069 2124 7075 2136
rect 6877 2104 6883 2116
rect 6781 1784 6787 1796
rect 6797 1784 6803 1856
rect 6925 1764 6931 1876
rect 6557 1684 6563 1696
rect 6285 1480 6300 1483
rect 6285 1477 6307 1480
rect 6205 1404 6211 1436
rect 6221 1384 6227 1416
rect 6157 1164 6163 1296
rect 6205 1184 6211 1256
rect 6237 1124 6243 1436
rect 6285 1364 6291 1477
rect 6333 1464 6339 1476
rect 6333 1384 6339 1456
rect 6349 1364 6355 1556
rect 6365 1524 6371 1536
rect 6381 1464 6387 1476
rect 6397 1444 6403 1496
rect 6477 1464 6483 1476
rect 6253 1204 6259 1316
rect 6365 1303 6371 1436
rect 6445 1364 6451 1396
rect 6477 1344 6483 1456
rect 6365 1297 6380 1303
rect 6397 1284 6403 1316
rect 6269 1163 6275 1236
rect 6253 1157 6275 1163
rect 6253 1104 6259 1157
rect 6093 1024 6099 1076
rect 6109 1023 6115 1094
rect 6109 1017 6131 1023
rect 6125 984 6131 1017
rect 6061 904 6067 916
rect 6013 704 6019 716
rect 6045 704 6051 836
rect 6077 784 6083 916
rect 6109 903 6115 936
rect 6173 924 6179 1096
rect 6221 1084 6227 1096
rect 6285 1084 6291 1236
rect 6205 944 6211 1076
rect 6221 984 6227 1076
rect 6237 1064 6243 1076
rect 6301 1063 6307 1096
rect 6397 1084 6403 1256
rect 6429 1124 6435 1296
rect 6477 1184 6483 1216
rect 6429 1084 6435 1116
rect 6285 1057 6307 1063
rect 6189 904 6195 916
rect 6093 897 6115 903
rect 6093 784 6099 897
rect 6157 884 6163 896
rect 6061 737 6076 743
rect 5946 614 5958 616
rect 5931 606 5933 614
rect 5941 606 5943 614
rect 5951 606 5953 614
rect 5961 606 5963 614
rect 5971 606 5973 614
rect 5946 604 5958 606
rect 5997 564 6003 596
rect 6029 584 6035 676
rect 5901 524 5907 556
rect 6061 524 6067 737
rect 6125 724 6131 776
rect 6077 697 6092 703
rect 6077 584 6083 697
rect 6109 703 6115 716
rect 6109 697 6131 703
rect 6125 644 6131 697
rect 5869 504 5875 516
rect 5876 477 5932 483
rect 5988 477 6012 483
rect 6029 463 6035 516
rect 6013 457 6035 463
rect 5981 304 5987 376
rect 6013 364 6019 457
rect 6045 324 6051 496
rect 6061 424 6067 456
rect 5805 184 5811 256
rect 5869 144 5875 176
rect 5517 97 5532 103
rect 5885 84 5891 236
rect 5901 224 5907 296
rect 5997 284 6003 316
rect 6029 284 6035 316
rect 6077 263 6083 556
rect 6109 544 6115 576
rect 6125 524 6131 636
rect 6141 564 6147 836
rect 6173 784 6179 816
rect 6205 704 6211 916
rect 6237 704 6243 1016
rect 6285 964 6291 1057
rect 6301 924 6307 1036
rect 6349 944 6355 1076
rect 6477 1064 6483 1096
rect 6493 1084 6499 1316
rect 6509 1303 6515 1436
rect 6525 1384 6531 1396
rect 6637 1384 6643 1494
rect 6669 1484 6675 1736
rect 6909 1724 6915 1756
rect 7005 1744 7011 1876
rect 7021 1864 7027 1916
rect 7037 1884 7043 2076
rect 7085 1884 7091 1936
rect 7117 1924 7123 2016
rect 7181 1944 7187 2516
rect 7213 2384 7219 2517
rect 7261 2503 7267 3296
rect 7277 3084 7283 3496
rect 7293 3304 7299 4076
rect 7309 3544 7315 4036
rect 7341 3584 7347 4216
rect 7389 3884 7395 5216
rect 7389 3744 7395 3876
rect 7357 3484 7363 3496
rect 7389 3464 7395 3516
rect 7293 3104 7299 3116
rect 7277 2584 7283 2936
rect 7293 2684 7299 3076
rect 7325 2804 7331 2916
rect 7277 2544 7283 2576
rect 7245 2497 7267 2503
rect 7245 2483 7251 2497
rect 7229 2477 7251 2483
rect 7197 2224 7203 2294
rect 7197 2104 7203 2176
rect 7197 2024 7203 2096
rect 7037 1724 7043 1876
rect 7117 1824 7123 1916
rect 7149 1884 7155 1896
rect 7181 1844 7187 1856
rect 7053 1724 7059 1736
rect 6861 1504 6867 1716
rect 7181 1704 7187 1816
rect 7213 1763 7219 2136
rect 7229 1784 7235 2477
rect 7261 2424 7267 2476
rect 7293 2344 7299 2436
rect 7309 2384 7315 2694
rect 7325 2524 7331 2536
rect 7261 2284 7267 2336
rect 7325 2324 7331 2496
rect 7277 2317 7292 2323
rect 7245 2184 7251 2236
rect 7261 2144 7267 2216
rect 7277 2184 7283 2317
rect 7293 2224 7299 2236
rect 7261 1884 7267 1896
rect 7213 1757 7235 1763
rect 7181 1684 7187 1696
rect 7005 1504 7011 1516
rect 7037 1504 7043 1516
rect 6749 1437 6764 1443
rect 6541 1344 6547 1376
rect 6541 1304 6547 1316
rect 6509 1297 6524 1303
rect 6381 1003 6387 1056
rect 6381 997 6403 1003
rect 6397 984 6403 997
rect 6381 964 6387 976
rect 6397 944 6403 976
rect 6429 924 6435 1036
rect 6461 924 6467 1016
rect 6493 984 6499 1076
rect 6509 984 6515 1276
rect 6605 1184 6611 1256
rect 6621 1204 6627 1356
rect 6653 1344 6659 1376
rect 6669 1344 6675 1396
rect 6669 1264 6675 1316
rect 6685 1304 6691 1316
rect 6685 1243 6691 1296
rect 6669 1237 6691 1243
rect 6557 1143 6563 1176
rect 6541 1137 6563 1143
rect 6525 1064 6531 1136
rect 6541 1104 6547 1137
rect 6557 1084 6563 1116
rect 6589 1084 6595 1136
rect 6605 1104 6611 1156
rect 6637 1124 6643 1136
rect 6605 1024 6611 1096
rect 6653 944 6659 956
rect 6621 924 6627 936
rect 6301 864 6307 896
rect 6317 844 6323 916
rect 6285 704 6291 716
rect 6381 704 6387 916
rect 6525 904 6531 918
rect 6637 884 6643 916
rect 6669 864 6675 1237
rect 6701 1104 6707 1296
rect 6733 1264 6739 1336
rect 6749 1324 6755 1437
rect 6788 1437 6803 1443
rect 6765 1363 6771 1436
rect 6797 1364 6803 1437
rect 6765 1357 6780 1363
rect 6797 1324 6803 1356
rect 6749 1184 6755 1316
rect 6765 1104 6771 1296
rect 6781 1144 6787 1276
rect 6781 1084 6787 1136
rect 6813 1084 6819 1236
rect 6861 1184 6867 1456
rect 6909 1424 6915 1494
rect 7069 1464 7075 1476
rect 6973 1444 6979 1456
rect 6957 1324 6963 1396
rect 6989 1384 6995 1416
rect 6877 1304 6883 1316
rect 6925 1284 6931 1296
rect 6829 1124 6835 1156
rect 6813 1064 6819 1076
rect 6461 684 6467 736
rect 6509 684 6515 696
rect 6157 524 6163 676
rect 6269 564 6275 656
rect 6237 544 6243 556
rect 6093 284 6099 496
rect 6125 343 6131 436
rect 6157 384 6163 496
rect 6173 444 6179 496
rect 6125 337 6147 343
rect 6141 304 6147 337
rect 6173 324 6179 436
rect 6221 424 6227 516
rect 6077 257 6099 263
rect 5901 184 5907 216
rect 5946 214 5958 216
rect 5931 206 5933 214
rect 5941 206 5943 214
rect 5951 206 5953 214
rect 5961 206 5963 214
rect 5971 206 5973 214
rect 5946 204 5958 206
rect 5997 204 6003 256
rect 5965 144 5971 156
rect 5933 104 5939 118
rect 6013 104 6019 236
rect 6077 104 6083 236
rect 6093 124 6099 257
rect 6109 244 6115 296
rect 6205 284 6211 376
rect 6285 364 6291 556
rect 6253 304 6259 356
rect 6109 124 6115 216
rect 6125 204 6131 276
rect 6189 177 6204 183
rect 6157 164 6163 176
rect 6189 163 6195 177
rect 6301 164 6307 656
rect 6333 524 6339 676
rect 6381 664 6387 676
rect 6429 604 6435 636
rect 6493 624 6499 676
rect 6525 663 6531 696
rect 6541 684 6547 716
rect 6605 704 6611 856
rect 6509 657 6531 663
rect 6477 524 6483 536
rect 6317 384 6323 496
rect 6381 484 6387 516
rect 6493 504 6499 616
rect 6365 384 6371 436
rect 6493 364 6499 436
rect 6509 384 6515 657
rect 6573 604 6579 656
rect 6589 644 6595 676
rect 6589 564 6595 636
rect 6541 544 6547 556
rect 6317 304 6323 356
rect 6349 284 6355 316
rect 6413 304 6419 356
rect 6493 324 6499 356
rect 6525 344 6531 376
rect 6381 284 6387 296
rect 6397 184 6403 236
rect 6429 164 6435 216
rect 6173 157 6195 163
rect 6173 84 6179 157
rect 6301 144 6307 156
rect 6189 104 6195 136
rect 6205 84 6211 116
rect 6269 104 6275 118
rect 6461 84 6467 256
rect 6493 104 6499 316
rect 6509 184 6515 196
rect 6541 164 6547 536
rect 6605 524 6611 696
rect 6653 584 6659 616
rect 6685 604 6691 956
rect 6717 924 6723 1016
rect 6740 937 6755 943
rect 6701 704 6707 716
rect 6717 684 6723 756
rect 6621 544 6627 576
rect 6653 544 6659 576
rect 6685 564 6691 596
rect 6717 564 6723 676
rect 6749 644 6755 937
rect 6781 904 6787 1036
rect 6877 944 6883 996
rect 6829 924 6835 936
rect 6877 904 6883 916
rect 6765 864 6771 876
rect 6813 784 6819 856
rect 6829 704 6835 896
rect 6845 884 6851 896
rect 6877 864 6883 896
rect 6893 724 6899 1116
rect 6909 943 6915 1256
rect 6941 1084 6947 1096
rect 6941 963 6947 1076
rect 6957 1044 6963 1316
rect 7005 1304 7011 1436
rect 7021 1264 7027 1296
rect 7005 1104 7011 1116
rect 6957 983 6963 1016
rect 6973 1004 6979 1096
rect 6989 1024 6995 1076
rect 7037 1024 7043 1276
rect 6957 977 6972 983
rect 6941 957 6956 963
rect 6989 944 6995 976
rect 7053 963 7059 1436
rect 7085 1404 7091 1496
rect 7117 1403 7123 1436
rect 7101 1397 7123 1403
rect 7101 1324 7107 1397
rect 7133 1324 7139 1676
rect 7165 1624 7171 1636
rect 7213 1624 7219 1736
rect 7229 1724 7235 1757
rect 7181 1524 7187 1556
rect 7245 1524 7251 1776
rect 7261 1744 7267 1856
rect 7293 1784 7299 2196
rect 7309 2164 7315 2256
rect 7309 2083 7315 2156
rect 7325 2124 7331 2216
rect 7341 2124 7347 2916
rect 7389 2543 7395 2956
rect 7405 2884 7411 2896
rect 7389 2537 7411 2543
rect 7357 2304 7363 2336
rect 7373 2284 7379 2516
rect 7309 2077 7331 2083
rect 7325 1844 7331 2077
rect 7325 1764 7331 1836
rect 7357 1743 7363 2276
rect 7389 2143 7395 2516
rect 7380 2137 7395 2143
rect 7373 2084 7379 2136
rect 7405 2104 7411 2537
rect 7341 1737 7363 1743
rect 7293 1724 7299 1736
rect 7069 1244 7075 1316
rect 7069 1104 7075 1236
rect 7133 1084 7139 1316
rect 7053 957 7075 963
rect 7069 944 7075 957
rect 6909 937 6924 943
rect 6909 784 6915 937
rect 6989 904 6995 916
rect 6717 524 6723 536
rect 6653 504 6659 516
rect 6573 363 6579 436
rect 6669 424 6675 516
rect 6733 444 6739 516
rect 6749 424 6755 436
rect 6557 357 6579 363
rect 6557 284 6563 357
rect 6573 304 6579 336
rect 6589 264 6595 276
rect 6621 244 6627 256
rect 6653 244 6659 276
rect 6701 244 6707 316
rect 6605 144 6611 156
rect 6669 124 6675 236
rect 6717 224 6723 296
rect 6749 224 6755 416
rect 6765 364 6771 556
rect 6781 484 6787 656
rect 6877 644 6883 656
rect 6909 544 6915 756
rect 6925 664 6931 696
rect 6957 564 6963 716
rect 6973 684 6979 796
rect 6989 704 6995 896
rect 6973 644 6979 656
rect 6861 524 6867 536
rect 6957 464 6963 536
rect 6989 524 6995 696
rect 7037 684 7043 936
rect 7053 924 7059 936
rect 7069 924 7075 936
rect 7085 924 7091 1016
rect 7069 784 7075 916
rect 7101 764 7107 1076
rect 7149 1003 7155 1436
rect 7165 1404 7171 1476
rect 7245 1464 7251 1496
rect 7261 1384 7267 1716
rect 7277 1684 7283 1716
rect 7277 1524 7283 1556
rect 7325 1524 7331 1536
rect 7309 1444 7315 1456
rect 7133 997 7155 1003
rect 7133 964 7139 997
rect 7165 983 7171 1096
rect 7156 977 7171 983
rect 7037 664 7043 676
rect 7005 584 7011 656
rect 7053 604 7059 736
rect 7117 724 7123 896
rect 7133 744 7139 956
rect 7165 944 7171 956
rect 7149 722 7155 916
rect 7005 544 7011 576
rect 7053 564 7059 596
rect 7005 444 7011 516
rect 7021 484 7027 536
rect 7069 484 7075 696
rect 7117 664 7123 696
rect 7085 584 7091 656
rect 7133 623 7139 716
rect 7117 617 7139 623
rect 6781 384 6787 436
rect 6765 324 6771 356
rect 6781 324 6787 336
rect 6765 184 6771 316
rect 6781 304 6787 316
rect 6829 304 6835 316
rect 6877 304 6883 376
rect 6701 164 6707 176
rect 6797 164 6803 216
rect 6733 144 6739 156
rect 6781 144 6787 156
rect 6829 144 6835 296
rect 6925 284 6931 296
rect 6637 104 6643 118
rect 6749 84 6755 116
rect 6893 104 6899 176
rect 6973 144 6979 196
rect 6989 184 6995 296
rect 7005 284 7011 436
rect 7021 384 7027 396
rect 7037 264 7043 276
rect 7053 204 7059 316
rect 7069 284 7075 296
rect 7085 284 7091 576
rect 7101 484 7107 516
rect 7117 504 7123 617
rect 7133 524 7139 536
rect 7149 504 7155 656
rect 7181 544 7187 1376
rect 7277 1144 7283 1416
rect 7293 1344 7299 1396
rect 7309 1323 7315 1356
rect 7293 1317 7315 1323
rect 7277 1064 7283 1136
rect 7229 944 7235 1056
rect 7245 964 7251 996
rect 7245 944 7251 956
rect 7261 944 7267 976
rect 7277 940 7283 1036
rect 7204 917 7219 923
rect 7197 884 7203 896
rect 7213 784 7219 917
rect 7229 904 7235 916
rect 7213 704 7219 716
rect 7117 304 7123 476
rect 7133 464 7139 476
rect 7165 304 7171 316
rect 7197 284 7203 636
rect 7245 524 7251 756
rect 7261 584 7267 676
rect 7277 664 7283 696
rect 7293 644 7299 1317
rect 7309 1164 7315 1296
rect 7325 1124 7331 1436
rect 7341 1364 7347 1737
rect 7373 1324 7379 1716
rect 7357 964 7363 1056
rect 7341 664 7347 936
rect 7357 784 7363 956
rect 7373 664 7379 776
rect 7069 184 7075 276
rect 7021 140 7027 176
rect 7085 124 7091 276
rect 7133 184 7139 276
rect 7213 203 7219 236
rect 7213 197 7235 203
rect 7117 164 7123 176
rect 7229 126 7235 197
rect 7245 144 7251 516
rect 7341 384 7347 636
rect 7293 304 7299 316
rect 7053 104 7059 116
rect 7101 84 7107 116
rect 7261 104 7267 256
rect 7357 144 7363 176
rect 7389 164 7395 1636
rect 6909 64 6915 76
rect 4845 -17 4851 36
rect 4845 -23 4867 -17
rect 4989 -23 4995 16
rect 5053 -17 5059 36
rect 5037 -23 5059 -17
rect 5069 -17 5075 36
rect 5245 -17 5251 36
rect 5357 -17 5363 36
rect 5405 -17 5411 36
rect 5581 -17 5587 36
rect 5629 -17 5635 36
rect 5069 -23 5091 -17
rect 5229 -23 5251 -17
rect 5341 -23 5363 -17
rect 5389 -23 5411 -17
rect 5565 -23 5587 -17
rect 5613 -23 5635 -17
rect 5709 -17 5715 36
rect 5757 -17 5763 36
rect 6061 -17 6067 36
rect 6141 -17 6147 36
rect 5709 -23 5731 -17
rect 5757 -23 5779 -17
rect 6061 -23 6083 -17
rect 6125 -23 6147 -17
rect 6413 -23 6419 16
<< m3contact >>
rect 2915 5406 2923 5414
rect 2925 5406 2933 5414
rect 2935 5406 2943 5414
rect 2945 5406 2953 5414
rect 2955 5406 2963 5414
rect 2965 5406 2973 5414
rect 620 5376 628 5384
rect 796 5376 804 5384
rect 1404 5376 1412 5384
rect 1548 5376 1556 5384
rect 524 5356 532 5364
rect 12 5336 20 5344
rect 140 5336 148 5344
rect 172 5336 180 5344
rect 252 5336 260 5344
rect 332 5336 340 5344
rect 172 5316 180 5324
rect 60 5296 68 5304
rect 156 5296 164 5304
rect 124 5256 132 5264
rect 236 5296 244 5304
rect 220 5276 228 5284
rect 284 5316 292 5324
rect 332 5316 340 5324
rect 524 5336 532 5344
rect 604 5336 612 5344
rect 316 5276 324 5284
rect 204 5236 212 5244
rect 268 5236 276 5244
rect 92 5216 100 5224
rect 140 5176 148 5184
rect 316 5156 324 5164
rect 508 5316 516 5324
rect 460 5216 468 5224
rect 476 5216 484 5224
rect 124 5136 132 5144
rect 220 5136 228 5144
rect 380 5136 388 5144
rect 108 5116 116 5124
rect 156 5116 164 5124
rect 316 5116 324 5124
rect 380 5116 388 5124
rect 28 5056 36 5064
rect 44 5016 52 5024
rect 172 5076 180 5084
rect 268 5076 276 5084
rect 204 5056 212 5064
rect 76 4956 84 4964
rect 124 4956 132 4964
rect 44 4936 52 4944
rect 12 4896 20 4904
rect 12 4556 20 4564
rect 12 4316 20 4324
rect 252 5056 260 5064
rect 236 5016 244 5024
rect 140 4936 148 4944
rect 124 4916 132 4924
rect 156 4916 164 4924
rect 76 4736 84 4744
rect 156 4696 164 4704
rect 204 4696 212 4704
rect 92 4676 100 4684
rect 332 5076 340 5084
rect 268 4916 276 4924
rect 252 4816 260 4824
rect 492 5196 500 5204
rect 444 5096 452 5104
rect 476 5076 484 5084
rect 348 5056 356 5064
rect 460 5056 468 5064
rect 508 5096 516 5104
rect 348 4996 356 5004
rect 460 4996 468 5004
rect 380 4956 388 4964
rect 508 4956 516 4964
rect 316 4936 324 4944
rect 364 4936 372 4944
rect 412 4936 420 4944
rect 444 4936 452 4944
rect 492 4936 500 4944
rect 300 4796 308 4804
rect 300 4696 308 4704
rect 364 4696 372 4704
rect 204 4676 212 4684
rect 236 4676 244 4684
rect 44 4556 52 4564
rect 428 4896 436 4904
rect 460 4896 468 4904
rect 988 5356 996 5364
rect 668 5336 676 5344
rect 636 5316 644 5324
rect 700 5316 708 5324
rect 588 5296 596 5304
rect 652 5296 660 5304
rect 668 5296 676 5304
rect 588 5276 596 5284
rect 636 5276 644 5284
rect 636 5176 644 5184
rect 540 4956 548 4964
rect 524 4936 532 4944
rect 412 4696 420 4704
rect 428 4696 436 4704
rect 268 4676 276 4684
rect 348 4680 356 4684
rect 348 4676 356 4680
rect 380 4676 388 4684
rect 252 4576 260 4584
rect 220 4556 228 4564
rect 332 4556 340 4564
rect 380 4556 388 4564
rect 76 4536 84 4544
rect 124 4536 132 4544
rect 396 4516 404 4524
rect 444 4676 452 4684
rect 604 5096 612 5104
rect 620 5076 628 5084
rect 572 5056 580 5064
rect 796 5336 804 5344
rect 876 5336 884 5344
rect 956 5336 964 5344
rect 764 5316 772 5324
rect 732 5276 740 5284
rect 748 5276 756 5284
rect 716 5256 724 5264
rect 956 5316 964 5324
rect 876 5296 884 5304
rect 908 5296 916 5304
rect 956 5236 964 5244
rect 876 5216 884 5224
rect 892 5216 900 5224
rect 844 5176 852 5184
rect 684 5156 692 5164
rect 748 5156 756 5164
rect 668 5116 676 5124
rect 716 5096 724 5104
rect 684 5076 692 5084
rect 732 5076 740 5084
rect 652 5036 660 5044
rect 844 5136 852 5144
rect 780 5116 788 5124
rect 812 5116 820 5124
rect 924 5116 932 5124
rect 796 5096 804 5104
rect 892 5096 900 5104
rect 812 5076 820 5084
rect 572 4976 580 4984
rect 604 4976 612 4984
rect 636 4976 644 4984
rect 748 4976 756 4984
rect 764 4976 772 4984
rect 588 4956 596 4964
rect 668 4936 676 4944
rect 636 4916 644 4924
rect 556 4896 564 4904
rect 588 4896 596 4904
rect 652 4896 660 4904
rect 588 4756 596 4764
rect 556 4696 564 4704
rect 572 4696 580 4704
rect 540 4676 548 4684
rect 524 4656 532 4664
rect 556 4656 564 4664
rect 508 4636 516 4644
rect 476 4556 484 4564
rect 684 4836 692 4844
rect 716 4916 724 4924
rect 876 5076 884 5084
rect 844 5056 852 5064
rect 940 5076 948 5084
rect 892 5056 900 5064
rect 876 5016 884 5024
rect 860 4996 868 5004
rect 780 4916 788 4924
rect 732 4896 740 4904
rect 780 4896 788 4904
rect 700 4736 708 4744
rect 620 4676 628 4684
rect 652 4636 660 4644
rect 588 4616 596 4624
rect 588 4556 596 4564
rect 124 4496 132 4504
rect 188 4496 196 4504
rect 76 4316 84 4324
rect 92 4316 100 4324
rect 284 4496 292 4504
rect 348 4496 356 4504
rect 252 4436 260 4444
rect 316 4356 324 4364
rect 348 4316 356 4324
rect 76 4296 84 4304
rect 108 4296 116 4304
rect 60 4256 68 4264
rect 12 4156 20 4164
rect 12 4116 20 4124
rect 332 4296 340 4304
rect 92 4276 100 4284
rect 316 4276 324 4284
rect 508 4516 516 4524
rect 636 4516 644 4524
rect 444 4356 452 4364
rect 428 4336 436 4344
rect 396 4296 404 4304
rect 156 4256 164 4264
rect 204 4256 212 4264
rect 396 4256 404 4264
rect 428 4256 436 4264
rect 108 4176 116 4184
rect 188 4176 196 4184
rect 348 4236 356 4244
rect 460 4236 468 4244
rect 124 4156 132 4164
rect 108 4136 116 4144
rect 172 4136 180 4144
rect 204 4156 212 4164
rect 284 4156 292 4164
rect 76 4116 84 4124
rect 236 4116 244 4124
rect 316 4116 324 4124
rect 268 4096 276 4104
rect 460 4156 468 4164
rect 412 4116 420 4124
rect 476 4116 484 4124
rect 364 4096 372 4104
rect 76 4076 84 4084
rect 284 4076 292 4084
rect 332 4076 340 4084
rect 60 3916 68 3924
rect 108 3916 116 3924
rect 124 3916 132 3924
rect 156 3896 164 3904
rect 12 3876 20 3884
rect 172 3876 180 3884
rect 236 4016 244 4024
rect 220 3896 228 3904
rect 300 3896 308 3904
rect 268 3876 276 3884
rect 300 3876 308 3884
rect 348 3876 356 3884
rect 268 3856 276 3864
rect 316 3856 324 3864
rect 332 3856 340 3864
rect 188 3776 196 3784
rect 524 4356 532 4364
rect 636 4356 644 4364
rect 556 4296 564 4304
rect 620 4296 628 4304
rect 684 4636 692 4644
rect 700 4636 708 4644
rect 780 4696 788 4704
rect 764 4676 772 4684
rect 732 4656 740 4664
rect 732 4636 740 4644
rect 716 4616 724 4624
rect 716 4556 724 4564
rect 684 4516 692 4524
rect 828 4936 836 4944
rect 812 4896 820 4904
rect 860 4896 868 4904
rect 924 4996 932 5004
rect 972 5076 980 5084
rect 1068 5296 1076 5304
rect 1004 5276 1012 5284
rect 1148 5336 1156 5344
rect 1116 5316 1124 5324
rect 1132 5236 1140 5244
rect 1100 5176 1108 5184
rect 1196 5316 1204 5324
rect 1196 5276 1204 5284
rect 1532 5356 1540 5364
rect 1628 5356 1636 5364
rect 2012 5356 2020 5364
rect 2204 5356 2212 5364
rect 2316 5356 2324 5364
rect 2508 5356 2516 5364
rect 1596 5336 1604 5344
rect 1932 5336 1940 5344
rect 1436 5316 1444 5324
rect 1196 5256 1204 5264
rect 1212 5256 1220 5264
rect 1148 5156 1156 5164
rect 1004 5136 1012 5144
rect 1036 5116 1044 5124
rect 1068 5116 1076 5124
rect 1132 5116 1140 5124
rect 1036 5096 1044 5104
rect 1148 5096 1156 5104
rect 1052 5076 1060 5084
rect 1116 5076 1124 5084
rect 1148 5076 1156 5084
rect 1020 5056 1028 5064
rect 956 4916 964 4924
rect 908 4876 916 4884
rect 892 4836 900 4844
rect 908 4736 916 4744
rect 828 4676 836 4684
rect 828 4616 836 4624
rect 812 4576 820 4584
rect 924 4656 932 4664
rect 892 4636 900 4644
rect 876 4576 884 4584
rect 812 4556 820 4564
rect 844 4556 852 4564
rect 860 4516 868 4524
rect 700 4476 708 4484
rect 748 4476 756 4484
rect 652 4336 660 4344
rect 684 4296 692 4304
rect 732 4296 740 4304
rect 524 4256 532 4264
rect 668 4236 676 4244
rect 668 4196 676 4204
rect 572 4156 580 4164
rect 540 4136 548 4144
rect 412 3916 420 3924
rect 476 3976 484 3984
rect 460 3936 468 3944
rect 476 3936 484 3944
rect 380 3896 388 3904
rect 380 3856 388 3864
rect 396 3856 404 3864
rect 364 3776 372 3784
rect 60 3756 68 3764
rect 124 3756 132 3764
rect 172 3756 180 3764
rect 188 3756 196 3764
rect 220 3756 228 3764
rect 300 3756 308 3764
rect 364 3756 372 3764
rect 396 3756 404 3764
rect 460 3916 468 3924
rect 444 3896 452 3904
rect 444 3876 452 3884
rect 460 3856 468 3864
rect 12 3716 20 3724
rect 108 3716 116 3724
rect 140 3696 148 3704
rect 60 3536 68 3544
rect 76 3496 84 3504
rect 60 3476 68 3484
rect 380 3736 388 3744
rect 284 3716 292 3724
rect 348 3716 356 3724
rect 428 3716 436 3724
rect 188 3696 196 3704
rect 220 3696 228 3704
rect 236 3616 244 3624
rect 172 3596 180 3604
rect 316 3696 324 3704
rect 364 3696 372 3704
rect 316 3596 324 3604
rect 300 3576 308 3584
rect 236 3556 244 3564
rect 268 3536 276 3544
rect 108 3516 116 3524
rect 156 3516 164 3524
rect 236 3496 244 3504
rect 108 3456 116 3464
rect 140 3456 148 3464
rect 12 3396 20 3404
rect 28 3396 36 3404
rect 44 3396 52 3404
rect 92 3396 100 3404
rect 12 3356 20 3364
rect 28 3216 36 3224
rect 92 3376 100 3384
rect 124 3376 132 3384
rect 76 3336 84 3344
rect 12 3096 20 3104
rect 28 2916 36 2924
rect 76 3216 84 3224
rect 76 3076 84 3084
rect 76 2936 84 2944
rect 204 3356 212 3364
rect 140 3336 148 3344
rect 252 3376 260 3384
rect 332 3496 340 3504
rect 316 3476 324 3484
rect 380 3616 388 3624
rect 412 3576 420 3584
rect 396 3496 404 3504
rect 444 3496 452 3504
rect 428 3476 436 3484
rect 316 3376 324 3384
rect 268 3336 276 3344
rect 156 3316 164 3324
rect 236 3316 244 3324
rect 124 3096 132 3104
rect 108 3076 116 3084
rect 204 3296 212 3304
rect 300 3296 308 3304
rect 412 3456 420 3464
rect 508 3936 516 3944
rect 636 4156 644 4164
rect 652 4136 660 4144
rect 700 4216 708 4224
rect 684 4136 692 4144
rect 748 4276 756 4284
rect 748 4196 756 4204
rect 748 4156 756 4164
rect 732 4136 740 4144
rect 748 4096 756 4104
rect 508 3916 516 3924
rect 540 3916 548 3924
rect 572 3916 580 3924
rect 492 3896 500 3904
rect 492 3856 500 3864
rect 492 3836 500 3844
rect 524 3876 532 3884
rect 556 3856 564 3864
rect 572 3856 580 3864
rect 604 3916 612 3924
rect 620 3896 628 3904
rect 636 3880 644 3884
rect 636 3876 644 3880
rect 780 4436 788 4444
rect 780 4336 788 4344
rect 796 4316 804 4324
rect 828 4316 836 4324
rect 860 4316 868 4324
rect 892 4556 900 4564
rect 988 4996 996 5004
rect 1020 4996 1028 5004
rect 1036 4996 1044 5004
rect 988 4936 996 4944
rect 988 4916 996 4924
rect 972 4856 980 4864
rect 1068 5036 1076 5044
rect 1052 4976 1060 4984
rect 1036 4956 1044 4964
rect 1052 4936 1060 4944
rect 1100 5036 1108 5044
rect 1244 5216 1252 5224
rect 1212 5136 1220 5144
rect 1196 5096 1204 5104
rect 1228 5116 1236 5124
rect 1276 5296 1284 5304
rect 1580 5296 1588 5304
rect 1580 5256 1588 5264
rect 1276 5216 1284 5224
rect 1564 5216 1572 5224
rect 1411 5206 1419 5214
rect 1421 5206 1429 5214
rect 1431 5206 1439 5214
rect 1441 5206 1449 5214
rect 1451 5206 1459 5214
rect 1461 5206 1469 5214
rect 1388 5196 1396 5204
rect 1276 5176 1284 5184
rect 1308 5156 1316 5164
rect 1260 5116 1268 5124
rect 1340 5136 1348 5144
rect 1324 5096 1332 5104
rect 1356 5056 1364 5064
rect 1388 5036 1396 5044
rect 1148 4976 1156 4984
rect 1164 4976 1172 4984
rect 1276 4956 1284 4964
rect 1100 4936 1108 4944
rect 1084 4916 1092 4924
rect 1116 4916 1124 4924
rect 1036 4896 1044 4904
rect 1068 4896 1076 4904
rect 988 4836 996 4844
rect 1020 4836 1028 4844
rect 972 4656 980 4664
rect 956 4616 964 4624
rect 1164 4876 1172 4884
rect 1196 4876 1204 4884
rect 1212 4856 1220 4864
rect 1068 4756 1076 4764
rect 1164 4736 1172 4744
rect 1116 4696 1124 4704
rect 1004 4676 1012 4684
rect 1020 4656 1028 4664
rect 1036 4656 1044 4664
rect 1084 4636 1092 4644
rect 988 4596 996 4604
rect 1068 4596 1076 4604
rect 956 4576 964 4584
rect 940 4556 948 4564
rect 1052 4556 1060 4564
rect 972 4536 980 4544
rect 924 4516 932 4524
rect 956 4516 964 4524
rect 988 4516 996 4524
rect 1036 4476 1044 4484
rect 892 4356 900 4364
rect 924 4356 932 4364
rect 940 4336 948 4344
rect 828 4296 836 4304
rect 876 4276 884 4284
rect 796 4256 804 4264
rect 860 4236 868 4244
rect 812 4156 820 4164
rect 764 3956 772 3964
rect 684 3916 692 3924
rect 668 3876 676 3884
rect 764 3896 772 3904
rect 700 3876 708 3884
rect 764 3856 772 3864
rect 700 3836 708 3844
rect 652 3796 660 3804
rect 620 3776 628 3784
rect 668 3776 676 3784
rect 1084 4576 1092 4584
rect 1116 4556 1124 4564
rect 1148 4556 1156 4564
rect 1228 4816 1236 4824
rect 1196 4716 1204 4724
rect 1180 4696 1188 4704
rect 1212 4676 1220 4684
rect 1212 4636 1220 4644
rect 1164 4536 1172 4544
rect 1068 4496 1076 4504
rect 1068 4476 1076 4484
rect 1372 4896 1380 4904
rect 1356 4876 1364 4884
rect 1308 4796 1316 4804
rect 1356 4736 1364 4744
rect 1420 5076 1428 5084
rect 1516 5136 1524 5144
rect 1660 5316 1668 5324
rect 1644 5296 1652 5304
rect 1964 5316 1972 5324
rect 2060 5276 2068 5284
rect 1804 5256 1812 5264
rect 1836 5236 1844 5244
rect 1612 5216 1620 5224
rect 1820 5156 1828 5164
rect 1708 5116 1716 5124
rect 1692 5096 1700 5104
rect 1724 5096 1732 5104
rect 1788 5096 1796 5104
rect 1820 5096 1828 5104
rect 1548 5076 1556 5084
rect 1596 5076 1604 5084
rect 1660 5076 1668 5084
rect 1596 5056 1604 5064
rect 1436 5036 1444 5044
rect 1612 5016 1620 5024
rect 1644 5016 1652 5024
rect 1548 4976 1556 4984
rect 1484 4956 1492 4964
rect 1468 4936 1476 4944
rect 1532 4936 1540 4944
rect 1516 4916 1524 4924
rect 1596 4936 1604 4944
rect 1580 4916 1588 4924
rect 1564 4856 1572 4864
rect 1484 4816 1492 4824
rect 1411 4806 1419 4814
rect 1421 4806 1429 4814
rect 1431 4806 1439 4814
rect 1441 4806 1449 4814
rect 1451 4806 1459 4814
rect 1461 4806 1469 4814
rect 1596 4836 1604 4844
rect 1580 4796 1588 4804
rect 1532 4716 1540 4724
rect 1372 4696 1380 4704
rect 1388 4696 1396 4704
rect 1580 4696 1588 4704
rect 1596 4676 1604 4684
rect 1644 4956 1652 4964
rect 1676 5036 1684 5044
rect 1756 5076 1764 5084
rect 1708 5056 1716 5064
rect 1708 5016 1716 5024
rect 1708 4976 1716 4984
rect 1692 4956 1700 4964
rect 1660 4936 1668 4944
rect 1628 4916 1636 4924
rect 1660 4916 1668 4924
rect 1628 4876 1636 4884
rect 1628 4836 1636 4844
rect 1660 4796 1668 4804
rect 1260 4656 1268 4664
rect 1388 4636 1396 4644
rect 1212 4536 1220 4544
rect 1244 4536 1252 4544
rect 1180 4476 1188 4484
rect 1148 4456 1156 4464
rect 1148 4436 1156 4444
rect 1276 4496 1284 4504
rect 1388 4616 1396 4624
rect 1356 4536 1364 4544
rect 1340 4516 1348 4524
rect 1452 4576 1460 4584
rect 1484 4556 1492 4564
rect 1468 4516 1476 4524
rect 1500 4516 1508 4524
rect 1420 4496 1428 4504
rect 1676 4736 1684 4744
rect 1740 4976 1748 4984
rect 1948 5176 1956 5184
rect 1900 5156 1908 5164
rect 1788 5016 1796 5024
rect 1772 4956 1780 4964
rect 1884 5036 1892 5044
rect 1820 5016 1828 5024
rect 1740 4916 1748 4924
rect 1756 4916 1764 4924
rect 1804 4916 1812 4924
rect 2268 5336 2276 5344
rect 2444 5336 2452 5344
rect 2572 5336 2580 5344
rect 2668 5336 2676 5344
rect 2748 5336 2756 5344
rect 2876 5336 2884 5344
rect 2892 5336 2900 5344
rect 2172 5316 2180 5324
rect 2220 5316 2228 5324
rect 2476 5316 2484 5324
rect 2524 5316 2532 5324
rect 2572 5316 2580 5324
rect 2716 5316 2724 5324
rect 2780 5316 2788 5324
rect 2140 5236 2148 5244
rect 2348 5296 2356 5304
rect 2316 5216 2324 5224
rect 2236 5136 2244 5144
rect 2172 5116 2180 5124
rect 1964 5096 1972 5104
rect 1996 5096 2004 5104
rect 2076 5096 2084 5104
rect 2092 5096 2100 5104
rect 2012 5076 2020 5084
rect 1996 5056 2004 5064
rect 2028 5056 2036 5064
rect 1948 5036 1956 5044
rect 2012 5016 2020 5024
rect 1948 4976 1956 4984
rect 1996 4976 2004 4984
rect 1964 4956 1972 4964
rect 1932 4916 1940 4924
rect 1852 4896 1860 4904
rect 1900 4896 1908 4904
rect 1820 4876 1828 4884
rect 1724 4856 1732 4864
rect 1804 4856 1812 4864
rect 1772 4776 1780 4784
rect 1756 4736 1764 4744
rect 1740 4716 1748 4724
rect 1708 4696 1716 4704
rect 1804 4736 1812 4744
rect 1820 4716 1828 4724
rect 1884 4856 1892 4864
rect 1852 4716 1860 4724
rect 1836 4696 1844 4704
rect 1660 4676 1668 4684
rect 1772 4676 1780 4684
rect 1644 4656 1652 4664
rect 1548 4576 1556 4584
rect 1580 4556 1588 4564
rect 1644 4556 1652 4564
rect 1532 4536 1540 4544
rect 1340 4476 1348 4484
rect 1388 4476 1396 4484
rect 1516 4476 1524 4484
rect 1244 4456 1252 4464
rect 1372 4456 1380 4464
rect 1196 4356 1204 4364
rect 1084 4336 1092 4344
rect 1228 4316 1236 4324
rect 1100 4296 1108 4304
rect 1132 4296 1140 4304
rect 1116 4276 1124 4284
rect 1164 4276 1172 4284
rect 1020 4256 1028 4264
rect 972 4216 980 4224
rect 956 4196 964 4204
rect 908 4176 916 4184
rect 892 4156 900 4164
rect 812 3996 820 4004
rect 844 3996 852 4004
rect 924 4136 932 4144
rect 908 4116 916 4124
rect 940 4116 948 4124
rect 1052 4196 1060 4204
rect 1004 4156 1012 4164
rect 988 4136 996 4144
rect 1004 4116 1012 4124
rect 1036 4116 1044 4124
rect 1100 4176 1108 4184
rect 1148 4256 1156 4264
rect 1196 4256 1204 4264
rect 1308 4336 1316 4344
rect 1292 4316 1300 4324
rect 1260 4296 1268 4304
rect 1676 4536 1684 4544
rect 1596 4516 1604 4524
rect 1612 4516 1620 4524
rect 1644 4516 1652 4524
rect 1580 4496 1588 4504
rect 1564 4476 1572 4484
rect 1532 4456 1540 4464
rect 1411 4406 1419 4414
rect 1421 4406 1429 4414
rect 1431 4406 1439 4414
rect 1441 4406 1449 4414
rect 1451 4406 1459 4414
rect 1461 4406 1469 4414
rect 1404 4376 1412 4384
rect 1356 4256 1364 4264
rect 1388 4256 1396 4264
rect 1244 4236 1252 4244
rect 1324 4236 1332 4244
rect 1324 4216 1332 4224
rect 1212 4196 1220 4204
rect 1132 4156 1140 4164
rect 1228 4156 1236 4164
rect 1340 4156 1348 4164
rect 1148 4136 1156 4144
rect 1212 4136 1220 4144
rect 1068 4116 1076 4124
rect 1116 4116 1124 4124
rect 1084 4076 1092 4084
rect 1100 4016 1108 4024
rect 1020 3976 1028 3984
rect 1068 3976 1076 3984
rect 972 3936 980 3944
rect 828 3876 836 3884
rect 892 3876 900 3884
rect 620 3756 628 3764
rect 684 3756 692 3764
rect 716 3756 724 3764
rect 748 3756 756 3764
rect 604 3736 612 3744
rect 668 3736 676 3744
rect 812 3736 820 3744
rect 652 3716 660 3724
rect 828 3716 836 3724
rect 764 3696 772 3704
rect 588 3656 596 3664
rect 652 3656 660 3664
rect 508 3536 516 3544
rect 556 3536 564 3544
rect 476 3476 484 3484
rect 364 3156 372 3164
rect 428 3416 436 3424
rect 412 3376 420 3384
rect 380 3116 388 3124
rect 476 3456 484 3464
rect 444 3376 452 3384
rect 476 3376 484 3384
rect 444 3296 452 3304
rect 460 3296 468 3304
rect 460 3276 468 3284
rect 444 3116 452 3124
rect 156 3096 164 3104
rect 268 3096 276 3104
rect 316 3096 324 3104
rect 396 3096 404 3104
rect 476 3096 484 3104
rect 124 3056 132 3064
rect 332 3076 340 3084
rect 380 3076 388 3084
rect 156 3056 164 3064
rect 172 3056 180 3064
rect 316 3056 324 3064
rect 364 3056 372 3064
rect 460 3056 468 3064
rect 156 3036 164 3044
rect 92 2916 100 2924
rect 140 2936 148 2944
rect 220 2936 228 2944
rect 540 3436 548 3444
rect 604 3516 612 3524
rect 636 3516 644 3524
rect 588 3416 596 3424
rect 604 3396 612 3404
rect 716 3516 724 3524
rect 668 3496 676 3504
rect 748 3476 756 3484
rect 908 3816 916 3824
rect 1036 3916 1044 3924
rect 1068 3916 1076 3924
rect 1068 3876 1076 3884
rect 940 3776 948 3784
rect 972 3776 980 3784
rect 860 3756 868 3764
rect 876 3716 884 3724
rect 908 3716 916 3724
rect 892 3596 900 3604
rect 844 3576 852 3584
rect 892 3516 900 3524
rect 876 3496 884 3504
rect 828 3476 836 3484
rect 652 3356 660 3364
rect 716 3456 724 3464
rect 780 3456 788 3464
rect 796 3456 804 3464
rect 748 3416 756 3424
rect 780 3416 788 3424
rect 700 3396 708 3404
rect 684 3376 692 3384
rect 668 3316 676 3324
rect 524 3296 532 3304
rect 540 3276 548 3284
rect 508 3216 516 3224
rect 508 3196 516 3204
rect 556 3156 564 3164
rect 540 3136 548 3144
rect 524 3096 532 3104
rect 492 3036 500 3044
rect 428 2940 436 2944
rect 428 2936 436 2940
rect 460 2936 468 2944
rect 236 2896 244 2904
rect 348 2896 356 2904
rect 300 2876 308 2884
rect 220 2856 228 2864
rect 380 2876 388 2884
rect 412 2876 420 2884
rect 380 2836 388 2844
rect 316 2796 324 2804
rect 252 2756 260 2764
rect 300 2756 308 2764
rect 60 2696 68 2704
rect 108 2696 116 2704
rect 156 2696 164 2704
rect 268 2736 276 2744
rect 300 2736 308 2744
rect 76 2656 84 2664
rect 60 2616 68 2624
rect 12 2516 20 2524
rect 156 2616 164 2624
rect 76 2556 84 2564
rect 44 2540 52 2544
rect 44 2536 52 2540
rect 76 2516 84 2524
rect 124 2516 132 2524
rect 156 2516 164 2524
rect 92 2496 100 2504
rect 44 2296 52 2304
rect 92 2296 100 2304
rect 124 2296 132 2304
rect 12 2256 20 2264
rect 76 2276 84 2284
rect 108 2276 116 2284
rect 140 2276 148 2284
rect 92 2256 100 2264
rect 60 2176 68 2184
rect 92 2156 100 2164
rect 28 2136 36 2144
rect 44 1896 52 1904
rect 12 1876 20 1884
rect 44 1876 52 1884
rect 156 2256 164 2264
rect 124 2176 132 2184
rect 284 2636 292 2644
rect 188 2616 196 2624
rect 220 2556 228 2564
rect 268 2516 276 2524
rect 204 2416 212 2424
rect 284 2496 292 2504
rect 396 2736 404 2744
rect 396 2716 404 2724
rect 332 2696 340 2704
rect 364 2696 372 2704
rect 380 2696 388 2704
rect 348 2676 356 2684
rect 380 2676 388 2684
rect 620 3156 628 3164
rect 796 3256 804 3264
rect 764 3156 772 3164
rect 780 3156 788 3164
rect 844 3416 852 3424
rect 860 3336 868 3344
rect 860 3316 868 3324
rect 988 3496 996 3504
rect 956 3456 964 3464
rect 908 3376 916 3384
rect 876 3256 884 3264
rect 860 3216 868 3224
rect 668 3136 676 3144
rect 732 3136 740 3144
rect 812 3136 820 3144
rect 636 3116 644 3124
rect 652 3096 660 3104
rect 572 3076 580 3084
rect 652 2976 660 2984
rect 604 2896 612 2904
rect 524 2876 532 2884
rect 444 2816 452 2824
rect 316 2476 324 2484
rect 252 2456 260 2464
rect 300 2456 308 2464
rect 236 2376 244 2384
rect 540 2856 548 2864
rect 620 2856 628 2864
rect 588 2796 596 2804
rect 508 2756 516 2764
rect 460 2736 468 2744
rect 508 2736 516 2744
rect 524 2736 532 2744
rect 460 2696 468 2704
rect 572 2716 580 2724
rect 700 3116 708 3124
rect 780 3116 788 3124
rect 700 3096 708 3104
rect 732 3096 740 3104
rect 780 3056 788 3064
rect 684 2976 692 2984
rect 796 2996 804 3004
rect 748 2916 756 2924
rect 700 2876 708 2884
rect 812 2976 820 2984
rect 796 2876 804 2884
rect 684 2856 692 2864
rect 716 2856 724 2864
rect 812 2856 820 2864
rect 716 2836 724 2844
rect 668 2796 676 2804
rect 668 2756 676 2764
rect 620 2716 628 2724
rect 524 2696 532 2704
rect 588 2656 596 2664
rect 700 2696 708 2704
rect 732 2696 740 2704
rect 796 2696 804 2704
rect 652 2556 660 2564
rect 604 2536 612 2544
rect 684 2536 692 2544
rect 364 2516 372 2524
rect 588 2516 596 2524
rect 620 2516 628 2524
rect 668 2516 676 2524
rect 556 2496 564 2504
rect 492 2476 500 2484
rect 460 2456 468 2464
rect 348 2436 356 2444
rect 348 2376 356 2384
rect 412 2376 420 2384
rect 332 2356 340 2364
rect 300 2336 308 2344
rect 364 2336 372 2344
rect 412 2336 420 2344
rect 204 2296 212 2304
rect 316 2276 324 2284
rect 220 2256 228 2264
rect 172 2176 180 2184
rect 396 2276 404 2284
rect 412 2236 420 2244
rect 348 2176 356 2184
rect 140 2156 148 2164
rect 364 2156 372 2164
rect 428 2156 436 2164
rect 124 2116 132 2124
rect 156 2136 164 2144
rect 428 2136 436 2144
rect 444 2136 452 2144
rect 172 2116 180 2124
rect 396 2116 404 2124
rect 236 2096 244 2104
rect 172 1916 180 1924
rect 108 1896 116 1904
rect 140 1876 148 1884
rect 92 1756 100 1764
rect 140 1756 148 1764
rect 76 1736 84 1744
rect 44 1496 52 1504
rect 12 1456 20 1464
rect 44 1456 52 1464
rect 60 1456 68 1464
rect 44 1316 52 1324
rect 172 1736 180 1744
rect 236 1896 244 1904
rect 204 1876 212 1884
rect 204 1856 212 1864
rect 364 2076 372 2084
rect 428 2076 436 2084
rect 380 2056 388 2064
rect 444 2056 452 2064
rect 940 3136 948 3144
rect 892 3116 900 3124
rect 972 3356 980 3364
rect 1068 3776 1076 3784
rect 1036 3756 1044 3764
rect 1660 4396 1668 4404
rect 1580 4356 1588 4364
rect 2108 4956 2116 4964
rect 2092 4936 2100 4944
rect 2396 5276 2404 5284
rect 2492 5116 2500 5124
rect 2188 5096 2196 5104
rect 2316 5096 2324 5104
rect 2236 5076 2244 5084
rect 2220 5016 2228 5024
rect 2396 5096 2404 5104
rect 2492 5096 2500 5104
rect 2364 5076 2372 5084
rect 2348 5016 2356 5024
rect 2172 4976 2180 4984
rect 2300 4976 2308 4984
rect 2316 4976 2324 4984
rect 2236 4956 2244 4964
rect 2300 4956 2308 4964
rect 2076 4916 2084 4924
rect 2092 4916 2100 4924
rect 1948 4896 1956 4904
rect 1980 4896 1988 4904
rect 2028 4896 2036 4904
rect 2060 4896 2068 4904
rect 1916 4836 1924 4844
rect 1964 4836 1972 4844
rect 1948 4776 1956 4784
rect 1932 4676 1940 4684
rect 1740 4636 1748 4644
rect 1868 4576 1876 4584
rect 1900 4636 1908 4644
rect 1836 4556 1844 4564
rect 1884 4556 1892 4564
rect 1740 4516 1748 4524
rect 1884 4516 1892 4524
rect 1772 4496 1780 4504
rect 1916 4496 1924 4504
rect 1772 4456 1780 4464
rect 1820 4456 1828 4464
rect 1756 4396 1764 4404
rect 1692 4336 1700 4344
rect 1740 4336 1748 4344
rect 1564 4276 1572 4284
rect 1612 4276 1620 4284
rect 1628 4256 1636 4264
rect 1676 4256 1684 4264
rect 1468 4176 1476 4184
rect 1516 4136 1524 4144
rect 1196 4116 1204 4124
rect 1244 4116 1252 4124
rect 1644 4196 1652 4204
rect 1740 4316 1748 4324
rect 1708 4296 1716 4304
rect 1724 4296 1732 4304
rect 1804 4336 1812 4344
rect 1852 4336 1860 4344
rect 1788 4296 1796 4304
rect 1820 4316 1828 4324
rect 2012 4816 2020 4824
rect 2012 4796 2020 4804
rect 2332 4936 2340 4944
rect 2364 4936 2372 4944
rect 2236 4916 2244 4924
rect 2124 4876 2132 4884
rect 2220 4876 2228 4884
rect 2012 4756 2020 4764
rect 2108 4756 2116 4764
rect 1980 4696 1988 4704
rect 1996 4636 2004 4644
rect 1964 4596 1972 4604
rect 1980 4596 1988 4604
rect 1948 4556 1956 4564
rect 1948 4516 1956 4524
rect 1980 4516 1988 4524
rect 1932 4376 1940 4384
rect 1948 4376 1956 4384
rect 2092 4716 2100 4724
rect 2140 4716 2148 4724
rect 2188 4716 2196 4724
rect 2412 5056 2420 5064
rect 2428 5036 2436 5044
rect 2460 5036 2468 5044
rect 2428 4996 2436 5004
rect 2428 4936 2436 4944
rect 2396 4916 2404 4924
rect 2348 4896 2356 4904
rect 2332 4856 2340 4864
rect 2284 4756 2292 4764
rect 2364 4756 2372 4764
rect 2252 4736 2260 4744
rect 2060 4596 2068 4604
rect 2044 4576 2052 4584
rect 2236 4676 2244 4684
rect 2156 4576 2164 4584
rect 2220 4576 2228 4584
rect 2028 4556 2036 4564
rect 2092 4556 2100 4564
rect 2492 4956 2500 4964
rect 2540 5216 2548 5224
rect 2556 5176 2564 5184
rect 2508 4936 2516 4944
rect 2524 4936 2532 4944
rect 2524 4916 2532 4924
rect 2524 4776 2532 4784
rect 2316 4736 2324 4744
rect 2412 4736 2420 4744
rect 2300 4676 2308 4684
rect 2380 4716 2388 4724
rect 2268 4636 2276 4644
rect 2316 4616 2324 4624
rect 2284 4556 2292 4564
rect 2108 4516 2116 4524
rect 2204 4516 2212 4524
rect 1996 4336 2004 4344
rect 1980 4316 1988 4324
rect 1996 4316 2004 4324
rect 1884 4296 1892 4304
rect 1900 4296 1908 4304
rect 1788 4276 1796 4284
rect 1868 4276 1876 4284
rect 1884 4276 1892 4284
rect 1548 4176 1556 4184
rect 1596 4176 1604 4184
rect 1708 4156 1716 4164
rect 1740 4156 1748 4164
rect 1564 4136 1572 4144
rect 1660 4136 1668 4144
rect 1676 4116 1684 4124
rect 1740 4116 1748 4124
rect 1180 4016 1188 4024
rect 1132 3896 1140 3904
rect 1228 3916 1236 3924
rect 1411 4006 1419 4014
rect 1421 4006 1429 4014
rect 1431 4006 1439 4014
rect 1441 4006 1449 4014
rect 1451 4006 1459 4014
rect 1461 4006 1469 4014
rect 1356 3976 1364 3984
rect 1212 3896 1220 3904
rect 1244 3896 1252 3904
rect 1164 3876 1172 3884
rect 1180 3876 1188 3884
rect 1196 3856 1204 3864
rect 1196 3756 1204 3764
rect 1052 3736 1060 3744
rect 1196 3736 1204 3744
rect 1228 3876 1236 3884
rect 1244 3796 1252 3804
rect 1276 3896 1284 3904
rect 1340 3896 1348 3904
rect 1404 3896 1412 3904
rect 1516 3896 1524 3904
rect 1548 3876 1556 3884
rect 1292 3856 1300 3864
rect 1308 3856 1316 3864
rect 1356 3856 1364 3864
rect 1388 3856 1396 3864
rect 1548 3856 1556 3864
rect 1308 3796 1316 3804
rect 1484 3776 1492 3784
rect 1356 3756 1364 3764
rect 1404 3756 1412 3764
rect 1388 3736 1396 3744
rect 1036 3596 1044 3604
rect 1068 3576 1076 3584
rect 1436 3716 1444 3724
rect 1292 3636 1300 3644
rect 1276 3596 1284 3604
rect 1084 3496 1092 3504
rect 1148 3496 1156 3504
rect 1164 3476 1172 3484
rect 1052 3456 1060 3464
rect 1020 3416 1028 3424
rect 1084 3416 1092 3424
rect 1020 3376 1028 3384
rect 1004 3336 1012 3344
rect 1068 3336 1076 3344
rect 1260 3516 1268 3524
rect 1196 3496 1204 3504
rect 1196 3456 1204 3464
rect 1411 3606 1419 3614
rect 1421 3606 1429 3614
rect 1431 3606 1439 3614
rect 1441 3606 1449 3614
rect 1451 3606 1459 3614
rect 1461 3606 1469 3614
rect 1388 3596 1396 3604
rect 1372 3556 1380 3564
rect 1404 3516 1412 3524
rect 1420 3516 1428 3524
rect 1228 3456 1236 3464
rect 1260 3456 1268 3464
rect 1116 3336 1124 3344
rect 972 3096 980 3104
rect 908 3056 916 3064
rect 908 2896 916 2904
rect 876 2876 884 2884
rect 908 2876 916 2884
rect 844 2736 852 2744
rect 828 2716 836 2724
rect 956 2936 964 2944
rect 924 2856 932 2864
rect 876 2776 884 2784
rect 908 2756 916 2764
rect 860 2696 868 2704
rect 764 2656 772 2664
rect 764 2556 772 2564
rect 748 2476 756 2484
rect 604 2436 612 2444
rect 636 2436 644 2444
rect 636 2376 644 2384
rect 732 2376 740 2384
rect 540 2356 548 2364
rect 556 2356 564 2364
rect 524 2316 532 2324
rect 476 2296 484 2304
rect 476 2276 484 2284
rect 508 2136 516 2144
rect 476 2116 484 2124
rect 460 2016 468 2024
rect 556 2336 564 2344
rect 620 2336 628 2344
rect 604 2296 612 2304
rect 556 2236 564 2244
rect 508 2076 516 2084
rect 556 2076 564 2084
rect 588 2156 596 2164
rect 572 2036 580 2044
rect 556 1996 564 2004
rect 524 1976 532 1984
rect 476 1956 484 1964
rect 364 1936 372 1944
rect 572 1936 580 1944
rect 300 1916 308 1924
rect 524 1916 532 1924
rect 268 1856 276 1864
rect 188 1716 196 1724
rect 172 1696 180 1704
rect 204 1696 212 1704
rect 108 1496 116 1504
rect 620 2156 628 2164
rect 604 2116 612 2124
rect 604 2096 612 2104
rect 652 2356 660 2364
rect 684 2336 692 2344
rect 940 2816 948 2824
rect 876 2636 884 2644
rect 908 2636 916 2644
rect 924 2636 932 2644
rect 780 2336 788 2344
rect 780 2316 788 2324
rect 732 2296 740 2304
rect 764 2296 772 2304
rect 844 2316 852 2324
rect 844 2236 852 2244
rect 748 2196 756 2204
rect 700 2156 708 2164
rect 700 2116 708 2124
rect 748 2116 756 2124
rect 828 2116 836 2124
rect 684 2076 692 2084
rect 812 2076 820 2084
rect 668 1936 676 1944
rect 636 1916 644 1924
rect 652 1916 660 1924
rect 556 1896 564 1904
rect 588 1896 596 1904
rect 652 1896 660 1904
rect 684 1896 692 1904
rect 332 1736 340 1744
rect 268 1716 276 1724
rect 348 1716 356 1724
rect 140 1456 148 1464
rect 204 1456 212 1464
rect 204 1436 212 1444
rect 92 1416 100 1424
rect 156 1416 164 1424
rect 156 1376 164 1384
rect 236 1436 244 1444
rect 220 1416 228 1424
rect 220 1396 228 1404
rect 412 1856 420 1864
rect 444 1856 452 1864
rect 428 1736 436 1744
rect 396 1716 404 1724
rect 412 1716 420 1724
rect 380 1696 388 1704
rect 316 1496 324 1504
rect 268 1396 276 1404
rect 252 1376 260 1384
rect 316 1476 324 1484
rect 796 1896 804 1904
rect 620 1876 628 1884
rect 716 1880 724 1884
rect 716 1876 724 1880
rect 780 1876 788 1884
rect 812 1876 820 1884
rect 828 1876 836 1884
rect 460 1836 468 1844
rect 524 1836 532 1844
rect 732 1816 740 1824
rect 700 1756 708 1764
rect 460 1740 468 1744
rect 460 1736 468 1740
rect 492 1736 500 1744
rect 604 1736 612 1744
rect 476 1696 484 1704
rect 588 1696 596 1704
rect 636 1696 644 1704
rect 668 1656 676 1664
rect 652 1636 660 1644
rect 492 1596 500 1604
rect 540 1596 548 1604
rect 380 1476 388 1484
rect 332 1436 340 1444
rect 492 1456 500 1464
rect 508 1456 516 1464
rect 476 1436 484 1444
rect 620 1556 628 1564
rect 556 1480 564 1484
rect 556 1476 564 1480
rect 524 1436 532 1444
rect 364 1396 372 1404
rect 268 1356 276 1364
rect 412 1356 420 1364
rect 524 1356 532 1364
rect 748 1756 756 1764
rect 796 1756 804 1764
rect 764 1736 772 1744
rect 748 1696 756 1704
rect 812 1716 820 1724
rect 748 1676 756 1684
rect 780 1676 788 1684
rect 780 1596 788 1604
rect 892 2276 900 2284
rect 860 2216 868 2224
rect 924 2516 932 2524
rect 988 2936 996 2944
rect 988 2916 996 2924
rect 1116 3256 1124 3264
rect 1308 3456 1316 3464
rect 1292 3416 1300 3424
rect 1292 3336 1300 3344
rect 1260 3296 1268 3304
rect 1276 3276 1284 3284
rect 1404 3376 1412 3384
rect 1420 3356 1428 3364
rect 1356 3316 1364 3324
rect 1324 3296 1332 3304
rect 1340 3276 1348 3284
rect 1196 3176 1204 3184
rect 1148 3136 1156 3144
rect 1164 3136 1172 3144
rect 1212 3136 1220 3144
rect 1052 3116 1060 3124
rect 1084 2996 1092 3004
rect 1148 3076 1156 3084
rect 1148 2996 1156 3004
rect 1100 2976 1108 2984
rect 1052 2956 1060 2964
rect 1084 2956 1092 2964
rect 1100 2956 1108 2964
rect 1132 2956 1140 2964
rect 1036 2916 1044 2924
rect 1180 2956 1188 2964
rect 1308 3256 1316 3264
rect 1308 3156 1316 3164
rect 1276 3116 1284 3124
rect 1260 3096 1268 3104
rect 1324 3136 1332 3144
rect 1324 3116 1332 3124
rect 1276 3076 1284 3084
rect 1244 2996 1252 3004
rect 1228 2976 1236 2984
rect 1260 2976 1268 2984
rect 1212 2936 1220 2944
rect 1244 2936 1252 2944
rect 1068 2876 1076 2884
rect 1132 2856 1140 2864
rect 1020 2796 1028 2804
rect 956 2756 964 2764
rect 956 2716 964 2724
rect 972 2656 980 2664
rect 956 2556 964 2564
rect 956 2436 964 2444
rect 940 2356 948 2364
rect 956 2336 964 2344
rect 1004 2756 1012 2764
rect 1036 2756 1044 2764
rect 1068 2796 1076 2804
rect 1116 2736 1124 2744
rect 1244 2876 1252 2884
rect 1212 2816 1220 2824
rect 1148 2796 1156 2804
rect 1196 2796 1204 2804
rect 1148 2736 1156 2744
rect 1292 2916 1300 2924
rect 1340 3096 1348 3104
rect 1411 3206 1419 3214
rect 1421 3206 1429 3214
rect 1431 3206 1439 3214
rect 1441 3206 1449 3214
rect 1451 3206 1459 3214
rect 1461 3206 1469 3214
rect 1388 3096 1396 3104
rect 1340 2956 1348 2964
rect 1340 2916 1348 2924
rect 1324 2896 1332 2904
rect 1292 2876 1300 2884
rect 1308 2816 1316 2824
rect 1276 2756 1284 2764
rect 1324 2796 1332 2804
rect 1532 3736 1540 3744
rect 1548 3716 1556 3724
rect 1628 3976 1636 3984
rect 1580 3936 1588 3944
rect 1580 3836 1588 3844
rect 1612 3836 1620 3844
rect 1596 3756 1604 3764
rect 1964 4276 1972 4284
rect 2012 4296 2020 4304
rect 1932 4256 1940 4264
rect 1916 4216 1924 4224
rect 1820 4156 1828 4164
rect 1900 4156 1908 4164
rect 1996 4196 2004 4204
rect 1836 4136 1844 4144
rect 1852 4116 1860 4124
rect 1756 4096 1764 4104
rect 1964 4116 1972 4124
rect 1948 4096 1956 4104
rect 1868 4076 1876 4084
rect 1900 3996 1908 4004
rect 1692 3976 1700 3984
rect 1836 3916 1844 3924
rect 1852 3916 1860 3924
rect 1708 3896 1716 3904
rect 1772 3896 1780 3904
rect 1804 3896 1812 3904
rect 1660 3756 1668 3764
rect 1660 3736 1668 3744
rect 1580 3696 1588 3704
rect 1564 3596 1572 3604
rect 1612 3696 1620 3704
rect 1628 3556 1636 3564
rect 1596 3516 1604 3524
rect 1644 3496 1652 3504
rect 1516 3476 1524 3484
rect 1500 3436 1508 3444
rect 1644 3436 1652 3444
rect 1532 3376 1540 3384
rect 1548 3356 1556 3364
rect 1612 3396 1620 3404
rect 1580 3356 1588 3364
rect 1564 3316 1572 3324
rect 1564 3276 1572 3284
rect 1516 3236 1524 3244
rect 1500 3176 1508 3184
rect 1548 3196 1556 3204
rect 1516 3096 1524 3104
rect 1484 3056 1492 3064
rect 1644 3336 1652 3344
rect 1676 3556 1684 3564
rect 1676 3476 1684 3484
rect 1724 3876 1732 3884
rect 1820 3876 1828 3884
rect 1836 3876 1844 3884
rect 1868 3876 1876 3884
rect 1980 3856 1988 3864
rect 1740 3756 1748 3764
rect 1708 3716 1716 3724
rect 1740 3716 1748 3724
rect 1692 3416 1700 3424
rect 1708 3396 1716 3404
rect 1692 3336 1700 3344
rect 1804 3796 1812 3804
rect 1852 3796 1860 3804
rect 1932 3776 1940 3784
rect 1836 3756 1844 3764
rect 1868 3756 1876 3764
rect 2044 4256 2052 4264
rect 2044 4216 2052 4224
rect 2108 4456 2116 4464
rect 2300 4496 2308 4504
rect 2348 4496 2356 4504
rect 2508 4702 2516 4704
rect 2508 4696 2516 4702
rect 2620 5156 2628 5164
rect 2700 5156 2708 5164
rect 2684 5096 2692 5104
rect 2732 5096 2740 5104
rect 2588 5076 2596 5084
rect 2556 5056 2564 5064
rect 2572 5016 2580 5024
rect 2556 4996 2564 5004
rect 2828 5296 2836 5304
rect 2908 5316 2916 5324
rect 3036 5296 3044 5304
rect 2988 5276 2996 5284
rect 2892 5216 2900 5224
rect 2908 5216 2916 5224
rect 2876 5116 2884 5124
rect 3020 5096 3028 5104
rect 2988 5076 2996 5084
rect 3004 5076 3012 5084
rect 2988 5016 2996 5024
rect 2915 5006 2923 5014
rect 2925 5006 2933 5014
rect 2935 5006 2943 5014
rect 2945 5006 2953 5014
rect 2955 5006 2963 5014
rect 2965 5006 2973 5014
rect 2812 4996 2820 5004
rect 2748 4976 2756 4984
rect 2748 4918 2756 4924
rect 2748 4916 2756 4918
rect 2812 4916 2820 4924
rect 2876 4916 2884 4924
rect 2572 4896 2580 4904
rect 2748 4896 2756 4904
rect 2844 4896 2852 4904
rect 2572 4876 2580 4884
rect 2620 4836 2628 4844
rect 2620 4796 2628 4804
rect 2604 4776 2612 4784
rect 2556 4756 2564 4764
rect 2668 4776 2676 4784
rect 2636 4736 2644 4744
rect 2732 4756 2740 4764
rect 2732 4716 2740 4724
rect 2940 4916 2948 4924
rect 3036 4916 3044 4924
rect 2924 4896 2932 4904
rect 2892 4876 2900 4884
rect 2860 4796 2868 4804
rect 2796 4736 2804 4744
rect 2572 4696 2580 4704
rect 2604 4696 2612 4704
rect 2700 4696 2708 4704
rect 2748 4696 2756 4704
rect 2652 4676 2660 4684
rect 2556 4576 2564 4584
rect 2492 4556 2500 4564
rect 2380 4456 2388 4464
rect 2172 4376 2180 4384
rect 2364 4356 2372 4364
rect 2092 4336 2100 4344
rect 2188 4336 2196 4344
rect 2076 4296 2084 4304
rect 2348 4316 2356 4324
rect 2124 4296 2132 4304
rect 2220 4296 2228 4304
rect 2124 4276 2132 4284
rect 2172 4276 2180 4284
rect 2140 4256 2148 4264
rect 2092 4196 2100 4204
rect 2172 4216 2180 4224
rect 2156 4196 2164 4204
rect 2044 4176 2052 4184
rect 2172 4176 2180 4184
rect 2092 4156 2100 4164
rect 2188 4156 2196 4164
rect 2348 4256 2356 4264
rect 2252 4216 2260 4224
rect 2300 4216 2308 4224
rect 2220 4136 2228 4144
rect 2284 4136 2292 4144
rect 2124 4116 2132 4124
rect 2252 4116 2260 4124
rect 2060 4096 2068 4104
rect 2220 4096 2228 4104
rect 2092 3976 2100 3984
rect 2236 3976 2244 3984
rect 2108 3936 2116 3944
rect 2140 3936 2148 3944
rect 2012 3896 2020 3904
rect 2028 3876 2036 3884
rect 2060 3876 2068 3884
rect 2108 3856 2116 3864
rect 2252 3896 2260 3904
rect 2684 4676 2692 4684
rect 2668 4656 2676 4664
rect 2732 4636 2740 4644
rect 2748 4556 2756 4564
rect 2684 4536 2692 4544
rect 2732 4536 2740 4544
rect 2572 4516 2580 4524
rect 2700 4516 2708 4524
rect 2556 4496 2564 4504
rect 2428 4296 2436 4304
rect 2476 4296 2484 4304
rect 2396 4276 2404 4284
rect 2444 4276 2452 4284
rect 2444 4216 2452 4224
rect 2460 4216 2468 4224
rect 2396 4196 2404 4204
rect 2380 4116 2388 4124
rect 2428 4116 2436 4124
rect 2316 4096 2324 4104
rect 2300 4036 2308 4044
rect 2444 4036 2452 4044
rect 2332 3936 2340 3944
rect 2348 3896 2356 3904
rect 2412 3896 2420 3904
rect 2188 3876 2196 3884
rect 2284 3876 2292 3884
rect 2316 3876 2324 3884
rect 2428 3876 2436 3884
rect 2220 3836 2228 3844
rect 2252 3836 2260 3844
rect 2140 3816 2148 3824
rect 2204 3776 2212 3784
rect 2172 3756 2180 3764
rect 2220 3756 2228 3764
rect 1948 3736 1956 3744
rect 1996 3736 2004 3744
rect 2044 3736 2052 3744
rect 1788 3716 1796 3724
rect 1820 3716 1828 3724
rect 1916 3716 1924 3724
rect 1964 3716 1972 3724
rect 1852 3596 1860 3604
rect 1900 3596 1908 3604
rect 1980 3596 1988 3604
rect 1740 3536 1748 3544
rect 1756 3536 1764 3544
rect 1740 3496 1748 3504
rect 1724 3316 1732 3324
rect 1660 3276 1668 3284
rect 1740 3216 1748 3224
rect 1724 3176 1732 3184
rect 1580 3076 1588 3084
rect 1708 3076 1716 3084
rect 1804 3476 1812 3484
rect 1788 3436 1796 3444
rect 1788 3356 1796 3364
rect 1836 3376 1844 3384
rect 1804 3316 1812 3324
rect 1820 3316 1828 3324
rect 1820 3296 1828 3304
rect 1948 3556 1956 3564
rect 1868 3536 1876 3544
rect 1932 3516 1940 3524
rect 1884 3496 1892 3504
rect 1916 3496 1924 3504
rect 1900 3456 1908 3464
rect 1964 3456 1972 3464
rect 1868 3356 1876 3364
rect 1964 3376 1972 3384
rect 2012 3556 2020 3564
rect 2348 3836 2356 3844
rect 2300 3796 2308 3804
rect 2300 3756 2308 3764
rect 2396 3736 2404 3744
rect 2300 3716 2308 3724
rect 2012 3536 2020 3544
rect 2044 3536 2052 3544
rect 2060 3536 2068 3544
rect 2172 3536 2180 3544
rect 2156 3496 2164 3504
rect 1996 3476 2004 3484
rect 2092 3476 2100 3484
rect 2140 3476 2148 3484
rect 2172 3476 2180 3484
rect 2012 3456 2020 3464
rect 2140 3456 2148 3464
rect 1996 3436 2004 3444
rect 2028 3416 2036 3424
rect 1996 3396 2004 3404
rect 1980 3356 1988 3364
rect 1932 3336 1940 3344
rect 1964 3340 1972 3344
rect 1964 3336 1972 3340
rect 1996 3336 2004 3344
rect 1868 3316 1876 3324
rect 2044 3316 2052 3324
rect 2076 3316 2084 3324
rect 1852 3276 1860 3284
rect 1852 3256 1860 3264
rect 1788 3216 1796 3224
rect 1804 3136 1812 3144
rect 1772 3116 1780 3124
rect 1564 3036 1572 3044
rect 1388 2956 1396 2964
rect 1404 2956 1412 2964
rect 1612 3036 1620 3044
rect 1724 3036 1732 3044
rect 1548 3016 1556 3024
rect 1596 2996 1604 3004
rect 1516 2956 1524 2964
rect 1516 2936 1524 2944
rect 1548 2936 1556 2944
rect 1516 2916 1524 2924
rect 1484 2856 1492 2864
rect 1532 2836 1540 2844
rect 1388 2816 1396 2824
rect 1500 2816 1508 2824
rect 1411 2806 1419 2814
rect 1421 2806 1429 2814
rect 1431 2806 1439 2814
rect 1441 2806 1449 2814
rect 1451 2806 1459 2814
rect 1461 2806 1469 2814
rect 1324 2756 1332 2764
rect 1372 2736 1380 2744
rect 1340 2716 1348 2724
rect 1004 2696 1012 2704
rect 1036 2696 1044 2704
rect 1212 2696 1220 2704
rect 1260 2696 1268 2704
rect 1036 2596 1044 2604
rect 1020 2556 1028 2564
rect 1116 2676 1124 2684
rect 1132 2556 1140 2564
rect 1148 2516 1156 2524
rect 1212 2516 1220 2524
rect 1164 2496 1172 2504
rect 1180 2496 1188 2504
rect 1116 2436 1124 2444
rect 1116 2376 1124 2384
rect 1004 2356 1012 2364
rect 924 2316 932 2324
rect 956 2316 964 2324
rect 940 2276 948 2284
rect 860 2116 868 2124
rect 972 2276 980 2284
rect 988 2256 996 2264
rect 972 2196 980 2204
rect 956 2136 964 2144
rect 988 2116 996 2124
rect 908 2096 916 2104
rect 940 2096 948 2104
rect 892 2016 900 2024
rect 860 1916 868 1924
rect 876 1876 884 1884
rect 844 1756 852 1764
rect 844 1736 852 1744
rect 828 1676 836 1684
rect 892 1696 900 1704
rect 892 1636 900 1644
rect 892 1616 900 1624
rect 860 1576 868 1584
rect 700 1556 708 1564
rect 732 1556 740 1564
rect 796 1556 804 1564
rect 860 1556 868 1564
rect 668 1516 676 1524
rect 764 1516 772 1524
rect 780 1516 788 1524
rect 828 1516 836 1524
rect 876 1516 884 1524
rect 700 1496 708 1504
rect 716 1496 724 1504
rect 780 1496 788 1504
rect 844 1496 852 1504
rect 652 1456 660 1464
rect 812 1476 820 1484
rect 588 1436 596 1444
rect 652 1436 660 1444
rect 684 1436 692 1444
rect 140 1316 148 1324
rect 188 1316 196 1324
rect 220 1316 228 1324
rect 12 1296 20 1304
rect 108 1236 116 1244
rect 844 1396 852 1404
rect 604 1356 612 1364
rect 700 1356 708 1364
rect 508 1336 516 1344
rect 668 1336 676 1344
rect 764 1336 772 1344
rect 364 1276 372 1284
rect 348 1176 356 1184
rect 220 1116 228 1124
rect 284 1116 292 1124
rect 348 1116 356 1124
rect 12 1096 20 1104
rect 300 1096 308 1104
rect 172 1076 180 1084
rect 236 1076 244 1084
rect 44 1056 52 1064
rect 108 1056 116 1064
rect 124 996 132 1004
rect 124 956 132 964
rect 12 896 20 904
rect 108 936 116 944
rect 92 916 100 924
rect 60 716 68 724
rect 44 696 52 704
rect 284 1076 292 1084
rect 316 1076 324 1084
rect 268 1056 276 1064
rect 236 996 244 1004
rect 204 936 212 944
rect 268 936 276 944
rect 300 916 308 924
rect 300 896 308 904
rect 268 876 276 884
rect 124 736 132 744
rect 204 736 212 744
rect 124 696 132 704
rect 332 1036 340 1044
rect 332 956 340 964
rect 428 1236 436 1244
rect 380 1156 388 1164
rect 380 1096 388 1104
rect 476 1116 484 1124
rect 396 1076 404 1084
rect 380 1056 388 1064
rect 460 1056 468 1064
rect 380 996 388 1004
rect 508 1076 516 1084
rect 492 1036 500 1044
rect 412 976 420 984
rect 396 956 404 964
rect 460 956 468 964
rect 508 956 516 964
rect 380 916 388 924
rect 428 916 436 924
rect 380 896 388 904
rect 556 1076 564 1084
rect 540 1036 548 1044
rect 556 976 564 984
rect 556 876 564 884
rect 524 856 532 864
rect 268 716 276 724
rect 396 716 404 724
rect 460 716 468 724
rect 492 716 500 724
rect 284 696 292 704
rect 412 696 420 704
rect 108 656 116 664
rect 188 656 196 664
rect 316 656 324 664
rect 76 576 84 584
rect 156 576 164 584
rect 252 576 260 584
rect 300 576 308 584
rect 364 656 372 664
rect 380 656 388 664
rect 444 676 452 684
rect 444 656 452 664
rect 364 636 372 644
rect 428 636 436 644
rect 332 616 340 624
rect 316 556 324 564
rect 412 556 420 564
rect 44 516 52 524
rect 172 516 180 524
rect 220 516 228 524
rect 284 516 292 524
rect 124 476 132 484
rect 124 316 132 324
rect 188 496 196 504
rect 92 296 100 304
rect 60 276 68 284
rect 108 276 116 284
rect 172 276 180 284
rect 220 276 228 284
rect 204 256 212 264
rect 12 216 20 224
rect 76 236 84 244
rect 332 516 340 524
rect 588 1316 596 1324
rect 620 1316 628 1324
rect 732 1256 740 1264
rect 684 1216 692 1224
rect 668 1116 676 1124
rect 588 1096 596 1104
rect 636 1076 644 1084
rect 812 1296 820 1304
rect 764 1136 772 1144
rect 700 1096 708 1104
rect 716 1096 724 1104
rect 588 1016 596 1024
rect 652 1056 660 1064
rect 652 996 660 1004
rect 636 976 644 984
rect 892 1316 900 1324
rect 956 2076 964 2084
rect 972 1976 980 1984
rect 1100 2336 1108 2344
rect 1052 2316 1060 2324
rect 1052 2236 1060 2244
rect 1100 2256 1108 2264
rect 1052 2216 1060 2224
rect 1132 2256 1140 2264
rect 1372 2696 1380 2704
rect 1484 2696 1492 2704
rect 1516 2776 1524 2784
rect 1564 2876 1572 2884
rect 1580 2836 1588 2844
rect 1564 2776 1572 2784
rect 1516 2656 1524 2664
rect 1292 2576 1300 2584
rect 1244 2556 1252 2564
rect 1500 2556 1508 2564
rect 1548 2736 1556 2744
rect 1628 2836 1636 2844
rect 1612 2756 1620 2764
rect 1612 2736 1620 2744
rect 1564 2696 1572 2704
rect 1628 2696 1636 2704
rect 1580 2656 1588 2664
rect 1628 2656 1636 2664
rect 1308 2516 1316 2524
rect 1356 2516 1364 2524
rect 1468 2516 1476 2524
rect 1500 2516 1508 2524
rect 1548 2516 1556 2524
rect 1228 2476 1236 2484
rect 1212 2436 1220 2444
rect 1180 2336 1188 2344
rect 1196 2336 1204 2344
rect 1180 2316 1188 2324
rect 1292 2316 1300 2324
rect 1356 2496 1364 2504
rect 1196 2296 1204 2304
rect 1212 2296 1220 2304
rect 1164 2216 1172 2224
rect 1148 2196 1156 2204
rect 1116 2156 1124 2164
rect 1148 2156 1156 2164
rect 1276 2236 1284 2244
rect 1228 2156 1236 2164
rect 1260 2156 1268 2164
rect 1260 2136 1268 2144
rect 1212 2116 1220 2124
rect 1052 2096 1060 2104
rect 1100 2096 1108 2104
rect 1180 2076 1188 2084
rect 1100 2036 1108 2044
rect 1020 1996 1028 2004
rect 1036 1936 1044 1944
rect 1068 1936 1076 1944
rect 1164 1936 1172 1944
rect 1036 1896 1044 1904
rect 1036 1876 1044 1884
rect 1068 1876 1076 1884
rect 940 1816 948 1824
rect 940 1756 948 1764
rect 1020 1756 1028 1764
rect 924 1576 932 1584
rect 924 1536 932 1544
rect 972 1716 980 1724
rect 1004 1696 1012 1704
rect 956 1676 964 1684
rect 956 1636 964 1644
rect 956 1596 964 1604
rect 988 1596 996 1604
rect 972 1536 980 1544
rect 1004 1536 1012 1544
rect 940 1516 948 1524
rect 956 1516 964 1524
rect 972 1496 980 1504
rect 972 1476 980 1484
rect 1068 1736 1076 1744
rect 1116 1896 1124 1904
rect 1164 1896 1172 1904
rect 1212 1916 1220 1924
rect 1212 1896 1220 1904
rect 1212 1876 1220 1884
rect 1180 1856 1188 1864
rect 1292 2136 1300 2144
rect 1411 2406 1419 2414
rect 1421 2406 1429 2414
rect 1431 2406 1439 2414
rect 1441 2406 1449 2414
rect 1451 2406 1459 2414
rect 1461 2406 1469 2414
rect 1468 2316 1476 2324
rect 1388 2296 1396 2304
rect 1388 2276 1396 2284
rect 1420 2276 1428 2284
rect 1372 2196 1380 2204
rect 1404 2256 1412 2264
rect 1388 2176 1396 2184
rect 1420 2156 1428 2164
rect 1388 2116 1396 2124
rect 1372 2096 1380 2104
rect 1340 2036 1348 2044
rect 1372 1976 1380 1984
rect 1324 1896 1332 1904
rect 1276 1876 1284 1884
rect 1276 1856 1284 1864
rect 1212 1776 1220 1784
rect 1484 2096 1492 2104
rect 1468 2076 1476 2084
rect 1420 2036 1428 2044
rect 1411 2006 1419 2014
rect 1421 2006 1429 2014
rect 1431 2006 1439 2014
rect 1441 2006 1449 2014
rect 1451 2006 1459 2014
rect 1461 2006 1469 2014
rect 1404 1936 1412 1944
rect 1548 2496 1556 2504
rect 1516 2476 1524 2484
rect 1676 2996 1684 3004
rect 1820 3096 1828 3104
rect 1852 3096 1860 3104
rect 1772 3056 1780 3064
rect 1788 3056 1796 3064
rect 1836 3056 1844 3064
rect 1852 3056 1860 3064
rect 1740 2936 1748 2944
rect 1660 2876 1668 2884
rect 1724 2876 1732 2884
rect 1692 2796 1700 2804
rect 1660 2756 1668 2764
rect 1612 2556 1620 2564
rect 1580 2396 1588 2404
rect 1532 2376 1540 2384
rect 1596 2376 1604 2384
rect 1564 2336 1572 2344
rect 1628 2356 1636 2364
rect 1612 2296 1620 2304
rect 1548 2256 1556 2264
rect 1564 2256 1572 2264
rect 1532 2176 1540 2184
rect 1548 2176 1556 2184
rect 1516 2156 1524 2164
rect 1500 2076 1508 2084
rect 1484 1896 1492 1904
rect 1596 2216 1604 2224
rect 1580 2196 1588 2204
rect 1516 1916 1524 1924
rect 1388 1776 1396 1784
rect 1132 1716 1140 1724
rect 1164 1716 1172 1724
rect 1116 1696 1124 1704
rect 1116 1656 1124 1664
rect 1084 1636 1092 1644
rect 1068 1596 1076 1604
rect 1068 1536 1076 1544
rect 1052 1516 1060 1524
rect 1084 1516 1092 1524
rect 1148 1636 1156 1644
rect 1292 1696 1300 1704
rect 1340 1736 1348 1744
rect 1484 1716 1492 1724
rect 1292 1656 1300 1664
rect 1276 1616 1284 1624
rect 1212 1556 1220 1564
rect 1228 1556 1236 1564
rect 1244 1516 1252 1524
rect 1164 1496 1172 1504
rect 1212 1496 1220 1504
rect 1036 1476 1044 1484
rect 1068 1476 1076 1484
rect 1132 1456 1140 1464
rect 1132 1436 1140 1444
rect 988 1416 996 1424
rect 1020 1416 1028 1424
rect 1068 1416 1076 1424
rect 1020 1396 1028 1404
rect 972 1376 980 1384
rect 924 1316 932 1324
rect 1036 1316 1044 1324
rect 1068 1316 1076 1324
rect 1100 1316 1108 1324
rect 1004 1216 1012 1224
rect 860 1196 868 1204
rect 924 1196 932 1204
rect 716 1076 724 1084
rect 764 1076 772 1084
rect 684 1056 692 1064
rect 732 1036 740 1044
rect 764 1016 772 1024
rect 620 956 628 964
rect 716 956 724 964
rect 796 956 804 964
rect 716 936 724 944
rect 796 936 804 944
rect 812 936 820 944
rect 780 916 788 924
rect 812 876 820 884
rect 748 836 756 844
rect 684 756 692 764
rect 540 736 548 744
rect 572 736 580 744
rect 636 716 644 724
rect 620 696 628 704
rect 556 676 564 684
rect 556 656 564 664
rect 636 656 644 664
rect 524 576 532 584
rect 556 576 564 584
rect 524 556 532 564
rect 380 496 388 504
rect 396 496 404 504
rect 348 476 356 484
rect 332 356 340 364
rect 620 636 628 644
rect 572 536 580 544
rect 604 516 612 524
rect 556 496 564 504
rect 508 356 516 364
rect 348 316 356 324
rect 380 316 388 324
rect 508 316 516 324
rect 348 296 356 304
rect 428 296 436 304
rect 476 296 484 304
rect 332 276 340 284
rect 396 276 404 284
rect 444 276 452 284
rect 492 276 500 284
rect 524 276 532 284
rect 204 216 212 224
rect 284 196 292 204
rect 60 176 68 184
rect 92 176 100 184
rect 268 176 276 184
rect 444 256 452 264
rect 476 236 484 244
rect 492 236 500 244
rect 316 216 324 224
rect 444 216 452 224
rect 396 196 404 204
rect 172 156 180 164
rect 316 156 324 164
rect 364 156 372 164
rect 60 136 68 144
rect 268 136 276 144
rect 284 136 292 144
rect 332 136 340 144
rect 428 136 436 144
rect 492 176 500 184
rect 476 156 484 164
rect 604 276 612 284
rect 668 696 676 704
rect 636 556 644 564
rect 748 736 756 744
rect 732 696 740 704
rect 700 636 708 644
rect 716 616 724 624
rect 732 576 740 584
rect 700 556 708 564
rect 812 816 820 824
rect 876 1116 884 1124
rect 972 1136 980 1144
rect 988 1136 996 1144
rect 956 1116 964 1124
rect 1004 1116 1012 1124
rect 892 1096 900 1104
rect 924 1096 932 1104
rect 940 1096 948 1104
rect 844 1076 852 1084
rect 876 1056 884 1064
rect 844 1036 852 1044
rect 844 976 852 984
rect 1084 1276 1092 1284
rect 1276 1496 1284 1504
rect 1308 1556 1316 1564
rect 1340 1656 1348 1664
rect 1411 1606 1419 1614
rect 1421 1606 1429 1614
rect 1431 1606 1439 1614
rect 1441 1606 1449 1614
rect 1451 1606 1459 1614
rect 1461 1606 1469 1614
rect 1516 1596 1524 1604
rect 1404 1496 1412 1504
rect 1372 1476 1380 1484
rect 1180 1456 1188 1464
rect 1260 1436 1268 1444
rect 1308 1436 1316 1444
rect 1180 1416 1188 1424
rect 1260 1376 1268 1384
rect 1372 1416 1380 1424
rect 1388 1416 1396 1424
rect 1324 1376 1332 1384
rect 1340 1356 1348 1364
rect 1148 1316 1156 1324
rect 1180 1316 1188 1324
rect 1148 1296 1156 1304
rect 1100 1196 1108 1204
rect 1132 1196 1140 1204
rect 988 1056 996 1064
rect 1036 1056 1044 1064
rect 1052 1056 1060 1064
rect 956 996 964 1004
rect 972 996 980 1004
rect 1068 1016 1076 1024
rect 940 956 948 964
rect 1020 956 1028 964
rect 860 936 868 944
rect 860 916 868 924
rect 908 756 916 764
rect 828 736 836 744
rect 908 736 916 744
rect 924 736 932 744
rect 892 696 900 704
rect 780 636 788 644
rect 780 576 788 584
rect 572 256 580 264
rect 620 256 628 264
rect 684 296 692 304
rect 844 656 852 664
rect 892 656 900 664
rect 764 536 772 544
rect 892 536 900 544
rect 1004 796 1012 804
rect 1020 696 1028 704
rect 1036 676 1044 684
rect 1116 1136 1124 1144
rect 1132 1136 1140 1144
rect 1116 1116 1124 1124
rect 1148 1116 1156 1124
rect 1164 1116 1172 1124
rect 1100 976 1108 984
rect 1100 956 1108 964
rect 1084 816 1092 824
rect 1084 696 1092 704
rect 1068 656 1076 664
rect 1052 596 1060 604
rect 1132 1036 1140 1044
rect 1164 1096 1172 1104
rect 1164 956 1172 964
rect 1196 1296 1204 1304
rect 1196 1236 1204 1244
rect 1212 1136 1220 1144
rect 1196 1036 1204 1044
rect 1228 1096 1236 1104
rect 1260 1236 1268 1244
rect 1244 1076 1252 1084
rect 1196 956 1204 964
rect 1292 1216 1300 1224
rect 1340 1156 1348 1164
rect 1500 1376 1508 1384
rect 1420 1356 1428 1364
rect 1548 2016 1556 2024
rect 1676 2736 1684 2744
rect 1692 2696 1700 2704
rect 1740 2696 1748 2704
rect 1724 2676 1732 2684
rect 1724 2576 1732 2584
rect 1740 2576 1748 2584
rect 1740 2516 1748 2524
rect 1708 2456 1716 2464
rect 1724 2456 1732 2464
rect 1692 2436 1700 2444
rect 1660 2376 1668 2384
rect 1644 2276 1652 2284
rect 1628 2236 1636 2244
rect 1612 2176 1620 2184
rect 1676 2236 1684 2244
rect 1820 2996 1828 3004
rect 1772 2956 1780 2964
rect 1836 2936 1844 2944
rect 2044 3296 2052 3304
rect 1900 3216 1908 3224
rect 1884 2936 1892 2944
rect 1820 2856 1828 2864
rect 1836 2856 1844 2864
rect 1772 2836 1780 2844
rect 1804 2776 1812 2784
rect 1788 2716 1796 2724
rect 1788 2696 1796 2704
rect 1836 2736 1844 2744
rect 1820 2716 1828 2724
rect 1820 2696 1828 2704
rect 1820 2656 1828 2664
rect 1804 2636 1812 2644
rect 2428 3796 2436 3804
rect 2524 4156 2532 4164
rect 2556 4216 2564 4224
rect 2604 4496 2612 4504
rect 2668 4496 2676 4504
rect 2620 4436 2628 4444
rect 2604 4216 2612 4224
rect 2588 4176 2596 4184
rect 2540 4136 2548 4144
rect 2556 4136 2564 4144
rect 2572 4136 2580 4144
rect 2492 4116 2500 4124
rect 2588 4096 2596 4104
rect 2476 4056 2484 4064
rect 2652 4336 2660 4344
rect 2636 4296 2644 4304
rect 2652 4176 2660 4184
rect 2652 4116 2660 4124
rect 2844 4716 2852 4724
rect 2924 4716 2932 4724
rect 5923 5406 5931 5414
rect 5933 5406 5941 5414
rect 5943 5406 5951 5414
rect 5953 5406 5961 5414
rect 5963 5406 5971 5414
rect 5973 5406 5981 5414
rect 6012 5396 6020 5404
rect 3804 5376 3812 5384
rect 3996 5376 4004 5384
rect 4284 5376 4292 5384
rect 4604 5376 4612 5384
rect 3676 5356 3684 5364
rect 3756 5356 3764 5364
rect 3884 5356 3892 5364
rect 3996 5356 4004 5364
rect 3212 5336 3220 5344
rect 3228 5336 3236 5344
rect 3324 5336 3332 5344
rect 3516 5336 3524 5344
rect 3212 5296 3220 5304
rect 3196 5236 3204 5244
rect 3100 5216 3108 5224
rect 3180 5176 3188 5184
rect 3164 5136 3172 5144
rect 3116 5116 3124 5124
rect 3100 5096 3108 5104
rect 3148 5096 3156 5104
rect 3180 5116 3188 5124
rect 3212 5176 3220 5184
rect 3292 5136 3300 5144
rect 3196 5096 3204 5104
rect 3148 5056 3156 5064
rect 3244 5076 3252 5084
rect 3276 5076 3284 5084
rect 3564 5316 3572 5324
rect 3692 5296 3700 5304
rect 3372 5276 3380 5284
rect 3404 5196 3412 5204
rect 3724 5316 3732 5324
rect 3708 5216 3716 5224
rect 3788 5216 3796 5224
rect 5276 5356 5284 5364
rect 3932 5336 3940 5344
rect 4028 5336 4036 5344
rect 4092 5336 4100 5344
rect 4348 5336 4356 5344
rect 4812 5336 4820 5344
rect 4908 5336 4916 5344
rect 5100 5336 5108 5344
rect 5132 5336 5140 5344
rect 5180 5336 5188 5344
rect 5212 5336 5220 5344
rect 3964 5316 3972 5324
rect 4108 5316 4116 5324
rect 4028 5296 4036 5304
rect 4076 5296 4084 5304
rect 4092 5276 4100 5284
rect 4108 5276 4116 5284
rect 3916 5216 3924 5224
rect 3884 5196 3892 5204
rect 3484 5156 3492 5164
rect 3548 5156 3556 5164
rect 3356 5116 3364 5124
rect 3340 5096 3348 5104
rect 3388 5096 3396 5104
rect 3436 5096 3444 5104
rect 3452 5096 3460 5104
rect 3180 4976 3188 4984
rect 3116 4956 3124 4964
rect 3164 4956 3172 4964
rect 3148 4936 3156 4944
rect 3164 4936 3172 4944
rect 3244 4936 3252 4944
rect 3068 4896 3076 4904
rect 3100 4916 3108 4924
rect 3084 4876 3092 4884
rect 3020 4856 3028 4864
rect 3052 4856 3060 4864
rect 3036 4776 3044 4784
rect 2812 4696 2820 4704
rect 2940 4696 2948 4704
rect 2908 4676 2916 4684
rect 2844 4656 2852 4664
rect 2860 4636 2868 4644
rect 2780 4596 2788 4604
rect 2812 4596 2820 4604
rect 2915 4606 2923 4614
rect 2925 4606 2933 4614
rect 2935 4606 2943 4614
rect 2945 4606 2953 4614
rect 2955 4606 2963 4614
rect 2965 4606 2973 4614
rect 2764 4516 2772 4524
rect 2716 4476 2724 4484
rect 2748 4236 2756 4244
rect 2796 4436 2804 4444
rect 2780 4336 2788 4344
rect 2812 4296 2820 4304
rect 2716 4136 2724 4144
rect 3052 4456 3060 4464
rect 3036 4296 3044 4304
rect 2860 4276 2868 4284
rect 3068 4276 3076 4284
rect 3036 4256 3044 4264
rect 2915 4206 2923 4214
rect 2925 4206 2933 4214
rect 2935 4206 2943 4214
rect 2945 4206 2953 4214
rect 2955 4206 2963 4214
rect 2965 4206 2973 4214
rect 2876 4176 2884 4184
rect 2780 4136 2788 4144
rect 2860 4136 2868 4144
rect 2892 4156 2900 4164
rect 2908 4136 2916 4144
rect 2764 4116 2772 4124
rect 2636 4096 2644 4104
rect 2684 4096 2692 4104
rect 2492 3976 2500 3984
rect 2620 3976 2628 3984
rect 2588 3956 2596 3964
rect 2700 4036 2708 4044
rect 2652 3956 2660 3964
rect 2572 3876 2580 3884
rect 2620 3856 2628 3864
rect 2636 3836 2644 3844
rect 2460 3796 2468 3804
rect 2684 3936 2692 3944
rect 2668 3896 2676 3904
rect 3180 4916 3188 4924
rect 3164 4702 3172 4704
rect 3164 4696 3172 4702
rect 3228 4696 3236 4704
rect 3260 4916 3268 4924
rect 3228 4656 3236 4664
rect 3324 5056 3332 5064
rect 3468 5076 3476 5084
rect 3436 5056 3444 5064
rect 3484 5056 3492 5064
rect 3500 5056 3508 5064
rect 3436 4956 3444 4964
rect 3452 4956 3460 4964
rect 3484 4956 3492 4964
rect 3356 4936 3364 4944
rect 3388 4916 3396 4924
rect 3404 4916 3412 4924
rect 3372 4896 3380 4904
rect 3420 4836 3428 4844
rect 3436 4836 3444 4844
rect 3372 4816 3380 4824
rect 3356 4716 3364 4724
rect 3276 4616 3284 4624
rect 3324 4576 3332 4584
rect 3468 4916 3476 4924
rect 3628 5136 3636 5144
rect 3532 4916 3540 4924
rect 3500 4876 3508 4884
rect 3580 4876 3588 4884
rect 3548 4856 3556 4864
rect 3660 5116 3668 5124
rect 3708 5116 3716 5124
rect 3804 5116 3812 5124
rect 3644 5076 3652 5084
rect 3724 5096 3732 5104
rect 3820 5076 3828 5084
rect 3612 5056 3620 5064
rect 3644 5036 3652 5044
rect 3660 5036 3668 5044
rect 3692 5056 3700 5064
rect 3740 5056 3748 5064
rect 3788 5056 3796 5064
rect 3724 5036 3732 5044
rect 3756 5036 3764 5044
rect 3852 5016 3860 5024
rect 3868 5016 3876 5024
rect 3660 4976 3668 4984
rect 3628 4956 3636 4964
rect 3644 4956 3652 4964
rect 3612 4936 3620 4944
rect 3724 4956 3732 4964
rect 3740 4956 3748 4964
rect 3900 4976 3908 4984
rect 3676 4916 3684 4924
rect 3708 4916 3716 4924
rect 3756 4916 3764 4924
rect 3644 4896 3652 4904
rect 3692 4896 3700 4904
rect 3596 4776 3604 4784
rect 3612 4736 3620 4744
rect 3660 4736 3668 4744
rect 3628 4716 3636 4724
rect 3564 4696 3572 4704
rect 3500 4676 3508 4684
rect 3484 4656 3492 4664
rect 3468 4636 3476 4644
rect 3452 4596 3460 4604
rect 3676 4716 3684 4724
rect 3708 4856 3716 4864
rect 3708 4816 3716 4824
rect 3692 4676 3700 4684
rect 3660 4656 3668 4664
rect 3580 4636 3588 4644
rect 3676 4596 3684 4604
rect 3580 4576 3588 4584
rect 3564 4556 3572 4564
rect 3676 4556 3684 4564
rect 3212 4536 3220 4544
rect 3308 4536 3316 4544
rect 3516 4536 3524 4544
rect 3276 4516 3284 4524
rect 3356 4516 3364 4524
rect 3148 4276 3156 4284
rect 3084 4156 3092 4164
rect 3292 4496 3300 4504
rect 3356 4496 3364 4504
rect 3164 4256 3172 4264
rect 3244 4236 3252 4244
rect 3180 4216 3188 4224
rect 3228 4216 3236 4224
rect 3276 4216 3284 4224
rect 3164 4156 3172 4164
rect 3052 4136 3060 4144
rect 3196 4116 3204 4124
rect 2812 4096 2820 4104
rect 2988 4096 2996 4104
rect 3068 4096 3076 4104
rect 3116 3976 3124 3984
rect 2748 3916 2756 3924
rect 2732 3896 2740 3904
rect 2780 3896 2788 3904
rect 2876 3896 2884 3904
rect 2892 3896 2900 3904
rect 3116 3896 3124 3904
rect 2620 3736 2628 3744
rect 2588 3718 2596 3724
rect 2588 3716 2596 3718
rect 2540 3696 2548 3704
rect 2380 3656 2388 3664
rect 2412 3656 2420 3664
rect 2524 3656 2532 3664
rect 2300 3596 2308 3604
rect 2252 3576 2260 3584
rect 2252 3556 2260 3564
rect 2284 3536 2292 3544
rect 2220 3476 2228 3484
rect 2236 3476 2244 3484
rect 2332 3516 2340 3524
rect 2300 3476 2308 3484
rect 2268 3456 2276 3464
rect 2252 3436 2260 3444
rect 2220 3316 2228 3324
rect 2188 3236 2196 3244
rect 2124 3176 2132 3184
rect 2156 3156 2164 3164
rect 2060 3136 2068 3144
rect 2156 3136 2164 3144
rect 1932 3116 1940 3124
rect 1980 3116 1988 3124
rect 1980 3056 1988 3064
rect 1932 2996 1940 3004
rect 1964 2996 1972 3004
rect 1932 2956 1940 2964
rect 1948 2936 1956 2944
rect 2092 3116 2100 3124
rect 2076 3056 2084 3064
rect 2060 3016 2068 3024
rect 1964 2856 1972 2864
rect 1900 2836 1908 2844
rect 1900 2736 1908 2744
rect 1884 2696 1892 2704
rect 2028 2936 2036 2944
rect 1996 2836 2004 2844
rect 1980 2796 1988 2804
rect 1932 2736 1940 2744
rect 1948 2696 1956 2704
rect 1852 2676 1860 2684
rect 1868 2676 1876 2684
rect 1916 2676 1924 2684
rect 1932 2676 1940 2684
rect 1836 2636 1844 2644
rect 1884 2556 1892 2564
rect 1772 2536 1780 2544
rect 1772 2516 1780 2524
rect 1788 2476 1796 2484
rect 1836 2476 1844 2484
rect 1852 2476 1860 2484
rect 1788 2396 1796 2404
rect 1772 2376 1780 2384
rect 1756 2336 1764 2344
rect 1724 2236 1732 2244
rect 1740 2236 1748 2244
rect 1548 1956 1556 1964
rect 1580 1936 1588 1944
rect 1596 1916 1604 1924
rect 1644 2076 1652 2084
rect 1660 2016 1668 2024
rect 1660 1936 1668 1944
rect 1692 2116 1700 2124
rect 1708 2016 1716 2024
rect 1692 1976 1700 1984
rect 1724 1976 1732 1984
rect 1708 1956 1716 1964
rect 1868 2416 1876 2424
rect 1916 2416 1924 2424
rect 1852 2396 1860 2404
rect 1948 2656 1956 2664
rect 1980 2696 1988 2704
rect 2220 3116 2228 3124
rect 2140 3056 2148 3064
rect 2108 3036 2116 3044
rect 2188 3036 2196 3044
rect 2156 2956 2164 2964
rect 2092 2916 2100 2924
rect 2060 2756 2068 2764
rect 2076 2736 2084 2744
rect 2012 2696 2020 2704
rect 2044 2676 2052 2684
rect 1996 2576 2004 2584
rect 2044 2576 2052 2584
rect 1964 2556 1972 2564
rect 1996 2536 2004 2544
rect 1980 2516 1988 2524
rect 2028 2516 2036 2524
rect 2060 2516 2068 2524
rect 1948 2476 1956 2484
rect 2044 2436 2052 2444
rect 1948 2416 1956 2424
rect 1804 2356 1812 2364
rect 1820 2336 1828 2344
rect 1932 2336 1940 2344
rect 2012 2336 2020 2344
rect 1820 2296 1828 2304
rect 1884 2296 1892 2304
rect 1820 2256 1828 2264
rect 1868 2256 1876 2264
rect 1916 2256 1924 2264
rect 1820 2236 1828 2244
rect 1788 2136 1796 2144
rect 1756 2016 1764 2024
rect 1628 1916 1636 1924
rect 1676 1916 1684 1924
rect 1692 1916 1700 1924
rect 1548 1856 1556 1864
rect 1612 1896 1620 1904
rect 1660 1896 1668 1904
rect 1596 1796 1604 1804
rect 1564 1756 1572 1764
rect 1548 1736 1556 1744
rect 1612 1736 1620 1744
rect 1644 1876 1652 1884
rect 1644 1776 1652 1784
rect 1628 1716 1636 1724
rect 1628 1696 1636 1704
rect 1628 1636 1636 1644
rect 1564 1556 1572 1564
rect 1596 1536 1604 1544
rect 1532 1516 1540 1524
rect 1756 1936 1764 1944
rect 1788 1916 1796 1924
rect 1804 1896 1812 1904
rect 1836 2196 1844 2204
rect 1900 2236 1908 2244
rect 1916 2236 1924 2244
rect 1884 2196 1892 2204
rect 1916 2156 1924 2164
rect 1852 2116 1860 2124
rect 1852 2096 1860 2104
rect 1836 1936 1844 1944
rect 1852 1936 1860 1944
rect 1836 1896 1844 1904
rect 1724 1816 1732 1824
rect 1692 1736 1700 1744
rect 1708 1736 1716 1744
rect 1692 1676 1700 1684
rect 1772 1856 1780 1864
rect 1756 1736 1764 1744
rect 1756 1676 1764 1684
rect 1564 1496 1572 1504
rect 1676 1496 1684 1504
rect 1740 1616 1748 1624
rect 1724 1516 1732 1524
rect 1580 1476 1588 1484
rect 1644 1476 1652 1484
rect 1708 1476 1716 1484
rect 1532 1456 1540 1464
rect 1596 1456 1604 1464
rect 1644 1456 1652 1464
rect 1548 1356 1556 1364
rect 1628 1336 1636 1344
rect 1484 1296 1492 1304
rect 1404 1236 1412 1244
rect 1411 1206 1419 1214
rect 1421 1206 1429 1214
rect 1431 1206 1439 1214
rect 1441 1206 1449 1214
rect 1451 1206 1459 1214
rect 1461 1206 1469 1214
rect 1612 1316 1620 1324
rect 1564 1236 1572 1244
rect 1388 1196 1396 1204
rect 1484 1196 1492 1204
rect 1580 1176 1588 1184
rect 1500 1156 1508 1164
rect 1516 1156 1524 1164
rect 1516 1116 1524 1124
rect 1532 1116 1540 1124
rect 1628 1216 1636 1224
rect 1692 1356 1700 1364
rect 1708 1356 1716 1364
rect 1676 1336 1684 1344
rect 1708 1336 1716 1344
rect 1660 1316 1668 1324
rect 1644 1136 1652 1144
rect 1292 1096 1300 1104
rect 1388 1096 1396 1104
rect 1484 1096 1492 1104
rect 1564 1096 1572 1104
rect 1612 1096 1620 1104
rect 1596 1076 1604 1084
rect 1388 1056 1396 1064
rect 1532 1056 1540 1064
rect 1612 1056 1620 1064
rect 1340 1036 1348 1044
rect 1292 1016 1300 1024
rect 1260 996 1268 1004
rect 1276 956 1284 964
rect 1324 996 1332 1004
rect 1372 976 1380 984
rect 1548 996 1556 1004
rect 1564 996 1572 1004
rect 1612 976 1620 984
rect 1500 956 1508 964
rect 1548 956 1556 964
rect 1580 956 1588 964
rect 1484 936 1492 944
rect 1564 936 1572 944
rect 1596 936 1604 944
rect 1228 916 1236 924
rect 1292 916 1300 924
rect 1308 916 1316 924
rect 1356 916 1364 924
rect 1468 916 1476 924
rect 1628 936 1636 944
rect 1132 756 1140 764
rect 1180 756 1188 764
rect 1148 736 1156 744
rect 1164 716 1172 724
rect 1212 796 1220 804
rect 1260 736 1268 744
rect 1212 716 1220 724
rect 1148 696 1156 704
rect 1196 696 1204 704
rect 1244 696 1252 704
rect 1116 656 1124 664
rect 1132 656 1140 664
rect 1132 596 1140 604
rect 924 556 932 564
rect 1100 556 1108 564
rect 796 516 804 524
rect 780 376 788 384
rect 908 436 916 444
rect 908 376 916 384
rect 700 276 708 284
rect 828 276 836 284
rect 860 276 868 284
rect 796 256 804 264
rect 828 256 836 264
rect 876 256 884 264
rect 604 236 612 244
rect 652 236 660 244
rect 556 216 564 224
rect 572 176 580 184
rect 524 136 532 144
rect 780 196 788 204
rect 700 176 708 184
rect 620 156 628 164
rect 636 156 644 164
rect 764 156 772 164
rect 892 176 900 184
rect 940 536 948 544
rect 1004 536 1012 544
rect 940 516 948 524
rect 1356 896 1364 904
rect 1532 896 1540 904
rect 1468 876 1476 884
rect 1516 876 1524 884
rect 1484 816 1492 824
rect 1411 806 1419 814
rect 1421 806 1429 814
rect 1431 806 1439 814
rect 1441 806 1449 814
rect 1451 806 1459 814
rect 1461 806 1469 814
rect 1308 696 1316 704
rect 1420 696 1428 704
rect 1180 656 1188 664
rect 1132 536 1140 544
rect 1084 516 1092 524
rect 1036 476 1044 484
rect 1132 476 1140 484
rect 1004 436 1012 444
rect 988 356 996 364
rect 1020 336 1028 344
rect 1084 336 1092 344
rect 1004 316 1012 324
rect 940 296 948 304
rect 1052 296 1060 304
rect 956 256 964 264
rect 988 256 996 264
rect 1036 256 1044 264
rect 1068 256 1076 264
rect 1116 256 1124 264
rect 988 236 996 244
rect 940 216 948 224
rect 972 216 980 224
rect 940 176 948 184
rect 1036 196 1044 204
rect 1148 356 1156 364
rect 1356 656 1364 664
rect 1340 636 1348 644
rect 1324 616 1332 624
rect 1292 556 1300 564
rect 1196 536 1204 544
rect 1228 516 1236 524
rect 1244 496 1252 504
rect 1292 496 1300 504
rect 1212 476 1220 484
rect 1196 436 1204 444
rect 1260 376 1268 384
rect 1340 596 1348 604
rect 1340 536 1348 544
rect 1340 516 1348 524
rect 1436 636 1444 644
rect 1372 556 1380 564
rect 1436 536 1444 544
rect 1372 516 1380 524
rect 1500 736 1508 744
rect 1516 696 1524 704
rect 1548 656 1556 664
rect 1468 596 1476 604
rect 1564 616 1572 624
rect 1516 536 1524 544
rect 1500 516 1508 524
rect 1564 516 1572 524
rect 1548 496 1556 504
rect 1484 476 1492 484
rect 1484 416 1492 424
rect 1411 406 1419 414
rect 1421 406 1429 414
rect 1431 406 1439 414
rect 1441 406 1449 414
rect 1451 406 1459 414
rect 1461 406 1469 414
rect 1436 336 1444 344
rect 1420 316 1428 324
rect 1388 296 1396 304
rect 1164 236 1172 244
rect 1196 176 1204 184
rect 1228 156 1236 164
rect 1292 276 1300 284
rect 1324 256 1332 264
rect 1388 276 1396 284
rect 1372 156 1380 164
rect 620 116 628 124
rect 668 116 676 124
rect 1052 136 1060 144
rect 1100 136 1108 144
rect 1244 136 1252 144
rect 716 116 724 124
rect 1132 116 1140 124
rect 1276 116 1284 124
rect 1388 136 1396 144
rect 1596 596 1604 604
rect 1692 1116 1700 1124
rect 1772 1556 1780 1564
rect 1756 1496 1764 1504
rect 1836 1856 1844 1864
rect 1836 1736 1844 1744
rect 1820 1676 1828 1684
rect 1804 1616 1812 1624
rect 1916 2116 1924 2124
rect 1916 2076 1924 2084
rect 1868 1876 1876 1884
rect 1916 1856 1924 1864
rect 1868 1776 1876 1784
rect 2060 2376 2068 2384
rect 2076 2356 2084 2364
rect 2044 2316 2052 2324
rect 1964 2296 1972 2304
rect 2012 2296 2020 2304
rect 2076 2296 2084 2304
rect 2028 2276 2036 2284
rect 1948 2236 1956 2244
rect 2012 2256 2020 2264
rect 1948 2176 1956 2184
rect 1964 2176 1972 2184
rect 1980 2136 1988 2144
rect 2044 2176 2052 2184
rect 2028 2156 2036 2164
rect 1996 2116 2004 2124
rect 2108 2876 2116 2884
rect 2204 3016 2212 3024
rect 2252 3376 2260 3384
rect 2236 2996 2244 3004
rect 2220 2956 2228 2964
rect 2284 3316 2292 3324
rect 2316 3456 2324 3464
rect 2300 3176 2308 3184
rect 2332 3156 2340 3164
rect 2460 3536 2468 3544
rect 2412 3496 2420 3504
rect 2636 3636 2644 3644
rect 2668 3576 2676 3584
rect 2636 3516 2644 3524
rect 2508 3476 2516 3484
rect 2508 3456 2516 3464
rect 2412 3436 2420 3444
rect 2396 3376 2404 3384
rect 2588 3396 2596 3404
rect 2572 3336 2580 3344
rect 2620 3376 2628 3384
rect 2604 3356 2612 3364
rect 2380 3316 2388 3324
rect 2364 3236 2372 3244
rect 2348 3076 2356 3084
rect 2300 2996 2308 3004
rect 2268 2936 2276 2944
rect 2284 2936 2292 2944
rect 2108 2736 2116 2744
rect 2124 2696 2132 2704
rect 2124 2516 2132 2524
rect 2252 2896 2260 2904
rect 2172 2876 2180 2884
rect 2236 2856 2244 2864
rect 2332 2976 2340 2984
rect 2460 3316 2468 3324
rect 2412 3176 2420 3184
rect 2524 3316 2532 3324
rect 2380 3116 2388 3124
rect 2444 3116 2452 3124
rect 2380 3096 2388 3104
rect 2572 3196 2580 3204
rect 2588 3176 2596 3184
rect 2524 3096 2532 3104
rect 2668 3476 2676 3484
rect 2700 3836 2708 3844
rect 2716 3716 2724 3724
rect 2764 3856 2772 3864
rect 2812 3756 2820 3764
rect 2844 3756 2852 3764
rect 3164 3976 3172 3984
rect 3132 3876 3140 3884
rect 3164 3876 3172 3884
rect 3020 3856 3028 3864
rect 2915 3806 2923 3814
rect 2925 3806 2933 3814
rect 2935 3806 2943 3814
rect 2945 3806 2953 3814
rect 2955 3806 2963 3814
rect 2965 3806 2973 3814
rect 3148 3776 3156 3784
rect 2812 3736 2820 3744
rect 2892 3736 2900 3744
rect 2780 3718 2788 3724
rect 2780 3716 2788 3718
rect 2844 3716 2852 3724
rect 2844 3696 2852 3704
rect 2748 3656 2756 3664
rect 2796 3576 2804 3584
rect 2700 3556 2708 3564
rect 2892 3716 2900 3724
rect 3020 3716 3028 3724
rect 2892 3676 2900 3684
rect 2732 3436 2740 3444
rect 2876 3436 2884 3444
rect 2780 3416 2788 3424
rect 2764 3376 2772 3384
rect 2684 3336 2692 3344
rect 2620 3256 2628 3264
rect 2684 3256 2692 3264
rect 2620 3136 2628 3144
rect 2668 3116 2676 3124
rect 2604 3096 2612 3104
rect 2668 3096 2676 3104
rect 2620 3076 2628 3084
rect 2396 3036 2404 3044
rect 2380 3016 2388 3024
rect 2460 2956 2468 2964
rect 2460 2936 2468 2944
rect 2316 2896 2324 2904
rect 2364 2896 2372 2904
rect 2268 2856 2276 2864
rect 2284 2856 2292 2864
rect 2348 2856 2356 2864
rect 2396 2856 2404 2864
rect 2284 2796 2292 2804
rect 2172 2736 2180 2744
rect 2236 2736 2244 2744
rect 2204 2716 2212 2724
rect 2556 3036 2564 3044
rect 2572 2976 2580 2984
rect 2508 2916 2516 2924
rect 2460 2896 2468 2904
rect 2572 2876 2580 2884
rect 2652 3056 2660 3064
rect 2796 3196 2804 3204
rect 2716 3176 2724 3184
rect 2764 3176 2772 3184
rect 2764 3136 2772 3144
rect 2780 3136 2788 3144
rect 2732 3076 2740 3084
rect 2732 2976 2740 2984
rect 2828 3116 2836 3124
rect 2796 3076 2804 3084
rect 2828 3056 2836 3064
rect 2812 3036 2820 3044
rect 2652 2940 2660 2944
rect 2652 2936 2660 2940
rect 2780 2936 2788 2944
rect 2828 2976 2836 2984
rect 2915 3406 2923 3414
rect 2925 3406 2933 3414
rect 2935 3406 2943 3414
rect 2945 3406 2953 3414
rect 2955 3406 2963 3414
rect 2965 3406 2973 3414
rect 2908 3376 2916 3384
rect 2940 3336 2948 3344
rect 2988 3336 2996 3344
rect 3036 3696 3044 3704
rect 3020 3296 3028 3304
rect 3180 3716 3188 3724
rect 3180 3696 3188 3704
rect 3260 3776 3268 3784
rect 3452 4518 3460 4524
rect 3452 4516 3460 4518
rect 3628 4516 3636 4524
rect 3548 4456 3556 4464
rect 3388 4396 3396 4404
rect 3372 4316 3380 4324
rect 3468 4316 3476 4324
rect 3404 4256 3412 4264
rect 3356 4176 3364 4184
rect 3452 4276 3460 4284
rect 3500 4236 3508 4244
rect 3468 4176 3476 4184
rect 3436 4156 3444 4164
rect 3324 4136 3332 4144
rect 3420 4136 3428 4144
rect 3436 4136 3444 4144
rect 3388 4116 3396 4124
rect 3484 4156 3492 4164
rect 3436 4096 3444 4104
rect 3372 3896 3380 3904
rect 3404 3896 3412 3904
rect 3404 3776 3412 3784
rect 3276 3736 3284 3744
rect 3228 3716 3236 3724
rect 3180 3496 3188 3504
rect 3180 3436 3188 3444
rect 3148 3376 3156 3384
rect 3084 3356 3092 3364
rect 3260 3596 3268 3604
rect 3276 3596 3284 3604
rect 3228 3396 3236 3404
rect 3116 3316 3124 3324
rect 3164 3316 3172 3324
rect 3052 3216 3060 3224
rect 3436 4076 3444 4084
rect 3484 4056 3492 4064
rect 3500 4016 3508 4024
rect 3580 4316 3588 4324
rect 3628 4356 3636 4364
rect 3660 4496 3668 4504
rect 3644 4316 3652 4324
rect 3596 4276 3604 4284
rect 3660 4296 3668 4304
rect 3612 4236 3620 4244
rect 3612 4136 3620 4144
rect 3564 4116 3572 4124
rect 3596 4116 3604 4124
rect 3724 4636 3732 4644
rect 3708 4556 3716 4564
rect 3708 4536 3716 4544
rect 3820 4896 3828 4904
rect 3772 4816 3780 4824
rect 3804 4776 3812 4784
rect 3868 4896 3876 4904
rect 3852 4876 3860 4884
rect 3836 4696 3844 4704
rect 3820 4676 3828 4684
rect 3836 4656 3844 4664
rect 3772 4636 3780 4644
rect 3836 4616 3844 4624
rect 3884 4616 3892 4624
rect 4044 5196 4052 5204
rect 3932 5096 3940 5104
rect 4012 5096 4020 5104
rect 4028 5096 4036 5104
rect 3932 5076 3940 5084
rect 3964 5076 3972 5084
rect 3980 5056 3988 5064
rect 4028 5076 4036 5084
rect 3996 5036 4004 5044
rect 4028 5016 4036 5024
rect 3932 4956 3940 4964
rect 3996 4956 4004 4964
rect 3964 4916 3972 4924
rect 3980 4876 3988 4884
rect 3964 4856 3972 4864
rect 3932 4836 3940 4844
rect 3916 4696 3924 4704
rect 3980 4836 3988 4844
rect 3980 4716 3988 4724
rect 3964 4696 3972 4704
rect 4316 5316 4324 5324
rect 4252 5296 4260 5304
rect 4396 5296 4404 5304
rect 4236 5256 4244 5264
rect 4236 5236 4244 5244
rect 4236 5196 4244 5204
rect 4300 5176 4308 5184
rect 4140 5156 4148 5164
rect 4156 5156 4164 5164
rect 4284 5156 4292 5164
rect 4204 5136 4212 5144
rect 4220 5136 4228 5144
rect 4156 5116 4164 5124
rect 4172 5096 4180 5104
rect 4092 5076 4100 5084
rect 4060 5056 4068 5064
rect 4060 4936 4068 4944
rect 4108 5056 4116 5064
rect 4188 5056 4196 5064
rect 4236 5116 4244 5124
rect 4268 5116 4276 5124
rect 4236 5096 4244 5104
rect 4300 5076 4308 5084
rect 4252 5056 4260 5064
rect 4284 5056 4292 5064
rect 4236 5016 4244 5024
rect 4092 4876 4100 4884
rect 4076 4836 4084 4844
rect 4044 4816 4052 4824
rect 4060 4816 4068 4824
rect 4124 4916 4132 4924
rect 4140 4896 4148 4904
rect 4172 4916 4180 4924
rect 4204 4916 4212 4924
rect 4220 4896 4228 4904
rect 4156 4876 4164 4884
rect 4124 4836 4132 4844
rect 4364 5036 4372 5044
rect 4332 4976 4340 4984
rect 4348 4976 4356 4984
rect 4316 4956 4324 4964
rect 4252 4916 4260 4924
rect 4236 4816 4244 4824
rect 4044 4756 4052 4764
rect 4172 4756 4180 4764
rect 4012 4716 4020 4724
rect 4060 4716 4068 4724
rect 4060 4696 4068 4704
rect 3996 4676 4004 4684
rect 4188 4696 4196 4704
rect 4204 4696 4212 4704
rect 3932 4616 3940 4624
rect 3852 4596 3860 4604
rect 3900 4596 3908 4604
rect 3772 4536 3780 4544
rect 3804 4536 3812 4544
rect 3756 4376 3764 4384
rect 3756 4356 3764 4364
rect 3724 4316 3732 4324
rect 3788 4376 3796 4384
rect 3772 4316 3780 4324
rect 3804 4356 3812 4364
rect 3916 4336 3924 4344
rect 3772 4296 3780 4304
rect 3708 4276 3716 4284
rect 3788 4276 3796 4284
rect 3692 4236 3700 4244
rect 3740 4236 3748 4244
rect 3692 4176 3700 4184
rect 3820 4196 3828 4204
rect 3804 4136 3812 4144
rect 3756 4116 3764 4124
rect 3644 4096 3652 4104
rect 3564 4016 3572 4024
rect 3612 4016 3620 4024
rect 3724 4076 3732 4084
rect 3788 4076 3796 4084
rect 3772 4036 3780 4044
rect 3676 3996 3684 4004
rect 3484 3896 3492 3904
rect 3452 3876 3460 3884
rect 3452 3736 3460 3744
rect 3548 3876 3556 3884
rect 3500 3776 3508 3784
rect 3548 3776 3556 3784
rect 3532 3756 3540 3764
rect 3548 3736 3556 3744
rect 3644 3896 3652 3904
rect 3580 3856 3588 3864
rect 3628 3856 3636 3864
rect 3644 3856 3652 3864
rect 3612 3796 3620 3804
rect 3420 3716 3428 3724
rect 3468 3716 3476 3724
rect 3580 3716 3588 3724
rect 3500 3676 3508 3684
rect 3564 3676 3572 3684
rect 3292 3576 3300 3584
rect 3324 3576 3332 3584
rect 3340 3576 3348 3584
rect 3372 3576 3380 3584
rect 3468 3536 3476 3544
rect 3436 3516 3444 3524
rect 3564 3616 3572 3624
rect 3548 3556 3556 3564
rect 3532 3516 3540 3524
rect 3340 3496 3348 3504
rect 3452 3496 3460 3504
rect 3484 3496 3492 3504
rect 3308 3436 3316 3444
rect 3292 3416 3300 3424
rect 3404 3416 3412 3424
rect 3484 3476 3492 3484
rect 3660 3796 3668 3804
rect 3660 3756 3668 3764
rect 3628 3736 3636 3744
rect 3612 3616 3620 3624
rect 3596 3556 3604 3564
rect 3612 3536 3620 3544
rect 3596 3516 3604 3524
rect 3580 3496 3588 3504
rect 3660 3636 3668 3644
rect 3660 3536 3668 3544
rect 3644 3516 3652 3524
rect 3452 3356 3460 3364
rect 3516 3456 3524 3464
rect 3612 3456 3620 3464
rect 3724 3916 3732 3924
rect 3740 3896 3748 3904
rect 3772 3896 3780 3904
rect 3692 3876 3700 3884
rect 3724 3776 3732 3784
rect 3740 3776 3748 3784
rect 3708 3736 3716 3744
rect 3708 3676 3716 3684
rect 3708 3556 3716 3564
rect 3692 3536 3700 3544
rect 3676 3496 3684 3504
rect 3724 3516 3732 3524
rect 3756 3696 3764 3704
rect 3900 4296 3908 4304
rect 3916 4296 3924 4304
rect 3884 4276 3892 4284
rect 3836 4056 3844 4064
rect 3820 3956 3828 3964
rect 3804 3816 3812 3824
rect 3948 4136 3956 4144
rect 3980 4196 3988 4204
rect 3964 4116 3972 4124
rect 3884 3976 3892 3984
rect 3852 3916 3860 3924
rect 3836 3876 3844 3884
rect 3836 3776 3844 3784
rect 3820 3756 3828 3764
rect 3804 3696 3812 3704
rect 3820 3696 3828 3704
rect 3804 3676 3812 3684
rect 3788 3656 3796 3664
rect 3820 3616 3828 3624
rect 3772 3536 3780 3544
rect 3500 3356 3508 3364
rect 3164 3176 3172 3184
rect 2924 3116 2932 3124
rect 3452 3276 3460 3284
rect 3276 3116 3284 3124
rect 3436 3196 3444 3204
rect 3212 3096 3220 3104
rect 3260 3096 3268 3104
rect 3372 3096 3380 3104
rect 2892 3076 2900 3084
rect 2972 3076 2980 3084
rect 2988 3076 2996 3084
rect 3068 3076 3076 3084
rect 3180 3076 3188 3084
rect 3244 3076 3252 3084
rect 3196 3056 3204 3064
rect 3276 3056 3284 3064
rect 3132 3036 3140 3044
rect 3260 3036 3268 3044
rect 2915 3006 2923 3014
rect 2925 3006 2933 3014
rect 2935 3006 2943 3014
rect 2945 3006 2953 3014
rect 2955 3006 2963 3014
rect 2965 3006 2973 3014
rect 2876 2916 2884 2924
rect 2828 2816 2836 2824
rect 2444 2756 2452 2764
rect 2588 2756 2596 2764
rect 2812 2736 2820 2744
rect 2348 2716 2356 2724
rect 2188 2696 2196 2704
rect 2252 2696 2260 2704
rect 2364 2696 2372 2704
rect 2476 2696 2484 2704
rect 2284 2656 2292 2664
rect 2252 2556 2260 2564
rect 2188 2516 2196 2524
rect 2348 2576 2356 2584
rect 2332 2556 2340 2564
rect 2220 2516 2228 2524
rect 2268 2496 2276 2504
rect 2220 2476 2228 2484
rect 2108 2456 2116 2464
rect 2092 2276 2100 2284
rect 2076 2256 2084 2264
rect 2124 2396 2132 2404
rect 2172 2336 2180 2344
rect 2156 2316 2164 2324
rect 2140 2296 2148 2304
rect 2108 2176 2116 2184
rect 2060 2156 2068 2164
rect 2236 2416 2244 2424
rect 2220 2396 2228 2404
rect 2204 2256 2212 2264
rect 2172 2156 2180 2164
rect 2156 2136 2164 2144
rect 2028 2096 2036 2104
rect 2140 2096 2148 2104
rect 2012 2016 2020 2024
rect 2236 2236 2244 2244
rect 2316 2496 2324 2504
rect 2300 2456 2308 2464
rect 2300 2416 2308 2424
rect 2412 2636 2420 2644
rect 2492 2656 2500 2664
rect 2540 2716 2548 2724
rect 2524 2696 2532 2704
rect 2556 2696 2564 2704
rect 2604 2696 2612 2704
rect 2716 2676 2724 2684
rect 2828 2676 2836 2684
rect 2556 2656 2564 2664
rect 2700 2656 2708 2664
rect 2700 2616 2708 2624
rect 2508 2596 2516 2604
rect 2684 2596 2692 2604
rect 2428 2576 2436 2584
rect 2476 2576 2484 2584
rect 2604 2576 2612 2584
rect 2668 2576 2676 2584
rect 2716 2576 2724 2584
rect 2412 2556 2420 2564
rect 2780 2576 2788 2584
rect 2844 2576 2852 2584
rect 2876 2556 2884 2564
rect 2540 2536 2548 2544
rect 2636 2536 2644 2544
rect 2652 2536 2660 2544
rect 2684 2536 2692 2544
rect 2748 2536 2756 2544
rect 2876 2536 2884 2544
rect 2364 2516 2372 2524
rect 2428 2516 2436 2524
rect 2348 2496 2356 2504
rect 2380 2496 2388 2504
rect 2524 2496 2532 2504
rect 2348 2476 2356 2484
rect 2268 2316 2276 2324
rect 2300 2316 2308 2324
rect 2252 2176 2260 2184
rect 2220 2156 2228 2164
rect 2204 2136 2212 2144
rect 2220 2076 2228 2084
rect 2092 2056 2100 2064
rect 2108 2056 2116 2064
rect 2188 2056 2196 2064
rect 1964 1916 1972 1924
rect 2012 1916 2020 1924
rect 2108 2036 2116 2044
rect 2364 2356 2372 2364
rect 2332 2276 2340 2284
rect 2316 2216 2324 2224
rect 2300 2136 2308 2144
rect 2348 2256 2356 2264
rect 2348 2236 2356 2244
rect 2348 2176 2356 2184
rect 2284 2096 2292 2104
rect 2188 1936 2196 1944
rect 2044 1896 2052 1904
rect 2076 1896 2084 1904
rect 1996 1856 2004 1864
rect 2060 1856 2068 1864
rect 2012 1836 2020 1844
rect 1964 1816 1972 1824
rect 1948 1796 1956 1804
rect 1932 1756 1940 1764
rect 1916 1716 1924 1724
rect 2012 1796 2020 1804
rect 2076 1796 2084 1804
rect 2060 1736 2068 1744
rect 2156 1916 2164 1924
rect 2300 1936 2308 1944
rect 2300 1916 2308 1924
rect 2380 2336 2388 2344
rect 2508 2376 2516 2384
rect 2508 2316 2516 2324
rect 2412 2296 2420 2304
rect 2444 2296 2452 2304
rect 2588 2516 2596 2524
rect 2604 2336 2612 2344
rect 2556 2316 2564 2324
rect 2588 2316 2596 2324
rect 2748 2516 2756 2524
rect 2876 2516 2884 2524
rect 2844 2476 2852 2484
rect 2700 2356 2708 2364
rect 2956 2676 2964 2684
rect 2988 2676 2996 2684
rect 3020 2676 3028 2684
rect 2915 2606 2923 2614
rect 2925 2606 2933 2614
rect 2935 2606 2943 2614
rect 2945 2606 2953 2614
rect 2955 2606 2963 2614
rect 2965 2606 2973 2614
rect 3180 2936 3188 2944
rect 3276 2916 3284 2924
rect 3212 2896 3220 2904
rect 3308 2896 3316 2904
rect 3676 3456 3684 3464
rect 3692 3456 3700 3464
rect 3756 3456 3764 3464
rect 3516 3276 3524 3284
rect 3500 3216 3508 3224
rect 3468 3196 3476 3204
rect 3484 3196 3492 3204
rect 3420 3056 3428 3064
rect 3388 3036 3396 3044
rect 3484 3056 3492 3064
rect 3548 3376 3556 3384
rect 3692 3416 3700 3424
rect 3724 3396 3732 3404
rect 3612 3356 3620 3364
rect 3596 3336 3604 3344
rect 3644 3336 3652 3344
rect 3692 3336 3700 3344
rect 3580 3316 3588 3324
rect 3628 3276 3636 3284
rect 3564 3216 3572 3224
rect 3564 3196 3572 3204
rect 3644 3196 3652 3204
rect 3516 3156 3524 3164
rect 3532 3156 3540 3164
rect 3516 3016 3524 3024
rect 3660 3156 3668 3164
rect 3676 3156 3684 3164
rect 3740 3116 3748 3124
rect 3692 3096 3700 3104
rect 3724 3096 3732 3104
rect 3596 3076 3604 3084
rect 3580 3036 3588 3044
rect 3452 2976 3460 2984
rect 3532 2976 3540 2984
rect 3564 2956 3572 2964
rect 3868 3596 3876 3604
rect 3852 3496 3860 3504
rect 3948 3936 3956 3944
rect 4172 4616 4180 4624
rect 4076 4596 4084 4604
rect 4060 4556 4068 4564
rect 4028 4516 4036 4524
rect 4364 4896 4372 4904
rect 4476 5318 4484 5324
rect 4476 5316 4484 5318
rect 4444 5276 4452 5284
rect 4636 5276 4644 5284
rect 4419 5206 4427 5214
rect 4429 5206 4437 5214
rect 4439 5206 4447 5214
rect 4449 5206 4457 5214
rect 4459 5206 4467 5214
rect 4469 5206 4477 5214
rect 4636 5176 4644 5184
rect 4412 5136 4420 5144
rect 4508 5136 4516 5144
rect 4604 5096 4612 5104
rect 4540 5016 4548 5024
rect 4492 4956 4500 4964
rect 4556 4976 4564 4984
rect 4572 4936 4580 4944
rect 4540 4916 4548 4924
rect 4508 4896 4516 4904
rect 4419 4806 4427 4814
rect 4429 4806 4437 4814
rect 4439 4806 4447 4814
rect 4449 4806 4457 4814
rect 4459 4806 4467 4814
rect 4469 4806 4477 4814
rect 4396 4736 4404 4744
rect 4492 4736 4500 4744
rect 4348 4702 4356 4704
rect 4348 4696 4356 4702
rect 4380 4616 4388 4624
rect 4252 4596 4260 4604
rect 4188 4556 4196 4564
rect 4236 4556 4244 4564
rect 4124 4536 4132 4544
rect 4156 4536 4164 4544
rect 4076 4516 4084 4524
rect 4060 4456 4068 4464
rect 4012 4276 4020 4284
rect 4060 4256 4068 4264
rect 4124 4456 4132 4464
rect 4236 4496 4244 4504
rect 4188 4476 4196 4484
rect 4172 4396 4180 4404
rect 4172 4356 4180 4364
rect 4092 4236 4100 4244
rect 4108 4236 4116 4244
rect 4124 4236 4132 4244
rect 4156 4236 4164 4244
rect 4140 4196 4148 4204
rect 4108 4136 4116 4144
rect 3996 3956 4004 3964
rect 4108 4016 4116 4024
rect 4044 3936 4052 3944
rect 4060 3936 4068 3944
rect 4044 3896 4052 3904
rect 3964 3856 3972 3864
rect 3964 3836 3972 3844
rect 3948 3736 3956 3744
rect 3932 3696 3940 3704
rect 3948 3676 3956 3684
rect 4028 3756 4036 3764
rect 4028 3736 4036 3744
rect 4028 3716 4036 3724
rect 3964 3596 3972 3604
rect 4044 3696 4052 3704
rect 4044 3676 4052 3684
rect 3916 3556 3924 3564
rect 3996 3556 4004 3564
rect 4028 3536 4036 3544
rect 3788 3456 3796 3464
rect 3948 3496 3956 3504
rect 3980 3496 3988 3504
rect 3900 3476 3908 3484
rect 3884 3456 3892 3464
rect 3868 3436 3876 3444
rect 3852 3376 3860 3384
rect 3788 3316 3796 3324
rect 3772 3216 3780 3224
rect 3772 3096 3780 3104
rect 3804 3276 3812 3284
rect 3948 3456 3956 3464
rect 3916 3416 3924 3424
rect 3948 3396 3956 3404
rect 3900 3356 3908 3364
rect 4204 4376 4212 4384
rect 4364 4576 4372 4584
rect 4268 4556 4276 4564
rect 4300 4556 4308 4564
rect 4284 4516 4292 4524
rect 4284 4336 4292 4344
rect 4332 4336 4340 4344
rect 4300 4276 4308 4284
rect 4188 4236 4196 4244
rect 4236 4236 4244 4244
rect 4284 4236 4292 4244
rect 4268 4176 4276 4184
rect 4188 4136 4196 4144
rect 4204 4116 4212 4124
rect 4220 4076 4228 4084
rect 4156 4036 4164 4044
rect 4252 4096 4260 4104
rect 4236 4056 4244 4064
rect 4236 4016 4244 4024
rect 4412 4576 4420 4584
rect 4444 4556 4452 4564
rect 4476 4556 4484 4564
rect 4460 4456 4468 4464
rect 4380 4416 4388 4424
rect 4364 4316 4372 4324
rect 4492 4436 4500 4444
rect 4419 4406 4427 4414
rect 4429 4406 4437 4414
rect 4439 4406 4447 4414
rect 4449 4406 4457 4414
rect 4459 4406 4467 4414
rect 4469 4406 4477 4414
rect 4492 4396 4500 4404
rect 4492 4356 4500 4364
rect 4348 4236 4356 4244
rect 4396 4236 4404 4244
rect 4348 4156 4356 4164
rect 4300 4136 4308 4144
rect 4396 4136 4404 4144
rect 4284 4076 4292 4084
rect 4268 4056 4276 4064
rect 4332 3996 4340 4004
rect 4316 3956 4324 3964
rect 4204 3916 4212 3924
rect 4092 3876 4100 3884
rect 4108 3876 4116 3884
rect 4108 3856 4116 3864
rect 4140 3856 4148 3864
rect 4092 3796 4100 3804
rect 4076 3776 4084 3784
rect 4172 3756 4180 3764
rect 4108 3736 4116 3744
rect 4188 3736 4196 3744
rect 4124 3716 4132 3724
rect 4252 3896 4260 3904
rect 4268 3896 4276 3904
rect 4268 3816 4276 3824
rect 4252 3796 4260 3804
rect 4300 3816 4308 3824
rect 4332 3816 4340 3824
rect 4252 3776 4260 3784
rect 4268 3776 4276 3784
rect 4284 3756 4292 3764
rect 4284 3736 4292 3744
rect 4236 3716 4244 3724
rect 4076 3656 4084 3664
rect 4012 3416 4020 3424
rect 4028 3416 4036 3424
rect 3980 3356 3988 3364
rect 4044 3356 4052 3364
rect 4140 3616 4148 3624
rect 4092 3556 4100 3564
rect 4124 3516 4132 3524
rect 4124 3436 4132 3444
rect 3964 3336 3972 3344
rect 4060 3336 4068 3344
rect 4028 3316 4036 3324
rect 4044 3316 4052 3324
rect 3852 3196 3860 3204
rect 3996 3296 4004 3304
rect 4012 3276 4020 3284
rect 4028 3276 4036 3284
rect 3964 3256 3972 3264
rect 3868 3176 3876 3184
rect 3852 3116 3860 3124
rect 3788 3076 3796 3084
rect 3612 3056 3620 3064
rect 3756 3056 3764 3064
rect 3804 3056 3812 3064
rect 3676 3036 3684 3044
rect 3836 3036 3844 3044
rect 3612 2956 3620 2964
rect 3340 2936 3348 2944
rect 3404 2936 3412 2944
rect 3500 2936 3508 2944
rect 3580 2936 3588 2944
rect 3388 2916 3396 2924
rect 3436 2916 3444 2924
rect 3468 2896 3476 2904
rect 3228 2876 3236 2884
rect 3292 2876 3300 2884
rect 3116 2716 3124 2724
rect 3164 2716 3172 2724
rect 3132 2696 3140 2704
rect 3004 2636 3012 2644
rect 2972 2536 2980 2544
rect 2988 2536 2996 2544
rect 2924 2476 2932 2484
rect 2540 2296 2548 2304
rect 2668 2296 2676 2304
rect 2844 2296 2852 2304
rect 2892 2296 2900 2304
rect 2524 2276 2532 2284
rect 2604 2276 2612 2284
rect 2652 2276 2660 2284
rect 2780 2276 2788 2284
rect 2828 2276 2836 2284
rect 2540 2236 2548 2244
rect 2652 2236 2660 2244
rect 2444 2196 2452 2204
rect 2492 2196 2500 2204
rect 2412 2156 2420 2164
rect 2716 2196 2724 2204
rect 3052 2636 3060 2644
rect 3292 2716 3300 2724
rect 3260 2676 3268 2684
rect 3164 2656 3172 2664
rect 3132 2556 3140 2564
rect 3132 2536 3140 2544
rect 3068 2516 3076 2524
rect 3036 2496 3044 2504
rect 3036 2476 3044 2484
rect 3020 2396 3028 2404
rect 2988 2316 2996 2324
rect 3020 2316 3028 2324
rect 3052 2416 3060 2424
rect 3116 2476 3124 2484
rect 3084 2416 3092 2424
rect 3052 2336 3060 2344
rect 3228 2516 3236 2524
rect 3276 2576 3284 2584
rect 3356 2736 3364 2744
rect 3340 2716 3348 2724
rect 3516 2916 3524 2924
rect 3580 2916 3588 2924
rect 3484 2736 3492 2744
rect 3420 2716 3428 2724
rect 3468 2716 3476 2724
rect 3388 2696 3396 2704
rect 3340 2676 3348 2684
rect 3324 2576 3332 2584
rect 3372 2556 3380 2564
rect 3308 2536 3316 2544
rect 3244 2476 3252 2484
rect 3164 2436 3172 2444
rect 3340 2436 3348 2444
rect 3148 2416 3156 2424
rect 3132 2376 3140 2384
rect 3132 2316 3140 2324
rect 2972 2236 2980 2244
rect 2860 2216 2868 2224
rect 2915 2206 2923 2214
rect 2925 2206 2933 2214
rect 2935 2206 2943 2214
rect 2945 2206 2953 2214
rect 2955 2206 2963 2214
rect 2965 2206 2973 2214
rect 2796 2176 2804 2184
rect 2508 2156 2516 2164
rect 2604 2136 2612 2144
rect 2636 2136 2644 2144
rect 2780 2136 2788 2144
rect 2572 2116 2580 2124
rect 2364 2096 2372 2104
rect 2396 2096 2404 2104
rect 2460 2096 2468 2104
rect 2524 2096 2532 2104
rect 2540 2096 2548 2104
rect 2572 2096 2580 2104
rect 2620 2096 2628 2104
rect 2428 2056 2436 2064
rect 2636 2036 2644 2044
rect 2444 2016 2452 2024
rect 2444 1996 2452 2004
rect 2348 1916 2356 1924
rect 2316 1896 2324 1904
rect 2268 1876 2276 1884
rect 2300 1876 2308 1884
rect 2332 1876 2340 1884
rect 2140 1836 2148 1844
rect 2284 1836 2292 1844
rect 2204 1816 2212 1824
rect 2204 1796 2212 1804
rect 2316 1796 2324 1804
rect 2108 1776 2116 1784
rect 2124 1776 2132 1784
rect 2284 1756 2292 1764
rect 2332 1756 2340 1764
rect 2252 1736 2260 1744
rect 2028 1716 2036 1724
rect 2108 1716 2116 1724
rect 2156 1716 2164 1724
rect 2220 1716 2228 1724
rect 2236 1716 2244 1724
rect 2108 1696 2116 1704
rect 1900 1676 1908 1684
rect 1932 1676 1940 1684
rect 1996 1676 2004 1684
rect 2060 1676 2068 1684
rect 1868 1556 1876 1564
rect 1852 1536 1860 1544
rect 1852 1516 1860 1524
rect 1836 1496 1844 1504
rect 1884 1496 1892 1504
rect 1980 1516 1988 1524
rect 2236 1676 2244 1684
rect 2204 1556 2212 1564
rect 2092 1516 2100 1524
rect 2172 1516 2180 1524
rect 1996 1496 2004 1504
rect 2060 1476 2068 1484
rect 1788 1456 1796 1464
rect 1788 1336 1796 1344
rect 1756 1296 1764 1304
rect 1900 1316 1908 1324
rect 1868 1296 1876 1304
rect 1932 1356 1940 1364
rect 1756 1256 1764 1264
rect 1724 1216 1732 1224
rect 1740 1216 1748 1224
rect 1772 1156 1780 1164
rect 1708 1096 1716 1104
rect 1676 1076 1684 1084
rect 1804 1096 1812 1104
rect 1692 1056 1700 1064
rect 1756 1056 1764 1064
rect 1884 1216 1892 1224
rect 1852 1136 1860 1144
rect 1836 1076 1844 1084
rect 1820 1056 1828 1064
rect 1724 956 1732 964
rect 1676 856 1684 864
rect 1740 816 1748 824
rect 1820 916 1828 924
rect 1852 916 1860 924
rect 1772 896 1780 904
rect 1788 896 1796 904
rect 1852 896 1860 904
rect 1980 1436 1988 1444
rect 2012 1436 2020 1444
rect 2076 1456 2084 1464
rect 2044 1376 2052 1384
rect 2060 1376 2068 1384
rect 1964 1336 1972 1344
rect 1980 1336 1988 1344
rect 2060 1336 2068 1344
rect 2188 1496 2196 1504
rect 2124 1436 2132 1444
rect 2220 1516 2228 1524
rect 2396 1936 2404 1944
rect 2460 1936 2468 1944
rect 2412 1916 2420 1924
rect 2380 1896 2388 1904
rect 2652 2016 2660 2024
rect 2668 1976 2676 1984
rect 2492 1896 2500 1904
rect 2524 1896 2532 1904
rect 2556 1896 2564 1904
rect 2652 1896 2660 1904
rect 2444 1876 2452 1884
rect 2460 1876 2468 1884
rect 2476 1876 2484 1884
rect 2364 1736 2372 1744
rect 2396 1736 2404 1744
rect 3148 2296 3156 2304
rect 3036 2256 3044 2264
rect 3020 2156 3028 2164
rect 3020 2136 3028 2144
rect 2892 2116 2900 2124
rect 2828 2096 2836 2104
rect 2796 2036 2804 2044
rect 3004 2096 3012 2104
rect 2892 2016 2900 2024
rect 2876 1996 2884 2004
rect 2780 1976 2788 1984
rect 2780 1956 2788 1964
rect 2796 1956 2804 1964
rect 2764 1916 2772 1924
rect 2780 1916 2788 1924
rect 2748 1896 2756 1904
rect 2796 1896 2804 1904
rect 2540 1876 2548 1884
rect 2588 1876 2596 1884
rect 2636 1876 2644 1884
rect 2716 1876 2724 1884
rect 2812 1876 2820 1884
rect 2492 1856 2500 1864
rect 2476 1816 2484 1824
rect 2492 1816 2500 1824
rect 2572 1816 2580 1824
rect 2476 1776 2484 1784
rect 2540 1776 2548 1784
rect 2604 1776 2612 1784
rect 2508 1756 2516 1764
rect 2732 1856 2740 1864
rect 2780 1856 2788 1864
rect 2716 1836 2724 1844
rect 2700 1816 2708 1824
rect 3100 2136 3108 2144
rect 3036 2016 3044 2024
rect 2924 1976 2932 1984
rect 3036 1976 3044 1984
rect 2908 1936 2916 1944
rect 2988 1956 2996 1964
rect 2924 1896 2932 1904
rect 3036 1916 3044 1924
rect 3324 2376 3332 2384
rect 3468 2696 3476 2704
rect 3436 2356 3444 2364
rect 3372 2316 3380 2324
rect 3420 2316 3428 2324
rect 3548 2896 3556 2904
rect 3564 2796 3572 2804
rect 3532 2616 3540 2624
rect 3580 2696 3588 2704
rect 3500 2536 3508 2544
rect 3580 2516 3588 2524
rect 3532 2316 3540 2324
rect 3564 2316 3572 2324
rect 3340 2296 3348 2304
rect 3388 2296 3396 2304
rect 3452 2296 3460 2304
rect 3468 2296 3476 2304
rect 3260 2276 3268 2284
rect 3372 2276 3380 2284
rect 3420 2276 3428 2284
rect 3292 2256 3300 2264
rect 3372 2256 3380 2264
rect 3388 2256 3396 2264
rect 3468 2256 3476 2264
rect 3292 2196 3300 2204
rect 3292 2176 3300 2184
rect 3532 2256 3540 2264
rect 3516 2196 3524 2204
rect 3436 2176 3444 2184
rect 3484 2176 3492 2184
rect 3500 2176 3508 2184
rect 3564 2196 3572 2204
rect 3196 2136 3204 2144
rect 3468 2156 3476 2164
rect 3500 2136 3508 2144
rect 3180 2116 3188 2124
rect 3260 2116 3268 2124
rect 3548 2176 3556 2184
rect 3164 2096 3172 2104
rect 3148 2056 3156 2064
rect 3212 2056 3220 2064
rect 3132 2036 3140 2044
rect 3308 2036 3316 2044
rect 3356 1996 3364 2004
rect 3292 1956 3300 1964
rect 3132 1936 3140 1944
rect 3084 1916 3092 1924
rect 3116 1916 3124 1924
rect 3052 1896 3060 1904
rect 3100 1896 3108 1904
rect 3084 1876 3092 1884
rect 3164 1916 3172 1924
rect 3180 1876 3188 1884
rect 2908 1856 2916 1864
rect 3084 1856 3092 1864
rect 3164 1856 3172 1864
rect 2876 1836 2884 1844
rect 2780 1816 2788 1824
rect 2915 1806 2923 1814
rect 2925 1806 2933 1814
rect 2935 1806 2943 1814
rect 2945 1806 2953 1814
rect 2955 1806 2963 1814
rect 2965 1806 2973 1814
rect 3068 1776 3076 1784
rect 2684 1756 2692 1764
rect 2732 1756 2740 1764
rect 2876 1756 2884 1764
rect 3004 1756 3012 1764
rect 2556 1736 2564 1744
rect 2732 1736 2740 1744
rect 2268 1716 2276 1724
rect 2444 1716 2452 1724
rect 2540 1716 2548 1724
rect 2316 1696 2324 1704
rect 2508 1696 2516 1704
rect 2252 1536 2260 1544
rect 2268 1536 2276 1544
rect 2236 1496 2244 1504
rect 2220 1456 2228 1464
rect 2204 1436 2212 1444
rect 2284 1496 2292 1504
rect 2268 1476 2276 1484
rect 2220 1336 2228 1344
rect 1964 1316 1972 1324
rect 1980 1316 1988 1324
rect 2044 1316 2052 1324
rect 2060 1316 2068 1324
rect 2076 1316 2084 1324
rect 2076 1296 2084 1304
rect 2092 1296 2100 1304
rect 1980 1216 1988 1224
rect 2012 1216 2020 1224
rect 1948 1096 1956 1104
rect 1900 1076 1908 1084
rect 1932 1076 1940 1084
rect 1996 1076 2004 1084
rect 1916 1056 1924 1064
rect 1948 1056 1956 1064
rect 1964 1056 1972 1064
rect 1996 1056 2004 1064
rect 1916 996 1924 1004
rect 1900 956 1908 964
rect 1980 936 1988 944
rect 1916 916 1924 924
rect 1948 916 1956 924
rect 1884 896 1892 904
rect 1932 896 1940 904
rect 1868 876 1876 884
rect 1804 776 1812 784
rect 1996 896 2004 904
rect 1852 736 1860 744
rect 1964 736 1972 744
rect 1708 716 1716 724
rect 1660 696 1668 704
rect 1756 696 1764 704
rect 1836 696 1844 704
rect 1884 696 1892 704
rect 1948 696 1956 704
rect 1612 556 1620 564
rect 1644 556 1652 564
rect 1628 536 1636 544
rect 1884 656 1892 664
rect 1980 716 1988 724
rect 2028 1156 2036 1164
rect 2044 1116 2052 1124
rect 2076 1216 2084 1224
rect 2044 1056 2052 1064
rect 2172 1316 2180 1324
rect 2220 1316 2228 1324
rect 2156 1216 2164 1224
rect 2124 1076 2132 1084
rect 2044 996 2052 1004
rect 2076 976 2084 984
rect 2060 876 2068 884
rect 2076 776 2084 784
rect 2252 1356 2260 1364
rect 2332 1656 2340 1664
rect 2348 1656 2356 1664
rect 2396 1656 2404 1664
rect 2332 1556 2340 1564
rect 2428 1556 2436 1564
rect 2380 1536 2388 1544
rect 2396 1536 2404 1544
rect 2364 1516 2372 1524
rect 2300 1456 2308 1464
rect 2316 1456 2324 1464
rect 2284 1436 2292 1444
rect 2300 1436 2308 1444
rect 2268 1316 2276 1324
rect 2252 1296 2260 1304
rect 2268 1296 2276 1304
rect 2188 1116 2196 1124
rect 2268 1056 2276 1064
rect 2300 1376 2308 1384
rect 2300 1356 2308 1364
rect 2300 1296 2308 1304
rect 2348 1416 2356 1424
rect 2364 1416 2372 1424
rect 2444 1516 2452 1524
rect 2396 1396 2404 1404
rect 2588 1676 2596 1684
rect 2652 1656 2660 1664
rect 2588 1516 2596 1524
rect 2460 1476 2468 1484
rect 2492 1476 2500 1484
rect 2604 1476 2612 1484
rect 2764 1716 2772 1724
rect 2812 1716 2820 1724
rect 3132 1756 3140 1764
rect 3052 1736 3060 1744
rect 3100 1736 3108 1744
rect 3004 1716 3012 1724
rect 3052 1716 3060 1724
rect 2716 1696 2724 1704
rect 2828 1696 2836 1704
rect 2844 1696 2852 1704
rect 2988 1696 2996 1704
rect 2764 1496 2772 1504
rect 2652 1456 2660 1464
rect 2668 1456 2676 1464
rect 2460 1436 2468 1444
rect 2508 1436 2516 1444
rect 2572 1436 2580 1444
rect 2636 1436 2644 1444
rect 2396 1376 2404 1384
rect 2428 1376 2436 1384
rect 2332 1356 2340 1364
rect 2396 1336 2404 1344
rect 2444 1336 2452 1344
rect 2380 1296 2388 1304
rect 2364 1236 2372 1244
rect 2316 1176 2324 1184
rect 2300 1056 2308 1064
rect 2316 996 2324 1004
rect 2348 1156 2356 1164
rect 2412 1316 2420 1324
rect 2444 1316 2452 1324
rect 2428 1196 2436 1204
rect 2220 976 2228 984
rect 2284 976 2292 984
rect 2332 976 2340 984
rect 2156 956 2164 964
rect 2188 956 2196 964
rect 2252 956 2260 964
rect 2268 956 2276 964
rect 2108 936 2116 944
rect 2156 936 2164 944
rect 2124 836 2132 844
rect 2060 696 2068 704
rect 2028 676 2036 684
rect 2140 696 2148 704
rect 2012 656 2020 664
rect 2060 656 2068 664
rect 2092 656 2100 664
rect 1964 556 1972 564
rect 2092 636 2100 644
rect 2092 576 2100 584
rect 2044 556 2052 564
rect 2140 556 2148 564
rect 2188 916 2196 924
rect 2220 916 2228 924
rect 2204 836 2212 844
rect 2172 716 2180 724
rect 2204 716 2212 724
rect 2204 676 2212 684
rect 2188 656 2196 664
rect 2300 896 2308 904
rect 2412 1056 2420 1064
rect 2396 1036 2404 1044
rect 2492 1416 2500 1424
rect 2476 1376 2484 1384
rect 2460 1196 2468 1204
rect 2556 1416 2564 1424
rect 2540 1376 2548 1384
rect 2700 1456 2708 1464
rect 2684 1436 2692 1444
rect 2668 1416 2676 1424
rect 2652 1396 2660 1404
rect 2828 1516 2836 1524
rect 2796 1496 2804 1504
rect 2796 1456 2804 1464
rect 2652 1376 2660 1384
rect 2588 1356 2596 1364
rect 2604 1356 2612 1364
rect 2524 1336 2532 1344
rect 2540 1336 2548 1344
rect 2588 1336 2596 1344
rect 2636 1336 2644 1344
rect 2700 1376 2708 1384
rect 2732 1356 2740 1364
rect 2764 1356 2772 1364
rect 2684 1336 2692 1344
rect 2716 1336 2724 1344
rect 2604 1316 2612 1324
rect 2620 1316 2628 1324
rect 2668 1316 2676 1324
rect 2588 1196 2596 1204
rect 2668 1196 2676 1204
rect 2492 1116 2500 1124
rect 2508 1116 2516 1124
rect 2524 1116 2532 1124
rect 2572 1116 2580 1124
rect 2636 1116 2644 1124
rect 2476 976 2484 984
rect 2492 976 2500 984
rect 2556 976 2564 984
rect 2572 976 2580 984
rect 2460 956 2468 964
rect 2428 936 2436 944
rect 2380 916 2388 924
rect 2412 916 2420 924
rect 2460 916 2468 924
rect 2348 836 2356 844
rect 2444 796 2452 804
rect 2316 756 2324 764
rect 2428 736 2436 744
rect 2252 716 2260 724
rect 2284 696 2292 704
rect 2316 696 2324 704
rect 2396 696 2404 704
rect 2460 736 2468 744
rect 2476 736 2484 744
rect 2540 716 2548 724
rect 2476 696 2484 704
rect 2492 696 2500 704
rect 2428 676 2436 684
rect 2524 676 2532 684
rect 2236 656 2244 664
rect 2284 656 2292 664
rect 2380 656 2388 664
rect 2444 656 2452 664
rect 2508 656 2516 664
rect 2300 576 2308 584
rect 2332 576 2340 584
rect 2284 536 2292 544
rect 2316 536 2324 544
rect 1900 516 1908 524
rect 2076 516 2084 524
rect 2124 516 2132 524
rect 2172 516 2180 524
rect 2188 516 2196 524
rect 2220 516 2228 524
rect 1708 496 1716 504
rect 1740 496 1748 504
rect 1788 496 1796 504
rect 1724 456 1732 464
rect 1580 436 1588 444
rect 1612 416 1620 424
rect 1692 336 1700 344
rect 1852 496 1860 504
rect 1804 416 1812 424
rect 1836 416 1844 424
rect 1676 256 1684 264
rect 1548 236 1556 244
rect 1692 176 1700 184
rect 1916 356 1924 364
rect 1820 256 1828 264
rect 1564 156 1572 164
rect 1644 156 1652 164
rect 1756 156 1764 164
rect 1532 136 1540 144
rect 1628 136 1636 144
rect 1660 116 1668 124
rect 2092 416 2100 424
rect 1980 356 1988 364
rect 1948 336 1956 344
rect 2076 336 2084 344
rect 2156 316 2164 324
rect 2172 316 2180 324
rect 2188 316 2196 324
rect 1996 276 2004 284
rect 2028 276 2036 284
rect 2044 276 2052 284
rect 2076 276 2084 284
rect 2156 276 2164 284
rect 2300 496 2308 504
rect 2300 456 2308 464
rect 2284 316 2292 324
rect 2220 296 2228 304
rect 2364 556 2372 564
rect 2348 516 2356 524
rect 2332 376 2340 384
rect 2428 556 2436 564
rect 2508 556 2516 564
rect 2524 556 2532 564
rect 2444 536 2452 544
rect 2508 536 2516 544
rect 2428 516 2436 524
rect 2524 516 2532 524
rect 2748 1316 2756 1324
rect 2780 1336 2788 1344
rect 2908 1516 2916 1524
rect 3180 1736 3188 1744
rect 3164 1696 3172 1704
rect 3052 1636 3060 1644
rect 3100 1576 3108 1584
rect 3084 1536 3092 1544
rect 3004 1516 3012 1524
rect 3052 1516 3060 1524
rect 2892 1456 2900 1464
rect 2876 1436 2884 1444
rect 2828 1356 2836 1364
rect 2812 1336 2820 1344
rect 2860 1396 2868 1404
rect 2876 1376 2884 1384
rect 2915 1406 2923 1414
rect 2925 1406 2933 1414
rect 2935 1406 2943 1414
rect 2945 1406 2953 1414
rect 2955 1406 2963 1414
rect 2965 1406 2973 1414
rect 2908 1376 2916 1384
rect 2860 1356 2868 1364
rect 2892 1356 2900 1364
rect 2924 1356 2932 1364
rect 2940 1356 2948 1364
rect 2924 1336 2932 1344
rect 2844 1316 2852 1324
rect 2860 1316 2868 1324
rect 2764 1196 2772 1204
rect 2812 1196 2820 1204
rect 2828 1196 2836 1204
rect 2876 1196 2884 1204
rect 2892 1196 2900 1204
rect 2860 1116 2868 1124
rect 2620 956 2628 964
rect 2684 956 2692 964
rect 2588 916 2596 924
rect 2604 916 2612 924
rect 2572 896 2580 904
rect 2636 896 2644 904
rect 2620 836 2628 844
rect 2652 836 2660 844
rect 2636 756 2644 764
rect 2620 736 2628 744
rect 2636 736 2644 744
rect 2684 796 2692 804
rect 2748 1056 2756 1064
rect 2764 1056 2772 1064
rect 2812 1056 2820 1064
rect 2844 1056 2852 1064
rect 2732 976 2740 984
rect 3068 1436 3076 1444
rect 3036 1416 3044 1424
rect 3228 1796 3236 1804
rect 3212 1756 3220 1764
rect 3244 1776 3252 1784
rect 3260 1756 3268 1764
rect 3196 1696 3204 1704
rect 3388 1916 3396 1924
rect 3468 1916 3476 1924
rect 3612 2896 3620 2904
rect 3884 3056 3892 3064
rect 3820 3016 3828 3024
rect 3868 3016 3876 3024
rect 3788 2996 3796 3004
rect 3884 2996 3892 3004
rect 3644 2916 3652 2924
rect 3660 2896 3668 2904
rect 3772 2916 3780 2924
rect 3708 2856 3716 2864
rect 3756 2856 3764 2864
rect 3628 2796 3636 2804
rect 3628 2716 3636 2724
rect 3724 2716 3732 2724
rect 3724 2676 3732 2684
rect 3772 2676 3780 2684
rect 3948 3176 3956 3184
rect 3932 3116 3940 3124
rect 4060 3216 4068 3224
rect 3964 3156 3972 3164
rect 4060 3156 4068 3164
rect 4044 3116 4052 3124
rect 4076 3116 4084 3124
rect 4012 3096 4020 3104
rect 4060 3096 4068 3104
rect 3948 3016 3956 3024
rect 3916 2736 3924 2744
rect 3868 2716 3876 2724
rect 4044 2996 4052 3004
rect 3996 2916 4004 2924
rect 4028 2776 4036 2784
rect 4044 2716 4052 2724
rect 3996 2696 4004 2704
rect 3948 2676 3956 2684
rect 3788 2636 3796 2644
rect 3692 2576 3700 2584
rect 3692 2556 3700 2564
rect 3660 2536 3668 2544
rect 3676 2516 3684 2524
rect 3676 2496 3684 2504
rect 3596 2476 3604 2484
rect 3596 2376 3604 2384
rect 3628 2316 3636 2324
rect 3676 2296 3684 2304
rect 3612 2276 3620 2284
rect 3644 2256 3652 2264
rect 3596 2116 3604 2124
rect 3548 2056 3556 2064
rect 3580 2056 3588 2064
rect 3324 1896 3332 1904
rect 3356 1896 3364 1904
rect 3452 1896 3460 1904
rect 3500 1896 3508 1904
rect 3516 1896 3524 1904
rect 3548 1896 3556 1904
rect 3340 1876 3348 1884
rect 3388 1876 3396 1884
rect 3372 1816 3380 1824
rect 3324 1796 3332 1804
rect 3452 1856 3460 1864
rect 3420 1816 3428 1824
rect 3436 1796 3444 1804
rect 3388 1736 3396 1744
rect 3260 1716 3268 1724
rect 3276 1716 3284 1724
rect 3196 1576 3204 1584
rect 3516 1816 3524 1824
rect 3580 1856 3588 1864
rect 3564 1816 3572 1824
rect 3532 1796 3540 1804
rect 3516 1776 3524 1784
rect 3612 2036 3620 2044
rect 3676 2156 3684 2164
rect 3788 2576 3796 2584
rect 3868 2556 3876 2564
rect 4060 2556 4068 2564
rect 4140 3336 4148 3344
rect 4188 3376 4196 3384
rect 4156 3316 4164 3324
rect 4156 3176 4164 3184
rect 4172 3096 4180 3104
rect 4140 3016 4148 3024
rect 4220 3116 4228 3124
rect 4220 3096 4228 3104
rect 4220 2996 4228 3004
rect 4204 2956 4212 2964
rect 4092 2936 4100 2944
rect 4188 2936 4196 2944
rect 4284 3676 4292 3684
rect 4348 3796 4356 3804
rect 4428 4296 4436 4304
rect 4460 4276 4468 4284
rect 4460 4236 4468 4244
rect 4444 4216 4452 4224
rect 4428 4156 4436 4164
rect 4380 4096 4388 4104
rect 4380 4076 4388 4084
rect 4364 3776 4372 3784
rect 4316 3736 4324 3744
rect 4460 4036 4468 4044
rect 4419 4006 4427 4014
rect 4429 4006 4437 4014
rect 4439 4006 4447 4014
rect 4449 4006 4457 4014
rect 4459 4006 4467 4014
rect 4469 4006 4477 4014
rect 4588 4916 4596 4924
rect 4588 4796 4596 4804
rect 4588 4716 4596 4724
rect 4588 4536 4596 4544
rect 4796 5156 4804 5164
rect 4684 5116 4692 5124
rect 4668 5096 4676 5104
rect 4764 5102 4772 5104
rect 4764 5096 4772 5102
rect 4684 5076 4692 5084
rect 4732 5076 4740 5084
rect 4636 5036 4644 5044
rect 4684 5036 4692 5044
rect 4620 5016 4628 5024
rect 4732 5016 4740 5024
rect 4700 4996 4708 5004
rect 4732 4956 4740 4964
rect 4764 4956 4772 4964
rect 4748 4916 4756 4924
rect 4620 4696 4628 4704
rect 4668 4816 4676 4824
rect 4668 4796 4676 4804
rect 4636 4636 4644 4644
rect 4748 4896 4756 4904
rect 4748 4876 4756 4884
rect 4732 4836 4740 4844
rect 4764 4816 4772 4824
rect 4764 4796 4772 4804
rect 4732 4676 4740 4684
rect 4684 4656 4692 4664
rect 4748 4636 4756 4644
rect 4636 4536 4644 4544
rect 4556 4516 4564 4524
rect 4604 4516 4612 4524
rect 4620 4516 4628 4524
rect 4588 4476 4596 4484
rect 4556 4456 4564 4464
rect 4540 4376 4548 4384
rect 4556 4356 4564 4364
rect 4540 4316 4548 4324
rect 4620 4376 4628 4384
rect 4668 4476 4676 4484
rect 4652 4396 4660 4404
rect 4588 4336 4596 4344
rect 4572 4156 4580 4164
rect 4876 5316 4884 5324
rect 4972 5318 4980 5324
rect 4972 5316 4980 5318
rect 4940 5276 4948 5284
rect 4828 5256 4836 5264
rect 4876 5256 4884 5264
rect 4892 5176 4900 5184
rect 4924 5176 4932 5184
rect 4908 5136 4916 5144
rect 5036 5102 5044 5104
rect 5036 5096 5044 5102
rect 5116 5316 5124 5324
rect 5164 5316 5172 5324
rect 5100 5216 5108 5224
rect 5180 5196 5188 5204
rect 5132 5176 5140 5184
rect 5180 5176 5188 5184
rect 5100 5136 5108 5144
rect 5148 5096 5156 5104
rect 5068 5056 5076 5064
rect 5228 5056 5236 5064
rect 5196 5036 5204 5044
rect 4812 4956 4820 4964
rect 4860 4936 4868 4944
rect 4828 4916 4836 4924
rect 4812 4896 4820 4904
rect 4828 4896 4836 4904
rect 4796 4836 4804 4844
rect 4796 4816 4804 4824
rect 4956 4916 4964 4924
rect 4988 4916 4996 4924
rect 5004 4916 5012 4924
rect 5036 4916 5044 4924
rect 5068 4916 5076 4924
rect 5116 4916 5124 4924
rect 4908 4896 4916 4904
rect 4892 4876 4900 4884
rect 4988 4876 4996 4884
rect 4892 4816 4900 4824
rect 4908 4816 4916 4824
rect 4876 4796 4884 4804
rect 4908 4776 4916 4784
rect 4780 4676 4788 4684
rect 4780 4636 4788 4644
rect 4764 4596 4772 4604
rect 4748 4516 4756 4524
rect 4748 4396 4756 4404
rect 4700 4376 4708 4384
rect 4636 4336 4644 4344
rect 4684 4336 4692 4344
rect 4732 4336 4740 4344
rect 4620 4116 4628 4124
rect 4524 4096 4532 4104
rect 4604 4056 4612 4064
rect 4588 3996 4596 4004
rect 4508 3976 4516 3984
rect 4492 3856 4500 3864
rect 4428 3816 4436 3824
rect 4412 3716 4420 3724
rect 4364 3636 4372 3644
rect 4380 3636 4388 3644
rect 4419 3606 4427 3614
rect 4429 3606 4437 3614
rect 4439 3606 4447 3614
rect 4449 3606 4457 3614
rect 4459 3606 4467 3614
rect 4469 3606 4477 3614
rect 4636 4016 4644 4024
rect 4620 3996 4628 4004
rect 4620 3976 4628 3984
rect 4604 3936 4612 3944
rect 4556 3796 4564 3804
rect 4540 3756 4548 3764
rect 4716 4256 4724 4264
rect 4668 4236 4676 4244
rect 4668 4136 4676 4144
rect 4652 3976 4660 3984
rect 4684 4116 4692 4124
rect 4716 4116 4724 4124
rect 4700 3956 4708 3964
rect 4748 4076 4756 4084
rect 4972 4756 4980 4764
rect 4924 4736 4932 4744
rect 4860 4696 4868 4704
rect 4796 4576 4804 4584
rect 4876 4576 4884 4584
rect 5052 4896 5060 4904
rect 5068 4896 5076 4904
rect 5180 4976 5188 4984
rect 5196 4956 5204 4964
rect 5132 4896 5140 4904
rect 5148 4876 5156 4884
rect 5148 4856 5156 4864
rect 5084 4836 5092 4844
rect 5084 4776 5092 4784
rect 5068 4736 5076 4744
rect 5020 4696 5028 4704
rect 5068 4696 5076 4704
rect 5132 4756 5140 4764
rect 5100 4696 5108 4704
rect 5052 4656 5060 4664
rect 5084 4656 5092 4664
rect 5004 4616 5012 4624
rect 5020 4616 5028 4624
rect 4924 4556 4932 4564
rect 4892 4316 4900 4324
rect 4940 4536 4948 4544
rect 5004 4376 5012 4384
rect 5036 4576 5044 4584
rect 5164 4716 5172 4724
rect 5228 4836 5236 4844
rect 6172 5376 6180 5384
rect 6252 5376 6260 5384
rect 5404 5336 5412 5344
rect 5292 5316 5300 5324
rect 5420 5316 5428 5324
rect 5404 5276 5412 5284
rect 5484 5336 5492 5344
rect 5580 5336 5588 5344
rect 5500 5316 5508 5324
rect 5452 5236 5460 5244
rect 5404 5196 5412 5204
rect 5500 5176 5508 5184
rect 5404 5136 5412 5144
rect 5292 5016 5300 5024
rect 5388 5036 5396 5044
rect 5372 4976 5380 4984
rect 5420 5096 5428 5104
rect 5484 5116 5492 5124
rect 5436 5076 5444 5084
rect 5452 5076 5460 5084
rect 5532 5116 5540 5124
rect 5548 5116 5556 5124
rect 5548 5076 5556 5084
rect 5516 5016 5524 5024
rect 5484 4996 5492 5004
rect 5500 4996 5508 5004
rect 5468 4976 5476 4984
rect 5404 4956 5412 4964
rect 5452 4956 5460 4964
rect 5436 4936 5444 4944
rect 5308 4876 5316 4884
rect 5420 4876 5428 4884
rect 5420 4756 5428 4764
rect 5276 4716 5284 4724
rect 5340 4716 5348 4724
rect 5164 4636 5172 4644
rect 5116 4596 5124 4604
rect 5116 4576 5124 4584
rect 5084 4536 5092 4544
rect 5148 4536 5156 4544
rect 5036 4516 5044 4524
rect 5020 4336 5028 4344
rect 4796 4296 4804 4304
rect 4876 4296 4884 4304
rect 4828 4256 4836 4264
rect 4860 4236 4868 4244
rect 5020 4316 5028 4324
rect 5036 4316 5044 4324
rect 4924 4216 4932 4224
rect 4876 4156 4884 4164
rect 4860 4116 4868 4124
rect 4748 3996 4756 4004
rect 4764 3936 4772 3944
rect 4716 3876 4724 3884
rect 4748 3856 4756 3864
rect 4732 3816 4740 3824
rect 4748 3816 4756 3824
rect 4668 3756 4676 3764
rect 4604 3716 4612 3724
rect 4540 3676 4548 3684
rect 4492 3596 4500 3604
rect 4396 3536 4404 3544
rect 4300 3476 4308 3484
rect 4252 3456 4260 3464
rect 4364 3456 4372 3464
rect 4284 3396 4292 3404
rect 4348 3396 4356 3404
rect 4252 3316 4260 3324
rect 4300 3336 4308 3344
rect 4380 3356 4388 3364
rect 4332 3316 4340 3324
rect 4364 3316 4372 3324
rect 4364 3256 4372 3264
rect 4268 3196 4276 3204
rect 4364 3176 4372 3184
rect 4252 3116 4260 3124
rect 4316 3102 4324 3104
rect 4316 3096 4324 3102
rect 4284 2976 4292 2984
rect 4252 2956 4260 2964
rect 4188 2876 4196 2884
rect 4236 2876 4244 2884
rect 4108 2796 4116 2804
rect 4092 2776 4100 2784
rect 4092 2636 4100 2644
rect 4140 2736 4148 2744
rect 4124 2716 4132 2724
rect 4156 2716 4164 2724
rect 4172 2676 4180 2684
rect 4348 2936 4356 2944
rect 4508 3516 4516 3524
rect 4636 3676 4644 3684
rect 4620 3616 4628 3624
rect 4716 3756 4724 3764
rect 4796 3976 4804 3984
rect 4796 3936 4804 3944
rect 4780 3916 4788 3924
rect 4892 4116 4900 4124
rect 4892 4096 4900 4104
rect 4876 3996 4884 4004
rect 4892 3996 4900 4004
rect 4828 3976 4836 3984
rect 4924 4096 4932 4104
rect 4908 3956 4916 3964
rect 4924 3956 4932 3964
rect 5020 4156 5028 4164
rect 4892 3936 4900 3944
rect 4908 3916 4916 3924
rect 4812 3896 4820 3904
rect 4860 3896 4868 3904
rect 4892 3896 4900 3904
rect 4924 3896 4932 3904
rect 4876 3876 4884 3884
rect 4796 3856 4804 3864
rect 4844 3816 4852 3824
rect 4700 3716 4708 3724
rect 4780 3796 4788 3804
rect 4828 3756 4836 3764
rect 4764 3696 4772 3704
rect 4812 3696 4820 3704
rect 4668 3676 4676 3684
rect 4748 3676 4756 3684
rect 4700 3636 4708 3644
rect 4668 3616 4676 3624
rect 4652 3596 4660 3604
rect 4556 3536 4564 3544
rect 4620 3536 4628 3544
rect 4588 3516 4596 3524
rect 4652 3516 4660 3524
rect 4684 3596 4692 3604
rect 4700 3596 4708 3604
rect 4556 3476 4564 3484
rect 4636 3476 4644 3484
rect 4668 3476 4676 3484
rect 4684 3476 4692 3484
rect 4620 3456 4628 3464
rect 4524 3436 4532 3444
rect 4556 3396 4564 3404
rect 4540 3376 4548 3384
rect 4492 3356 4500 3364
rect 4508 3356 4516 3364
rect 4428 3336 4436 3344
rect 4444 3336 4452 3344
rect 4444 3296 4452 3304
rect 4412 3256 4420 3264
rect 4396 3216 4404 3224
rect 4524 3256 4532 3264
rect 4419 3206 4427 3214
rect 4429 3206 4437 3214
rect 4439 3206 4447 3214
rect 4449 3206 4457 3214
rect 4459 3206 4467 3214
rect 4469 3206 4477 3214
rect 4492 3196 4500 3204
rect 4444 3116 4452 3124
rect 4492 3076 4500 3084
rect 4380 3036 4388 3044
rect 4236 2816 4244 2824
rect 4268 2816 4276 2824
rect 4220 2716 4228 2724
rect 4172 2596 4180 2604
rect 4188 2596 4196 2604
rect 3996 2536 4004 2544
rect 4204 2536 4212 2544
rect 4252 2716 4260 2724
rect 4268 2676 4276 2684
rect 4236 2636 4244 2644
rect 3756 2516 3764 2524
rect 4028 2516 4036 2524
rect 4076 2516 4084 2524
rect 4172 2516 4180 2524
rect 4076 2476 4084 2484
rect 4108 2476 4116 2484
rect 4060 2356 4068 2364
rect 3948 2316 3956 2324
rect 3868 2296 3876 2304
rect 3820 2276 3828 2284
rect 3772 2136 3780 2144
rect 3660 1916 3668 1924
rect 3628 1896 3636 1904
rect 3596 1736 3604 1744
rect 3420 1716 3428 1724
rect 3468 1716 3476 1724
rect 3596 1716 3604 1724
rect 3308 1536 3316 1544
rect 3212 1516 3220 1524
rect 3116 1496 3124 1504
rect 3148 1496 3156 1504
rect 3180 1496 3188 1504
rect 3244 1496 3252 1504
rect 3132 1456 3140 1464
rect 3116 1396 3124 1404
rect 3036 1316 3044 1324
rect 3068 1336 3076 1344
rect 3100 1336 3108 1344
rect 3036 1296 3044 1304
rect 3052 1296 3060 1304
rect 3020 1236 3028 1244
rect 3036 1236 3044 1244
rect 2972 1116 2980 1124
rect 2940 1076 2948 1084
rect 2988 1076 2996 1084
rect 2892 1016 2900 1024
rect 2915 1006 2923 1014
rect 2925 1006 2933 1014
rect 2935 1006 2943 1014
rect 2945 1006 2953 1014
rect 2955 1006 2963 1014
rect 2965 1006 2973 1014
rect 2844 996 2852 1004
rect 2892 996 2900 1004
rect 2828 976 2836 984
rect 2716 956 2724 964
rect 2764 956 2772 964
rect 2924 976 2932 984
rect 2716 916 2724 924
rect 2796 916 2804 924
rect 2860 956 2868 964
rect 2892 956 2900 964
rect 2892 936 2900 944
rect 2844 916 2852 924
rect 2860 916 2868 924
rect 2796 836 2804 844
rect 2812 836 2820 844
rect 2700 776 2708 784
rect 2700 756 2708 764
rect 2572 696 2580 704
rect 2604 696 2612 704
rect 2668 696 2676 704
rect 2636 676 2644 684
rect 2604 656 2612 664
rect 2796 796 2804 804
rect 2828 756 2836 764
rect 2876 896 2884 904
rect 2892 896 2900 904
rect 2860 836 2868 844
rect 2892 836 2900 844
rect 2940 836 2948 844
rect 2908 796 2916 804
rect 2876 776 2884 784
rect 2876 736 2884 744
rect 2844 696 2852 704
rect 2684 676 2692 684
rect 2716 676 2724 684
rect 2892 676 2900 684
rect 2668 596 2676 604
rect 2796 656 2804 664
rect 2732 596 2740 604
rect 2620 556 2628 564
rect 2684 556 2692 564
rect 2748 556 2756 564
rect 2812 556 2820 564
rect 2588 516 2596 524
rect 2556 496 2564 504
rect 2604 456 2612 464
rect 2492 436 2500 444
rect 2540 436 2548 444
rect 2204 276 2212 284
rect 1916 256 1924 264
rect 1980 256 1988 264
rect 2012 256 2020 264
rect 1932 236 1940 244
rect 1868 176 1876 184
rect 1820 136 1828 144
rect 2012 236 2020 244
rect 2124 256 2132 264
rect 2300 256 2308 264
rect 2108 196 2116 204
rect 2172 196 2180 204
rect 2092 176 2100 184
rect 2108 156 2116 164
rect 1868 116 1876 124
rect 2012 116 2020 124
rect 12 96 20 104
rect 556 96 564 104
rect 652 96 660 104
rect 684 96 692 104
rect 1724 96 1732 104
rect 2204 176 2212 184
rect 2380 236 2388 244
rect 2332 136 2340 144
rect 2140 116 2148 124
rect 2268 116 2276 124
rect 2284 116 2292 124
rect 2460 236 2468 244
rect 2540 236 2548 244
rect 2412 176 2420 184
rect 2508 176 2516 184
rect 2396 156 2404 164
rect 2428 156 2436 164
rect 2476 136 2484 144
rect 2572 256 2580 264
rect 2876 616 2884 624
rect 2940 656 2948 664
rect 2915 606 2923 614
rect 2925 606 2933 614
rect 2935 606 2943 614
rect 2945 606 2953 614
rect 2955 606 2963 614
rect 2965 606 2973 614
rect 2892 596 2900 604
rect 2876 576 2884 584
rect 2876 556 2884 564
rect 2748 536 2756 544
rect 2844 536 2852 544
rect 2636 516 2644 524
rect 2780 516 2788 524
rect 2828 496 2836 504
rect 2860 476 2868 484
rect 2652 456 2660 464
rect 2796 456 2804 464
rect 3020 996 3028 1004
rect 3100 1196 3108 1204
rect 3148 1416 3156 1424
rect 3388 1476 3396 1484
rect 3260 1456 3268 1464
rect 3276 1396 3284 1404
rect 3308 1396 3316 1404
rect 3196 1376 3204 1384
rect 3292 1376 3300 1384
rect 3260 1336 3268 1344
rect 3148 1296 3156 1304
rect 3148 1196 3156 1204
rect 3228 1296 3236 1304
rect 3180 1196 3188 1204
rect 3164 1116 3172 1124
rect 3132 1096 3140 1104
rect 3084 1076 3092 1084
rect 3116 1056 3124 1064
rect 3052 1016 3060 1024
rect 3116 1016 3124 1024
rect 3020 956 3028 964
rect 3052 956 3060 964
rect 3004 936 3012 944
rect 3052 936 3060 944
rect 3068 936 3076 944
rect 3148 936 3156 944
rect 3020 916 3028 924
rect 3036 916 3044 924
rect 3084 916 3092 924
rect 3148 916 3156 924
rect 3228 1116 3236 1124
rect 3196 1056 3204 1064
rect 3228 1056 3236 1064
rect 3244 1056 3252 1064
rect 3196 1016 3204 1024
rect 3228 976 3236 984
rect 3276 1296 3284 1304
rect 3276 1016 3284 1024
rect 3260 956 3268 964
rect 3196 916 3204 924
rect 3244 916 3252 924
rect 3180 876 3188 884
rect 3004 836 3012 844
rect 3004 796 3012 804
rect 3036 796 3044 804
rect 3196 796 3204 804
rect 3276 796 3284 804
rect 3020 736 3028 744
rect 3004 696 3012 704
rect 3004 616 3012 624
rect 3052 716 3060 724
rect 3100 716 3108 724
rect 3244 756 3252 764
rect 3212 736 3220 744
rect 3276 736 3284 744
rect 3324 1316 3332 1324
rect 3420 1476 3428 1484
rect 3420 1436 3428 1444
rect 3628 1776 3636 1784
rect 3724 2116 3732 2124
rect 3692 1956 3700 1964
rect 3804 1956 3812 1964
rect 3724 1896 3732 1904
rect 3708 1876 3716 1884
rect 3692 1736 3700 1744
rect 3660 1676 3668 1684
rect 3676 1656 3684 1664
rect 3660 1636 3668 1644
rect 3644 1556 3652 1564
rect 3676 1596 3684 1604
rect 3788 1896 3796 1904
rect 3724 1856 3732 1864
rect 3756 1856 3764 1864
rect 3756 1796 3764 1804
rect 3772 1776 3780 1784
rect 3740 1756 3748 1764
rect 3740 1716 3748 1724
rect 3788 1716 3796 1724
rect 3724 1636 3732 1644
rect 3772 1616 3780 1624
rect 3724 1596 3732 1604
rect 3724 1536 3732 1544
rect 3548 1502 3556 1504
rect 3548 1496 3556 1502
rect 3612 1496 3620 1504
rect 3628 1496 3636 1504
rect 3708 1496 3716 1504
rect 3756 1496 3764 1504
rect 3612 1456 3620 1464
rect 3484 1416 3492 1424
rect 3500 1416 3508 1424
rect 3388 1376 3396 1384
rect 3404 1356 3412 1364
rect 3356 1336 3364 1344
rect 3468 1336 3476 1344
rect 3468 1276 3476 1284
rect 3372 1196 3380 1204
rect 3340 1156 3348 1164
rect 3308 1116 3316 1124
rect 3596 1436 3604 1444
rect 3724 1436 3732 1444
rect 3788 1596 3796 1604
rect 4204 2496 4212 2504
rect 4220 2496 4228 2504
rect 4188 2436 4196 2444
rect 4172 2356 4180 2364
rect 4092 2316 4100 2324
rect 4124 2316 4132 2324
rect 4092 2296 4100 2304
rect 4140 2296 4148 2304
rect 3948 2196 3956 2204
rect 4044 2156 4052 2164
rect 3932 2136 3940 2144
rect 3980 2116 3988 2124
rect 3948 2096 3956 2104
rect 3884 1996 3892 2004
rect 3868 1936 3876 1944
rect 3900 1916 3908 1924
rect 3836 1896 3844 1904
rect 3916 1896 3924 1904
rect 3964 1896 3972 1904
rect 3884 1876 3892 1884
rect 3820 1856 3828 1864
rect 3996 2096 4004 2104
rect 3948 1776 3956 1784
rect 3980 1776 3988 1784
rect 3868 1696 3876 1704
rect 3804 1536 3812 1544
rect 3916 1516 3924 1524
rect 3980 1756 3988 1764
rect 3964 1636 3972 1644
rect 3836 1496 3844 1504
rect 3852 1496 3860 1504
rect 3820 1476 3828 1484
rect 3612 1356 3620 1364
rect 3692 1356 3700 1364
rect 3772 1356 3780 1364
rect 3596 1336 3604 1344
rect 3548 1316 3556 1324
rect 3564 1316 3572 1324
rect 3548 1276 3556 1284
rect 3500 1196 3508 1204
rect 3532 1196 3540 1204
rect 3564 1196 3572 1204
rect 3580 1196 3588 1204
rect 3484 1116 3492 1124
rect 3644 1336 3652 1344
rect 3628 1236 3636 1244
rect 3676 1236 3684 1244
rect 3612 1116 3620 1124
rect 3372 1096 3380 1104
rect 3404 1096 3412 1104
rect 3452 1096 3460 1104
rect 3324 1056 3332 1064
rect 3340 1056 3348 1064
rect 3388 1056 3396 1064
rect 3340 1016 3348 1024
rect 3340 976 3348 984
rect 3372 956 3380 964
rect 3356 936 3364 944
rect 3420 956 3428 964
rect 3436 936 3444 944
rect 3324 896 3332 904
rect 3340 896 3348 904
rect 3372 896 3380 904
rect 3388 896 3396 904
rect 3404 876 3412 884
rect 3436 876 3444 884
rect 3500 1016 3508 1024
rect 3580 1036 3588 1044
rect 3516 996 3524 1004
rect 3548 976 3556 984
rect 3532 956 3540 964
rect 3484 816 3492 824
rect 3452 756 3460 764
rect 3292 716 3300 724
rect 3356 716 3364 724
rect 3388 716 3396 724
rect 3484 716 3492 724
rect 3148 696 3156 704
rect 3196 696 3204 704
rect 3292 696 3300 704
rect 3084 676 3092 684
rect 3100 676 3108 684
rect 3116 616 3124 624
rect 3084 576 3092 584
rect 3084 556 3092 564
rect 3132 556 3140 564
rect 3004 536 3012 544
rect 2892 336 2900 344
rect 2812 296 2820 304
rect 2844 296 2852 304
rect 2780 276 2788 284
rect 2828 276 2836 284
rect 2668 256 2676 264
rect 2604 216 2612 224
rect 2556 176 2564 184
rect 2604 176 2612 184
rect 2876 296 2884 304
rect 2652 236 2660 244
rect 2700 236 2708 244
rect 2860 236 2868 244
rect 2716 216 2724 224
rect 2796 196 2804 204
rect 2588 156 2596 164
rect 2620 156 2628 164
rect 2652 156 2660 164
rect 2716 156 2724 164
rect 2828 156 2836 164
rect 2588 136 2596 144
rect 2636 136 2644 144
rect 2732 136 2740 144
rect 2892 276 2900 284
rect 2988 456 2996 464
rect 3068 536 3076 544
rect 3116 536 3124 544
rect 3052 496 3060 504
rect 3132 496 3140 504
rect 3116 476 3124 484
rect 3228 676 3236 684
rect 3276 676 3284 684
rect 3260 616 3268 624
rect 3180 556 3188 564
rect 3196 536 3204 544
rect 3180 496 3188 504
rect 3164 456 3172 464
rect 3164 436 3172 444
rect 3036 336 3044 344
rect 3308 676 3316 684
rect 3340 676 3348 684
rect 3308 656 3316 664
rect 3276 556 3284 564
rect 3324 556 3332 564
rect 3372 676 3380 684
rect 3420 696 3428 704
rect 3404 676 3412 684
rect 3452 676 3460 684
rect 3388 616 3396 624
rect 3372 556 3380 564
rect 3452 656 3460 664
rect 3468 656 3476 664
rect 3436 556 3444 564
rect 3276 536 3284 544
rect 3356 536 3364 544
rect 3276 516 3284 524
rect 3308 516 3316 524
rect 3356 516 3364 524
rect 3404 516 3412 524
rect 3260 336 3268 344
rect 3212 316 3220 324
rect 3084 296 3092 304
rect 3180 296 3188 304
rect 3404 316 3412 324
rect 3260 296 3268 304
rect 3308 296 3316 304
rect 3340 296 3348 304
rect 3180 276 3188 284
rect 3212 276 3220 284
rect 3292 276 3300 284
rect 3004 256 3012 264
rect 3100 256 3108 264
rect 3132 256 3140 264
rect 3260 256 3268 264
rect 2915 206 2923 214
rect 2925 206 2933 214
rect 2935 206 2943 214
rect 2945 206 2953 214
rect 2955 206 2963 214
rect 2965 206 2973 214
rect 2892 196 2900 204
rect 3100 236 3108 244
rect 2924 176 2932 184
rect 2940 156 2948 164
rect 3052 136 3060 144
rect 2524 116 2532 124
rect 2620 116 2628 124
rect 2716 116 2724 124
rect 2908 116 2916 124
rect 3020 116 3028 124
rect 3180 176 3188 184
rect 3244 156 3252 164
rect 3260 156 3268 164
rect 3436 316 3444 324
rect 3484 636 3492 644
rect 3484 536 3492 544
rect 3468 496 3476 504
rect 3596 898 3604 904
rect 3596 896 3604 898
rect 3644 1216 3652 1224
rect 3900 1456 3908 1464
rect 3916 1436 3924 1444
rect 3868 1396 3876 1404
rect 4124 2136 4132 2144
rect 4060 2076 4068 2084
rect 4332 2896 4340 2904
rect 4348 2896 4356 2904
rect 4364 2856 4372 2864
rect 4316 2736 4324 2744
rect 4508 2956 4516 2964
rect 4492 2916 4500 2924
rect 4508 2916 4516 2924
rect 4492 2816 4500 2824
rect 4419 2806 4427 2814
rect 4429 2806 4437 2814
rect 4439 2806 4447 2814
rect 4449 2806 4457 2814
rect 4459 2806 4467 2814
rect 4469 2806 4477 2814
rect 4508 2796 4516 2804
rect 4588 3356 4596 3364
rect 4652 3356 4660 3364
rect 4652 3296 4660 3304
rect 4636 3256 4644 3264
rect 4748 3596 4756 3604
rect 4780 3596 4788 3604
rect 4732 3476 4740 3484
rect 4748 3396 4756 3404
rect 4700 3376 4708 3384
rect 4844 3616 4852 3624
rect 4860 3616 4868 3624
rect 4828 3596 4836 3604
rect 4908 3856 4916 3864
rect 4876 3536 4884 3544
rect 4956 3936 4964 3944
rect 5020 4076 5028 4084
rect 5004 3956 5012 3964
rect 5020 3956 5028 3964
rect 4988 3916 4996 3924
rect 5068 4496 5076 4504
rect 5148 4496 5156 4504
rect 5212 4596 5220 4604
rect 5196 4576 5204 4584
rect 5340 4676 5348 4684
rect 5404 4676 5412 4684
rect 5308 4616 5316 4624
rect 5324 4556 5332 4564
rect 5388 4616 5396 4624
rect 5244 4536 5252 4544
rect 5260 4536 5268 4544
rect 5180 4436 5188 4444
rect 5132 4356 5140 4364
rect 5084 4316 5092 4324
rect 5100 4236 5108 4244
rect 5084 4216 5092 4224
rect 5116 4176 5124 4184
rect 5068 4116 5076 4124
rect 5068 3996 5076 4004
rect 5052 3976 5060 3984
rect 5036 3936 5044 3944
rect 4972 3876 4980 3884
rect 4940 3856 4948 3864
rect 5036 3856 5044 3864
rect 5164 4256 5172 4264
rect 5228 4516 5236 4524
rect 5324 4518 5332 4524
rect 5324 4516 5332 4518
rect 5356 4496 5364 4504
rect 5260 4436 5268 4444
rect 5244 4416 5252 4424
rect 5196 4316 5204 4324
rect 5212 4296 5220 4304
rect 5372 4476 5380 4484
rect 5356 4456 5364 4464
rect 5292 4396 5300 4404
rect 5356 4396 5364 4404
rect 5276 4256 5284 4264
rect 5212 4236 5220 4244
rect 5324 4236 5332 4244
rect 5180 4176 5188 4184
rect 5180 4136 5188 4144
rect 5228 4136 5236 4144
rect 5340 4196 5348 4204
rect 5276 4156 5284 4164
rect 5148 4116 5156 4124
rect 5260 4116 5268 4124
rect 5180 4056 5188 4064
rect 5196 4056 5204 4064
rect 5116 4036 5124 4044
rect 5084 3936 5092 3944
rect 5164 3896 5172 3904
rect 5116 3876 5124 3884
rect 5164 3876 5172 3884
rect 5100 3856 5108 3864
rect 4940 3756 4948 3764
rect 4972 3756 4980 3764
rect 5068 3756 5076 3764
rect 4924 3616 4932 3624
rect 5052 3736 5060 3744
rect 5100 3796 5108 3804
rect 5116 3776 5124 3784
rect 5132 3736 5140 3744
rect 5100 3716 5108 3724
rect 4972 3676 4980 3684
rect 5164 3676 5172 3684
rect 4924 3536 4932 3544
rect 4940 3536 4948 3544
rect 4908 3516 4916 3524
rect 4812 3476 4820 3484
rect 4860 3476 4868 3484
rect 4956 3476 4964 3484
rect 4796 3396 4804 3404
rect 4732 3356 4740 3364
rect 4748 3336 4756 3344
rect 4780 3316 4788 3324
rect 4764 3296 4772 3304
rect 4988 3616 4996 3624
rect 5116 3616 5124 3624
rect 5164 3596 5172 3604
rect 5004 3476 5012 3484
rect 4828 3436 4836 3444
rect 4812 3356 4820 3364
rect 4828 3316 4836 3324
rect 4716 3276 4724 3284
rect 4796 3276 4804 3284
rect 4700 3256 4708 3264
rect 4716 3256 4724 3264
rect 4668 3176 4676 3184
rect 4604 3156 4612 3164
rect 4716 3156 4724 3164
rect 4636 3116 4644 3124
rect 4716 3116 4724 3124
rect 4748 3116 4756 3124
rect 4572 3096 4580 3104
rect 4700 3096 4708 3104
rect 4732 3076 4740 3084
rect 4796 3076 4804 3084
rect 4588 3056 4596 3064
rect 4684 3056 4692 3064
rect 4716 3056 4724 3064
rect 4764 2976 4772 2984
rect 4556 2936 4564 2944
rect 4700 2956 4708 2964
rect 4732 2956 4740 2964
rect 4924 3436 4932 3444
rect 4940 3436 4948 3444
rect 4876 3376 4884 3384
rect 4860 3176 4868 3184
rect 4908 3376 4916 3384
rect 4940 3376 4948 3384
rect 4924 3336 4932 3344
rect 4892 3316 4900 3324
rect 4924 3316 4932 3324
rect 4892 3296 4900 3304
rect 4892 3276 4900 3284
rect 4908 3036 4916 3044
rect 4892 3016 4900 3024
rect 4876 2976 4884 2984
rect 4844 2956 4852 2964
rect 4940 3296 4948 3304
rect 5004 3456 5012 3464
rect 4972 3376 4980 3384
rect 4956 3276 4964 3284
rect 4972 3276 4980 3284
rect 5020 3436 5028 3444
rect 5036 3436 5044 3444
rect 5068 3436 5076 3444
rect 5100 3436 5108 3444
rect 5036 3376 5044 3384
rect 5020 3316 5028 3324
rect 5100 3396 5108 3404
rect 5116 3376 5124 3384
rect 5084 3356 5092 3364
rect 5116 3336 5124 3344
rect 5180 3396 5188 3404
rect 5244 3996 5252 4004
rect 5212 3976 5220 3984
rect 5388 4376 5396 4384
rect 5372 4276 5380 4284
rect 5532 4976 5540 4984
rect 5500 4876 5508 4884
rect 5548 4876 5556 4884
rect 5580 5036 5588 5044
rect 5596 5036 5604 5044
rect 5564 4836 5572 4844
rect 5564 4716 5572 4724
rect 5500 4636 5508 4644
rect 5452 4576 5460 4584
rect 5532 4636 5540 4644
rect 5484 4536 5492 4544
rect 5468 4516 5476 4524
rect 5452 4456 5460 4464
rect 5468 4436 5476 4444
rect 5468 4316 5476 4324
rect 5532 4516 5540 4524
rect 5548 4516 5556 4524
rect 5500 4436 5508 4444
rect 5500 4416 5508 4424
rect 5548 4396 5556 4404
rect 5580 4636 5588 4644
rect 5580 4596 5588 4604
rect 5596 4576 5604 4584
rect 5644 5316 5652 5324
rect 5724 5316 5732 5324
rect 5852 5256 5860 5264
rect 5708 5236 5716 5244
rect 5868 5196 5876 5204
rect 5724 5076 5732 5084
rect 5756 5076 5764 5084
rect 5660 5056 5668 5064
rect 5644 4916 5652 4924
rect 5644 4896 5652 4904
rect 5772 5036 5780 5044
rect 5708 5016 5716 5024
rect 5676 4956 5684 4964
rect 5788 4996 5796 5004
rect 5740 4956 5748 4964
rect 5756 4916 5764 4924
rect 5724 4896 5732 4904
rect 5740 4896 5748 4904
rect 5676 4876 5684 4884
rect 5692 4776 5700 4784
rect 5740 4776 5748 4784
rect 5628 4636 5636 4644
rect 5612 4536 5620 4544
rect 5676 4576 5684 4584
rect 5580 4436 5588 4444
rect 5596 4436 5604 4444
rect 5580 4416 5588 4424
rect 5564 4376 5572 4384
rect 5516 4356 5524 4364
rect 5516 4336 5524 4344
rect 5548 4336 5556 4344
rect 5532 4316 5540 4324
rect 5500 4296 5508 4304
rect 5420 4276 5428 4284
rect 5404 4256 5412 4264
rect 5436 4256 5444 4264
rect 5388 4196 5396 4204
rect 5372 4116 5380 4124
rect 5276 4076 5284 4084
rect 5308 4076 5316 4084
rect 5420 4136 5428 4144
rect 5404 3936 5412 3944
rect 5260 3896 5268 3904
rect 5324 3896 5332 3904
rect 5372 3896 5380 3904
rect 5228 3876 5236 3884
rect 5324 3876 5332 3884
rect 5212 3856 5220 3864
rect 5292 3856 5300 3864
rect 5372 3856 5380 3864
rect 5388 3836 5396 3844
rect 5228 3796 5236 3804
rect 5260 3776 5268 3784
rect 5340 3776 5348 3784
rect 5404 3776 5412 3784
rect 5308 3716 5316 3724
rect 5228 3616 5236 3624
rect 5292 3696 5300 3704
rect 5324 3696 5332 3704
rect 5228 3596 5236 3604
rect 5244 3596 5252 3604
rect 5276 3556 5284 3564
rect 5260 3516 5268 3524
rect 5212 3456 5220 3464
rect 5196 3336 5204 3344
rect 5068 3316 5076 3324
rect 5164 3316 5172 3324
rect 5036 3296 5044 3304
rect 5084 3276 5092 3284
rect 5212 3276 5220 3284
rect 4988 3216 4996 3224
rect 4956 3196 4964 3204
rect 5068 3176 5076 3184
rect 5020 3136 5028 3144
rect 5036 3136 5044 3144
rect 5052 3136 5060 3144
rect 4940 3076 4948 3084
rect 4940 3036 4948 3044
rect 4828 2936 4836 2944
rect 4620 2916 4628 2924
rect 4652 2916 4660 2924
rect 4716 2916 4724 2924
rect 4844 2916 4852 2924
rect 4540 2876 4548 2884
rect 4636 2876 4644 2884
rect 4556 2796 4564 2804
rect 4540 2736 4548 2744
rect 4524 2716 4532 2724
rect 4412 2696 4420 2704
rect 4588 2696 4596 2704
rect 4604 2696 4612 2704
rect 4300 2656 4308 2664
rect 4332 2656 4340 2664
rect 4348 2656 4356 2664
rect 4284 2556 4292 2564
rect 4316 2556 4324 2564
rect 4300 2536 4308 2544
rect 4252 2516 4260 2524
rect 4268 2516 4276 2524
rect 4380 2656 4388 2664
rect 4524 2576 4532 2584
rect 4412 2556 4420 2564
rect 4556 2556 4564 2564
rect 4380 2496 4388 2504
rect 4332 2416 4340 2424
rect 4316 2356 4324 2364
rect 4252 2296 4260 2304
rect 4300 2296 4308 2304
rect 4188 2076 4196 2084
rect 4012 2036 4020 2044
rect 4140 2036 4148 2044
rect 4028 1976 4036 1984
rect 4044 1976 4052 1984
rect 4012 1916 4020 1924
rect 4060 1936 4068 1944
rect 4140 1936 4148 1944
rect 4028 1896 4036 1904
rect 4028 1876 4036 1884
rect 4012 1816 4020 1824
rect 4092 1916 4100 1924
rect 4268 2156 4276 2164
rect 4300 2156 4308 2164
rect 4268 2136 4276 2144
rect 4316 1956 4324 1964
rect 4236 1936 4244 1944
rect 4220 1896 4228 1904
rect 4092 1876 4100 1884
rect 4156 1876 4164 1884
rect 4060 1856 4068 1864
rect 4092 1836 4100 1844
rect 4028 1716 4036 1724
rect 4204 1856 4212 1864
rect 4236 1856 4244 1864
rect 4188 1836 4196 1844
rect 4124 1716 4132 1724
rect 4108 1696 4116 1704
rect 4044 1676 4052 1684
rect 4092 1676 4100 1684
rect 3996 1636 4004 1644
rect 3980 1576 3988 1584
rect 3884 1376 3892 1384
rect 3836 1336 3844 1344
rect 3980 1456 3988 1464
rect 3916 1336 3924 1344
rect 3964 1336 3972 1344
rect 3932 1256 3940 1264
rect 3932 1236 3940 1244
rect 3660 1136 3668 1144
rect 3708 1096 3716 1104
rect 3756 1096 3764 1104
rect 3884 1096 3892 1104
rect 3900 1102 3908 1104
rect 3900 1096 3908 1102
rect 3692 1076 3700 1084
rect 3756 1076 3764 1084
rect 3724 1056 3732 1064
rect 3644 1036 3652 1044
rect 3692 1036 3700 1044
rect 3740 1036 3748 1044
rect 3660 996 3668 1004
rect 3628 956 3636 964
rect 3516 856 3524 864
rect 3612 856 3620 864
rect 3548 836 3556 844
rect 3564 716 3572 724
rect 3644 796 3652 804
rect 3644 736 3652 744
rect 3804 976 3812 984
rect 3708 936 3716 944
rect 3772 936 3780 944
rect 3708 916 3716 924
rect 3756 916 3764 924
rect 3724 836 3732 844
rect 3692 756 3700 764
rect 3692 716 3700 724
rect 3756 676 3764 684
rect 3676 656 3684 664
rect 3564 636 3572 644
rect 3532 616 3540 624
rect 3548 516 3556 524
rect 3516 496 3524 504
rect 3532 476 3540 484
rect 3532 436 3540 444
rect 3468 316 3476 324
rect 3516 316 3524 324
rect 3452 296 3460 304
rect 3372 256 3380 264
rect 3356 176 3364 184
rect 3340 156 3348 164
rect 3132 136 3140 144
rect 3308 136 3316 144
rect 3500 276 3508 284
rect 3580 536 3588 544
rect 3676 636 3684 644
rect 3772 576 3780 584
rect 3708 556 3716 564
rect 3612 516 3620 524
rect 3628 516 3636 524
rect 3836 956 3844 964
rect 3836 936 3844 944
rect 3900 1016 3908 1024
rect 3996 1356 4004 1364
rect 4012 1296 4020 1304
rect 4012 1196 4020 1204
rect 3980 1116 3988 1124
rect 3996 1116 4004 1124
rect 4028 1116 4036 1124
rect 4156 1596 4164 1604
rect 4092 1556 4100 1564
rect 4076 1476 4084 1484
rect 4076 1356 4084 1364
rect 4108 1516 4116 1524
rect 4172 1516 4180 1524
rect 4172 1436 4180 1444
rect 4284 1916 4292 1924
rect 4268 1876 4276 1884
rect 4220 1836 4228 1844
rect 4252 1836 4260 1844
rect 4204 1776 4212 1784
rect 4220 1756 4228 1764
rect 4204 1716 4212 1724
rect 4236 1616 4244 1624
rect 4252 1576 4260 1584
rect 4236 1476 4244 1484
rect 4236 1436 4244 1444
rect 4140 1296 4148 1304
rect 4076 1256 4084 1264
rect 4092 1256 4100 1264
rect 4060 1136 4068 1144
rect 4044 1096 4052 1104
rect 3964 1076 3972 1084
rect 3964 976 3972 984
rect 3900 936 3908 944
rect 3820 916 3828 924
rect 3884 916 3892 924
rect 3852 896 3860 904
rect 3916 896 3924 904
rect 3948 896 3956 904
rect 3820 856 3828 864
rect 3884 816 3892 824
rect 3884 796 3892 804
rect 3820 702 3828 704
rect 3820 696 3828 702
rect 3852 656 3860 664
rect 3820 636 3828 644
rect 3788 536 3796 544
rect 3740 516 3748 524
rect 3804 516 3812 524
rect 3852 576 3860 584
rect 3868 556 3876 564
rect 3836 536 3844 544
rect 3644 476 3652 484
rect 3676 476 3684 484
rect 3692 396 3700 404
rect 3660 376 3668 384
rect 3580 356 3588 364
rect 3644 356 3652 364
rect 3660 356 3668 364
rect 3580 316 3588 324
rect 3692 316 3700 324
rect 3628 276 3636 284
rect 3708 276 3716 284
rect 3724 276 3732 284
rect 3580 256 3588 264
rect 3452 216 3460 224
rect 3484 156 3492 164
rect 3692 156 3700 164
rect 3436 136 3444 144
rect 3884 436 3892 444
rect 3836 396 3844 404
rect 3852 396 3860 404
rect 3772 256 3780 264
rect 3324 116 3332 124
rect 3660 118 3668 124
rect 3660 116 3668 118
rect 3756 116 3764 124
rect 2316 96 2324 104
rect 2348 96 2356 104
rect 2364 96 2372 104
rect 2444 96 2452 104
rect 2476 96 2484 104
rect 2556 96 2564 104
rect 2636 96 2644 104
rect 3068 96 3076 104
rect 3132 96 3140 104
rect 3212 96 3220 104
rect 3308 96 3316 104
rect 3356 96 3364 104
rect 1772 76 1780 84
rect 2540 76 2548 84
rect 3820 316 3828 324
rect 3916 876 3924 884
rect 3916 716 3924 724
rect 3916 696 3924 704
rect 3932 676 3940 684
rect 3932 636 3940 644
rect 3916 596 3924 604
rect 3964 676 3972 684
rect 3964 656 3972 664
rect 3916 396 3924 404
rect 3900 356 3908 364
rect 3900 276 3908 284
rect 3852 256 3860 264
rect 3868 176 3876 184
rect 3948 316 3956 324
rect 4028 956 4036 964
rect 3996 876 4004 884
rect 3996 836 4004 844
rect 4028 756 4036 764
rect 4172 1196 4180 1204
rect 4204 1176 4212 1184
rect 4284 1836 4292 1844
rect 4300 1816 4308 1824
rect 4316 1816 4324 1824
rect 4348 2376 4356 2384
rect 4364 2316 4372 2324
rect 4380 2316 4388 2324
rect 4652 2796 4660 2804
rect 4652 2736 4660 2744
rect 4908 2796 4916 2804
rect 4860 2736 4868 2744
rect 4636 2696 4644 2704
rect 4668 2696 4676 2704
rect 4748 2696 4756 2704
rect 4620 2656 4628 2664
rect 4572 2536 4580 2544
rect 4492 2456 4500 2464
rect 4524 2456 4532 2464
rect 4419 2406 4427 2414
rect 4429 2406 4437 2414
rect 4439 2406 4447 2414
rect 4449 2406 4457 2414
rect 4459 2406 4467 2414
rect 4469 2406 4477 2414
rect 4460 2376 4468 2384
rect 4428 2276 4436 2284
rect 4380 2256 4388 2264
rect 4396 2176 4404 2184
rect 4428 2176 4436 2184
rect 4652 2576 4660 2584
rect 4780 2716 4788 2724
rect 4844 2716 4852 2724
rect 4796 2696 4804 2704
rect 4764 2656 4772 2664
rect 4700 2616 4708 2624
rect 4732 2616 4740 2624
rect 4732 2596 4740 2604
rect 4764 2536 4772 2544
rect 4604 2516 4612 2524
rect 4668 2516 4676 2524
rect 4780 2496 4788 2504
rect 4588 2456 4596 2464
rect 4732 2456 4740 2464
rect 4700 2376 4708 2384
rect 4716 2376 4724 2384
rect 4492 2356 4500 2364
rect 4572 2336 4580 2344
rect 4620 2336 4628 2344
rect 4492 2296 4500 2304
rect 4476 2276 4484 2284
rect 4492 2256 4500 2264
rect 4492 2176 4500 2184
rect 4364 2096 4372 2104
rect 4364 2076 4372 2084
rect 4396 2076 4404 2084
rect 4396 2016 4404 2024
rect 4419 2006 4427 2014
rect 4429 2006 4437 2014
rect 4439 2006 4447 2014
rect 4449 2006 4457 2014
rect 4459 2006 4467 2014
rect 4469 2006 4477 2014
rect 4524 2156 4532 2164
rect 4556 2136 4564 2144
rect 4524 2116 4532 2124
rect 4540 2116 4548 2124
rect 4348 1956 4356 1964
rect 4348 1916 4356 1924
rect 4492 1956 4500 1964
rect 4508 1956 4516 1964
rect 4540 2076 4548 2084
rect 4572 1996 4580 2004
rect 4556 1936 4564 1944
rect 4508 1896 4516 1904
rect 4524 1896 4532 1904
rect 4348 1816 4356 1824
rect 4332 1796 4340 1804
rect 4540 1876 4548 1884
rect 4604 2016 4612 2024
rect 4636 2296 4644 2304
rect 4684 2296 4692 2304
rect 4636 2276 4644 2284
rect 4700 2276 4708 2284
rect 4748 2436 4756 2444
rect 4652 2136 4660 2144
rect 4716 2136 4724 2144
rect 4636 2116 4644 2124
rect 4620 1976 4628 1984
rect 4588 1916 4596 1924
rect 4620 1916 4628 1924
rect 4636 1916 4644 1924
rect 4588 1896 4596 1904
rect 4652 1896 4660 1904
rect 4604 1876 4612 1884
rect 4572 1856 4580 1864
rect 4620 1836 4628 1844
rect 4396 1816 4404 1824
rect 4316 1776 4324 1784
rect 4332 1776 4340 1784
rect 4284 1456 4292 1464
rect 4396 1736 4404 1744
rect 4620 1816 4628 1824
rect 4588 1796 4596 1804
rect 4556 1756 4564 1764
rect 4636 1776 4644 1784
rect 4492 1716 4500 1724
rect 4556 1716 4564 1724
rect 4716 2096 4724 2104
rect 4732 2096 4740 2104
rect 4828 2656 4836 2664
rect 4876 2716 4884 2724
rect 4908 2716 4916 2724
rect 4956 2996 4964 3004
rect 5004 2996 5012 3004
rect 5004 2956 5012 2964
rect 4988 2916 4996 2924
rect 4988 2896 4996 2904
rect 4972 2776 4980 2784
rect 4940 2696 4948 2704
rect 4972 2696 4980 2704
rect 4860 2656 4868 2664
rect 4924 2656 4932 2664
rect 4972 2656 4980 2664
rect 4828 2596 4836 2604
rect 4844 2596 4852 2604
rect 4876 2596 4884 2604
rect 4908 2596 4916 2604
rect 4844 2576 4852 2584
rect 4828 2536 4836 2544
rect 4860 2536 4868 2544
rect 4988 2576 4996 2584
rect 4940 2556 4948 2564
rect 4892 2536 4900 2544
rect 4988 2536 4996 2544
rect 4892 2516 4900 2524
rect 4972 2516 4980 2524
rect 5052 2936 5060 2944
rect 5036 2896 5044 2904
rect 5052 2816 5060 2824
rect 5036 2796 5044 2804
rect 5020 2736 5028 2744
rect 5036 2716 5044 2724
rect 5228 3216 5236 3224
rect 5164 3176 5172 3184
rect 5148 3136 5156 3144
rect 5276 3396 5284 3404
rect 5260 3136 5268 3144
rect 5228 3056 5236 3064
rect 5116 3036 5124 3044
rect 5132 3036 5140 3044
rect 5100 3016 5108 3024
rect 5100 2916 5108 2924
rect 5132 2816 5140 2824
rect 5244 3036 5252 3044
rect 5260 2996 5268 3004
rect 5164 2916 5172 2924
rect 5180 2876 5188 2884
rect 5212 2876 5220 2884
rect 5116 2796 5124 2804
rect 5148 2796 5156 2804
rect 5068 2736 5076 2744
rect 5084 2736 5092 2744
rect 5084 2716 5092 2724
rect 5036 2696 5044 2704
rect 5020 2676 5028 2684
rect 4796 2456 4804 2464
rect 4908 2456 4916 2464
rect 4876 2436 4884 2444
rect 4780 2396 4788 2404
rect 4796 2356 4804 2364
rect 4844 2302 4852 2304
rect 4844 2296 4852 2302
rect 4844 2276 4852 2284
rect 4844 2236 4852 2244
rect 4908 2396 4916 2404
rect 4972 2376 4980 2384
rect 4924 2356 4932 2364
rect 4940 2316 4948 2324
rect 4956 2316 4964 2324
rect 4908 2276 4916 2284
rect 4908 2176 4916 2184
rect 4764 2116 4772 2124
rect 4860 2116 4868 2124
rect 4828 2096 4836 2104
rect 4812 2016 4820 2024
rect 4748 1976 4756 1984
rect 4860 1976 4868 1984
rect 4780 1956 4788 1964
rect 4668 1876 4676 1884
rect 4652 1736 4660 1744
rect 4716 1916 4724 1924
rect 4732 1896 4740 1904
rect 4764 1896 4772 1904
rect 4716 1836 4724 1844
rect 4700 1776 4708 1784
rect 4540 1696 4548 1704
rect 4572 1696 4580 1704
rect 4636 1676 4644 1684
rect 4556 1656 4564 1664
rect 4588 1656 4596 1664
rect 4668 1716 4676 1724
rect 4668 1676 4676 1684
rect 4492 1616 4500 1624
rect 4419 1606 4427 1614
rect 4429 1606 4437 1614
rect 4439 1606 4447 1614
rect 4449 1606 4457 1614
rect 4459 1606 4467 1614
rect 4469 1606 4477 1614
rect 4364 1596 4372 1604
rect 4460 1536 4468 1544
rect 4380 1516 4388 1524
rect 4412 1516 4420 1524
rect 4332 1496 4340 1504
rect 4364 1496 4372 1504
rect 4316 1396 4324 1404
rect 4300 1356 4308 1364
rect 4268 1236 4276 1244
rect 4156 1136 4164 1144
rect 4236 1136 4244 1144
rect 4172 1116 4180 1124
rect 4140 1096 4148 1104
rect 4156 1076 4164 1084
rect 4108 996 4116 1004
rect 4348 1236 4356 1244
rect 4428 1416 4436 1424
rect 4396 1356 4404 1364
rect 4700 1676 4708 1684
rect 4716 1616 4724 1624
rect 4604 1576 4612 1584
rect 4652 1576 4660 1584
rect 4684 1576 4692 1584
rect 4524 1496 4532 1504
rect 4540 1496 4548 1504
rect 4604 1496 4612 1504
rect 4508 1476 4516 1484
rect 4524 1476 4532 1484
rect 4508 1456 4516 1464
rect 4492 1436 4500 1444
rect 4716 1476 4724 1484
rect 4620 1436 4628 1444
rect 4652 1436 4660 1444
rect 4668 1436 4676 1444
rect 4700 1456 4708 1464
rect 4812 1936 4820 1944
rect 4796 1836 4804 1844
rect 4828 1916 4836 1924
rect 4892 2116 4900 2124
rect 4892 1976 4900 1984
rect 4940 2156 4948 2164
rect 4972 2276 4980 2284
rect 4972 2236 4980 2244
rect 4956 2136 4964 2144
rect 4908 1956 4916 1964
rect 4876 1936 4884 1944
rect 4972 2096 4980 2104
rect 5004 2416 5012 2424
rect 5052 2656 5060 2664
rect 5084 2676 5092 2684
rect 5148 2716 5156 2724
rect 5212 2716 5220 2724
rect 5244 2916 5252 2924
rect 5372 3676 5380 3684
rect 5356 3596 5364 3604
rect 5340 3536 5348 3544
rect 5356 3536 5364 3544
rect 5340 3436 5348 3444
rect 5388 3536 5396 3544
rect 5388 3476 5396 3484
rect 5452 4196 5460 4204
rect 5596 4396 5604 4404
rect 5628 4456 5636 4464
rect 5628 4436 5636 4444
rect 5612 4356 5620 4364
rect 5628 4356 5636 4364
rect 5612 4296 5620 4304
rect 5628 4296 5636 4304
rect 5564 4276 5572 4284
rect 5580 4276 5588 4284
rect 5532 4236 5540 4244
rect 5516 4176 5524 4184
rect 5468 4136 5476 4144
rect 5468 4096 5476 4104
rect 5484 4076 5492 4084
rect 5548 4096 5556 4104
rect 5532 3936 5540 3944
rect 5516 3896 5524 3904
rect 5468 3836 5476 3844
rect 5452 3736 5460 3744
rect 5532 3816 5540 3824
rect 5532 3776 5540 3784
rect 5660 4516 5668 4524
rect 5676 4516 5684 4524
rect 5660 4436 5668 4444
rect 5724 4676 5732 4684
rect 5852 5096 5860 5104
rect 5852 4976 5860 4984
rect 5852 4936 5860 4944
rect 5836 4876 5844 4884
rect 5852 4876 5860 4884
rect 5820 4776 5828 4784
rect 5820 4716 5828 4724
rect 5820 4676 5828 4684
rect 5756 4616 5764 4624
rect 5772 4616 5780 4624
rect 5756 4576 5764 4584
rect 5708 4536 5716 4544
rect 5724 4456 5732 4464
rect 5868 4816 5876 4824
rect 5852 4736 5860 4744
rect 5804 4596 5812 4604
rect 5836 4596 5844 4604
rect 5820 4536 5828 4544
rect 5788 4516 5796 4524
rect 5820 4456 5828 4464
rect 5756 4396 5764 4404
rect 5772 4396 5780 4404
rect 5692 4336 5700 4344
rect 5756 4336 5764 4344
rect 5788 4336 5796 4344
rect 5708 4296 5716 4304
rect 5788 4296 5796 4304
rect 5676 4276 5684 4284
rect 5740 4256 5748 4264
rect 5788 4256 5796 4264
rect 5900 5356 5908 5364
rect 6060 5336 6068 5344
rect 5916 5316 5924 5324
rect 5932 5296 5940 5304
rect 6028 5296 6036 5304
rect 6140 5256 6148 5264
rect 6044 5196 6052 5204
rect 6028 5156 6036 5164
rect 6060 5156 6068 5164
rect 5900 5096 5908 5104
rect 6012 5096 6020 5104
rect 5980 5076 5988 5084
rect 5923 5006 5931 5014
rect 5933 5006 5941 5014
rect 5943 5006 5951 5014
rect 5953 5006 5961 5014
rect 5963 5006 5971 5014
rect 5973 5006 5981 5014
rect 5900 4936 5908 4944
rect 6012 4996 6020 5004
rect 6140 5116 6148 5124
rect 6476 5356 6484 5364
rect 6364 5336 6372 5344
rect 6428 5336 6436 5344
rect 6076 5096 6084 5104
rect 6172 5096 6180 5104
rect 6092 5036 6100 5044
rect 6060 4996 6068 5004
rect 6076 4996 6084 5004
rect 6012 4956 6020 4964
rect 6044 4956 6052 4964
rect 5916 4916 5924 4924
rect 5932 4896 5940 4904
rect 5980 4856 5988 4864
rect 5996 4816 6004 4824
rect 5868 4716 5876 4724
rect 5884 4716 5892 4724
rect 5900 4696 5908 4704
rect 5884 4656 5892 4664
rect 5868 4616 5876 4624
rect 5868 4596 5876 4604
rect 5923 4606 5931 4614
rect 5933 4606 5941 4614
rect 5943 4606 5951 4614
rect 5953 4606 5961 4614
rect 5963 4606 5971 4614
rect 5973 4606 5981 4614
rect 5900 4576 5908 4584
rect 5916 4576 5924 4584
rect 5884 4556 5892 4564
rect 5852 4516 5860 4524
rect 5884 4476 5892 4484
rect 6076 4916 6084 4924
rect 6108 4896 6116 4904
rect 6044 4776 6052 4784
rect 6012 4676 6020 4684
rect 6012 4616 6020 4624
rect 5932 4456 5940 4464
rect 5996 4456 6004 4464
rect 6172 5056 6180 5064
rect 6140 4836 6148 4844
rect 6156 4796 6164 4804
rect 6124 4756 6132 4764
rect 6204 5116 6212 5124
rect 6236 5116 6244 5124
rect 6252 5056 6260 5064
rect 6220 4996 6228 5004
rect 6236 4996 6244 5004
rect 6284 5096 6292 5104
rect 6332 5096 6340 5104
rect 6300 5036 6308 5044
rect 6316 5036 6324 5044
rect 6348 5036 6356 5044
rect 6268 4956 6276 4964
rect 6332 4956 6340 4964
rect 6268 4916 6276 4924
rect 6284 4916 6292 4924
rect 6284 4896 6292 4904
rect 6252 4856 6260 4864
rect 6236 4836 6244 4844
rect 6188 4796 6196 4804
rect 6300 4776 6308 4784
rect 6172 4736 6180 4744
rect 6252 4716 6260 4724
rect 6268 4676 6276 4684
rect 6300 4676 6308 4684
rect 6108 4596 6116 4604
rect 6140 4596 6148 4604
rect 6108 4556 6116 4564
rect 6044 4536 6052 4544
rect 5916 4336 5924 4344
rect 5932 4336 5940 4344
rect 6012 4336 6020 4344
rect 6028 4336 6036 4344
rect 5836 4276 5844 4284
rect 5724 4236 5732 4244
rect 5788 4236 5796 4244
rect 5612 4136 5620 4144
rect 5644 4136 5652 4144
rect 5596 4036 5604 4044
rect 5596 3996 5604 4004
rect 5644 3936 5652 3944
rect 5628 3856 5636 3864
rect 5628 3796 5636 3804
rect 5676 4196 5684 4204
rect 5740 4196 5748 4204
rect 5804 4196 5812 4204
rect 5772 4156 5780 4164
rect 5740 4136 5748 4144
rect 5724 4036 5732 4044
rect 5708 3996 5716 4004
rect 5692 3956 5700 3964
rect 5692 3856 5700 3864
rect 5532 3716 5540 3724
rect 5484 3696 5492 3704
rect 5484 3676 5492 3684
rect 5436 3576 5444 3584
rect 5484 3576 5492 3584
rect 5500 3576 5508 3584
rect 5468 3536 5476 3544
rect 5452 3476 5460 3484
rect 5420 3456 5428 3464
rect 5404 3436 5412 3444
rect 5324 3376 5332 3384
rect 5356 3376 5364 3384
rect 5292 3116 5300 3124
rect 5420 3336 5428 3344
rect 5388 3316 5396 3324
rect 5404 3296 5412 3304
rect 5436 3276 5444 3284
rect 5356 3256 5364 3264
rect 5468 3436 5476 3444
rect 5468 3256 5476 3264
rect 5468 3196 5476 3204
rect 5516 3336 5524 3344
rect 5564 3676 5572 3684
rect 5548 3616 5556 3624
rect 5500 3296 5508 3304
rect 5532 3296 5540 3304
rect 5500 3256 5508 3264
rect 5484 3176 5492 3184
rect 5500 3136 5508 3144
rect 5516 3136 5524 3144
rect 5500 3116 5508 3124
rect 5324 3056 5332 3064
rect 5372 3076 5380 3084
rect 5372 2936 5380 2944
rect 5356 2916 5364 2924
rect 5276 2816 5284 2824
rect 5276 2736 5284 2744
rect 5084 2616 5092 2624
rect 5132 2616 5140 2624
rect 5164 2676 5172 2684
rect 5196 2676 5204 2684
rect 5212 2656 5220 2664
rect 5164 2616 5172 2624
rect 5180 2616 5188 2624
rect 5036 2536 5044 2544
rect 5068 2556 5076 2564
rect 5148 2576 5156 2584
rect 5100 2536 5108 2544
rect 5036 2496 5044 2504
rect 5036 2436 5044 2444
rect 5036 2376 5044 2384
rect 5020 2296 5028 2304
rect 5004 2276 5012 2284
rect 4844 1896 4852 1904
rect 4940 1896 4948 1904
rect 4828 1796 4836 1804
rect 4748 1696 4756 1704
rect 4780 1696 4788 1704
rect 4764 1676 4772 1684
rect 4748 1616 4756 1624
rect 4764 1556 4772 1564
rect 4748 1516 4756 1524
rect 4796 1676 4804 1684
rect 4876 1856 4884 1864
rect 5004 1796 5012 1804
rect 4908 1756 4916 1764
rect 4988 1716 4996 1724
rect 4892 1696 4900 1704
rect 4844 1676 4852 1684
rect 4924 1676 4932 1684
rect 4812 1616 4820 1624
rect 4812 1536 4820 1544
rect 4796 1476 4804 1484
rect 4812 1476 4820 1484
rect 4508 1416 4516 1424
rect 4556 1416 4564 1424
rect 4572 1416 4580 1424
rect 4444 1296 4452 1304
rect 4492 1296 4500 1304
rect 4412 1256 4420 1264
rect 4419 1206 4427 1214
rect 4429 1206 4437 1214
rect 4439 1206 4447 1214
rect 4449 1206 4457 1214
rect 4459 1206 4467 1214
rect 4469 1206 4477 1214
rect 4364 1176 4372 1184
rect 4364 1156 4372 1164
rect 4348 1136 4356 1144
rect 4380 1136 4388 1144
rect 4428 1136 4436 1144
rect 4220 1096 4228 1104
rect 4332 1096 4340 1104
rect 4412 1096 4420 1104
rect 4364 1076 4372 1084
rect 4252 1016 4260 1024
rect 4172 996 4180 1004
rect 4092 976 4100 984
rect 4124 976 4132 984
rect 4140 976 4148 984
rect 4188 976 4196 984
rect 4076 796 4084 804
rect 4060 756 4068 764
rect 3996 716 4004 724
rect 4044 716 4052 724
rect 4124 896 4132 904
rect 4140 896 4148 904
rect 4172 896 4180 904
rect 4172 836 4180 844
rect 4044 676 4052 684
rect 4076 676 4084 684
rect 4076 576 4084 584
rect 3996 518 4004 524
rect 3996 516 4004 518
rect 4060 396 4068 404
rect 3948 276 3956 284
rect 3980 276 3988 284
rect 3852 136 3860 144
rect 3884 136 3892 144
rect 3836 116 3844 124
rect 3868 116 3876 124
rect 3932 116 3940 124
rect 3852 96 3860 104
rect 3884 96 3892 104
rect 3804 56 3812 64
rect 3836 56 3844 64
rect 1411 6 1419 14
rect 1421 6 1429 14
rect 1431 6 1439 14
rect 1441 6 1449 14
rect 1451 6 1459 14
rect 1461 6 1469 14
rect 4172 696 4180 704
rect 4124 676 4132 684
rect 4204 956 4212 964
rect 4236 836 4244 844
rect 4364 1016 4372 1024
rect 4428 1016 4436 1024
rect 4284 976 4292 984
rect 4300 936 4308 944
rect 4284 916 4292 924
rect 4284 896 4292 904
rect 4492 976 4500 984
rect 4364 816 4372 824
rect 4236 696 4244 704
rect 4252 676 4260 684
rect 4188 636 4196 644
rect 4140 556 4148 564
rect 4236 536 4244 544
rect 4204 516 4212 524
rect 4252 476 4260 484
rect 4124 436 4132 444
rect 4108 396 4116 404
rect 4156 376 4164 384
rect 4172 276 4180 284
rect 4284 676 4292 684
rect 4396 916 4404 924
rect 4492 816 4500 824
rect 4419 806 4427 814
rect 4429 806 4437 814
rect 4439 806 4447 814
rect 4449 806 4457 814
rect 4459 806 4467 814
rect 4469 806 4477 814
rect 4652 1376 4660 1384
rect 4572 1336 4580 1344
rect 4588 1336 4596 1344
rect 4604 1316 4612 1324
rect 4636 1296 4644 1304
rect 4572 1236 4580 1244
rect 4588 1236 4596 1244
rect 4556 1216 4564 1224
rect 4572 1136 4580 1144
rect 4732 1376 4740 1384
rect 4764 1376 4772 1384
rect 4780 1376 4788 1384
rect 4732 1316 4740 1324
rect 4716 1276 4724 1284
rect 4668 1256 4676 1264
rect 4636 1196 4644 1204
rect 4636 1156 4644 1164
rect 4588 1096 4596 1104
rect 4588 1076 4596 1084
rect 4780 1336 4788 1344
rect 4796 1296 4804 1304
rect 4828 1436 4836 1444
rect 4972 1616 4980 1624
rect 4876 1556 4884 1564
rect 4940 1516 4948 1524
rect 4892 1496 4900 1504
rect 4844 1396 4852 1404
rect 4764 1216 4772 1224
rect 4780 1216 4788 1224
rect 4764 1196 4772 1204
rect 4684 1156 4692 1164
rect 4732 1156 4740 1164
rect 4748 1156 4756 1164
rect 4668 1136 4676 1144
rect 4540 1056 4548 1064
rect 4620 1056 4628 1064
rect 4556 956 4564 964
rect 4572 956 4580 964
rect 4524 916 4532 924
rect 4508 716 4516 724
rect 4540 676 4548 684
rect 4300 536 4308 544
rect 4316 536 4324 544
rect 4492 536 4500 544
rect 4604 716 4612 724
rect 4636 856 4644 864
rect 4668 1096 4676 1104
rect 4668 976 4676 984
rect 4588 616 4596 624
rect 4572 536 4580 544
rect 4284 516 4292 524
rect 4508 516 4516 524
rect 4300 456 4308 464
rect 4348 436 4356 444
rect 4419 406 4427 414
rect 4429 406 4437 414
rect 4439 406 4447 414
rect 4449 406 4457 414
rect 4459 406 4467 414
rect 4469 406 4477 414
rect 4268 356 4276 364
rect 4348 316 4356 324
rect 4252 276 4260 284
rect 4268 276 4276 284
rect 4300 276 4308 284
rect 4204 256 4212 264
rect 4236 256 4244 264
rect 4092 236 4100 244
rect 4204 236 4212 244
rect 4236 236 4244 244
rect 4284 256 4292 264
rect 4428 316 4436 324
rect 4396 276 4404 284
rect 4476 276 4484 284
rect 4556 276 4564 284
rect 4364 256 4372 264
rect 4412 256 4420 264
rect 4332 236 4340 244
rect 4284 196 4292 204
rect 4540 256 4548 264
rect 4076 156 4084 164
rect 4108 136 4116 144
rect 4380 136 4388 144
rect 4140 116 4148 124
rect 4188 116 4196 124
rect 4252 116 4260 124
rect 4348 118 4356 124
rect 4348 116 4356 118
rect 4076 96 4084 104
rect 4156 96 4164 104
rect 4060 36 4068 44
rect 4092 36 4100 44
rect 4060 16 4068 24
rect 4252 16 4260 24
rect 4419 6 4427 14
rect 4429 6 4437 14
rect 4439 6 4447 14
rect 4449 6 4457 14
rect 4459 6 4467 14
rect 4469 6 4477 14
rect 4620 616 4628 624
rect 4604 576 4612 584
rect 4620 496 4628 504
rect 4604 236 4612 244
rect 4572 136 4580 144
rect 4668 536 4676 544
rect 4652 496 4660 504
rect 4668 316 4676 324
rect 4636 256 4644 264
rect 4652 256 4660 264
rect 4668 236 4676 244
rect 4700 1096 4708 1104
rect 4732 1096 4740 1104
rect 4732 1076 4740 1084
rect 4780 1096 4788 1104
rect 4764 1076 4772 1084
rect 4748 1016 4756 1024
rect 4828 1256 4836 1264
rect 4844 1236 4852 1244
rect 4892 1416 4900 1424
rect 4940 1356 4948 1364
rect 5116 2496 5124 2504
rect 5068 2476 5076 2484
rect 5052 2356 5060 2364
rect 5084 2396 5092 2404
rect 5100 2396 5108 2404
rect 5052 2276 5060 2284
rect 5084 2236 5092 2244
rect 5084 2196 5092 2204
rect 5196 2596 5204 2604
rect 5164 2536 5172 2544
rect 5180 2496 5188 2504
rect 5308 2676 5316 2684
rect 5260 2596 5268 2604
rect 5244 2576 5252 2584
rect 5260 2576 5268 2584
rect 5132 2316 5140 2324
rect 5164 2316 5172 2324
rect 5228 2316 5236 2324
rect 5116 2296 5124 2304
rect 5132 2276 5140 2284
rect 5116 2196 5124 2204
rect 5308 2636 5316 2644
rect 5276 2456 5284 2464
rect 5260 2376 5268 2384
rect 5260 2336 5268 2344
rect 5244 2236 5252 2244
rect 5260 2236 5268 2244
rect 5212 2176 5220 2184
rect 5260 2176 5268 2184
rect 5100 2136 5108 2144
rect 5180 2136 5188 2144
rect 5132 2116 5140 2124
rect 5148 2116 5156 2124
rect 5068 2096 5076 2104
rect 5052 2076 5060 2084
rect 5100 2076 5108 2084
rect 5148 2076 5156 2084
rect 5164 2016 5172 2024
rect 5244 2096 5252 2104
rect 5228 2076 5236 2084
rect 5180 1976 5188 1984
rect 5212 1976 5220 1984
rect 5148 1896 5156 1904
rect 5292 2376 5300 2384
rect 5452 3076 5460 3084
rect 5420 3036 5428 3044
rect 5452 3036 5460 3044
rect 5436 2956 5444 2964
rect 5404 2916 5412 2924
rect 5420 2876 5428 2884
rect 5388 2736 5396 2744
rect 5516 3076 5524 3084
rect 5500 2916 5508 2924
rect 5676 3736 5684 3744
rect 5660 3716 5668 3724
rect 5676 3716 5684 3724
rect 5644 3656 5652 3664
rect 5580 3576 5588 3584
rect 5612 3576 5620 3584
rect 5596 3536 5604 3544
rect 5564 3496 5572 3504
rect 5580 3476 5588 3484
rect 5916 4296 5924 4304
rect 5948 4316 5956 4324
rect 5932 4256 5940 4264
rect 5948 4256 5956 4264
rect 5852 4156 5860 4164
rect 5868 4136 5876 4144
rect 5772 3896 5780 3904
rect 5756 3756 5764 3764
rect 5724 3696 5732 3704
rect 5692 3616 5700 3624
rect 5724 3616 5732 3624
rect 5660 3576 5668 3584
rect 5628 3496 5636 3504
rect 5628 3476 5636 3484
rect 5596 3436 5604 3444
rect 5756 3576 5764 3584
rect 5772 3556 5780 3564
rect 5820 3936 5828 3944
rect 5836 3936 5844 3944
rect 5820 3816 5828 3824
rect 5804 3776 5812 3784
rect 5804 3736 5812 3744
rect 5923 4206 5931 4214
rect 5933 4206 5941 4214
rect 5943 4206 5951 4214
rect 5953 4206 5961 4214
rect 5963 4206 5971 4214
rect 5973 4206 5981 4214
rect 6012 4216 6020 4224
rect 5996 4196 6004 4204
rect 6124 4516 6132 4524
rect 6092 4496 6100 4504
rect 6172 4616 6180 4624
rect 6076 4356 6084 4364
rect 6092 4356 6100 4364
rect 6140 4456 6148 4464
rect 6204 4576 6212 4584
rect 6220 4536 6228 4544
rect 6268 4536 6276 4544
rect 6220 4496 6228 4504
rect 6204 4456 6212 4464
rect 6044 4236 6052 4244
rect 6124 4296 6132 4304
rect 6188 4296 6196 4304
rect 6108 4256 6116 4264
rect 6156 4256 6164 4264
rect 6188 4256 6196 4264
rect 6092 4236 6100 4244
rect 6156 4236 6164 4244
rect 6172 4236 6180 4244
rect 6060 4216 6068 4224
rect 6092 4176 6100 4184
rect 5916 4156 5924 4164
rect 6028 4156 6036 4164
rect 6012 4136 6020 4144
rect 6044 4136 6052 4144
rect 5996 4116 6004 4124
rect 6124 4136 6132 4144
rect 6156 4116 6164 4124
rect 6124 4096 6132 4104
rect 6188 4076 6196 4084
rect 6156 4036 6164 4044
rect 6012 3996 6020 4004
rect 5900 3936 5908 3944
rect 5868 3916 5876 3924
rect 6012 3896 6020 3904
rect 5868 3856 5876 3864
rect 5884 3776 5892 3784
rect 5923 3806 5931 3814
rect 5933 3806 5941 3814
rect 5943 3806 5951 3814
rect 5953 3806 5961 3814
rect 5963 3806 5971 3814
rect 5973 3806 5981 3814
rect 5884 3696 5892 3704
rect 5900 3696 5908 3704
rect 5820 3616 5828 3624
rect 5852 3576 5860 3584
rect 5820 3536 5828 3544
rect 5756 3516 5764 3524
rect 5788 3516 5796 3524
rect 5852 3516 5860 3524
rect 5660 3416 5668 3424
rect 5692 3456 5700 3464
rect 5756 3496 5764 3504
rect 5724 3456 5732 3464
rect 5740 3456 5748 3464
rect 5804 3456 5812 3464
rect 5708 3436 5716 3444
rect 5676 3336 5684 3344
rect 5708 3336 5716 3344
rect 5580 3296 5588 3304
rect 5580 3276 5588 3284
rect 5612 3276 5620 3284
rect 5756 3436 5764 3444
rect 5772 3436 5780 3444
rect 5740 3416 5748 3424
rect 5772 3396 5780 3404
rect 5788 3396 5796 3404
rect 5788 3336 5796 3344
rect 5644 3316 5652 3324
rect 5660 3316 5668 3324
rect 5772 3316 5780 3324
rect 5580 3196 5588 3204
rect 5628 3196 5636 3204
rect 5644 3196 5652 3204
rect 5564 3116 5572 3124
rect 5612 3176 5620 3184
rect 5596 3076 5604 3084
rect 5596 3056 5604 3064
rect 5628 2956 5636 2964
rect 5564 2936 5572 2944
rect 5628 2916 5636 2924
rect 5532 2876 5540 2884
rect 5532 2736 5540 2744
rect 5468 2716 5476 2724
rect 5452 2696 5460 2704
rect 5356 2676 5364 2684
rect 5356 2576 5364 2584
rect 5356 2516 5364 2524
rect 5340 2456 5348 2464
rect 5324 2436 5332 2444
rect 5308 2356 5316 2364
rect 5404 2676 5412 2684
rect 5372 2476 5380 2484
rect 5436 2596 5444 2604
rect 5516 2676 5524 2684
rect 5516 2616 5524 2624
rect 5548 2696 5556 2704
rect 5532 2596 5540 2604
rect 5452 2556 5460 2564
rect 5436 2536 5444 2544
rect 5548 2556 5556 2564
rect 5452 2516 5460 2524
rect 5500 2516 5508 2524
rect 5532 2516 5540 2524
rect 5452 2496 5460 2504
rect 5484 2496 5492 2504
rect 5404 2456 5412 2464
rect 5468 2456 5476 2464
rect 5388 2436 5396 2444
rect 5356 2396 5364 2404
rect 5388 2356 5396 2364
rect 5452 2356 5460 2364
rect 5356 2296 5364 2304
rect 5436 2296 5444 2304
rect 5324 2236 5332 2244
rect 5372 2236 5380 2244
rect 5324 2156 5332 2164
rect 5516 2376 5524 2384
rect 5500 2296 5508 2304
rect 5548 2496 5556 2504
rect 5532 2356 5540 2364
rect 5836 3436 5844 3444
rect 5836 3416 5844 3424
rect 5852 3396 5860 3404
rect 5852 3356 5860 3364
rect 5916 3676 5924 3684
rect 5900 3516 5908 3524
rect 5916 3516 5924 3524
rect 5900 3476 5908 3484
rect 5820 3316 5828 3324
rect 5820 3276 5828 3284
rect 5836 3236 5844 3244
rect 5820 3176 5828 3184
rect 5724 3136 5732 3144
rect 5692 3096 5700 3104
rect 5788 3056 5796 3064
rect 5884 3336 5892 3344
rect 5884 3316 5892 3324
rect 5868 3256 5876 3264
rect 6012 3716 6020 3724
rect 6124 3936 6132 3944
rect 6076 3896 6084 3904
rect 6076 3856 6084 3864
rect 6092 3816 6100 3824
rect 6108 3776 6116 3784
rect 6060 3716 6068 3724
rect 6092 3716 6100 3724
rect 6028 3696 6036 3704
rect 5996 3676 6004 3684
rect 6028 3656 6036 3664
rect 6012 3496 6020 3504
rect 5932 3456 5940 3464
rect 5996 3416 6004 3424
rect 5923 3406 5931 3414
rect 5933 3406 5941 3414
rect 5943 3406 5951 3414
rect 5953 3406 5961 3414
rect 5963 3406 5971 3414
rect 5973 3406 5981 3414
rect 5964 3336 5972 3344
rect 6044 3616 6052 3624
rect 6060 3616 6068 3624
rect 6188 3996 6196 4004
rect 6188 3976 6196 3984
rect 6300 4496 6308 4504
rect 6236 4476 6244 4484
rect 6284 4316 6292 4324
rect 6348 4816 6356 4824
rect 6332 4756 6340 4764
rect 6332 4696 6340 4704
rect 6380 5276 6388 5284
rect 6396 5256 6404 5264
rect 6428 5236 6436 5244
rect 6396 5216 6404 5224
rect 6380 5116 6388 5124
rect 6460 5036 6468 5044
rect 6396 5016 6404 5024
rect 6444 4956 6452 4964
rect 6428 4936 6436 4944
rect 6460 4876 6468 4884
rect 6428 4856 6436 4864
rect 6620 5336 6628 5344
rect 6812 5336 6820 5344
rect 7228 5336 7236 5344
rect 6588 5276 6596 5284
rect 6620 5196 6628 5204
rect 6492 5156 6500 5164
rect 6652 5156 6660 5164
rect 6556 5136 6564 5144
rect 6524 5116 6532 5124
rect 6620 5116 6628 5124
rect 6716 5116 6724 5124
rect 6556 5076 6564 5084
rect 6636 5076 6644 5084
rect 6540 5056 6548 5064
rect 6572 5056 6580 5064
rect 6524 4956 6532 4964
rect 6492 4936 6500 4944
rect 6508 4896 6516 4904
rect 6524 4896 6532 4904
rect 6604 5016 6612 5024
rect 6588 4996 6596 5004
rect 6668 5016 6676 5024
rect 6652 4976 6660 4984
rect 6620 4956 6628 4964
rect 6588 4916 6596 4924
rect 6540 4856 6548 4864
rect 6476 4816 6484 4824
rect 6540 4816 6548 4824
rect 6380 4776 6388 4784
rect 6444 4736 6452 4744
rect 6332 4676 6340 4684
rect 6332 4596 6340 4604
rect 6364 4676 6372 4684
rect 6348 4516 6356 4524
rect 6492 4696 6500 4704
rect 6492 4656 6500 4664
rect 6476 4636 6484 4644
rect 6428 4616 6436 4624
rect 6396 4536 6404 4544
rect 6332 4476 6340 4484
rect 6332 4336 6340 4344
rect 6236 4296 6244 4304
rect 6268 4296 6276 4304
rect 6316 4296 6324 4304
rect 6316 4276 6324 4284
rect 6332 4256 6340 4264
rect 6316 4236 6324 4244
rect 6300 4196 6308 4204
rect 6332 4196 6340 4204
rect 6252 4176 6260 4184
rect 6316 4136 6324 4144
rect 6268 4116 6276 4124
rect 6236 4056 6244 4064
rect 6220 4016 6228 4024
rect 6252 4016 6260 4024
rect 6220 3996 6228 4004
rect 6236 3976 6244 3984
rect 6220 3936 6228 3944
rect 6172 3896 6180 3904
rect 6204 3896 6212 3904
rect 6156 3856 6164 3864
rect 6236 3856 6244 3864
rect 6172 3816 6180 3824
rect 6156 3796 6164 3804
rect 6172 3796 6180 3804
rect 6284 4096 6292 4104
rect 6300 4056 6308 4064
rect 6396 4516 6404 4524
rect 6380 4496 6388 4504
rect 6412 4476 6420 4484
rect 6396 4136 6404 4144
rect 6300 4036 6308 4044
rect 6316 4036 6324 4044
rect 6284 4016 6292 4024
rect 6332 3996 6340 4004
rect 6332 3896 6340 3904
rect 6268 3876 6276 3884
rect 6284 3876 6292 3884
rect 6300 3876 6308 3884
rect 6396 4116 6404 4124
rect 6364 4096 6372 4104
rect 6364 3916 6372 3924
rect 6268 3756 6276 3764
rect 6300 3756 6308 3764
rect 6348 3756 6356 3764
rect 6364 3756 6372 3764
rect 6140 3716 6148 3724
rect 6300 3736 6308 3744
rect 6236 3716 6244 3724
rect 6284 3716 6292 3724
rect 6124 3676 6132 3684
rect 6156 3616 6164 3624
rect 6092 3536 6100 3544
rect 6044 3456 6052 3464
rect 6028 3396 6036 3404
rect 6028 3336 6036 3344
rect 6172 3576 6180 3584
rect 6220 3676 6228 3684
rect 6252 3636 6260 3644
rect 6236 3576 6244 3584
rect 6220 3496 6228 3504
rect 6140 3456 6148 3464
rect 6204 3456 6212 3464
rect 6140 3416 6148 3424
rect 6076 3396 6084 3404
rect 6204 3396 6212 3404
rect 6188 3376 6196 3384
rect 6124 3336 6132 3344
rect 6172 3336 6180 3344
rect 6044 3296 6052 3304
rect 5996 3276 6004 3284
rect 6028 3276 6036 3284
rect 5996 3216 6004 3224
rect 5980 3176 5988 3184
rect 6028 3116 6036 3124
rect 5996 3096 6004 3104
rect 6284 3616 6292 3624
rect 6460 4336 6468 4344
rect 6460 4156 6468 4164
rect 6428 4116 6436 4124
rect 6476 4116 6484 4124
rect 6428 4076 6436 4084
rect 6460 4076 6468 4084
rect 6412 4056 6420 4064
rect 6412 3996 6420 4004
rect 6444 3976 6452 3984
rect 6396 3896 6404 3904
rect 6396 3876 6404 3884
rect 6380 3736 6388 3744
rect 6316 3676 6324 3684
rect 6332 3656 6340 3664
rect 6300 3536 6308 3544
rect 6428 3856 6436 3864
rect 6412 3736 6420 3744
rect 6332 3516 6340 3524
rect 6396 3516 6404 3524
rect 6476 3836 6484 3844
rect 6460 3756 6468 3764
rect 6428 3716 6436 3724
rect 6476 3716 6484 3724
rect 6428 3676 6436 3684
rect 6460 3676 6468 3684
rect 6460 3656 6468 3664
rect 6380 3496 6388 3504
rect 6348 3476 6356 3484
rect 6316 3396 6324 3404
rect 6428 3476 6436 3484
rect 6396 3456 6404 3464
rect 6300 3376 6308 3384
rect 6380 3376 6388 3384
rect 6396 3336 6404 3344
rect 6236 3316 6244 3324
rect 6140 3296 6148 3304
rect 6156 3296 6164 3304
rect 6076 3276 6084 3284
rect 5932 3076 5940 3084
rect 5852 3056 5860 3064
rect 5900 3056 5908 3064
rect 5836 3016 5844 3024
rect 5772 2956 5780 2964
rect 5660 2936 5668 2944
rect 5724 2936 5732 2944
rect 5772 2936 5780 2944
rect 5820 2936 5828 2944
rect 5660 2896 5668 2904
rect 5708 2896 5716 2904
rect 5628 2876 5636 2884
rect 5740 2876 5748 2884
rect 5580 2796 5588 2804
rect 5708 2716 5716 2724
rect 5932 3036 5940 3044
rect 6012 3036 6020 3044
rect 5996 3016 6004 3024
rect 5923 3006 5931 3014
rect 5933 3006 5941 3014
rect 5943 3006 5951 3014
rect 5953 3006 5961 3014
rect 5963 3006 5971 3014
rect 5973 3006 5981 3014
rect 5884 2956 5892 2964
rect 5836 2896 5844 2904
rect 5788 2796 5796 2804
rect 5788 2716 5796 2724
rect 5788 2696 5796 2704
rect 5740 2676 5748 2684
rect 5852 2676 5860 2684
rect 5644 2636 5652 2644
rect 5564 2476 5572 2484
rect 5612 2336 5620 2344
rect 5772 2636 5780 2644
rect 5836 2636 5844 2644
rect 5740 2556 5748 2564
rect 5852 2536 5860 2544
rect 5676 2518 5684 2524
rect 5676 2516 5684 2518
rect 5772 2516 5780 2524
rect 5772 2496 5780 2504
rect 5740 2456 5748 2464
rect 5660 2356 5668 2364
rect 5676 2356 5684 2364
rect 5660 2336 5668 2344
rect 5500 2256 5508 2264
rect 5564 2256 5572 2264
rect 5612 2276 5620 2284
rect 5484 2196 5492 2204
rect 5468 2176 5476 2184
rect 5420 2156 5428 2164
rect 5308 2096 5316 2104
rect 5388 2096 5396 2104
rect 5452 2116 5460 2124
rect 5340 2076 5348 2084
rect 5372 2076 5380 2084
rect 5404 2076 5412 2084
rect 5340 2016 5348 2024
rect 5436 2016 5444 2024
rect 5324 1976 5332 1984
rect 5372 1976 5380 1984
rect 5276 1796 5284 1804
rect 5292 1796 5300 1804
rect 5084 1756 5092 1764
rect 5148 1756 5156 1764
rect 5132 1736 5140 1744
rect 5068 1696 5076 1704
rect 5132 1676 5140 1684
rect 5052 1596 5060 1604
rect 5036 1536 5044 1544
rect 5020 1516 5028 1524
rect 5020 1496 5028 1504
rect 5180 1656 5188 1664
rect 5116 1536 5124 1544
rect 5084 1516 5092 1524
rect 5068 1496 5076 1504
rect 5004 1476 5012 1484
rect 5020 1456 5028 1464
rect 5084 1436 5092 1444
rect 5020 1376 5028 1384
rect 5052 1376 5060 1384
rect 4876 1296 4884 1304
rect 4892 1296 4900 1304
rect 4924 1216 4932 1224
rect 4908 1116 4916 1124
rect 4812 996 4820 1004
rect 4748 896 4756 904
rect 4764 896 4772 904
rect 4716 876 4724 884
rect 4716 736 4724 744
rect 4812 736 4820 744
rect 4700 696 4708 704
rect 4796 696 4804 704
rect 4700 656 4708 664
rect 4716 536 4724 544
rect 4700 516 4708 524
rect 4700 416 4708 424
rect 4700 396 4708 404
rect 4844 976 4852 984
rect 4892 916 4900 924
rect 4908 896 4916 904
rect 4860 856 4868 864
rect 4956 1336 4964 1344
rect 4988 1336 4996 1344
rect 5036 1336 5044 1344
rect 5084 1336 5092 1344
rect 4956 1316 4964 1324
rect 4972 1316 4980 1324
rect 4988 1296 4996 1304
rect 5004 1296 5012 1304
rect 4940 1136 4948 1144
rect 4972 1076 4980 1084
rect 4956 1056 4964 1064
rect 4940 956 4948 964
rect 4972 996 4980 1004
rect 4956 916 4964 924
rect 4940 896 4948 904
rect 4924 816 4932 824
rect 4892 796 4900 804
rect 4844 716 4852 724
rect 4876 716 4884 724
rect 4844 696 4852 704
rect 4924 736 4932 744
rect 4956 696 4964 704
rect 5260 1716 5268 1724
rect 5292 1676 5300 1684
rect 5628 2256 5636 2264
rect 5692 2336 5700 2344
rect 5724 2296 5732 2304
rect 6012 2996 6020 3004
rect 5996 2916 6004 2924
rect 5996 2896 6004 2904
rect 5980 2856 5988 2864
rect 6060 3076 6068 3084
rect 6060 3036 6068 3044
rect 6028 2916 6036 2924
rect 6012 2816 6020 2824
rect 6060 2796 6068 2804
rect 6012 2656 6020 2664
rect 5900 2636 5908 2644
rect 5923 2606 5931 2614
rect 5933 2606 5941 2614
rect 5943 2606 5951 2614
rect 5953 2606 5961 2614
rect 5963 2606 5971 2614
rect 5973 2606 5981 2614
rect 5932 2536 5940 2544
rect 5996 2516 6004 2524
rect 5884 2496 5892 2504
rect 5996 2496 6004 2504
rect 5884 2456 5892 2464
rect 5836 2436 5844 2444
rect 5756 2416 5764 2424
rect 5836 2356 5844 2364
rect 5788 2336 5796 2344
rect 5804 2336 5812 2344
rect 5708 2276 5716 2284
rect 5756 2276 5764 2284
rect 5692 2256 5700 2264
rect 5596 2196 5604 2204
rect 5660 2196 5668 2204
rect 5580 2136 5588 2144
rect 5468 2096 5476 2104
rect 5868 2316 5876 2324
rect 5820 2256 5828 2264
rect 5676 2176 5684 2184
rect 5788 2176 5796 2184
rect 5788 2156 5796 2164
rect 5532 2116 5540 2124
rect 5644 2096 5652 2104
rect 5516 2056 5524 2064
rect 5564 2056 5572 2064
rect 5532 1996 5540 2004
rect 5468 1936 5476 1944
rect 5356 1916 5364 1924
rect 5452 1916 5460 1924
rect 5404 1896 5412 1904
rect 5340 1756 5348 1764
rect 5532 1916 5540 1924
rect 5516 1876 5524 1884
rect 5532 1876 5540 1884
rect 5468 1856 5476 1864
rect 5516 1856 5524 1864
rect 5388 1776 5396 1784
rect 5436 1776 5444 1784
rect 5340 1736 5348 1744
rect 5356 1736 5364 1744
rect 5404 1756 5412 1764
rect 5372 1696 5380 1704
rect 5388 1696 5396 1704
rect 5356 1676 5364 1684
rect 5324 1656 5332 1664
rect 5212 1596 5220 1604
rect 5276 1576 5284 1584
rect 5292 1556 5300 1564
rect 5324 1536 5332 1544
rect 5420 1736 5428 1744
rect 5484 1736 5492 1744
rect 5452 1716 5460 1724
rect 5404 1596 5412 1604
rect 5404 1556 5412 1564
rect 5132 1496 5140 1504
rect 5308 1496 5316 1504
rect 5116 1256 5124 1264
rect 5180 1476 5188 1484
rect 5228 1476 5236 1484
rect 5212 1456 5220 1464
rect 5292 1476 5300 1484
rect 5324 1476 5332 1484
rect 5372 1476 5380 1484
rect 5180 1416 5188 1424
rect 5196 1416 5204 1424
rect 5308 1416 5316 1424
rect 5244 1356 5252 1364
rect 5260 1356 5268 1364
rect 5212 1336 5220 1344
rect 5196 1316 5204 1324
rect 5244 1316 5252 1324
rect 5180 1296 5188 1304
rect 5228 1296 5236 1304
rect 5148 1256 5156 1264
rect 5132 1236 5140 1244
rect 5196 1236 5204 1244
rect 5052 1196 5060 1204
rect 5084 1176 5092 1184
rect 5004 1156 5012 1164
rect 5100 1096 5108 1104
rect 5052 1076 5060 1084
rect 5132 1096 5140 1104
rect 5148 1076 5156 1084
rect 5116 1056 5124 1064
rect 5004 1016 5012 1024
rect 5068 976 5076 984
rect 5036 956 5044 964
rect 5196 1076 5204 1084
rect 5164 1056 5172 1064
rect 5100 956 5108 964
rect 5212 1056 5220 1064
rect 5068 916 5076 924
rect 5084 916 5092 924
rect 5148 916 5156 924
rect 5020 896 5028 904
rect 4988 856 4996 864
rect 4988 716 4996 724
rect 5036 716 5044 724
rect 5132 896 5140 904
rect 5164 836 5172 844
rect 5100 816 5108 824
rect 5276 1296 5284 1304
rect 5260 1216 5268 1224
rect 5308 1236 5316 1244
rect 5308 1216 5316 1224
rect 5292 1096 5300 1104
rect 5276 1076 5284 1084
rect 5260 1016 5268 1024
rect 5260 956 5268 964
rect 5420 1536 5428 1544
rect 5452 1656 5460 1664
rect 5452 1596 5460 1604
rect 5436 1496 5444 1504
rect 5420 1436 5428 1444
rect 5356 1376 5364 1384
rect 5340 1336 5348 1344
rect 5388 1336 5396 1344
rect 5340 1236 5348 1244
rect 5372 1196 5380 1204
rect 5372 1156 5380 1164
rect 5356 1096 5364 1104
rect 5356 1076 5364 1084
rect 5372 1016 5380 1024
rect 5372 976 5380 984
rect 5324 936 5332 944
rect 5356 936 5364 944
rect 5340 916 5348 924
rect 5212 796 5220 804
rect 5260 896 5268 904
rect 5308 896 5316 904
rect 5324 876 5332 884
rect 5324 796 5332 804
rect 5308 776 5316 784
rect 5276 736 5284 744
rect 5228 716 5236 724
rect 5100 702 5108 704
rect 5100 696 5108 702
rect 5276 696 5284 704
rect 5068 676 5076 684
rect 5260 676 5268 684
rect 5292 676 5300 684
rect 4796 596 4804 604
rect 4828 596 4836 604
rect 4748 516 4756 524
rect 4764 516 4772 524
rect 4748 496 4756 504
rect 4732 396 4740 404
rect 4716 276 4724 284
rect 4972 656 4980 664
rect 4876 576 4884 584
rect 4812 556 4820 564
rect 4844 556 4852 564
rect 4812 496 4820 504
rect 4748 376 4756 384
rect 4796 376 4804 384
rect 4764 356 4772 364
rect 4764 276 4772 284
rect 4796 276 4804 284
rect 4764 256 4772 264
rect 4748 156 4756 164
rect 4796 136 4804 144
rect 4828 316 4836 324
rect 4908 616 4916 624
rect 4892 516 4900 524
rect 4876 496 4884 504
rect 4860 376 4868 384
rect 5068 596 5076 604
rect 5004 576 5012 584
rect 4940 556 4948 564
rect 5228 556 5236 564
rect 5100 536 5108 544
rect 5196 536 5204 544
rect 5228 536 5236 544
rect 5020 516 5028 524
rect 5020 376 5028 384
rect 5100 376 5108 384
rect 4972 356 4980 364
rect 5116 336 5124 344
rect 5164 416 5172 424
rect 5324 736 5332 744
rect 5308 636 5316 644
rect 5276 576 5284 584
rect 5308 540 5316 544
rect 5308 536 5316 540
rect 5292 516 5300 524
rect 5292 456 5300 464
rect 5260 396 5268 404
rect 5244 336 5252 344
rect 5196 296 5204 304
rect 4988 276 4996 284
rect 4844 256 4852 264
rect 4828 216 4836 224
rect 4716 76 4724 84
rect 4748 16 4756 24
rect 4876 136 4884 144
rect 4924 176 4932 184
rect 4940 136 4948 144
rect 5276 276 5284 284
rect 5036 236 5044 244
rect 5004 136 5012 144
rect 4972 116 4980 124
rect 5004 116 5012 124
rect 5308 436 5316 444
rect 5372 816 5380 824
rect 5548 1836 5556 1844
rect 5516 1696 5524 1704
rect 5532 1696 5540 1704
rect 5548 1656 5556 1664
rect 5596 2016 5604 2024
rect 5612 1936 5620 1944
rect 5596 1896 5604 1904
rect 5660 1902 5668 1904
rect 5660 1896 5668 1902
rect 5852 2196 5860 2204
rect 5884 2196 5892 2204
rect 5868 2176 5876 2184
rect 5804 2096 5812 2104
rect 5932 2236 5940 2244
rect 5923 2206 5931 2214
rect 5933 2206 5941 2214
rect 5943 2206 5951 2214
rect 5953 2206 5961 2214
rect 5963 2206 5971 2214
rect 5973 2206 5981 2214
rect 5916 2156 5924 2164
rect 5932 2156 5940 2164
rect 5948 2136 5956 2144
rect 5948 2096 5956 2104
rect 5900 2056 5908 2064
rect 5916 2016 5924 2024
rect 6012 2436 6020 2444
rect 6028 2396 6036 2404
rect 6108 3156 6116 3164
rect 6092 2996 6100 3004
rect 6092 2976 6100 2984
rect 6108 2916 6116 2924
rect 6108 2876 6116 2884
rect 6124 2856 6132 2864
rect 6236 3296 6244 3304
rect 6316 3296 6324 3304
rect 6284 3256 6292 3264
rect 6172 3216 6180 3224
rect 6156 3196 6164 3204
rect 6188 3196 6196 3204
rect 6156 3076 6164 3084
rect 6156 2976 6164 2984
rect 6284 3096 6292 3104
rect 6348 3176 6356 3184
rect 6396 3176 6404 3184
rect 6332 3136 6340 3144
rect 6252 3056 6260 3064
rect 6300 3056 6308 3064
rect 6220 3036 6228 3044
rect 6332 3036 6340 3044
rect 6316 3016 6324 3024
rect 6268 2996 6276 3004
rect 6092 2656 6100 2664
rect 6108 2556 6116 2564
rect 6140 2516 6148 2524
rect 6140 2496 6148 2504
rect 6124 2436 6132 2444
rect 6108 2376 6116 2384
rect 6124 2376 6132 2384
rect 6092 2356 6100 2364
rect 6028 2176 6036 2184
rect 6060 2236 6068 2244
rect 6060 2216 6068 2224
rect 6076 2156 6084 2164
rect 6060 2136 6068 2144
rect 6124 2096 6132 2104
rect 6028 2056 6036 2064
rect 6012 2016 6020 2024
rect 6028 1956 6036 1964
rect 5788 1936 5796 1944
rect 5932 1936 5940 1944
rect 5996 1936 6004 1944
rect 5804 1896 5812 1904
rect 5900 1896 5908 1904
rect 5660 1816 5668 1824
rect 5708 1796 5716 1804
rect 5836 1876 5844 1884
rect 5916 1876 5924 1884
rect 5932 1876 5940 1884
rect 5740 1776 5748 1784
rect 5756 1776 5764 1784
rect 5708 1756 5716 1764
rect 5580 1696 5588 1704
rect 5644 1696 5652 1704
rect 5692 1696 5700 1704
rect 5596 1676 5604 1684
rect 5580 1656 5588 1664
rect 5532 1576 5540 1584
rect 5484 1396 5492 1404
rect 5484 1376 5492 1384
rect 5516 1376 5524 1384
rect 5468 1356 5476 1364
rect 5500 1356 5508 1364
rect 5436 1336 5444 1344
rect 5484 1336 5492 1344
rect 5420 1256 5428 1264
rect 5436 1096 5444 1104
rect 5420 1076 5428 1084
rect 5468 1316 5476 1324
rect 5564 1456 5572 1464
rect 5628 1656 5636 1664
rect 5612 1636 5620 1644
rect 5596 1516 5604 1524
rect 5596 1336 5604 1344
rect 5532 1316 5540 1324
rect 5580 1316 5588 1324
rect 5532 1276 5540 1284
rect 5596 1176 5604 1184
rect 5628 1596 5636 1604
rect 5740 1736 5748 1744
rect 5708 1616 5716 1624
rect 5692 1596 5700 1604
rect 5724 1556 5732 1564
rect 5740 1516 5748 1524
rect 5660 1496 5668 1504
rect 5724 1456 5732 1464
rect 5660 1376 5668 1384
rect 5708 1376 5716 1384
rect 5628 1336 5636 1344
rect 5692 1318 5700 1324
rect 5692 1316 5700 1318
rect 5708 1236 5716 1244
rect 5644 1176 5652 1184
rect 5692 1176 5700 1184
rect 5468 1116 5476 1124
rect 5484 1116 5492 1124
rect 5612 1116 5620 1124
rect 5532 1096 5540 1104
rect 5516 1076 5524 1084
rect 5564 1076 5572 1084
rect 5468 1056 5476 1064
rect 5532 1016 5540 1024
rect 5452 996 5460 1004
rect 5468 976 5476 984
rect 5484 976 5492 984
rect 5436 936 5444 944
rect 5500 936 5508 944
rect 5452 916 5460 924
rect 5468 916 5476 924
rect 5404 896 5412 904
rect 5548 956 5556 964
rect 5564 956 5572 964
rect 5580 936 5588 944
rect 5564 916 5572 924
rect 5468 816 5476 824
rect 5388 796 5396 804
rect 5420 796 5428 804
rect 5356 776 5364 784
rect 5340 716 5348 724
rect 5404 696 5412 704
rect 5452 756 5460 764
rect 5436 696 5444 704
rect 5404 656 5412 664
rect 5420 636 5428 644
rect 5404 556 5412 564
rect 5484 716 5492 724
rect 5628 1016 5636 1024
rect 5676 1076 5684 1084
rect 5644 976 5652 984
rect 5724 1136 5732 1144
rect 5772 1756 5780 1764
rect 5788 1716 5796 1724
rect 5900 1816 5908 1824
rect 5923 1806 5931 1814
rect 5933 1806 5941 1814
rect 5943 1806 5951 1814
rect 5953 1806 5961 1814
rect 5963 1806 5971 1814
rect 5973 1806 5981 1814
rect 6012 1916 6020 1924
rect 6076 1996 6084 2004
rect 6140 1976 6148 1984
rect 6060 1956 6068 1964
rect 6076 1956 6084 1964
rect 6076 1936 6084 1944
rect 6140 1936 6148 1944
rect 6092 1916 6100 1924
rect 6348 2976 6356 2984
rect 6380 2976 6388 2984
rect 6316 2956 6324 2964
rect 6444 3096 6452 3104
rect 6524 4516 6532 4524
rect 6524 4256 6532 4264
rect 6524 3896 6532 3904
rect 6508 3836 6516 3844
rect 6572 4716 6580 4724
rect 6572 4676 6580 4684
rect 6636 4896 6644 4904
rect 6604 4876 6612 4884
rect 6652 4836 6660 4844
rect 6668 4836 6676 4844
rect 6604 4756 6612 4764
rect 6652 4736 6660 4744
rect 6652 4716 6660 4724
rect 6668 4696 6676 4704
rect 6716 5056 6724 5064
rect 6748 4996 6756 5004
rect 6716 4956 6724 4964
rect 6764 4936 6772 4944
rect 6732 4916 6740 4924
rect 6700 4856 6708 4864
rect 6684 4676 6692 4684
rect 6684 4656 6692 4664
rect 6684 4616 6692 4624
rect 6620 4536 6628 4544
rect 6588 4476 6596 4484
rect 6572 4336 6580 4344
rect 6556 4316 6564 4324
rect 6604 4376 6612 4384
rect 6604 4316 6612 4324
rect 6972 5318 6980 5324
rect 6972 5316 6980 5318
rect 7004 5316 7012 5324
rect 7164 5318 7172 5324
rect 7164 5316 7172 5318
rect 7244 5316 7252 5324
rect 6908 5196 6916 5204
rect 6924 5176 6932 5184
rect 6844 5156 6852 5164
rect 6892 5096 6900 5104
rect 6844 4996 6852 5004
rect 6812 4916 6820 4924
rect 6828 4856 6836 4864
rect 6892 5056 6900 5064
rect 6828 4836 6836 4844
rect 6860 4836 6868 4844
rect 6796 4736 6804 4744
rect 6780 4696 6788 4704
rect 6748 4676 6756 4684
rect 6780 4656 6788 4664
rect 6748 4596 6756 4604
rect 6732 4576 6740 4584
rect 6716 4536 6724 4544
rect 6636 4516 6644 4524
rect 6700 4516 6708 4524
rect 6652 4496 6660 4504
rect 6652 4476 6660 4484
rect 6684 4376 6692 4384
rect 6636 4316 6644 4324
rect 6652 4316 6660 4324
rect 6716 4476 6724 4484
rect 6748 4476 6756 4484
rect 6716 4436 6724 4444
rect 6684 4296 6692 4304
rect 6588 4196 6596 4204
rect 6620 4276 6628 4284
rect 6636 4156 6644 4164
rect 6732 4356 6740 4364
rect 6748 4356 6756 4364
rect 6764 4356 6772 4364
rect 6860 4576 6868 4584
rect 6828 4556 6836 4564
rect 6812 4536 6820 4544
rect 6796 4396 6804 4404
rect 6684 4196 6692 4204
rect 6716 4196 6724 4204
rect 6748 4196 6756 4204
rect 6732 4176 6740 4184
rect 6668 4116 6676 4124
rect 6700 4116 6708 4124
rect 6668 4076 6676 4084
rect 6604 3896 6612 3904
rect 6588 3796 6596 3804
rect 6540 3776 6548 3784
rect 6524 3756 6532 3764
rect 6572 3756 6580 3764
rect 6540 3716 6548 3724
rect 6508 3696 6516 3704
rect 6492 3656 6500 3664
rect 6476 3496 6484 3504
rect 6492 3336 6500 3344
rect 6476 3256 6484 3264
rect 6556 3616 6564 3624
rect 6524 3516 6532 3524
rect 6540 3516 6548 3524
rect 6636 3916 6644 3924
rect 6716 3956 6724 3964
rect 6732 3896 6740 3904
rect 6652 3836 6660 3844
rect 6652 3816 6660 3824
rect 6620 3676 6628 3684
rect 6700 3816 6708 3824
rect 6716 3776 6724 3784
rect 6684 3656 6692 3664
rect 6572 3536 6580 3544
rect 6604 3536 6612 3544
rect 6652 3516 6660 3524
rect 6668 3516 6676 3524
rect 6604 3496 6612 3504
rect 6588 3476 6596 3484
rect 6540 3456 6548 3464
rect 6556 3456 6564 3464
rect 6588 3456 6596 3464
rect 6556 3336 6564 3344
rect 6620 3436 6628 3444
rect 6684 3476 6692 3484
rect 6796 4316 6804 4324
rect 6780 4236 6788 4244
rect 6796 4116 6804 4124
rect 6908 4976 6916 4984
rect 6892 4916 6900 4924
rect 6972 5056 6980 5064
rect 6940 5036 6948 5044
rect 6956 4916 6964 4924
rect 6908 4896 6916 4904
rect 6908 4756 6916 4764
rect 6988 4636 6996 4644
rect 6908 4616 6916 4624
rect 6988 4616 6996 4624
rect 6924 4576 6932 4584
rect 6956 4576 6964 4584
rect 6940 4516 6948 4524
rect 6908 4476 6916 4484
rect 6876 4416 6884 4424
rect 6844 4376 6852 4384
rect 6844 4316 6852 4324
rect 6844 4296 6852 4304
rect 6876 4256 6884 4264
rect 6828 4156 6836 4164
rect 6796 3956 6804 3964
rect 6812 3956 6820 3964
rect 6780 3896 6788 3904
rect 6860 4118 6868 4124
rect 6860 4116 6868 4118
rect 6876 3936 6884 3944
rect 6764 3856 6772 3864
rect 6780 3836 6788 3844
rect 6860 3896 6868 3904
rect 6812 3736 6820 3744
rect 6860 3856 6868 3864
rect 6844 3716 6852 3724
rect 6780 3656 6788 3664
rect 6748 3616 6756 3624
rect 6732 3596 6740 3604
rect 6732 3556 6740 3564
rect 6716 3456 6724 3464
rect 6716 3376 6724 3384
rect 6700 3296 6708 3304
rect 6508 3236 6516 3244
rect 6620 3216 6628 3224
rect 6668 3176 6676 3184
rect 6668 3156 6676 3164
rect 6604 3136 6612 3144
rect 6572 3116 6580 3124
rect 6524 3096 6532 3104
rect 6620 3116 6628 3124
rect 6636 3096 6644 3104
rect 6652 3096 6660 3104
rect 6268 2896 6276 2904
rect 6284 2896 6292 2904
rect 6236 2816 6244 2824
rect 6300 2816 6308 2824
rect 6220 2676 6228 2684
rect 6204 2616 6212 2624
rect 6204 2556 6212 2564
rect 6268 2676 6276 2684
rect 6252 2636 6260 2644
rect 6268 2636 6276 2644
rect 6236 2536 6244 2544
rect 6220 2516 6228 2524
rect 6188 2496 6196 2504
rect 6204 2476 6212 2484
rect 6332 2716 6340 2724
rect 6332 2676 6340 2684
rect 6316 2656 6324 2664
rect 6348 2636 6356 2644
rect 6284 2556 6292 2564
rect 6284 2536 6292 2544
rect 6412 2896 6420 2904
rect 6428 2896 6436 2904
rect 6588 3076 6596 3084
rect 6556 3056 6564 3064
rect 6492 2996 6500 3004
rect 6508 2976 6516 2984
rect 6460 2956 6468 2964
rect 6492 2956 6500 2964
rect 6572 3016 6580 3024
rect 6492 2916 6500 2924
rect 6556 2916 6564 2924
rect 6476 2896 6484 2904
rect 6556 2896 6564 2904
rect 6476 2876 6484 2884
rect 6460 2776 6468 2784
rect 6460 2716 6468 2724
rect 6444 2636 6452 2644
rect 6412 2536 6420 2544
rect 6444 2516 6452 2524
rect 6268 2456 6276 2464
rect 6284 2436 6292 2444
rect 6508 2776 6516 2784
rect 6588 2976 6596 2984
rect 6668 2976 6676 2984
rect 6620 2936 6628 2944
rect 6604 2716 6612 2724
rect 6556 2676 6564 2684
rect 6588 2676 6596 2684
rect 6636 2916 6644 2924
rect 6636 2896 6644 2904
rect 6636 2796 6644 2804
rect 6540 2656 6548 2664
rect 6508 2596 6516 2604
rect 6524 2536 6532 2544
rect 6380 2496 6388 2504
rect 6460 2496 6468 2504
rect 6396 2396 6404 2404
rect 6332 2336 6340 2344
rect 6220 2296 6228 2304
rect 6252 2296 6260 2304
rect 6220 2276 6228 2284
rect 6252 2256 6260 2264
rect 6332 2256 6340 2264
rect 6348 2256 6356 2264
rect 6252 2136 6260 2144
rect 6316 2236 6324 2244
rect 6300 2176 6308 2184
rect 6316 2176 6324 2184
rect 6284 2096 6292 2104
rect 6332 2136 6340 2144
rect 6380 2136 6388 2144
rect 6428 2336 6436 2344
rect 6444 2336 6452 2344
rect 6364 2116 6372 2124
rect 6476 2456 6484 2464
rect 6476 2416 6484 2424
rect 6492 2396 6500 2404
rect 6524 2376 6532 2384
rect 6508 2316 6516 2324
rect 6508 2276 6516 2284
rect 6444 2256 6452 2264
rect 6460 2256 6468 2264
rect 6492 2256 6500 2264
rect 6460 2196 6468 2204
rect 6492 2156 6500 2164
rect 6364 2056 6372 2064
rect 6444 2056 6452 2064
rect 6204 1996 6212 2004
rect 6172 1976 6180 1984
rect 6300 1936 6308 1944
rect 6412 2036 6420 2044
rect 6476 2136 6484 2144
rect 6460 1976 6468 1984
rect 6396 1936 6404 1944
rect 6508 2136 6516 2144
rect 6508 2116 6516 2124
rect 6588 2656 6596 2664
rect 6556 2596 6564 2604
rect 6588 2576 6596 2584
rect 6556 2416 6564 2424
rect 6572 2356 6580 2364
rect 6572 2336 6580 2344
rect 6620 2616 6628 2624
rect 6604 2536 6612 2544
rect 6700 3236 6708 3244
rect 6748 3536 6756 3544
rect 6748 3456 6756 3464
rect 6876 3776 6884 3784
rect 6876 3756 6884 3764
rect 6876 3736 6884 3744
rect 6860 3596 6868 3604
rect 6796 3416 6804 3424
rect 6796 3376 6804 3384
rect 6796 3356 6804 3364
rect 6780 3316 6788 3324
rect 6764 3296 6772 3304
rect 6748 3236 6756 3244
rect 6972 4456 6980 4464
rect 6972 4296 6980 4304
rect 6924 4176 6932 4184
rect 6956 4136 6964 4144
rect 6972 4116 6980 4124
rect 6924 3936 6932 3944
rect 6924 3916 6932 3924
rect 6956 3916 6964 3924
rect 6908 3816 6916 3824
rect 6972 3796 6980 3804
rect 6956 3776 6964 3784
rect 6924 3716 6932 3724
rect 6940 3696 6948 3704
rect 6924 3536 6932 3544
rect 6892 3476 6900 3484
rect 7036 5196 7044 5204
rect 7100 5096 7108 5104
rect 7228 5096 7236 5104
rect 7052 5036 7060 5044
rect 7036 4956 7044 4964
rect 7068 4876 7076 4884
rect 7020 4636 7028 4644
rect 7004 4536 7012 4544
rect 7004 4516 7012 4524
rect 7004 4476 7012 4484
rect 7148 4876 7156 4884
rect 7132 4696 7140 4704
rect 7084 4676 7092 4684
rect 7356 5216 7364 5224
rect 7388 5216 7396 5224
rect 7356 5196 7364 5204
rect 7324 5156 7332 5164
rect 7212 4976 7220 4984
rect 7196 4876 7204 4884
rect 7180 4856 7188 4864
rect 7212 4856 7220 4864
rect 7180 4756 7188 4764
rect 7164 4736 7172 4744
rect 7180 4736 7188 4744
rect 7164 4716 7172 4724
rect 7164 4696 7172 4704
rect 7100 4576 7108 4584
rect 7052 4556 7060 4564
rect 7132 4556 7140 4564
rect 7036 4496 7044 4504
rect 7116 4496 7124 4504
rect 7100 4396 7108 4404
rect 7084 4356 7092 4364
rect 7004 4256 7012 4264
rect 7020 4236 7028 4244
rect 7052 4236 7060 4244
rect 7004 4136 7012 4144
rect 7132 4376 7140 4384
rect 7116 4336 7124 4344
rect 7116 4296 7124 4304
rect 7084 4156 7092 4164
rect 7084 4116 7092 4124
rect 7100 4056 7108 4064
rect 7052 4036 7060 4044
rect 7052 3956 7060 3964
rect 7004 3896 7012 3904
rect 7020 3776 7028 3784
rect 7004 3636 7012 3644
rect 6988 3556 6996 3564
rect 7004 3476 7012 3484
rect 6972 3416 6980 3424
rect 7004 3416 7012 3424
rect 6988 3396 6996 3404
rect 6876 3336 6884 3344
rect 6876 3316 6884 3324
rect 6908 3296 6916 3304
rect 6748 3136 6756 3144
rect 6908 3136 6916 3144
rect 6844 3116 6852 3124
rect 6972 3116 6980 3124
rect 6812 3096 6820 3104
rect 6764 3056 6772 3064
rect 6828 3056 6836 3064
rect 6684 2916 6692 2924
rect 6652 2756 6660 2764
rect 6684 2756 6692 2764
rect 6716 3016 6724 3024
rect 6892 3056 6900 3064
rect 6844 3036 6852 3044
rect 6876 3036 6884 3044
rect 6892 3036 6900 3044
rect 6860 2956 6868 2964
rect 6956 3036 6964 3044
rect 6908 2996 6916 3004
rect 6940 2996 6948 3004
rect 6956 2976 6964 2984
rect 6988 3056 6996 3064
rect 6988 3016 6996 3024
rect 6780 2916 6788 2924
rect 6748 2896 6756 2904
rect 6764 2896 6772 2904
rect 6764 2856 6772 2864
rect 6700 2696 6708 2704
rect 6668 2676 6676 2684
rect 6668 2656 6676 2664
rect 6652 2636 6660 2644
rect 6716 2656 6724 2664
rect 6716 2636 6724 2644
rect 6684 2556 6692 2564
rect 6700 2556 6708 2564
rect 6668 2516 6676 2524
rect 6604 2496 6612 2504
rect 6636 2496 6644 2504
rect 6748 2596 6756 2604
rect 6620 2476 6628 2484
rect 6604 2316 6612 2324
rect 6652 2316 6660 2324
rect 6684 2336 6692 2344
rect 6636 2256 6644 2264
rect 6556 2236 6564 2244
rect 6572 2156 6580 2164
rect 6556 2116 6564 2124
rect 6636 2116 6644 2124
rect 6652 2116 6660 2124
rect 6620 2096 6628 2104
rect 6540 2076 6548 2084
rect 6476 1916 6484 1924
rect 6540 1916 6548 1924
rect 6620 1916 6628 1924
rect 6668 1916 6676 1924
rect 6076 1876 6084 1884
rect 6076 1816 6084 1824
rect 6012 1796 6020 1804
rect 6044 1796 6052 1804
rect 5900 1736 5908 1744
rect 5852 1716 5860 1724
rect 5820 1676 5828 1684
rect 5852 1676 5860 1684
rect 6044 1776 6052 1784
rect 5996 1736 6004 1744
rect 5980 1656 5988 1664
rect 5884 1636 5892 1644
rect 5804 1536 5812 1544
rect 5900 1516 5908 1524
rect 6076 1676 6084 1684
rect 6044 1536 6052 1544
rect 5996 1516 6004 1524
rect 5788 1496 5796 1504
rect 5900 1496 5908 1504
rect 5852 1476 5860 1484
rect 5772 1456 5780 1464
rect 5820 1456 5828 1464
rect 5868 1456 5876 1464
rect 5820 1376 5828 1384
rect 5916 1476 5924 1484
rect 6060 1456 6068 1464
rect 5923 1406 5931 1414
rect 5933 1406 5941 1414
rect 5943 1406 5951 1414
rect 5953 1406 5961 1414
rect 5963 1406 5971 1414
rect 5973 1406 5981 1414
rect 6076 1436 6084 1444
rect 6060 1416 6068 1424
rect 5932 1376 5940 1384
rect 6012 1376 6020 1384
rect 5868 1336 5876 1344
rect 5916 1296 5924 1304
rect 5852 1276 5860 1284
rect 6028 1236 6036 1244
rect 6076 1236 6084 1244
rect 5836 1176 5844 1184
rect 5772 1116 5780 1124
rect 5868 1116 5876 1124
rect 5756 1096 5764 1104
rect 5852 1096 5860 1104
rect 5820 1076 5828 1084
rect 5900 1076 5908 1084
rect 5740 1056 5748 1064
rect 5756 1056 5764 1064
rect 5692 936 5700 944
rect 5532 796 5540 804
rect 5516 696 5524 704
rect 5500 656 5508 664
rect 5468 596 5476 604
rect 5500 596 5508 604
rect 5580 756 5588 764
rect 5660 916 5668 924
rect 5564 736 5572 744
rect 5644 736 5652 744
rect 5548 716 5556 724
rect 5644 716 5652 724
rect 5724 916 5732 924
rect 5756 996 5764 1004
rect 5772 976 5780 984
rect 5772 936 5780 944
rect 5772 916 5780 924
rect 5756 896 5764 904
rect 5740 876 5748 884
rect 5804 976 5812 984
rect 5820 936 5828 944
rect 5884 996 5892 1004
rect 5923 1006 5931 1014
rect 5933 1006 5941 1014
rect 5943 1006 5951 1014
rect 5953 1006 5961 1014
rect 5963 1006 5971 1014
rect 5973 1006 5981 1014
rect 5900 976 5908 984
rect 5916 976 5924 984
rect 5932 956 5940 964
rect 5820 916 5828 924
rect 5788 856 5796 864
rect 5708 756 5716 764
rect 5884 936 5892 944
rect 5916 936 5924 944
rect 5868 916 5876 924
rect 5900 916 5908 924
rect 5820 856 5828 864
rect 5852 856 5860 864
rect 5836 836 5844 844
rect 5756 716 5764 724
rect 5772 716 5780 724
rect 5564 696 5572 704
rect 5612 696 5620 704
rect 5692 696 5700 704
rect 5804 696 5812 704
rect 5548 656 5556 664
rect 5532 576 5540 584
rect 5372 516 5380 524
rect 5356 396 5364 404
rect 5388 336 5396 344
rect 5340 276 5348 284
rect 5260 256 5268 264
rect 5196 196 5204 204
rect 5164 136 5172 144
rect 5276 136 5284 144
rect 5388 276 5396 284
rect 5596 676 5604 684
rect 5660 676 5668 684
rect 5724 676 5732 684
rect 5852 756 5860 764
rect 5884 696 5892 704
rect 5612 616 5620 624
rect 5452 536 5460 544
rect 5596 536 5604 544
rect 5500 516 5508 524
rect 5532 516 5540 524
rect 5468 496 5476 504
rect 5500 496 5508 504
rect 5580 496 5588 504
rect 5692 596 5700 604
rect 5644 576 5652 584
rect 5660 556 5668 564
rect 5676 516 5684 524
rect 5628 456 5636 464
rect 5644 456 5652 464
rect 5596 436 5604 444
rect 5484 356 5492 364
rect 5468 336 5476 344
rect 5548 336 5556 344
rect 5532 316 5540 324
rect 5580 296 5588 304
rect 5468 256 5476 264
rect 5404 196 5412 204
rect 5356 156 5364 164
rect 5404 156 5412 164
rect 5372 116 5380 124
rect 5420 116 5428 124
rect 4812 96 4820 104
rect 4956 96 4964 104
rect 5452 196 5460 204
rect 5500 156 5508 164
rect 5532 136 5540 144
rect 5644 396 5652 404
rect 5612 356 5620 364
rect 5660 356 5668 364
rect 5660 296 5668 304
rect 5788 616 5796 624
rect 5820 616 5828 624
rect 5836 616 5844 624
rect 5708 496 5716 504
rect 5708 416 5716 424
rect 5692 296 5700 304
rect 5772 556 5780 564
rect 5740 536 5748 544
rect 5772 536 5780 544
rect 5756 516 5764 524
rect 5772 496 5780 504
rect 5740 416 5748 424
rect 5740 336 5748 344
rect 5724 316 5732 324
rect 5772 316 5780 324
rect 5740 276 5748 284
rect 5756 256 5764 264
rect 5676 236 5684 244
rect 5692 236 5700 244
rect 5596 216 5604 224
rect 5660 216 5668 224
rect 5644 176 5652 184
rect 5676 176 5684 184
rect 5740 196 5748 204
rect 5772 196 5780 204
rect 5676 156 5684 164
rect 5596 136 5604 144
rect 5804 576 5812 584
rect 5820 576 5828 584
rect 5820 556 5828 564
rect 5804 496 5812 504
rect 5804 396 5812 404
rect 5820 376 5828 384
rect 5836 296 5844 304
rect 5868 676 5876 684
rect 5916 836 5924 844
rect 5932 816 5940 824
rect 5916 796 5924 804
rect 5932 796 5940 804
rect 6012 976 6020 984
rect 6108 1676 6116 1684
rect 6124 1576 6132 1584
rect 6172 1896 6180 1904
rect 6284 1896 6292 1904
rect 6188 1816 6196 1824
rect 6748 2496 6756 2504
rect 6748 2296 6756 2304
rect 6860 2896 6868 2904
rect 6940 2876 6948 2884
rect 6972 2796 6980 2804
rect 6828 2776 6836 2784
rect 6796 2716 6804 2724
rect 6780 2696 6788 2704
rect 6876 2696 6884 2704
rect 6796 2596 6804 2604
rect 6812 2596 6820 2604
rect 6812 2536 6820 2544
rect 6860 2536 6868 2544
rect 6796 2396 6804 2404
rect 6908 2656 6916 2664
rect 6956 2676 6964 2684
rect 6924 2616 6932 2624
rect 6988 2636 6996 2644
rect 7036 3756 7044 3764
rect 7116 3916 7124 3924
rect 7084 3876 7092 3884
rect 7068 3816 7076 3824
rect 7084 3736 7092 3744
rect 7068 3696 7076 3704
rect 7036 3676 7044 3684
rect 7052 3676 7060 3684
rect 7036 3496 7044 3504
rect 7052 3496 7060 3504
rect 7084 3656 7092 3664
rect 7180 4536 7188 4544
rect 7164 4336 7172 4344
rect 7276 4956 7284 4964
rect 7340 4956 7348 4964
rect 7276 4876 7284 4884
rect 7324 4876 7332 4884
rect 7260 4736 7268 4744
rect 7244 4676 7252 4684
rect 7212 4596 7220 4604
rect 7292 4696 7300 4704
rect 7276 4616 7284 4624
rect 7244 4576 7252 4584
rect 7276 4576 7284 4584
rect 7244 4556 7252 4564
rect 7196 4356 7204 4364
rect 7164 4316 7172 4324
rect 7164 4296 7172 4304
rect 7148 4276 7156 4284
rect 7148 4036 7156 4044
rect 7196 4176 7204 4184
rect 7180 4076 7188 4084
rect 7180 4016 7188 4024
rect 7132 3776 7140 3784
rect 7164 3836 7172 3844
rect 7212 4156 7220 4164
rect 7212 4116 7220 4124
rect 7212 4076 7220 4084
rect 7228 3876 7236 3884
rect 7244 3836 7252 3844
rect 7212 3756 7220 3764
rect 7164 3716 7172 3724
rect 7148 3696 7156 3704
rect 7132 3676 7140 3684
rect 7052 3316 7060 3324
rect 7116 3616 7124 3624
rect 7148 3656 7156 3664
rect 7100 3356 7108 3364
rect 7132 3396 7140 3404
rect 7068 3256 7076 3264
rect 7052 3196 7060 3204
rect 7068 3136 7076 3144
rect 7036 3096 7044 3104
rect 7116 3076 7124 3084
rect 7100 3056 7108 3064
rect 7052 3036 7060 3044
rect 7116 3036 7124 3044
rect 7132 3036 7140 3044
rect 7100 2996 7108 3004
rect 7052 2976 7060 2984
rect 7036 2936 7044 2944
rect 7292 4496 7300 4504
rect 7308 4376 7316 4384
rect 7308 4316 7316 4324
rect 7340 4216 7348 4224
rect 7308 4116 7316 4124
rect 7292 4096 7300 4104
rect 7292 4076 7300 4084
rect 7324 4076 7332 4084
rect 7276 3576 7284 3584
rect 7260 3496 7268 3504
rect 7244 3476 7252 3484
rect 7260 3456 7268 3464
rect 7212 3436 7220 3444
rect 7196 3396 7204 3404
rect 7180 3376 7188 3384
rect 7212 3376 7220 3384
rect 7244 3316 7252 3324
rect 7260 3296 7268 3304
rect 7196 3176 7204 3184
rect 7180 3136 7188 3144
rect 7164 3116 7172 3124
rect 7164 3056 7172 3064
rect 7164 3036 7172 3044
rect 7148 2976 7156 2984
rect 7244 3096 7252 3104
rect 7244 3016 7252 3024
rect 7212 2996 7220 3004
rect 7116 2956 7124 2964
rect 7148 2956 7156 2964
rect 7084 2936 7092 2944
rect 7116 2916 7124 2924
rect 7052 2856 7060 2864
rect 7020 2656 7028 2664
rect 7068 2636 7076 2644
rect 7020 2576 7028 2584
rect 6988 2536 6996 2544
rect 7004 2536 7012 2544
rect 6908 2476 6916 2484
rect 6844 2276 6852 2284
rect 6796 2256 6804 2264
rect 6844 2256 6852 2264
rect 6828 2216 6836 2224
rect 6764 2196 6772 2204
rect 6764 2176 6772 2184
rect 6876 2196 6884 2204
rect 6732 2136 6740 2144
rect 6844 2136 6852 2144
rect 6796 2116 6804 2124
rect 6700 2096 6708 2104
rect 6684 1896 6692 1904
rect 6572 1876 6580 1884
rect 6300 1856 6308 1864
rect 6348 1856 6356 1864
rect 6444 1856 6452 1864
rect 6588 1856 6596 1864
rect 6460 1836 6468 1844
rect 6492 1836 6500 1844
rect 6188 1736 6196 1744
rect 6252 1736 6260 1744
rect 6172 1656 6180 1664
rect 6172 1516 6180 1524
rect 6140 1496 6148 1504
rect 6140 1436 6148 1444
rect 6156 1416 6164 1424
rect 6156 1396 6164 1404
rect 6252 1696 6260 1704
rect 6204 1656 6212 1664
rect 6364 1776 6372 1784
rect 6316 1716 6324 1724
rect 6428 1718 6436 1724
rect 6428 1716 6436 1718
rect 6284 1656 6292 1664
rect 6220 1616 6228 1624
rect 6300 1616 6308 1624
rect 6204 1596 6212 1604
rect 6268 1556 6276 1564
rect 6252 1516 6260 1524
rect 6508 1796 6516 1804
rect 6492 1756 6500 1764
rect 6492 1716 6500 1724
rect 6620 1776 6628 1784
rect 6748 2096 6756 2104
rect 6764 2096 6772 2104
rect 6716 2056 6724 2064
rect 6764 2016 6772 2024
rect 6796 1936 6804 1944
rect 6716 1916 6724 1924
rect 6764 1916 6772 1924
rect 6764 1896 6772 1904
rect 7100 2736 7108 2744
rect 7116 2676 7124 2684
rect 7100 2616 7108 2624
rect 7084 2596 7092 2604
rect 7116 2576 7124 2584
rect 7036 2556 7044 2564
rect 7020 2496 7028 2504
rect 7084 2496 7092 2504
rect 7132 2476 7140 2484
rect 7164 2816 7172 2824
rect 7180 2576 7188 2584
rect 7180 2536 7188 2544
rect 7164 2516 7172 2524
rect 7180 2516 7188 2524
rect 7228 2916 7236 2924
rect 7212 2876 7220 2884
rect 7212 2796 7220 2804
rect 7228 2596 7236 2604
rect 7068 2336 7076 2344
rect 7148 2336 7156 2344
rect 6956 2276 6964 2284
rect 7132 2276 7140 2284
rect 7004 2236 7012 2244
rect 7164 2156 7172 2164
rect 6908 2136 6916 2144
rect 6924 2136 6932 2144
rect 7068 2136 7076 2144
rect 6956 2116 6964 2124
rect 6876 2096 6884 2104
rect 6924 2096 6932 2104
rect 7036 2076 7044 2084
rect 7004 1956 7012 1964
rect 7020 1916 7028 1924
rect 6908 1896 6916 1904
rect 6844 1876 6852 1884
rect 6972 1876 6980 1884
rect 7004 1876 7012 1884
rect 6796 1856 6804 1864
rect 6700 1796 6708 1804
rect 6780 1796 6788 1804
rect 6652 1756 6660 1764
rect 6908 1756 6916 1764
rect 6588 1736 6596 1744
rect 6540 1716 6548 1724
rect 6652 1718 6660 1724
rect 6652 1716 6660 1718
rect 6556 1676 6564 1684
rect 6524 1636 6532 1644
rect 6348 1556 6356 1564
rect 6460 1556 6468 1564
rect 6220 1476 6228 1484
rect 6220 1416 6228 1424
rect 6204 1396 6212 1404
rect 6108 1336 6116 1344
rect 6172 1336 6180 1344
rect 6204 1276 6212 1284
rect 6204 1256 6212 1264
rect 6156 1156 6164 1164
rect 6332 1456 6340 1464
rect 6364 1536 6372 1544
rect 6444 1516 6452 1524
rect 6524 1516 6532 1524
rect 6572 1516 6580 1524
rect 6572 1496 6580 1504
rect 6380 1456 6388 1464
rect 6540 1476 6548 1484
rect 6476 1456 6484 1464
rect 6396 1436 6404 1444
rect 6428 1436 6436 1444
rect 6252 1316 6260 1324
rect 6300 1316 6308 1324
rect 6444 1396 6452 1404
rect 6428 1336 6436 1344
rect 6476 1336 6484 1344
rect 6380 1316 6388 1324
rect 6412 1316 6420 1324
rect 6492 1316 6500 1324
rect 6428 1296 6436 1304
rect 6396 1276 6404 1284
rect 6396 1256 6404 1264
rect 6284 1236 6292 1244
rect 6252 1196 6260 1204
rect 6236 1116 6244 1124
rect 6268 1136 6276 1144
rect 6252 1096 6260 1104
rect 6092 1016 6100 1024
rect 6140 956 6148 964
rect 6076 936 6084 944
rect 6156 936 6164 944
rect 6012 916 6020 924
rect 6060 916 6068 924
rect 6092 916 6100 924
rect 6044 836 6052 844
rect 5996 776 6004 784
rect 6012 716 6020 724
rect 6300 1116 6308 1124
rect 6300 1096 6308 1104
rect 6204 1076 6212 1084
rect 6220 1076 6228 1084
rect 6236 1056 6244 1064
rect 6476 1216 6484 1224
rect 6444 1116 6452 1124
rect 6428 1076 6436 1084
rect 6236 1016 6244 1024
rect 6220 976 6228 984
rect 6204 936 6212 944
rect 6172 916 6180 924
rect 6204 916 6212 924
rect 6188 896 6196 904
rect 6156 876 6164 884
rect 6140 836 6148 844
rect 6076 776 6084 784
rect 6124 776 6132 784
rect 5932 656 5940 664
rect 5996 656 6004 664
rect 5900 616 5908 624
rect 5923 606 5931 614
rect 5933 606 5941 614
rect 5943 606 5951 614
rect 5953 606 5961 614
rect 5963 606 5971 614
rect 5973 606 5981 614
rect 5996 596 6004 604
rect 5868 556 5876 564
rect 5996 556 6004 564
rect 5948 536 5956 544
rect 6108 576 6116 584
rect 6076 556 6084 564
rect 5900 516 5908 524
rect 5868 496 5876 504
rect 6060 496 6068 504
rect 5980 376 5988 384
rect 6012 356 6020 364
rect 6060 456 6068 464
rect 6060 416 6068 424
rect 5996 316 6004 324
rect 6028 316 6036 324
rect 6044 316 6052 324
rect 5884 276 5892 284
rect 5804 256 5812 264
rect 5868 176 5876 184
rect 6044 296 6052 304
rect 5996 256 6004 264
rect 6028 256 6036 264
rect 6092 536 6100 544
rect 6172 816 6180 824
rect 6252 936 6260 944
rect 6524 1396 6532 1404
rect 7116 2016 7124 2024
rect 7084 1936 7092 1944
rect 7068 1916 7076 1924
rect 7068 1896 7076 1904
rect 7196 2496 7204 2504
rect 7244 2516 7252 2524
rect 7228 2496 7236 2504
rect 7404 4536 7412 4544
rect 7388 3736 7396 3744
rect 7308 3536 7316 3544
rect 7388 3516 7396 3524
rect 7308 3476 7316 3484
rect 7356 3476 7364 3484
rect 7292 3296 7300 3304
rect 7292 3116 7300 3124
rect 7276 3076 7284 3084
rect 7276 2956 7284 2964
rect 7276 2936 7284 2944
rect 7388 2956 7396 2964
rect 7308 2916 7316 2924
rect 7324 2796 7332 2804
rect 7292 2676 7300 2684
rect 7276 2576 7284 2584
rect 7212 2376 7220 2384
rect 7196 2216 7204 2224
rect 7196 2176 7204 2184
rect 7196 2016 7204 2024
rect 7180 1936 7188 1944
rect 7196 1936 7204 1944
rect 7148 1896 7156 1904
rect 7180 1896 7188 1904
rect 7180 1836 7188 1844
rect 7116 1816 7124 1824
rect 7180 1816 7188 1824
rect 7052 1736 7060 1744
rect 7036 1716 7044 1724
rect 7260 2416 7268 2424
rect 7324 2516 7332 2524
rect 7260 2336 7268 2344
rect 7292 2336 7300 2344
rect 7244 2236 7252 2244
rect 7260 2216 7268 2224
rect 7292 2316 7300 2324
rect 7324 2316 7332 2324
rect 7292 2216 7300 2224
rect 7292 2196 7300 2204
rect 7276 2176 7284 2184
rect 7276 2156 7284 2164
rect 7260 1876 7268 1884
rect 7260 1856 7268 1864
rect 7244 1776 7252 1784
rect 7180 1676 7188 1684
rect 7196 1676 7204 1684
rect 6988 1516 6996 1524
rect 7036 1516 7044 1524
rect 7004 1496 7012 1504
rect 7020 1496 7028 1504
rect 6860 1456 6868 1464
rect 6668 1396 6676 1404
rect 6540 1376 6548 1384
rect 6652 1376 6660 1384
rect 6588 1336 6596 1344
rect 6604 1316 6612 1324
rect 6540 1296 6548 1304
rect 6508 1276 6516 1284
rect 6588 1276 6596 1284
rect 6492 1076 6500 1084
rect 6476 1056 6484 1064
rect 6380 976 6388 984
rect 6348 936 6356 944
rect 6396 936 6404 944
rect 6460 1016 6468 1024
rect 6604 1256 6612 1264
rect 6716 1376 6724 1384
rect 6732 1336 6740 1344
rect 6684 1296 6692 1304
rect 6700 1296 6708 1304
rect 6668 1256 6676 1264
rect 6620 1196 6628 1204
rect 6556 1176 6564 1184
rect 6540 1156 6548 1164
rect 6604 1156 6612 1164
rect 6636 1136 6644 1144
rect 6620 1116 6628 1124
rect 6556 1076 6564 1084
rect 6588 1076 6596 1084
rect 6524 1056 6532 1064
rect 6636 1076 6644 1084
rect 6604 1016 6612 1024
rect 6492 976 6500 984
rect 6508 976 6516 984
rect 6588 956 6596 964
rect 6652 936 6660 944
rect 6300 916 6308 924
rect 6380 916 6388 924
rect 6428 916 6436 924
rect 6268 896 6276 904
rect 6300 856 6308 864
rect 6316 836 6324 844
rect 6364 756 6372 764
rect 6284 716 6292 724
rect 6620 916 6628 924
rect 6524 896 6532 904
rect 6588 896 6596 904
rect 6636 876 6644 884
rect 6764 1436 6772 1444
rect 6796 1316 6804 1324
rect 6844 1316 6852 1324
rect 6732 1256 6740 1264
rect 6764 1296 6772 1304
rect 6748 1176 6756 1184
rect 6780 1136 6788 1144
rect 7052 1476 7060 1484
rect 7068 1456 7076 1464
rect 6972 1436 6980 1444
rect 7004 1436 7012 1444
rect 7052 1436 7060 1444
rect 6908 1416 6916 1424
rect 6988 1416 6996 1424
rect 6956 1396 6964 1404
rect 6876 1336 6884 1344
rect 6892 1316 6900 1324
rect 6876 1296 6884 1304
rect 6924 1276 6932 1284
rect 6908 1256 6916 1264
rect 6828 1156 6836 1164
rect 6892 1116 6900 1124
rect 6684 1076 6692 1084
rect 6812 1076 6820 1084
rect 6876 1076 6884 1084
rect 6716 1016 6724 1024
rect 6684 956 6692 964
rect 6604 856 6612 864
rect 6668 856 6676 864
rect 6460 736 6468 744
rect 6204 696 6212 704
rect 6444 696 6452 704
rect 6492 716 6500 724
rect 6540 716 6548 724
rect 6572 716 6580 724
rect 6332 676 6340 684
rect 6380 676 6388 684
rect 6508 676 6516 684
rect 6140 556 6148 564
rect 6268 656 6276 664
rect 6188 556 6196 564
rect 6236 556 6244 564
rect 6204 536 6212 544
rect 6268 536 6276 544
rect 6156 516 6164 524
rect 6092 496 6100 504
rect 6172 436 6180 444
rect 6140 376 6148 384
rect 6156 376 6164 384
rect 6124 316 6132 324
rect 6156 336 6164 344
rect 6220 416 6228 424
rect 6188 376 6196 384
rect 6204 376 6212 384
rect 6172 316 6180 324
rect 6092 276 6100 284
rect 5900 216 5908 224
rect 5923 206 5931 214
rect 5933 206 5941 214
rect 5943 206 5951 214
rect 5953 206 5961 214
rect 5963 206 5971 214
rect 5973 206 5981 214
rect 5996 196 6004 204
rect 5900 176 5908 184
rect 5964 156 5972 164
rect 6252 356 6260 364
rect 6284 356 6292 364
rect 6220 336 6228 344
rect 6124 276 6132 284
rect 6204 276 6212 284
rect 6108 236 6116 244
rect 6108 216 6116 224
rect 6188 256 6196 264
rect 6284 256 6292 264
rect 6124 196 6132 204
rect 6156 176 6164 184
rect 6172 176 6180 184
rect 6204 176 6212 184
rect 6604 696 6612 704
rect 6588 676 6596 684
rect 6492 616 6500 624
rect 6428 596 6436 604
rect 6476 536 6484 544
rect 6380 516 6388 524
rect 6492 496 6500 504
rect 6492 436 6500 444
rect 6316 376 6324 384
rect 6364 376 6372 384
rect 6572 656 6580 664
rect 6572 596 6580 604
rect 6540 556 6548 564
rect 6524 376 6532 384
rect 6316 356 6324 364
rect 6412 356 6420 364
rect 6492 356 6500 364
rect 6476 316 6484 324
rect 6380 296 6388 304
rect 6348 276 6356 284
rect 6396 276 6404 284
rect 6380 256 6388 264
rect 6460 256 6468 264
rect 6396 236 6404 244
rect 6428 216 6436 224
rect 5932 96 5940 104
rect 6012 96 6020 104
rect 6076 96 6084 104
rect 6300 156 6308 164
rect 6188 96 6196 104
rect 6412 116 6420 124
rect 6268 96 6276 104
rect 6476 116 6484 124
rect 6508 296 6516 304
rect 6508 196 6516 204
rect 6652 616 6660 624
rect 6700 916 6708 924
rect 6716 756 6724 764
rect 6700 716 6708 724
rect 6684 596 6692 604
rect 6620 576 6628 584
rect 6652 576 6660 584
rect 6764 916 6772 924
rect 6876 996 6884 1004
rect 6828 936 6836 944
rect 6764 896 6772 904
rect 6780 896 6788 904
rect 6844 896 6852 904
rect 6876 896 6884 904
rect 6764 876 6772 884
rect 6780 876 6788 884
rect 6812 856 6820 864
rect 6860 876 6868 884
rect 6876 856 6884 864
rect 6940 1096 6948 1104
rect 7020 1316 7028 1324
rect 7020 1296 7028 1304
rect 7004 1116 7012 1124
rect 6956 1036 6964 1044
rect 6956 1016 6964 1024
rect 7020 1076 7028 1084
rect 7004 1056 7012 1064
rect 6988 1016 6996 1024
rect 7036 1016 7044 1024
rect 6972 996 6980 1004
rect 6988 976 6996 984
rect 7036 956 7044 964
rect 7084 1396 7092 1404
rect 7228 1716 7236 1724
rect 7228 1696 7236 1704
rect 7164 1616 7172 1624
rect 7212 1616 7220 1624
rect 7180 1556 7188 1564
rect 7196 1556 7204 1564
rect 7324 2216 7332 2224
rect 7308 2156 7316 2164
rect 7404 2896 7412 2904
rect 7388 2516 7396 2524
rect 7356 2496 7364 2504
rect 7356 2336 7364 2344
rect 7356 2276 7364 2284
rect 7340 2116 7348 2124
rect 7340 2096 7348 2104
rect 7308 1896 7316 1904
rect 7324 1836 7332 1844
rect 7292 1776 7300 1784
rect 7340 1756 7348 1764
rect 7308 1736 7316 1744
rect 7404 2096 7412 2104
rect 7372 2076 7380 2084
rect 7260 1716 7268 1724
rect 7292 1716 7300 1724
rect 7244 1516 7252 1524
rect 7212 1476 7220 1484
rect 7068 1316 7076 1324
rect 7100 1316 7108 1324
rect 7068 1096 7076 1104
rect 7084 1016 7092 1024
rect 6924 936 6932 944
rect 7036 936 7044 944
rect 7052 936 7060 944
rect 6940 916 6948 924
rect 6988 896 6996 904
rect 6924 876 6932 884
rect 6972 796 6980 804
rect 6908 756 6916 764
rect 6892 716 6900 724
rect 6812 696 6820 704
rect 6828 696 6836 704
rect 6860 696 6868 704
rect 6780 656 6788 664
rect 6828 656 6836 664
rect 6844 656 6852 664
rect 6748 636 6756 644
rect 6716 556 6724 564
rect 6764 556 6772 564
rect 6700 536 6708 544
rect 6652 516 6660 524
rect 6716 516 6724 524
rect 6732 436 6740 444
rect 6668 416 6676 424
rect 6748 416 6756 424
rect 6572 336 6580 344
rect 6684 316 6692 324
rect 6556 276 6564 284
rect 6636 276 6644 284
rect 6588 256 6596 264
rect 6620 236 6628 244
rect 6652 236 6660 244
rect 6700 236 6708 244
rect 6540 156 6548 164
rect 6604 156 6612 164
rect 6876 636 6884 644
rect 6956 716 6964 724
rect 6924 656 6932 664
rect 6972 636 6980 644
rect 6956 556 6964 564
rect 6860 536 6868 544
rect 6940 516 6948 524
rect 6780 476 6788 484
rect 7068 916 7076 924
rect 7084 916 7092 924
rect 7084 896 7092 904
rect 7068 776 7076 784
rect 7244 1456 7252 1464
rect 7164 1396 7172 1404
rect 7276 1676 7284 1684
rect 7276 1556 7284 1564
rect 7324 1536 7332 1544
rect 7276 1496 7284 1504
rect 7292 1456 7300 1464
rect 7308 1436 7316 1444
rect 7276 1416 7284 1424
rect 7180 1376 7188 1384
rect 7164 1316 7172 1324
rect 7164 956 7172 964
rect 7100 756 7108 764
rect 7052 736 7060 744
rect 7004 656 7012 664
rect 7036 656 7044 664
rect 7036 636 7044 644
rect 7148 916 7156 924
rect 7132 736 7140 744
rect 7116 716 7124 724
rect 7132 716 7140 724
rect 7068 696 7076 704
rect 7052 596 7060 604
rect 7004 576 7012 584
rect 7036 576 7044 584
rect 6988 516 6996 524
rect 6988 496 6996 504
rect 6956 456 6964 464
rect 7052 516 7060 524
rect 7100 676 7108 684
rect 7116 656 7124 664
rect 7148 656 7156 664
rect 7084 576 7092 584
rect 7020 476 7028 484
rect 7068 476 7076 484
rect 6780 436 6788 444
rect 7004 436 7012 444
rect 6876 376 6884 384
rect 6764 356 6772 364
rect 6796 336 6804 344
rect 6860 336 6868 344
rect 6780 316 6788 324
rect 6716 216 6724 224
rect 6748 216 6756 224
rect 6988 336 6996 344
rect 6828 296 6836 304
rect 6924 296 6932 304
rect 6988 296 6996 304
rect 6796 216 6804 224
rect 6700 176 6708 184
rect 6764 176 6772 184
rect 6732 156 6740 164
rect 6876 276 6884 284
rect 6972 196 6980 204
rect 6892 176 6900 184
rect 6748 136 6756 144
rect 6780 136 6788 144
rect 6668 116 6676 124
rect 6844 116 6852 124
rect 6876 116 6884 124
rect 6636 96 6644 104
rect 6700 96 6708 104
rect 7020 396 7028 404
rect 7036 336 7044 344
rect 7004 276 7012 284
rect 7036 276 7044 284
rect 7100 536 7108 544
rect 7132 536 7140 544
rect 7260 1296 7268 1304
rect 7292 1396 7300 1404
rect 7308 1376 7316 1384
rect 7308 1356 7316 1364
rect 7196 976 7204 984
rect 7276 1036 7284 1044
rect 7244 996 7252 1004
rect 7260 976 7268 984
rect 7244 956 7252 964
rect 7228 936 7236 944
rect 7196 876 7204 884
rect 7228 896 7236 904
rect 7244 756 7252 764
rect 7228 736 7236 744
rect 7196 716 7204 724
rect 7212 716 7220 724
rect 7196 636 7204 644
rect 7180 536 7188 544
rect 7100 476 7108 484
rect 7132 476 7140 484
rect 7180 436 7188 444
rect 7164 296 7172 304
rect 7276 736 7284 744
rect 7276 656 7284 664
rect 7308 1156 7316 1164
rect 7356 1476 7364 1484
rect 7340 1356 7348 1364
rect 7356 1336 7364 1344
rect 7340 1316 7348 1324
rect 7372 1316 7380 1324
rect 7324 1116 7332 1124
rect 7356 1116 7364 1124
rect 7340 1096 7348 1104
rect 7308 1076 7316 1084
rect 7356 1056 7364 1064
rect 7324 956 7332 964
rect 7340 936 7348 944
rect 7324 916 7332 924
rect 7308 836 7316 844
rect 7324 676 7332 684
rect 7372 776 7380 784
rect 7292 636 7300 644
rect 7340 636 7348 644
rect 7260 576 7268 584
rect 7292 516 7300 524
rect 7068 276 7076 284
rect 7084 276 7092 284
rect 7116 276 7124 284
rect 7132 276 7140 284
rect 7052 196 7060 204
rect 7020 176 7028 184
rect 7068 176 7076 184
rect 7228 256 7236 264
rect 7116 176 7124 184
rect 7164 156 7172 164
rect 7292 316 7300 324
rect 7276 276 7284 284
rect 6908 116 6916 124
rect 7052 116 7060 124
rect 7084 116 7092 124
rect 7100 116 7108 124
rect 7148 116 7156 124
rect 6876 96 6884 104
rect 6956 96 6964 104
rect 7388 156 7396 164
rect 7356 136 7364 144
rect 7260 96 7268 104
rect 5884 76 5892 84
rect 6172 76 6180 84
rect 6204 76 6212 84
rect 6428 76 6436 84
rect 6748 76 6756 84
rect 6908 76 6916 84
rect 6924 76 6932 84
rect 7100 76 7108 84
rect 4988 16 4996 24
rect 6412 16 6420 24
<< metal3 >>
rect 2914 5414 2974 5416
rect 2914 5406 2915 5414
rect 2924 5406 2925 5414
rect 2963 5406 2964 5414
rect 2973 5406 2974 5414
rect 2914 5404 2974 5406
rect 5922 5414 5982 5416
rect 5922 5406 5923 5414
rect 5932 5406 5933 5414
rect 5971 5406 5972 5414
rect 5981 5406 5982 5414
rect 5922 5404 5982 5406
rect 6020 5397 7340 5403
rect 628 5377 796 5383
rect 1412 5377 1548 5383
rect 3812 5377 3996 5383
rect 4292 5377 4604 5383
rect 4612 5377 6172 5383
rect 6260 5377 6988 5383
rect 532 5357 988 5363
rect 1540 5357 1628 5363
rect 2020 5357 2204 5363
rect 2324 5357 2508 5363
rect 3684 5357 3756 5363
rect 3764 5357 3884 5363
rect 4004 5357 5276 5363
rect 5908 5357 6476 5363
rect -35 5337 12 5343
rect 148 5337 172 5343
rect 260 5337 332 5343
rect 340 5337 524 5343
rect 612 5337 668 5343
rect 804 5337 876 5343
rect 964 5337 1148 5343
rect 1197 5337 1596 5343
rect 1197 5324 1203 5337
rect 1940 5337 2268 5343
rect 2452 5337 2572 5343
rect 2676 5337 2748 5343
rect 2756 5337 2876 5343
rect 2900 5337 3212 5343
rect 3236 5337 3324 5343
rect 3332 5337 3516 5343
rect 3940 5337 4028 5343
rect 4100 5337 4108 5343
rect 4356 5337 4812 5343
rect 4916 5337 5100 5343
rect 5140 5337 5180 5343
rect 5220 5337 5404 5343
rect 5492 5337 5580 5343
rect 6068 5337 6364 5343
rect 6436 5337 6620 5343
rect 6820 5337 7228 5343
rect 7236 5337 7308 5343
rect 180 5317 284 5323
rect 292 5317 332 5323
rect 516 5317 636 5323
rect 708 5317 764 5323
rect 772 5317 956 5323
rect 1124 5317 1196 5323
rect 1444 5317 1660 5323
rect 1668 5317 1964 5323
rect 2180 5317 2220 5323
rect 2228 5317 2476 5323
rect 2484 5317 2524 5323
rect 2580 5317 2716 5323
rect 2788 5317 2908 5323
rect 3572 5317 3724 5323
rect 3972 5317 4108 5323
rect 4324 5317 4476 5323
rect 4884 5317 4972 5323
rect 5124 5317 5132 5323
rect 5172 5317 5292 5323
rect 5428 5317 5500 5323
rect 5652 5317 5724 5323
rect 5924 5317 6412 5323
rect 6980 5317 7004 5323
rect 7172 5317 7244 5323
rect -35 5297 60 5303
rect 164 5297 236 5303
rect 596 5297 652 5303
rect 676 5297 876 5303
rect 884 5297 908 5303
rect 916 5297 972 5303
rect 1076 5297 1276 5303
rect 1652 5297 2348 5303
rect 2836 5297 3036 5303
rect 3220 5297 3692 5303
rect 3700 5297 3980 5303
rect 4036 5297 4076 5303
rect 4084 5297 4252 5303
rect 4260 5297 4396 5303
rect 5300 5297 5932 5303
rect 6036 5297 6604 5303
rect 228 5277 316 5283
rect 324 5277 588 5283
rect 644 5277 732 5283
rect 756 5277 1004 5283
rect 1204 5277 2060 5283
rect 2404 5277 2988 5283
rect 3380 5277 4092 5283
rect 4116 5277 4444 5283
rect 4452 5277 4636 5283
rect 4644 5277 4940 5283
rect 5412 5277 6380 5283
rect 6596 5277 7244 5283
rect 132 5257 268 5263
rect 724 5257 1196 5263
rect 1220 5257 1580 5263
rect 1812 5257 4236 5263
rect 4836 5257 4876 5263
rect 4884 5257 4940 5263
rect 5117 5257 5852 5263
rect 212 5237 268 5243
rect 276 5237 956 5243
rect 1140 5237 1836 5243
rect 2148 5237 3196 5243
rect 5117 5243 5123 5257
rect 5860 5257 6124 5263
rect 6148 5257 6220 5263
rect 6404 5257 6444 5263
rect 4244 5237 5123 5243
rect 5460 5237 5708 5243
rect 5716 5237 6428 5243
rect 100 5217 460 5223
rect 484 5217 876 5223
rect 900 5217 1244 5223
rect 1284 5217 1324 5223
rect 1572 5217 1612 5223
rect 1620 5217 2316 5223
rect 2548 5217 2892 5223
rect 2916 5217 3100 5223
rect 3716 5217 3788 5223
rect 3796 5217 3916 5223
rect 5108 5217 6396 5223
rect 6605 5217 7356 5223
rect 1410 5214 1470 5216
rect 1410 5206 1411 5214
rect 1420 5206 1421 5214
rect 1459 5206 1460 5214
rect 1469 5206 1470 5214
rect 1410 5204 1470 5206
rect 4418 5214 4478 5216
rect 4418 5206 4419 5214
rect 4428 5206 4429 5214
rect 4467 5206 4468 5214
rect 4477 5206 4478 5214
rect 4418 5204 4478 5206
rect 500 5197 1388 5203
rect 1588 5197 3404 5203
rect 3892 5197 4044 5203
rect 5188 5197 5404 5203
rect 5780 5197 5868 5203
rect 6052 5197 6092 5203
rect 6605 5203 6611 5217
rect 7364 5217 7388 5223
rect 6132 5197 6611 5203
rect 6628 5197 6892 5203
rect 6900 5197 6908 5203
rect 7044 5197 7356 5203
rect 148 5177 636 5183
rect 852 5177 1100 5183
rect 1108 5177 1276 5183
rect 1284 5177 1948 5183
rect 2564 5177 3180 5183
rect 3220 5177 4300 5183
rect 4644 5177 4892 5183
rect 4900 5177 4924 5183
rect 5140 5177 5180 5183
rect 5188 5177 5500 5183
rect 5508 5177 6924 5183
rect 324 5157 684 5163
rect 692 5157 748 5163
rect 1156 5157 1308 5163
rect 1316 5157 1820 5163
rect 1908 5157 2060 5163
rect 2068 5157 2620 5163
rect 2708 5157 3468 5163
rect 3492 5157 3548 5163
rect 3556 5157 3756 5163
rect 3764 5157 4140 5163
rect 4164 5157 4284 5163
rect 4804 5157 6028 5163
rect 6068 5157 6492 5163
rect 6660 5157 6700 5163
rect 6740 5157 6844 5163
rect 6852 5157 7324 5163
rect 132 5137 220 5143
rect 388 5137 844 5143
rect 1012 5137 1212 5143
rect 1220 5137 1340 5143
rect 1348 5137 1516 5143
rect 1524 5137 1644 5143
rect 2244 5137 3164 5143
rect 3300 5137 3628 5143
rect 3636 5137 3948 5143
rect 3956 5137 4204 5143
rect 4228 5137 4412 5143
rect 4516 5137 4908 5143
rect 4916 5137 5100 5143
rect 5412 5137 6556 5143
rect 116 5117 156 5123
rect 324 5117 380 5123
rect 676 5117 764 5123
rect 788 5117 812 5123
rect 932 5117 1036 5123
rect 1076 5117 1132 5123
rect 1140 5117 1228 5123
rect 1268 5117 1708 5123
rect 1716 5117 2172 5123
rect 2189 5117 2492 5123
rect 2189 5104 2195 5117
rect 2884 5117 3116 5123
rect 3188 5117 3356 5123
rect 3476 5117 3660 5123
rect 3716 5117 3804 5123
rect 3828 5117 4156 5123
rect 4244 5117 4268 5123
rect 4692 5117 5443 5123
rect 452 5097 508 5103
rect 612 5097 716 5103
rect 724 5097 796 5103
rect 820 5097 892 5103
rect 1044 5097 1148 5103
rect 1204 5097 1324 5103
rect 1332 5097 1692 5103
rect 1732 5097 1788 5103
rect 1828 5097 1868 5103
rect 2004 5097 2076 5103
rect 2100 5097 2188 5103
rect 2324 5097 2396 5103
rect 2500 5097 2684 5103
rect 2740 5097 3020 5103
rect 3108 5097 3148 5103
rect 3204 5097 3340 5103
rect 3380 5097 3388 5103
rect 3460 5097 3724 5103
rect 3940 5097 4012 5103
rect 4036 5097 4044 5103
rect 4180 5097 4236 5103
rect 4244 5097 4604 5103
rect 4676 5097 4764 5103
rect 5044 5097 5148 5103
rect 5437 5103 5443 5117
rect 5492 5117 5532 5123
rect 5556 5117 6067 5123
rect 6061 5104 6067 5117
rect 6148 5117 6204 5123
rect 6244 5117 6339 5123
rect 6333 5104 6339 5117
rect 6388 5117 6524 5123
rect 6628 5117 6716 5123
rect 5437 5097 5852 5103
rect 5908 5097 6012 5103
rect 6068 5097 6076 5103
rect 6180 5097 6284 5103
rect 6340 5097 6892 5103
rect 7108 5097 7228 5103
rect 180 5077 268 5083
rect 340 5077 476 5083
rect 628 5077 684 5083
rect 740 5077 812 5083
rect 884 5077 940 5083
rect 980 5077 1052 5083
rect 1124 5077 1148 5083
rect 1428 5077 1548 5083
rect 1604 5077 1660 5083
rect 1764 5077 1804 5083
rect 1821 5077 2012 5083
rect 36 5057 204 5063
rect 260 5057 348 5063
rect 468 5057 572 5063
rect 852 5057 892 5063
rect 1028 5057 1356 5063
rect 1604 5057 1708 5063
rect 1821 5063 1827 5077
rect 2020 5077 2028 5083
rect 2244 5077 2364 5083
rect 2596 5077 2988 5083
rect 3012 5077 3244 5083
rect 3284 5077 3459 5083
rect 1748 5057 1827 5063
rect 2004 5057 2028 5063
rect 2420 5057 2483 5063
rect 660 5037 1068 5043
rect 1108 5037 1388 5043
rect 1444 5037 1676 5043
rect 1693 5037 1884 5043
rect 52 5017 236 5023
rect 276 5017 876 5023
rect 980 5017 1612 5023
rect 1693 5023 1699 5037
rect 1956 5037 1996 5043
rect 2436 5037 2460 5043
rect 2477 5043 2483 5057
rect 2564 5057 3148 5063
rect 3332 5057 3436 5063
rect 3453 5063 3459 5077
rect 3476 5077 3644 5083
rect 3652 5077 3660 5083
rect 3668 5077 3820 5083
rect 3828 5077 3932 5083
rect 3972 5077 4028 5083
rect 4100 5077 4300 5083
rect 4308 5077 4684 5083
rect 4740 5077 5436 5083
rect 5460 5077 5548 5083
rect 5732 5077 5756 5083
rect 5988 5077 6188 5083
rect 6564 5077 6636 5083
rect 3453 5057 3484 5063
rect 3620 5057 3692 5063
rect 3709 5057 3740 5063
rect 2477 5037 3644 5043
rect 3709 5043 3715 5057
rect 3796 5057 3980 5063
rect 4068 5057 4108 5063
rect 4196 5057 4252 5063
rect 4292 5057 4908 5063
rect 5076 5057 5228 5063
rect 5236 5057 5660 5063
rect 5668 5057 6172 5063
rect 6260 5057 6540 5063
rect 6580 5057 6716 5063
rect 6900 5057 6972 5063
rect 3668 5037 3715 5043
rect 3732 5037 3756 5043
rect 4004 5037 4364 5043
rect 4644 5037 4684 5043
rect 4724 5037 5196 5043
rect 5396 5037 5580 5043
rect 5604 5037 5772 5043
rect 5789 5037 6003 5043
rect 1652 5017 1699 5023
rect 1716 5017 1740 5023
rect 1796 5017 1820 5023
rect 2020 5017 2220 5023
rect 2356 5017 2572 5023
rect 2996 5017 3852 5023
rect 3876 5017 4028 5023
rect 4036 5017 4236 5023
rect 4244 5017 4540 5023
rect 4628 5017 4732 5023
rect 5300 5017 5516 5023
rect 5789 5023 5795 5037
rect 5716 5017 5795 5023
rect 5997 5023 6003 5037
rect 6100 5037 6300 5043
rect 6324 5037 6348 5043
rect 6468 5037 6828 5043
rect 6948 5037 7052 5043
rect 5997 5017 6396 5023
rect 6612 5017 6668 5023
rect 2914 5014 2974 5016
rect 2914 5006 2915 5014
rect 2924 5006 2925 5014
rect 2963 5006 2964 5014
rect 2973 5006 2974 5014
rect 2914 5004 2974 5006
rect 5922 5014 5982 5016
rect 5922 5006 5923 5014
rect 5932 5006 5933 5014
rect 5971 5006 5972 5014
rect 5981 5006 5982 5014
rect 5922 5004 5982 5006
rect 356 4997 460 5003
rect 868 4997 924 5003
rect 996 4997 1020 5003
rect 1044 4997 2428 5003
rect 2564 4997 2812 5003
rect 3188 4997 3820 5003
rect 4116 4997 4700 5003
rect 4708 4997 5132 5003
rect 5140 4997 5484 5003
rect 5492 4997 5500 5003
rect 5508 4997 5788 5003
rect 6020 4997 6060 5003
rect 6084 4997 6220 5003
rect 6244 4997 6540 5003
rect 6596 4997 6748 5003
rect 6756 4997 6844 5003
rect 580 4977 604 4983
rect 644 4977 748 4983
rect 772 4977 1036 4983
rect 1060 4977 1148 4983
rect 1172 4977 1548 4983
rect 1652 4977 1708 4983
rect 1748 4977 1948 4983
rect 1956 4977 1996 4983
rect 2180 4977 2300 4983
rect 2308 4977 2316 4983
rect 2756 4977 3180 4983
rect 3188 4977 3660 4983
rect 3668 4977 3900 4983
rect 3908 4977 4332 4983
rect 4356 4977 4556 4983
rect 4564 4977 5180 4983
rect 5188 4977 5372 4983
rect 5389 4977 5468 4983
rect 84 4957 124 4963
rect 388 4957 508 4963
rect 548 4957 588 4963
rect 596 4957 1036 4963
rect 1284 4957 1484 4963
rect 1652 4957 1692 4963
rect 1780 4957 1964 4963
rect 1972 4957 2108 4963
rect 2244 4957 2300 4963
rect 2500 4957 2508 4963
rect 2516 4957 3116 4963
rect 3172 4957 3436 4963
rect 3460 4957 3484 4963
rect 3492 4957 3628 4963
rect 3652 4957 3724 4963
rect 3748 4957 3756 4963
rect 3940 4957 3948 4963
rect 3988 4957 3996 4963
rect 4004 4957 4316 4963
rect 4324 4957 4492 4963
rect 4500 4957 4716 4963
rect 4740 4957 4764 4963
rect 4820 4957 5123 4963
rect 52 4937 140 4943
rect 324 4937 364 4943
rect 372 4937 412 4943
rect 452 4937 492 4943
rect 532 4937 668 4943
rect 676 4937 828 4943
rect 836 4937 988 4943
rect 1044 4937 1052 4943
rect 1060 4937 1100 4943
rect 1476 4937 1532 4943
rect 1540 4937 1596 4943
rect 1668 4937 2092 4943
rect 2100 4937 2316 4943
rect 2340 4937 2364 4943
rect 2381 4937 2428 4943
rect 132 4917 156 4923
rect 276 4917 636 4923
rect 724 4917 780 4923
rect 797 4917 956 4923
rect -35 4897 12 4903
rect 436 4897 460 4903
rect 564 4897 588 4903
rect 660 4897 732 4903
rect 797 4903 803 4917
rect 996 4917 1084 4923
rect 1092 4917 1116 4923
rect 1524 4917 1580 4923
rect 1636 4917 1660 4923
rect 1668 4917 1740 4923
rect 1764 4917 1804 4923
rect 1940 4917 2076 4923
rect 2100 4917 2236 4923
rect 2381 4923 2387 4937
rect 2452 4937 2508 4943
rect 2532 4937 3148 4943
rect 3172 4937 3244 4943
rect 3364 4937 3612 4943
rect 3620 4937 4060 4943
rect 4068 4937 4572 4943
rect 4580 4937 4860 4943
rect 4868 4937 5100 4943
rect 5117 4943 5123 4957
rect 5389 4963 5395 4977
rect 5540 4977 5763 4983
rect 5204 4957 5395 4963
rect 5412 4957 5452 4963
rect 5684 4957 5740 4963
rect 5757 4963 5763 4977
rect 5860 4977 6652 4983
rect 6660 4977 6668 4983
rect 6676 4977 6908 4983
rect 6916 4977 7052 4983
rect 7060 4977 7212 4983
rect 5757 4957 6012 4963
rect 6052 4957 6156 4963
rect 6276 4957 6332 4963
rect 6452 4957 6524 4963
rect 6548 4957 6620 4963
rect 6724 4957 7036 4963
rect 7284 4957 7340 4963
rect 5117 4937 5436 4943
rect 5444 4937 5852 4943
rect 5908 4937 5939 4943
rect 2244 4917 2387 4923
rect 2404 4917 2524 4923
rect 2756 4917 2812 4923
rect 2884 4917 2940 4923
rect 2948 4917 3036 4923
rect 3044 4917 3100 4923
rect 3165 4923 3171 4936
rect 3108 4917 3171 4923
rect 3268 4917 3388 4923
rect 3412 4917 3468 4923
rect 3540 4917 3676 4923
rect 3716 4917 3756 4923
rect 3764 4917 3964 4923
rect 3972 4917 4124 4923
rect 4180 4917 4204 4923
rect 4260 4917 4540 4923
rect 4548 4917 4588 4923
rect 4756 4917 4828 4923
rect 4964 4917 4988 4923
rect 5044 4917 5068 4923
rect 5124 4917 5484 4923
rect 5492 4917 5644 4923
rect 5764 4917 5916 4923
rect 5933 4923 5939 4937
rect 6068 4937 6428 4943
rect 6500 4937 6764 4943
rect 5933 4917 6076 4923
rect 6164 4917 6268 4923
rect 6292 4917 6540 4923
rect 6596 4917 6732 4923
rect 6820 4917 6892 4923
rect 6900 4917 6956 4923
rect 788 4897 803 4903
rect 820 4897 860 4903
rect 868 4897 1036 4903
rect 1076 4897 1372 4903
rect 1380 4897 1804 4903
rect 1860 4897 1900 4903
rect 1956 4897 1980 4903
rect 2036 4897 2060 4903
rect 2356 4897 2572 4903
rect 2756 4897 2844 4903
rect 2932 4897 3068 4903
rect 3389 4897 3644 4903
rect 916 4877 1164 4883
rect 1364 4877 1628 4883
rect 1828 4877 2124 4883
rect 2132 4877 2220 4883
rect 2349 4883 2355 4896
rect 2228 4877 2355 4883
rect 2580 4877 2892 4883
rect 3389 4883 3395 4897
rect 3668 4897 3692 4903
rect 3828 4897 3868 4903
rect 4148 4897 4220 4903
rect 4372 4897 4508 4903
rect 4756 4897 4812 4903
rect 4820 4897 4828 4903
rect 4916 4897 5052 4903
rect 5140 4897 5571 4903
rect 3092 4877 3395 4883
rect 3508 4877 3580 4883
rect 3588 4877 3852 4883
rect 3860 4877 3980 4883
rect 3988 4877 4092 4883
rect 4100 4877 4156 4883
rect 4164 4877 4748 4883
rect 4900 4877 4988 4883
rect 4996 4877 5148 4883
rect 5316 4877 5420 4883
rect 5508 4877 5548 4883
rect 5565 4883 5571 4897
rect 5652 4897 5724 4903
rect 5748 4897 5932 4903
rect 6116 4897 6284 4903
rect 6292 4897 6508 4903
rect 6516 4897 6524 4903
rect 6644 4897 6908 4903
rect 5565 4877 5676 4883
rect 5725 4883 5731 4896
rect 5725 4877 5836 4883
rect 5860 4877 6460 4883
rect 6525 4877 6604 4883
rect 980 4857 1212 4863
rect 1572 4857 1724 4863
rect 1812 4857 1884 4863
rect 2004 4857 2332 4863
rect 3028 4857 3052 4863
rect 3556 4857 3708 4863
rect 3972 4857 5148 4863
rect 5428 4857 5980 4863
rect 5988 4857 6252 4863
rect 6525 4863 6531 4877
rect 7076 4877 7148 4883
rect 7188 4877 7196 4883
rect 7204 4877 7276 4883
rect 7284 4877 7324 4883
rect 6436 4857 6531 4863
rect 6548 4857 6700 4863
rect 6708 4857 6828 4863
rect 7188 4857 7212 4863
rect 692 4837 892 4843
rect 900 4837 988 4843
rect 1028 4837 1596 4843
rect 1636 4837 1916 4843
rect 1972 4837 2620 4843
rect 3380 4837 3420 4843
rect 3444 4837 3932 4843
rect 3988 4837 4076 4843
rect 4132 4837 4732 4843
rect 4804 4837 5004 4843
rect 5092 4837 5228 4843
rect 5572 4837 5868 4843
rect 5876 4837 6140 4843
rect 6148 4837 6236 4843
rect 6244 4837 6652 4843
rect 6660 4837 6668 4843
rect 6836 4837 6860 4843
rect 260 4817 1228 4823
rect 1492 4817 2012 4823
rect 3380 4817 3708 4823
rect 3780 4817 4044 4823
rect 4068 4817 4236 4823
rect 4676 4817 4764 4823
rect 4804 4817 4892 4823
rect 4916 4817 5868 4823
rect 6004 4817 6348 4823
rect 6484 4817 6540 4823
rect 1410 4814 1470 4816
rect 1410 4806 1411 4814
rect 1420 4806 1421 4814
rect 1459 4806 1460 4814
rect 1469 4806 1470 4814
rect 1410 4804 1470 4806
rect 4418 4814 4478 4816
rect 4418 4806 4419 4814
rect 4428 4806 4429 4814
rect 4467 4806 4468 4814
rect 4477 4806 4478 4814
rect 4418 4804 4478 4806
rect 308 4797 1308 4803
rect 1588 4797 1660 4803
rect 1972 4797 2012 4803
rect 2628 4797 2764 4803
rect 2868 4797 4131 4803
rect 1780 4777 1948 4783
rect 2532 4777 2604 4783
rect 2676 4777 3036 4783
rect 3604 4777 3804 4783
rect 3812 4777 4044 4783
rect 4052 4777 4108 4783
rect 4125 4783 4131 4797
rect 4596 4797 4668 4803
rect 4772 4797 4876 4803
rect 4916 4797 6156 4803
rect 6196 4797 6956 4803
rect 4125 4777 4908 4783
rect 5092 4777 5132 4783
rect 5700 4777 5740 4783
rect 5828 4777 6028 4783
rect 6052 4777 6300 4783
rect 6308 4777 6380 4783
rect 596 4757 1068 4763
rect 2020 4757 2108 4763
rect 2292 4757 2364 4763
rect 2564 4757 2732 4763
rect 2772 4757 4035 4763
rect 84 4737 700 4743
rect 916 4737 1164 4743
rect 1268 4737 1356 4743
rect 1684 4737 1756 4743
rect 1764 4737 1804 4743
rect 2036 4737 2188 4743
rect 2260 4737 2316 4743
rect 2324 4737 2412 4743
rect 2420 4737 2636 4743
rect 2644 4737 2796 4743
rect 3620 4737 3660 4743
rect 4029 4743 4035 4757
rect 4052 4757 4172 4763
rect 4189 4757 4972 4763
rect 4189 4743 4195 4757
rect 5012 4757 5132 4763
rect 5428 4757 6124 4763
rect 6340 4757 6604 4763
rect 6612 4757 6908 4763
rect 7092 4757 7180 4763
rect 3668 4737 4019 4743
rect 4029 4737 4195 4743
rect 4013 4724 4019 4737
rect 4404 4737 4492 4743
rect 4932 4737 5068 4743
rect 5332 4737 5852 4743
rect 6180 4737 6444 4743
rect 6660 4737 6796 4743
rect 7156 4737 7164 4743
rect 7188 4737 7260 4743
rect 1204 4717 1532 4723
rect 1748 4717 1820 4723
rect 1828 4717 1852 4723
rect 2100 4717 2140 4723
rect 2164 4717 2188 4723
rect 2196 4717 2380 4723
rect 2740 4717 2844 4723
rect 2852 4717 2924 4723
rect 3364 4717 3628 4723
rect 3684 4717 3980 4723
rect 4020 4717 4060 4723
rect 4596 4717 5123 4723
rect 164 4697 204 4703
rect 372 4697 412 4703
rect 436 4697 556 4703
rect 580 4697 780 4703
rect 1124 4697 1180 4703
rect 1213 4697 1372 4703
rect 1213 4684 1219 4697
rect 1396 4697 1580 4703
rect 1716 4697 1836 4703
rect 1988 4697 1996 4703
rect 2516 4697 2572 4703
rect 2612 4697 2700 4703
rect 2708 4697 2748 4703
rect 2820 4697 2940 4703
rect 3172 4697 3228 4703
rect 3572 4697 3836 4703
rect 3924 4697 3964 4703
rect 4068 4697 4188 4703
rect 4212 4697 4348 4703
rect 4628 4697 4860 4703
rect 5028 4697 5068 4703
rect 5117 4703 5123 4717
rect 5172 4717 5276 4723
rect 5348 4717 5564 4723
rect 5828 4717 5868 4723
rect 5892 4717 5923 4723
rect 5117 4697 5836 4703
rect 5844 4697 5900 4703
rect 5917 4703 5923 4717
rect 6196 4717 6252 4723
rect 6580 4717 6652 4723
rect 7172 4717 7276 4723
rect 5917 4697 6252 4703
rect 6340 4697 6492 4703
rect 6772 4697 6780 4703
rect 7124 4697 7132 4703
rect 7172 4697 7292 4703
rect 100 4677 204 4683
rect 212 4677 236 4683
rect 244 4677 268 4683
rect 356 4677 380 4683
rect 452 4677 540 4683
rect 548 4677 620 4683
rect 628 4677 764 4683
rect 772 4677 828 4683
rect 1012 4677 1212 4683
rect 1604 4677 1612 4683
rect 1668 4677 1772 4683
rect 1940 4677 2156 4683
rect 2244 4677 2300 4683
rect 2660 4677 2684 4683
rect 2916 4677 3500 4683
rect 3700 4677 3820 4683
rect 4004 4677 4076 4683
rect 4244 4677 4732 4683
rect 4740 4677 4748 4683
rect 4788 4677 4876 4683
rect 4916 4677 5123 4683
rect 532 4657 556 4663
rect 740 4657 924 4663
rect 932 4657 972 4663
rect 980 4657 1020 4663
rect 1044 4657 1260 4663
rect 1652 4657 1923 4663
rect 516 4637 652 4643
rect 660 4637 684 4643
rect 708 4637 732 4643
rect 740 4637 892 4643
rect 1021 4643 1027 4656
rect 1021 4637 1084 4643
rect 1220 4637 1388 4643
rect 1748 4637 1804 4643
rect 1812 4637 1900 4643
rect 1917 4643 1923 4657
rect 2004 4657 2668 4663
rect 2852 4657 3228 4663
rect 3492 4657 3660 4663
rect 3844 4657 4684 4663
rect 4692 4657 5004 4663
rect 5060 4657 5084 4663
rect 5117 4663 5123 4677
rect 5204 4677 5292 4683
rect 5348 4677 5404 4683
rect 5732 4677 5820 4683
rect 6020 4677 6268 4683
rect 6276 4677 6300 4683
rect 6340 4677 6364 4683
rect 6580 4677 6684 4683
rect 6692 4677 6748 4683
rect 7092 4677 7244 4683
rect 5117 4657 5324 4663
rect 5892 4657 6188 4663
rect 6228 4657 6492 4663
rect 6644 4657 6684 4663
rect 6708 4657 6780 4663
rect 1917 4637 1996 4643
rect 2004 4637 2268 4643
rect 2740 4637 2860 4643
rect 3476 4637 3580 4643
rect 3588 4637 3724 4643
rect 3732 4637 3772 4643
rect 3789 4637 4636 4643
rect 724 4617 828 4623
rect 964 4617 1388 4623
rect 1876 4617 2316 4623
rect 3789 4623 3795 4637
rect 4756 4637 4780 4643
rect 5172 4637 5500 4643
rect 5540 4637 5580 4643
rect 5636 4637 6476 4643
rect 6484 4637 6988 4643
rect 6996 4637 7020 4643
rect 3284 4617 3795 4623
rect 3844 4617 3884 4623
rect 3940 4617 4172 4623
rect 4388 4617 5004 4623
rect 5028 4617 5308 4623
rect 5396 4617 5756 4623
rect 5780 4617 5868 4623
rect 6020 4617 6172 4623
rect 6420 4617 6428 4623
rect 6692 4617 6908 4623
rect 7220 4617 7276 4623
rect 2914 4614 2974 4616
rect 2914 4606 2915 4614
rect 2924 4606 2925 4614
rect 2963 4606 2964 4614
rect 2973 4606 2974 4614
rect 2914 4604 2974 4606
rect 5922 4614 5982 4616
rect 5922 4606 5923 4614
rect 5932 4606 5933 4614
rect 5971 4606 5972 4614
rect 5981 4606 5982 4614
rect 5922 4604 5982 4606
rect 733 4597 988 4603
rect 733 4583 739 4597
rect 996 4597 1004 4603
rect 1076 4597 1964 4603
rect 1988 4597 2060 4603
rect 2788 4597 2812 4603
rect 3460 4597 3676 4603
rect 3860 4597 3900 4603
rect 3908 4597 4076 4603
rect 4116 4597 4252 4603
rect 4260 4597 4764 4603
rect 5124 4597 5212 4603
rect 5588 4597 5804 4603
rect 5844 4597 5868 4603
rect 6116 4597 6140 4603
rect 6196 4597 6332 4603
rect 6340 4597 6380 4603
rect 6756 4597 7212 4603
rect 260 4577 739 4583
rect 820 4577 876 4583
rect 964 4577 1084 4583
rect 1092 4577 1452 4583
rect 1556 4577 1580 4583
rect 1876 4577 2044 4583
rect 2164 4577 2220 4583
rect 2228 4577 2556 4583
rect 3332 4577 3580 4583
rect 3588 4577 4364 4583
rect 4420 4577 4796 4583
rect 4804 4577 4876 4583
rect 5044 4577 5116 4583
rect 5204 4577 5452 4583
rect 5604 4577 5676 4583
rect 5764 4577 5900 4583
rect 5924 4577 6204 4583
rect 6292 4577 6732 4583
rect 6868 4577 6924 4583
rect 6932 4577 6956 4583
rect 6964 4577 7100 4583
rect 7252 4577 7276 4583
rect 20 4557 44 4563
rect 52 4557 220 4563
rect 340 4557 380 4563
rect 484 4557 588 4563
rect 596 4557 716 4563
rect 820 4557 844 4563
rect 900 4557 940 4563
rect 948 4557 1052 4563
rect 1060 4557 1116 4563
rect 1124 4557 1148 4563
rect 1492 4557 1571 4563
rect 84 4537 124 4543
rect 845 4543 851 4556
rect 845 4537 972 4543
rect 1172 4537 1212 4543
rect 1252 4537 1292 4543
rect 1364 4537 1532 4543
rect 1565 4543 1571 4557
rect 1588 4557 1644 4563
rect 1661 4557 1836 4563
rect 1661 4543 1667 4557
rect 1892 4557 1948 4563
rect 1956 4557 2028 4563
rect 2100 4557 2284 4563
rect 2500 4557 2748 4563
rect 3572 4557 3676 4563
rect 3693 4557 3708 4563
rect 1565 4537 1667 4543
rect 1684 4537 2508 4543
rect 2692 4537 2732 4543
rect 3220 4537 3308 4543
rect 3693 4543 3699 4557
rect 4068 4557 4188 4563
rect 4196 4557 4236 4563
rect 4276 4557 4300 4563
rect 4308 4557 4444 4563
rect 4452 4557 4476 4563
rect 4932 4557 5324 4563
rect 5469 4557 5884 4563
rect 3524 4537 3699 4543
rect 3716 4537 3772 4543
rect 3812 4537 4124 4543
rect 4164 4537 4588 4543
rect 4644 4537 4684 4543
rect 4692 4537 4908 4543
rect 4948 4537 5084 4543
rect 5156 4537 5244 4543
rect 5469 4543 5475 4557
rect 6116 4557 6156 4563
rect 6164 4557 6700 4563
rect 6836 4557 7020 4563
rect 7028 4557 7052 4563
rect 7060 4557 7132 4563
rect 7140 4557 7244 4563
rect 5268 4537 5475 4543
rect 5492 4537 5612 4543
rect 5620 4537 5708 4543
rect 5716 4537 5820 4543
rect 5828 4537 6044 4543
rect 6228 4537 6268 4543
rect 6404 4537 6620 4543
rect 6724 4537 6812 4543
rect 7012 4537 7180 4543
rect 7412 4537 7443 4543
rect 404 4517 508 4523
rect 644 4517 684 4523
rect 868 4517 924 4523
rect 964 4517 988 4523
rect 1204 4517 1228 4523
rect 1348 4517 1468 4523
rect 1508 4517 1596 4523
rect 1620 4517 1644 4523
rect 1748 4517 1884 4523
rect 1956 4517 1980 4523
rect 2116 4517 2204 4523
rect 2580 4517 2700 4523
rect 2772 4517 3276 4523
rect 3364 4517 3452 4523
rect 3636 4517 3948 4523
rect 3956 4517 4028 4523
rect 4084 4517 4284 4523
rect 4564 4517 4604 4523
rect 4628 4517 4748 4523
rect 4948 4517 5036 4523
rect 5236 4517 5324 4523
rect 5476 4517 5532 4523
rect 5556 4517 5660 4523
rect 5684 4517 5788 4523
rect 5860 4517 6124 4523
rect 6132 4517 6348 4523
rect 6356 4517 6396 4523
rect 6461 4517 6524 4523
rect 132 4497 188 4503
rect 292 4497 348 4503
rect 1076 4497 1132 4503
rect 1284 4497 1420 4503
rect 1556 4497 1580 4503
rect 1780 4497 1916 4503
rect 2308 4497 2348 4503
rect 2356 4497 2556 4503
rect 2612 4497 2668 4503
rect 3156 4497 3292 4503
rect 3300 4497 3356 4503
rect 3540 4497 3660 4503
rect 4244 4497 5068 4503
rect 5076 4497 5148 4503
rect 5364 4497 6051 4503
rect 708 4477 748 4483
rect 1044 4477 1068 4483
rect 1188 4477 1340 4483
rect 1396 4477 1516 4483
rect 1572 4477 2572 4483
rect 2580 4477 2716 4483
rect 4196 4477 4556 4483
rect 4596 4477 4668 4483
rect 5380 4477 5884 4483
rect 6045 4483 6051 4497
rect 6068 4497 6092 4503
rect 6228 4497 6300 4503
rect 6461 4503 6467 4517
rect 6708 4517 6940 4523
rect 7012 4517 7084 4523
rect 6388 4497 6467 4503
rect 6484 4497 6652 4503
rect 6708 4497 7036 4503
rect 7044 4497 7116 4503
rect 7300 4497 7443 4503
rect 6045 4477 6236 4483
rect 6340 4477 6412 4483
rect 6548 4477 6588 4483
rect 6612 4477 6652 4483
rect 6724 4477 6748 4483
rect 6916 4477 7004 4483
rect 308 4457 556 4463
rect 564 4457 1148 4463
rect 1252 4457 1372 4463
rect 1380 4457 1532 4463
rect 1780 4457 1820 4463
rect 1828 4457 2108 4463
rect 2388 4457 3052 4463
rect 3556 4457 4060 4463
rect 4132 4457 4460 4463
rect 4468 4457 4556 4463
rect 4724 4457 5356 4463
rect 5460 4457 5628 4463
rect 5636 4457 5724 4463
rect 5828 4457 5932 4463
rect 6004 4457 6140 4463
rect 6212 4457 6972 4463
rect 260 4437 460 4443
rect 468 4437 780 4443
rect 1156 4437 2156 4443
rect 2628 4437 2796 4443
rect 4500 4437 5180 4443
rect 5268 4437 5468 4443
rect 5508 4437 5580 4443
rect 5604 4437 5628 4443
rect 5668 4437 5811 4443
rect 3732 4417 4380 4423
rect 5252 4417 5484 4423
rect 5492 4417 5500 4423
rect 5508 4417 5580 4423
rect 5805 4423 5811 4437
rect 6100 4437 6716 4443
rect 5805 4417 6876 4423
rect 1410 4414 1470 4416
rect 1410 4406 1411 4414
rect 1420 4406 1421 4414
rect 1459 4406 1460 4414
rect 1469 4406 1470 4414
rect 1410 4404 1470 4406
rect 4418 4414 4478 4416
rect 4418 4406 4419 4414
rect 4428 4406 4429 4414
rect 4467 4406 4468 4414
rect 4477 4406 4478 4414
rect 4418 4404 4478 4406
rect 1668 4397 1756 4403
rect 3396 4397 4172 4403
rect 4500 4397 4652 4403
rect 4660 4397 4748 4403
rect 4884 4397 5292 4403
rect 5364 4397 5548 4403
rect 5604 4397 5756 4403
rect 5780 4397 6668 4403
rect 7108 4397 7148 4403
rect 1412 4377 1868 4383
rect 1876 4377 1932 4383
rect 1956 4377 2172 4383
rect 3700 4377 3756 4383
rect 3764 4377 3788 4383
rect 4212 4377 4540 4383
rect 4628 4377 4700 4383
rect 5012 4377 5388 4383
rect 5492 4377 5564 4383
rect 5572 4377 6572 4383
rect 6612 4377 6684 4383
rect 6692 4377 6844 4383
rect 7140 4377 7308 4383
rect 324 4357 444 4363
rect 452 4357 524 4363
rect 644 4357 892 4363
rect 932 4357 1196 4363
rect 1204 4357 1580 4363
rect 1588 4357 2364 4363
rect 3636 4357 3756 4363
rect 3764 4357 3804 4363
rect 4180 4357 4492 4363
rect 4564 4357 5132 4363
rect 5140 4357 5516 4363
rect 5524 4357 5612 4363
rect 5636 4357 6076 4363
rect 6132 4357 6732 4363
rect 6756 4357 6764 4363
rect 6772 4357 7084 4363
rect 7092 4357 7196 4363
rect 660 4337 780 4343
rect 788 4337 940 4343
rect 1092 4337 1308 4343
rect 1700 4337 1740 4343
rect 1812 4337 1852 4343
rect 1860 4337 1996 4343
rect 2004 4337 2092 4343
rect 2196 4337 2652 4343
rect 2788 4337 3916 4343
rect 4292 4337 4332 4343
rect 4340 4337 4588 4343
rect 4644 4337 4684 4343
rect 4692 4337 4732 4343
rect 4740 4337 5020 4343
rect 5044 4337 5516 4343
rect 5556 4337 5692 4343
rect 5764 4337 5788 4343
rect 5812 4337 5916 4343
rect 5940 4337 6012 4343
rect 6036 4337 6332 4343
rect 6468 4337 6572 4343
rect 6676 4337 7116 4343
rect 7156 4337 7164 4343
rect 20 4317 76 4323
rect 100 4317 108 4323
rect 116 4317 348 4323
rect 804 4317 828 4323
rect 868 4317 1228 4323
rect 1300 4317 1740 4323
rect 1757 4317 1820 4323
rect 84 4297 108 4303
rect 340 4297 396 4303
rect 564 4297 620 4303
rect 692 4297 732 4303
rect 740 4297 828 4303
rect 1108 4297 1132 4303
rect 1268 4297 1708 4303
rect 1757 4303 1763 4317
rect 1988 4317 1996 4323
rect 2004 4317 2348 4323
rect 3380 4317 3468 4323
rect 3588 4317 3635 4323
rect 1732 4297 1763 4303
rect 1796 4297 1884 4303
rect 1908 4297 2012 4303
rect 2084 4297 2124 4303
rect 2228 4297 2428 4303
rect 2484 4297 2636 4303
rect 2644 4297 2812 4303
rect 3044 4297 3596 4303
rect 3629 4303 3635 4317
rect 3652 4317 3724 4323
rect 3732 4317 3772 4323
rect 4372 4317 4540 4323
rect 4548 4317 4684 4323
rect 4900 4317 5020 4323
rect 5044 4317 5084 4323
rect 5204 4317 5468 4323
rect 5540 4317 5948 4323
rect 6068 4317 6284 4323
rect 6564 4317 6572 4323
rect 6580 4317 6604 4323
rect 6612 4317 6636 4323
rect 6660 4317 6796 4323
rect 6804 4317 6844 4323
rect 7172 4317 7308 4323
rect 3629 4297 3660 4303
rect 3780 4297 3900 4303
rect 3924 4297 4428 4303
rect 4804 4297 4876 4303
rect 4884 4297 5036 4303
rect 5220 4297 5491 4303
rect 100 4277 316 4283
rect 756 4277 876 4283
rect 1124 4277 1164 4283
rect 1572 4277 1612 4283
rect 1796 4277 1868 4283
rect 1892 4277 1964 4283
rect 2132 4277 2172 4283
rect 2404 4277 2444 4283
rect 2868 4277 3068 4283
rect 3156 4277 3452 4283
rect 3460 4277 3596 4283
rect 3716 4277 3788 4283
rect 3892 4277 4012 4283
rect 4308 4277 4460 4283
rect 5012 4277 5372 4283
rect 5380 4277 5420 4283
rect 5485 4283 5491 4297
rect 5508 4297 5612 4303
rect 5636 4297 5708 4303
rect 5796 4297 5916 4303
rect 5924 4297 6124 4303
rect 6196 4297 6236 4303
rect 6276 4297 6316 4303
rect 6324 4297 6684 4303
rect 6852 4297 6972 4303
rect 7124 4297 7164 4303
rect 5485 4277 5564 4283
rect 5588 4277 5676 4283
rect 5844 4277 6195 4283
rect 6189 4264 6195 4277
rect 6324 4277 6547 4283
rect 68 4257 156 4263
rect 212 4257 396 4263
rect 404 4257 428 4263
rect 532 4257 588 4263
rect 804 4257 1020 4263
rect 1037 4257 1148 4263
rect 356 4237 460 4243
rect 468 4237 668 4243
rect 1037 4243 1043 4257
rect 1364 4257 1388 4263
rect 1636 4257 1676 4263
rect 1684 4257 1932 4263
rect 2052 4257 2140 4263
rect 2324 4257 2348 4263
rect 3044 4257 3164 4263
rect 3412 4257 4060 4263
rect 4068 4257 4716 4263
rect 4724 4257 4828 4263
rect 4836 4257 4972 4263
rect 5085 4257 5164 4263
rect 868 4237 1043 4243
rect 1108 4237 1244 4243
rect 1332 4237 2748 4243
rect 2605 4224 2611 4237
rect 3252 4237 3500 4243
rect 3508 4237 3612 4243
rect 3700 4237 3740 4243
rect 3748 4237 4092 4243
rect 4132 4237 4140 4243
rect 4164 4237 4188 4243
rect 4244 4237 4284 4243
rect 4356 4237 4396 4243
rect 4468 4237 4668 4243
rect 5085 4243 5091 4257
rect 5284 4257 5292 4263
rect 5412 4257 5436 4263
rect 5620 4257 5740 4263
rect 5796 4257 5932 4263
rect 5956 4257 6092 4263
rect 6116 4257 6156 4263
rect 6196 4257 6332 4263
rect 6340 4257 6524 4263
rect 6541 4263 6547 4277
rect 6628 4277 7148 4283
rect 6541 4257 6876 4263
rect 7012 4257 7116 4263
rect 4868 4237 5091 4243
rect 5172 4237 5212 4243
rect 5332 4237 5532 4243
rect 5732 4237 5788 4243
rect 5805 4237 6028 4243
rect 708 4217 972 4223
rect 980 4217 1324 4223
rect 1924 4217 2044 4223
rect 2180 4217 2252 4223
rect 2260 4217 2300 4223
rect 2308 4217 2444 4223
rect 2468 4217 2556 4223
rect 3188 4217 3228 4223
rect 3236 4217 3276 4223
rect 3316 4217 4163 4223
rect 2914 4214 2974 4216
rect 2914 4206 2915 4214
rect 2924 4206 2925 4214
rect 2963 4206 2964 4214
rect 2973 4206 2974 4214
rect 2914 4204 2974 4206
rect 676 4197 748 4203
rect 964 4197 1052 4203
rect 1060 4197 1212 4203
rect 1220 4197 1644 4203
rect 2004 4197 2092 4203
rect 2164 4197 2396 4203
rect 2989 4197 3715 4203
rect 116 4177 188 4183
rect 756 4177 908 4183
rect 916 4177 1100 4183
rect 1140 4177 1468 4183
rect 1556 4177 1596 4183
rect 2052 4177 2172 4183
rect 2596 4177 2652 4183
rect 2989 4183 2995 4197
rect 2884 4177 2995 4183
rect 3364 4177 3468 4183
rect 3476 4177 3692 4183
rect 3709 4183 3715 4197
rect 3828 4197 3980 4203
rect 3988 4197 4140 4203
rect 4157 4203 4163 4217
rect 4452 4217 4924 4223
rect 5805 4223 5811 4237
rect 6052 4237 6083 4243
rect 5092 4217 5811 4223
rect 6020 4217 6060 4223
rect 6077 4223 6083 4237
rect 6100 4237 6156 4243
rect 6180 4237 6316 4243
rect 6388 4237 6412 4243
rect 6420 4237 6780 4243
rect 6788 4237 7020 4243
rect 7060 4237 7180 4243
rect 6077 4217 6316 4223
rect 7252 4217 7340 4223
rect 5922 4214 5982 4216
rect 5922 4206 5923 4214
rect 5932 4206 5933 4214
rect 5971 4206 5972 4214
rect 5981 4206 5982 4214
rect 5922 4204 5982 4206
rect 4157 4197 5340 4203
rect 5396 4197 5452 4203
rect 5460 4197 5676 4203
rect 5748 4197 5804 4203
rect 6004 4197 6124 4203
rect 6141 4197 6284 4203
rect 3709 4177 4268 4183
rect 5124 4177 5132 4183
rect 5188 4177 5324 4183
rect 5533 4177 6051 4183
rect 20 4157 108 4163
rect 132 4157 204 4163
rect 292 4157 460 4163
rect 580 4157 636 4163
rect 756 4157 812 4163
rect 900 4157 1004 4163
rect 1012 4157 1132 4163
rect 1236 4157 1340 4163
rect 1716 4157 1740 4163
rect 1828 4157 1900 4163
rect 2100 4157 2188 4163
rect 2532 4157 2540 4163
rect 2548 4157 2892 4163
rect 3092 4157 3164 4163
rect 3444 4157 3484 4163
rect 4356 4157 4428 4163
rect 4580 4157 4876 4163
rect 5028 4157 5276 4163
rect 5533 4163 5539 4177
rect 5284 4157 5539 4163
rect 5812 4157 5852 4163
rect 5924 4157 6028 4163
rect 6045 4163 6051 4177
rect 6141 4183 6147 4197
rect 6308 4197 6332 4203
rect 6596 4197 6684 4203
rect 6724 4197 6748 4203
rect 6100 4177 6147 4183
rect 6260 4177 6732 4183
rect 6740 4177 6924 4183
rect 7204 4177 7212 4183
rect 6045 4157 6460 4163
rect 6644 4157 6828 4163
rect 6836 4157 6892 4163
rect 7092 4157 7212 4163
rect 116 4137 172 4143
rect 548 4137 652 4143
rect 660 4137 684 4143
rect 740 4137 924 4143
rect 932 4137 988 4143
rect 1156 4137 1212 4143
rect 1524 4137 1548 4143
rect 1556 4137 1564 4143
rect 1668 4137 1676 4143
rect 1844 4137 2220 4143
rect 2292 4137 2540 4143
rect 2564 4137 2572 4143
rect 2580 4137 2716 4143
rect 2724 4137 2780 4143
rect 2788 4137 2860 4143
rect 2868 4137 2908 4143
rect 2916 4137 3052 4143
rect 3332 4137 3420 4143
rect 3444 4137 3612 4143
rect 3812 4137 3948 4143
rect 4116 4137 4188 4143
rect 4308 4137 4396 4143
rect 4676 4137 5164 4143
rect 5188 4137 5228 4143
rect 5428 4137 5468 4143
rect 5476 4137 5484 4143
rect 5620 4137 5644 4143
rect 5748 4137 5868 4143
rect 6020 4137 6028 4143
rect 6052 4137 6124 4143
rect 6260 4137 6316 4143
rect 6404 4137 6668 4143
rect 6964 4137 7004 4143
rect 7245 4137 7308 4143
rect 7245 4124 7251 4137
rect 20 4117 76 4123
rect 84 4117 236 4123
rect 324 4117 412 4123
rect 420 4117 476 4123
rect 916 4117 940 4123
rect 948 4117 1004 4123
rect 1044 4117 1068 4123
rect 1124 4117 1196 4123
rect 1204 4117 1244 4123
rect 1252 4117 1676 4123
rect 1748 4117 1852 4123
rect 1972 4117 2124 4123
rect 2132 4117 2252 4123
rect 2388 4117 2428 4123
rect 2436 4117 2492 4123
rect 2644 4117 2652 4123
rect 2660 4117 2764 4123
rect 3204 4117 3388 4123
rect 3396 4117 3564 4123
rect 3604 4117 3756 4123
rect 3924 4117 3964 4123
rect 4052 4117 4204 4123
rect 4212 4117 4268 4123
rect 4276 4117 4620 4123
rect 4628 4117 4684 4123
rect 4724 4117 4860 4123
rect 4900 4117 5068 4123
rect 5156 4117 5260 4123
rect 5380 4117 5804 4123
rect 6004 4117 6060 4123
rect 6164 4117 6268 4123
rect 6276 4117 6396 4123
rect 6436 4117 6476 4123
rect 6708 4117 6796 4123
rect 6868 4117 6972 4123
rect 7092 4117 7212 4123
rect 7316 4117 7372 4123
rect 276 4097 364 4103
rect 1764 4097 1932 4103
rect 1956 4097 2060 4103
rect 2228 4097 2316 4103
rect 2596 4097 2636 4103
rect 2644 4097 2684 4103
rect 2692 4097 2812 4103
rect 2820 4097 2988 4103
rect 3076 4097 3436 4103
rect 3652 4097 4252 4103
rect 4260 4097 4380 4103
rect 4388 4097 4524 4103
rect 4532 4097 4892 4103
rect 4932 4097 4940 4103
rect 5476 4097 5548 4103
rect 6132 4097 6284 4103
rect 6292 4097 6364 4103
rect 6669 4103 6675 4116
rect 6548 4097 6675 4103
rect 7092 4097 7292 4103
rect 84 4077 284 4083
rect 292 4077 332 4083
rect 1076 4077 1084 4083
rect 1332 4077 1836 4083
rect 1876 4077 1964 4083
rect 3444 4077 3532 4083
rect 3732 4077 3788 4083
rect 4084 4077 4220 4083
rect 4292 4077 4380 4083
rect 4388 4077 4716 4083
rect 4756 4077 5020 4083
rect 5037 4077 5276 4083
rect 1556 4057 2444 4063
rect 2452 4057 2476 4063
rect 3492 4057 3836 4063
rect 3844 4057 4236 4063
rect 4276 4057 4483 4063
rect 468 4037 2300 4043
rect 2308 4037 2444 4043
rect 2708 4037 3772 4043
rect 4148 4037 4156 4043
rect 4164 4037 4460 4043
rect 4477 4043 4483 4057
rect 5037 4063 5043 4077
rect 5316 4077 5347 4083
rect 4612 4057 5043 4063
rect 5053 4057 5180 4063
rect 5053 4043 5059 4057
rect 5341 4063 5347 4077
rect 5492 4077 6156 4083
rect 6196 4077 6428 4083
rect 6468 4077 6668 4083
rect 7188 4077 7212 4083
rect 7284 4077 7292 4083
rect 7316 4077 7324 4083
rect 5341 4057 6179 4063
rect 4477 4037 5059 4043
rect 5124 4037 5596 4043
rect 5732 4037 6156 4043
rect 6173 4043 6179 4057
rect 6244 4057 6300 4063
rect 6324 4057 6412 4063
rect 6420 4057 7100 4063
rect 6173 4037 6300 4043
rect 6324 4037 6924 4043
rect 7060 4037 7148 4043
rect 244 4017 1100 4023
rect 1108 4017 1180 4023
rect 3508 4017 3564 4023
rect 3620 4017 4108 4023
rect 4212 4017 4236 4023
rect 4564 4017 4636 4023
rect 4644 4017 6220 4023
rect 6260 4017 6284 4023
rect 6452 4017 7180 4023
rect 1410 4014 1470 4016
rect 1410 4006 1411 4014
rect 1420 4006 1421 4014
rect 1459 4006 1460 4014
rect 1469 4006 1470 4014
rect 1410 4004 1470 4006
rect 4418 4014 4478 4016
rect 4418 4006 4419 4014
rect 4428 4006 4429 4014
rect 4467 4006 4468 4014
rect 4477 4006 4478 4014
rect 4418 4004 4478 4006
rect 820 3997 844 4003
rect 1908 3997 2092 4003
rect 3684 3997 4332 4003
rect 4596 3997 4620 4003
rect 4756 3997 4844 4003
rect 4852 3997 4876 4003
rect 4900 3997 5068 4003
rect 5252 3997 5260 4003
rect 5604 3997 5708 4003
rect 6020 3997 6188 4003
rect 6340 3997 6412 4003
rect 484 3977 812 3983
rect 1028 3977 1068 3983
rect 1364 3977 1628 3983
rect 1700 3977 1996 3983
rect 2100 3977 2236 3983
rect 2500 3977 2620 3983
rect 2628 3977 2700 3983
rect 3124 3977 3164 3983
rect 3172 3977 3372 3983
rect 3380 3977 3884 3983
rect 3892 3977 4508 3983
rect 4516 3977 4620 3983
rect 4660 3977 4796 3983
rect 4836 3977 5052 3983
rect 5220 3977 6188 3983
rect 6244 3977 6444 3983
rect 6452 3977 6732 3983
rect 772 3957 2588 3963
rect 2596 3957 2652 3963
rect 3828 3957 3996 3963
rect 4004 3957 4316 3963
rect 4692 3957 4700 3963
rect 4708 3957 4780 3963
rect 4788 3957 4908 3963
rect 4932 3957 5004 3963
rect 5028 3957 5196 3963
rect 5204 3957 5692 3963
rect 5700 3957 6716 3963
rect 6724 3957 6796 3963
rect 6820 3957 7052 3963
rect 180 3937 460 3943
rect 484 3937 508 3943
rect 980 3937 1100 3943
rect 1588 3937 2108 3943
rect 2148 3937 2332 3943
rect 2340 3937 2684 3943
rect 3956 3937 4044 3943
rect 4068 3937 4604 3943
rect 4772 3937 4796 3943
rect 4820 3937 4892 3943
rect 4909 3943 4915 3956
rect 4909 3937 4956 3943
rect 4964 3937 5036 3943
rect 5092 3937 5164 3943
rect 5412 3937 5532 3943
rect 5652 3937 5820 3943
rect 5844 3937 5900 3943
rect 6132 3937 6220 3943
rect 6228 3937 6876 3943
rect 6884 3937 6924 3943
rect 68 3917 108 3923
rect 132 3917 412 3923
rect 468 3917 508 3923
rect 548 3917 572 3923
rect 580 3917 604 3923
rect 612 3917 684 3923
rect 1044 3917 1068 3923
rect 1236 3917 1836 3923
rect 1860 3917 2060 3923
rect 2068 3917 2348 3923
rect 2756 3917 2764 3923
rect 3732 3917 3852 3923
rect 3860 3917 4204 3923
rect 4212 3917 4780 3923
rect 4788 3917 4908 3923
rect 4916 3917 4988 3923
rect 4996 3917 5868 3923
rect 6372 3917 6467 3923
rect 164 3897 220 3903
rect 228 3897 300 3903
rect 388 3897 444 3903
rect 452 3897 492 3903
rect 500 3897 620 3903
rect 692 3897 764 3903
rect 884 3897 1132 3903
rect 1140 3897 1212 3903
rect 1220 3897 1244 3903
rect 1284 3897 1340 3903
rect 1348 3897 1404 3903
rect 1412 3897 1516 3903
rect 1524 3897 1708 3903
rect 1716 3897 1772 3903
rect 1812 3897 2012 3903
rect 2020 3897 2252 3903
rect 2356 3897 2412 3903
rect 2676 3897 2732 3903
rect 2740 3897 2780 3903
rect 2788 3897 2876 3903
rect 2900 3897 3116 3903
rect 3380 3897 3404 3903
rect 3412 3897 3484 3903
rect 3652 3897 3692 3903
rect 3732 3897 3740 3903
rect 3748 3897 3772 3903
rect 4084 3897 4252 3903
rect 4276 3897 4739 3903
rect 20 3877 140 3883
rect 180 3877 268 3883
rect 308 3877 348 3883
rect 356 3877 428 3883
rect 436 3877 444 3883
rect 452 3877 524 3883
rect 532 3877 636 3883
rect 676 3877 700 3883
rect 836 3877 892 3883
rect 1076 3877 1164 3883
rect 1188 3877 1228 3883
rect 1236 3877 1548 3883
rect 1732 3877 1820 3883
rect 1844 3877 1868 3883
rect 1876 3877 2028 3883
rect 2068 3877 2188 3883
rect 2292 3877 2316 3883
rect 2324 3877 2428 3883
rect 2516 3877 2572 3883
rect 3140 3877 3164 3883
rect 3460 3877 3548 3883
rect 3700 3877 3836 3883
rect 3844 3877 4092 3883
rect 4116 3877 4515 3883
rect 276 3857 316 3863
rect 340 3857 380 3863
rect 404 3857 460 3863
rect 500 3857 556 3863
rect 669 3863 675 3876
rect 580 3857 675 3863
rect 772 3857 1196 3863
rect 1300 3857 1308 3863
rect 1316 3857 1356 3863
rect 1396 3857 1548 3863
rect 1725 3863 1731 3876
rect 1556 3857 1731 3863
rect 1988 3857 2108 3863
rect 2628 3857 2764 3863
rect 2772 3857 2828 3863
rect 3028 3857 3580 3863
rect 3636 3857 3644 3863
rect 3652 3857 3964 3863
rect 3972 3857 4108 3863
rect 4148 3857 4492 3863
rect 4509 3863 4515 3877
rect 4733 3883 4739 3897
rect 4820 3897 4851 3903
rect 4733 3877 4812 3883
rect 4845 3883 4851 3897
rect 4868 3897 4876 3903
rect 4900 3897 4924 3903
rect 4980 3897 5164 3903
rect 5181 3897 5260 3903
rect 4845 3877 4876 3883
rect 4980 3877 5116 3883
rect 5181 3883 5187 3897
rect 5332 3897 5372 3903
rect 5524 3897 5772 3903
rect 5812 3897 6012 3903
rect 6084 3897 6172 3903
rect 6212 3897 6332 3903
rect 6404 3897 6412 3903
rect 6461 3903 6467 3917
rect 6484 3917 6636 3923
rect 6932 3917 6956 3923
rect 7124 3917 7180 3923
rect 6461 3897 6524 3903
rect 6612 3897 6732 3903
rect 6740 3897 6780 3903
rect 6868 3897 7004 3903
rect 5172 3877 5187 3883
rect 5236 3877 5324 3883
rect 5588 3877 6268 3883
rect 6276 3877 6284 3883
rect 6308 3877 6396 3883
rect 7092 3877 7228 3883
rect 4509 3857 4748 3863
rect 4804 3857 4908 3863
rect 4948 3857 5036 3863
rect 5108 3857 5212 3863
rect 5220 3857 5292 3863
rect 5380 3857 5628 3863
rect 5636 3857 5692 3863
rect 5876 3857 6076 3863
rect 6164 3857 6236 3863
rect 6244 3857 6428 3863
rect 6772 3857 6860 3863
rect 500 3837 684 3843
rect 708 3837 1580 3843
rect 1981 3843 1987 3856
rect 1620 3837 1987 3843
rect 2228 3837 2252 3843
rect 2260 3837 2348 3843
rect 2644 3837 2700 3843
rect 3956 3837 3964 3843
rect 4212 3837 5100 3843
rect 5108 3837 5388 3843
rect 5396 3837 5468 3843
rect 5485 3837 6003 3843
rect 916 3817 1196 3823
rect 1204 3817 2140 3823
rect 3812 3817 4268 3823
rect 4308 3817 4332 3823
rect 4340 3817 4428 3823
rect 4436 3817 4732 3823
rect 4756 3817 4803 3823
rect 2914 3814 2974 3816
rect 2914 3806 2915 3814
rect 2924 3806 2925 3814
rect 2963 3806 2964 3814
rect 2973 3806 2974 3814
rect 2914 3804 2974 3806
rect 628 3797 652 3803
rect 1252 3797 1308 3803
rect 1812 3797 1852 3803
rect 1860 3797 2300 3803
rect 2436 3797 2460 3803
rect 3620 3797 3660 3803
rect 4100 3797 4252 3803
rect 4356 3797 4364 3803
rect 4564 3797 4780 3803
rect 4797 3803 4803 3817
rect 4852 3817 4908 3823
rect 5485 3823 5491 3837
rect 4948 3817 5491 3823
rect 5540 3817 5820 3823
rect 5997 3823 6003 3837
rect 6420 3837 6476 3843
rect 6516 3837 6652 3843
rect 6788 3837 7164 3843
rect 7172 3837 7244 3843
rect 5997 3817 6092 3823
rect 6180 3817 6652 3823
rect 6660 3817 6700 3823
rect 6916 3817 7068 3823
rect 5922 3814 5982 3816
rect 5922 3806 5923 3814
rect 5932 3806 5933 3814
rect 5971 3806 5972 3814
rect 5981 3806 5982 3814
rect 5922 3804 5982 3806
rect 4797 3797 5100 3803
rect 5172 3797 5228 3803
rect 5332 3797 5628 3803
rect 5997 3797 6156 3803
rect 196 3777 204 3783
rect 372 3777 620 3783
rect 676 3777 684 3783
rect 980 3777 1068 3783
rect 1300 3777 1484 3783
rect 1940 3777 2204 3783
rect 3156 3777 3260 3783
rect 3268 3777 3404 3783
rect 3412 3777 3500 3783
rect 3556 3777 3692 3783
rect 3732 3777 3740 3783
rect 3748 3777 3836 3783
rect 4084 3777 4252 3783
rect 4276 3777 4364 3783
rect 4372 3777 5075 3783
rect 68 3757 124 3763
rect 196 3757 220 3763
rect 308 3757 364 3763
rect 372 3757 396 3763
rect 628 3757 684 3763
rect 724 3757 748 3763
rect 868 3757 876 3763
rect 941 3763 947 3776
rect 5069 3764 5075 3777
rect 5124 3777 5260 3783
rect 5348 3777 5404 3783
rect 5412 3777 5532 3783
rect 5812 3777 5868 3783
rect 5997 3783 6003 3797
rect 6180 3797 6588 3803
rect 6772 3797 6972 3803
rect 5892 3777 6003 3783
rect 6116 3777 6307 3783
rect 6301 3764 6307 3777
rect 6548 3777 6716 3783
rect 6884 3777 6956 3783
rect 7028 3777 7132 3783
rect 941 3757 972 3763
rect 1044 3757 1196 3763
rect 1364 3757 1404 3763
rect 1604 3757 1660 3763
rect 1748 3757 1836 3763
rect 2180 3757 2220 3763
rect 2308 3757 2316 3763
rect 2820 3757 2844 3763
rect 3540 3757 3660 3763
rect 3828 3757 4028 3763
rect 4180 3757 4284 3763
rect 4548 3757 4668 3763
rect 4724 3757 4828 3763
rect 4836 3757 4940 3763
rect 5076 3757 5260 3763
rect 5268 3757 5756 3763
rect 5764 3757 6268 3763
rect 6308 3757 6348 3763
rect 6372 3757 6460 3763
rect 6532 3757 6572 3763
rect 6580 3757 6876 3763
rect 7044 3757 7212 3763
rect 388 3737 460 3743
rect 596 3737 604 3743
rect 612 3737 668 3743
rect 820 3737 1052 3743
rect 1060 3737 1196 3743
rect 1396 3737 1532 3743
rect 1620 3737 1660 3743
rect 1956 3737 1996 3743
rect 2004 3737 2044 3743
rect 2404 3737 2540 3743
rect 2548 3737 2604 3743
rect 2628 3737 2812 3743
rect 2820 3737 2892 3743
rect 3284 3737 3452 3743
rect 3460 3737 3548 3743
rect 3636 3737 3708 3743
rect 4036 3737 4076 3743
rect 4116 3737 4188 3743
rect 4196 3737 4284 3743
rect 4324 3737 4844 3743
rect 5060 3737 5132 3743
rect 5236 3737 5452 3743
rect 5460 3737 5676 3743
rect 5812 3737 6300 3743
rect 6388 3737 6412 3743
rect 6820 3737 6876 3743
rect 6884 3737 7084 3743
rect 7396 3737 7443 3743
rect 20 3717 108 3723
rect 292 3717 348 3723
rect 356 3717 428 3723
rect 660 3717 828 3723
rect 884 3717 908 3723
rect 1444 3717 1548 3723
rect 1716 3717 1740 3723
rect 1796 3717 1820 3723
rect 1844 3717 1916 3723
rect 1924 3717 1964 3723
rect 2164 3717 2300 3723
rect 2596 3717 2716 3723
rect 2788 3717 2844 3723
rect 2900 3717 3020 3723
rect 3188 3717 3228 3723
rect 3236 3717 3420 3723
rect 3476 3717 3580 3723
rect 4036 3717 4124 3723
rect 4244 3717 4412 3723
rect 4420 3717 4604 3723
rect 4660 3717 4700 3723
rect 4756 3717 4940 3723
rect 5108 3717 5308 3723
rect 5524 3717 5532 3723
rect 5620 3717 5660 3723
rect 5684 3717 5836 3723
rect 6020 3717 6060 3723
rect 6100 3717 6140 3723
rect 6148 3717 6236 3723
rect 6244 3717 6284 3723
rect 6436 3717 6476 3723
rect 6484 3717 6540 3723
rect 6852 3717 6924 3723
rect 6932 3717 7164 3723
rect 148 3697 188 3703
rect 228 3697 316 3703
rect 372 3697 764 3703
rect 772 3697 1004 3703
rect 1012 3697 1571 3703
rect 948 3677 972 3683
rect 1565 3683 1571 3697
rect 1588 3697 1612 3703
rect 2548 3697 2844 3703
rect 3044 3697 3180 3703
rect 3764 3697 3804 3703
rect 3940 3697 4044 3703
rect 4116 3697 4716 3703
rect 4772 3697 4812 3703
rect 4893 3697 5292 3703
rect 1565 3677 2892 3683
rect 3508 3677 3564 3683
rect 3572 3677 3708 3683
rect 3812 3677 3948 3683
rect 3988 3677 4044 3683
rect 4292 3677 4540 3683
rect 4644 3677 4668 3683
rect 4893 3683 4899 3697
rect 5332 3697 5484 3703
rect 5732 3697 5884 3703
rect 5892 3697 5900 3703
rect 6036 3697 6508 3703
rect 6948 3697 7068 3703
rect 7076 3697 7148 3703
rect 4756 3677 4899 3683
rect 4916 3677 4972 3683
rect 5108 3677 5132 3683
rect 5172 3677 5372 3683
rect 5492 3677 5564 3683
rect 5572 3677 5916 3683
rect 6004 3677 6051 3683
rect 596 3657 652 3663
rect 2388 3657 2412 3663
rect 2420 3657 2524 3663
rect 2756 3657 3683 3663
rect 1332 3637 2636 3643
rect 3677 3643 3683 3657
rect 3796 3657 4076 3663
rect 4084 3657 5612 3663
rect 5652 3657 6028 3663
rect 6045 3663 6051 3677
rect 6132 3677 6220 3683
rect 6324 3677 6428 3683
rect 6468 3677 6620 3683
rect 6628 3677 7036 3683
rect 7060 3677 7132 3683
rect 6045 3657 6332 3663
rect 6468 3657 6492 3663
rect 6692 3657 6780 3663
rect 6788 3657 7084 3663
rect 7124 3657 7148 3663
rect 3677 3637 4364 3643
rect 4388 3637 4700 3643
rect 4724 3637 5548 3643
rect 5556 3637 6252 3643
rect 6260 3637 6636 3643
rect 6644 3637 6860 3643
rect 7012 3637 7148 3643
rect 244 3617 380 3623
rect 3572 3617 3612 3623
rect 3700 3617 3820 3623
rect 3828 3617 4140 3623
rect 4532 3617 4620 3623
rect 4676 3617 4844 3623
rect 4868 3617 4924 3623
rect 4996 3617 5116 3623
rect 5172 3617 5228 3623
rect 5300 3617 5548 3623
rect 5700 3617 5724 3623
rect 5828 3617 6044 3623
rect 6068 3617 6156 3623
rect 6292 3617 6556 3623
rect 6756 3617 7116 3623
rect 1410 3614 1470 3616
rect 1410 3606 1411 3614
rect 1420 3606 1421 3614
rect 1459 3606 1460 3614
rect 1469 3606 1470 3614
rect 1410 3604 1470 3606
rect 4418 3614 4478 3616
rect 4418 3606 4419 3614
rect 4428 3606 4429 3614
rect 4467 3606 4468 3614
rect 4477 3606 4478 3614
rect 4418 3604 4478 3606
rect 180 3597 316 3603
rect 900 3597 1036 3603
rect 1284 3597 1388 3603
rect 1572 3597 1852 3603
rect 1908 3597 1980 3603
rect 2308 3597 3260 3603
rect 3284 3597 3868 3603
rect 3876 3597 3916 3603
rect 3972 3597 4012 3603
rect 4020 3597 4259 3603
rect 308 3577 412 3583
rect 852 3577 972 3583
rect 980 3577 1068 3583
rect 1076 3577 2252 3583
rect 2644 3577 2668 3583
rect 2676 3577 2796 3583
rect 2804 3577 3020 3583
rect 3300 3577 3324 3583
rect 3332 3577 3340 3583
rect 3348 3577 3372 3583
rect 4253 3583 4259 3597
rect 4500 3597 4652 3603
rect 4660 3597 4684 3603
rect 4708 3597 4748 3603
rect 4788 3597 4828 3603
rect 5172 3597 5228 3603
rect 5252 3597 5356 3603
rect 5373 3597 6732 3603
rect 5373 3583 5379 3597
rect 6868 3597 6892 3603
rect 3380 3577 4243 3583
rect 4253 3577 5379 3583
rect 4237 3564 4243 3577
rect 5444 3577 5484 3583
rect 5508 3577 5580 3583
rect 5668 3577 5676 3583
rect 5764 3577 5852 3583
rect 5876 3577 6172 3583
rect 6228 3577 6236 3583
rect 6964 3577 7276 3583
rect 244 3557 1372 3563
rect 1380 3557 1628 3563
rect 1636 3557 1676 3563
rect 1956 3557 2012 3563
rect 2260 3557 2476 3563
rect 2580 3557 2700 3563
rect 3556 3557 3596 3563
rect 3716 3557 3916 3563
rect 3924 3557 3996 3563
rect 4004 3557 4092 3563
rect 4244 3557 5276 3563
rect 5284 3557 5772 3563
rect 6740 3557 6796 3563
rect 68 3537 268 3543
rect 276 3537 508 3543
rect 564 3537 1740 3543
rect 1764 3537 1868 3543
rect 2020 3537 2044 3543
rect 2068 3537 2172 3543
rect 2180 3537 2284 3543
rect 2292 3537 2460 3543
rect 3476 3537 3612 3543
rect 3668 3537 3692 3543
rect 3780 3537 4028 3543
rect 4404 3537 4556 3543
rect 4628 3537 4780 3543
rect 4884 3537 4924 3543
rect 4948 3537 5340 3543
rect 5364 3537 5388 3543
rect 5396 3537 5468 3543
rect 5604 3537 5820 3543
rect 5844 3537 6092 3543
rect 6308 3537 6476 3543
rect 6580 3537 6604 3543
rect 6756 3537 6924 3543
rect 7220 3537 7308 3543
rect 116 3517 156 3523
rect 612 3517 636 3523
rect 644 3517 716 3523
rect 724 3517 892 3523
rect 900 3517 1203 3523
rect 1197 3504 1203 3517
rect 1268 3517 1404 3523
rect 1428 3517 1596 3523
rect 1940 3517 2332 3523
rect 2356 3517 2636 3523
rect 3444 3517 3532 3523
rect 3604 3517 3644 3523
rect 3652 3517 3724 3523
rect 4116 3517 4124 3523
rect 4516 3517 4588 3523
rect 4660 3517 4844 3523
rect 4916 3517 5260 3523
rect 5764 3517 5772 3523
rect 5796 3517 5804 3523
rect 5860 3517 5900 3523
rect 5924 3517 6332 3523
rect 6340 3517 6396 3523
rect 6404 3517 6524 3523
rect 6548 3517 6652 3523
rect 6676 3517 6828 3523
rect 6836 3517 7388 3523
rect 84 3497 236 3503
rect 301 3497 332 3503
rect 301 3483 307 3497
rect 340 3497 396 3503
rect 452 3497 668 3503
rect 884 3497 988 3503
rect 1092 3497 1148 3503
rect 1204 3497 1516 3503
rect 1652 3497 1740 3503
rect 1892 3497 1916 3503
rect 2388 3497 2412 3503
rect 3188 3497 3340 3503
rect 3460 3497 3484 3503
rect 3684 3497 3692 3503
rect 3860 3497 3948 3503
rect 3988 3497 5036 3503
rect 5076 3497 5564 3503
rect 5636 3497 5644 3503
rect 5764 3497 6012 3503
rect 6228 3497 6380 3503
rect 6484 3497 6604 3503
rect 7028 3497 7036 3503
rect 7268 3497 7276 3503
rect 68 3477 307 3483
rect 324 3477 428 3483
rect 484 3477 492 3483
rect 756 3477 828 3483
rect 884 3477 1164 3483
rect 1172 3477 1516 3483
rect 1684 3477 1804 3483
rect 2004 3477 2092 3483
rect 2100 3477 2140 3483
rect 2180 3477 2220 3483
rect 2244 3477 2300 3483
rect 2516 3477 2668 3483
rect 2676 3477 2700 3483
rect 3581 3483 3587 3496
rect 3492 3477 3900 3483
rect 3908 3477 4108 3483
rect 4116 3477 4300 3483
rect 4564 3477 4588 3483
rect 4644 3477 4668 3483
rect 4692 3477 4732 3483
rect 4820 3477 4860 3483
rect 4964 3477 5004 3483
rect 5012 3477 5388 3483
rect 5396 3477 5452 3483
rect 5476 3477 5580 3483
rect 5636 3477 5900 3483
rect 6356 3477 6428 3483
rect 6452 3477 6476 3483
rect 6596 3477 6604 3483
rect 6612 3477 6684 3483
rect 6900 3477 7004 3483
rect 7252 3477 7308 3483
rect 7316 3477 7356 3483
rect 116 3457 140 3463
rect 420 3457 476 3463
rect 724 3457 780 3463
rect 804 3457 956 3463
rect 964 3457 1052 3463
rect 1204 3457 1228 3463
rect 1268 3457 1308 3463
rect 1652 3457 1900 3463
rect 1908 3457 1964 3463
rect 1972 3457 2012 3463
rect 2148 3457 2268 3463
rect 2276 3457 2316 3463
rect 2324 3457 2508 3463
rect 3524 3457 3612 3463
rect 3636 3457 3676 3463
rect 3700 3457 3756 3463
rect 3796 3457 3884 3463
rect 3956 3457 4252 3463
rect 4372 3457 4524 3463
rect 4628 3457 5004 3463
rect 5012 3457 5212 3463
rect 5220 3457 5420 3463
rect 5428 3457 5692 3463
rect 5700 3457 5724 3463
rect 5748 3457 5804 3463
rect 5821 3457 5932 3463
rect 548 3437 1500 3443
rect 1508 3437 1644 3443
rect 1796 3437 1996 3443
rect 2260 3437 2412 3443
rect 2740 3437 2876 3443
rect 3188 3437 3308 3443
rect 3316 3437 3820 3443
rect 3876 3437 4124 3443
rect 4532 3437 4812 3443
rect 4836 3437 4924 3443
rect 4948 3437 5020 3443
rect 5044 3437 5068 3443
rect 5108 3437 5219 3443
rect 436 3417 556 3423
rect 596 3417 748 3423
rect 788 3417 844 3423
rect 852 3417 1020 3423
rect 1028 3417 1084 3423
rect 1092 3417 1292 3423
rect 1300 3417 1612 3423
rect 1700 3417 2028 3423
rect 2036 3417 2780 3423
rect 3300 3417 3404 3423
rect 3700 3417 3916 3423
rect 3924 3417 4012 3423
rect 4525 3423 4531 3436
rect 5213 3423 5219 3437
rect 5332 3437 5340 3443
rect 5412 3437 5452 3443
rect 5476 3437 5596 3443
rect 5716 3437 5756 3443
rect 5821 3443 5827 3457
rect 6052 3457 6140 3463
rect 6148 3457 6204 3463
rect 6404 3457 6540 3463
rect 6564 3457 6588 3463
rect 6724 3457 6748 3463
rect 6756 3457 7260 3463
rect 5780 3437 5827 3443
rect 5844 3437 6563 3443
rect 4036 3417 4531 3423
rect 4541 3417 5203 3423
rect 5213 3417 5660 3423
rect 2914 3414 2974 3416
rect 2914 3406 2915 3414
rect 2924 3406 2925 3414
rect 2963 3406 2964 3414
rect 2973 3406 2974 3414
rect 2914 3404 2974 3406
rect 20 3397 28 3403
rect 36 3397 44 3403
rect 100 3397 595 3403
rect 100 3377 124 3383
rect 260 3377 316 3383
rect 324 3377 412 3383
rect 420 3377 444 3383
rect 452 3377 476 3383
rect 589 3383 595 3397
rect 612 3397 700 3403
rect 1620 3397 1708 3403
rect 2004 3397 2588 3403
rect 3236 3397 3724 3403
rect 3956 3397 3980 3403
rect 4276 3397 4284 3403
rect 4541 3403 4547 3417
rect 4356 3397 4547 3403
rect 4564 3397 4748 3403
rect 4804 3397 5100 3403
rect 5172 3397 5180 3403
rect 5197 3403 5203 3417
rect 5748 3417 5836 3423
rect 6004 3417 6140 3423
rect 6516 3417 6540 3423
rect 6557 3423 6563 3437
rect 6628 3437 7212 3443
rect 6557 3417 6796 3423
rect 6980 3417 7004 3423
rect 5922 3414 5982 3416
rect 5922 3406 5923 3414
rect 5932 3406 5933 3414
rect 5971 3406 5972 3414
rect 5981 3406 5982 3414
rect 5922 3404 5982 3406
rect 5197 3397 5260 3403
rect 5284 3397 5772 3403
rect 5796 3397 5852 3403
rect 6036 3397 6076 3403
rect 6212 3397 6316 3403
rect 6356 3397 6988 3403
rect 7140 3397 7196 3403
rect 589 3377 684 3383
rect 916 3377 1020 3383
rect 1412 3377 1532 3383
rect 1540 3377 1836 3383
rect 1844 3377 1964 3383
rect 2260 3377 2396 3383
rect 2404 3377 2620 3383
rect 2916 3377 3148 3383
rect 3556 3377 3660 3383
rect 3860 3377 3948 3383
rect 3956 3377 4188 3383
rect 4372 3377 4524 3383
rect 4548 3377 4700 3383
rect 4708 3377 4876 3383
rect 4916 3377 4940 3383
rect 4980 3377 5036 3383
rect 5124 3377 5324 3383
rect 5364 3377 6188 3383
rect 6308 3377 6380 3383
rect 6388 3377 6716 3383
rect 6724 3377 6796 3383
rect 7188 3377 7212 3383
rect 20 3357 204 3363
rect 660 3357 972 3363
rect 1428 3357 1548 3363
rect 1588 3357 1788 3363
rect 1876 3357 1980 3363
rect 1988 3357 2211 3363
rect 84 3337 140 3343
rect 148 3337 268 3343
rect 820 3337 860 3343
rect 1076 3337 1116 3343
rect 1700 3337 1932 3343
rect 1972 3337 1996 3343
rect 2205 3343 2211 3357
rect 2484 3357 2604 3363
rect 3092 3357 3452 3363
rect 3508 3357 3612 3363
rect 3908 3357 3980 3363
rect 4388 3357 4492 3363
rect 4516 3357 4588 3363
rect 4660 3357 4732 3363
rect 4740 3357 4748 3363
rect 4756 3357 4812 3363
rect 4829 3357 5084 3363
rect 2205 3337 2572 3343
rect 2692 3337 2732 3343
rect 2948 3337 2988 3343
rect 3604 3337 3644 3343
rect 3700 3337 3964 3343
rect 3972 3337 4060 3343
rect 4148 3337 4300 3343
rect 4333 3337 4428 3343
rect 4333 3324 4339 3337
rect 4452 3337 4739 3343
rect 116 3317 156 3323
rect 164 3317 236 3323
rect 676 3317 860 3323
rect 868 3317 876 3323
rect 1364 3317 1564 3323
rect 1581 3317 1724 3323
rect 212 3297 300 3303
rect 308 3297 444 3303
rect 468 3297 524 3303
rect 1268 3297 1324 3303
rect 1581 3303 1587 3317
rect 1732 3317 1804 3323
rect 1828 3317 1868 3323
rect 2052 3317 2076 3323
rect 2228 3317 2284 3323
rect 2292 3317 2380 3323
rect 2468 3317 2524 3323
rect 3124 3317 3164 3323
rect 3588 3317 3788 3323
rect 3805 3317 4028 3323
rect 1332 3297 1587 3303
rect 1828 3297 2044 3303
rect 3805 3303 3811 3317
rect 4052 3317 4156 3323
rect 4260 3317 4332 3323
rect 4372 3317 4716 3323
rect 4733 3323 4739 3337
rect 4756 3337 4780 3343
rect 4829 3343 4835 3357
rect 5108 3357 5852 3363
rect 5860 3357 6796 3363
rect 6804 3357 7100 3363
rect 4797 3337 4835 3343
rect 4733 3317 4780 3323
rect 3028 3297 3811 3303
rect 4004 3297 4444 3303
rect 4596 3297 4652 3303
rect 4797 3303 4803 3337
rect 4932 3337 5068 3343
rect 5124 3337 5196 3343
rect 5428 3337 5516 3343
rect 5684 3337 5708 3343
rect 5796 3337 5884 3343
rect 5972 3337 6028 3343
rect 6132 3337 6172 3343
rect 6205 3337 6396 3343
rect 4820 3317 4828 3323
rect 4836 3317 4892 3323
rect 4900 3317 4924 3323
rect 5028 3317 5068 3323
rect 5076 3317 5164 3323
rect 5396 3317 5644 3323
rect 5668 3317 5772 3323
rect 5828 3317 5836 3323
rect 6205 3323 6211 3337
rect 6404 3337 6492 3343
rect 6564 3337 6876 3343
rect 5892 3317 6211 3323
rect 6228 3317 6236 3323
rect 6708 3317 6780 3323
rect 6884 3317 7052 3323
rect 7060 3317 7244 3323
rect 4772 3297 4803 3303
rect 4900 3297 4940 3303
rect 5044 3297 5404 3303
rect 5508 3297 5532 3303
rect 5588 3297 5612 3303
rect 5620 3297 6044 3303
rect 6052 3297 6140 3303
rect 6148 3297 6156 3303
rect 6164 3297 6236 3303
rect 6324 3297 6604 3303
rect 6621 3297 6700 3303
rect 468 3277 540 3283
rect 548 3277 1276 3283
rect 1284 3277 1340 3283
rect 1572 3277 1660 3283
rect 1860 3277 1868 3283
rect 3460 3277 3516 3283
rect 3636 3277 3804 3283
rect 3821 3277 4012 3283
rect 804 3257 876 3263
rect 884 3257 1116 3263
rect 1124 3257 1308 3263
rect 1316 3257 1852 3263
rect 1972 3257 1996 3263
rect 2628 3257 2684 3263
rect 3821 3263 3827 3277
rect 4036 3277 4716 3283
rect 4765 3277 4796 3283
rect 3412 3257 3827 3263
rect 3972 3257 4364 3263
rect 4420 3257 4524 3263
rect 4644 3257 4700 3263
rect 4765 3263 4771 3277
rect 4900 3277 4956 3283
rect 4980 3277 5036 3283
rect 5092 3277 5212 3283
rect 5444 3277 5580 3283
rect 5620 3277 5820 3283
rect 6004 3277 6028 3283
rect 6621 3283 6627 3297
rect 6772 3297 6908 3303
rect 7156 3297 7180 3303
rect 7268 3297 7292 3303
rect 6084 3277 6627 3283
rect 4724 3257 4771 3263
rect 4788 3257 5356 3263
rect 5428 3257 5468 3263
rect 5508 3257 5868 3263
rect 6292 3257 6476 3263
rect 6484 3257 7068 3263
rect 1524 3237 2188 3243
rect 2196 3237 2364 3243
rect 2516 3237 5740 3243
rect 5844 3237 6508 3243
rect 6708 3237 6748 3243
rect 36 3217 76 3223
rect 516 3217 860 3223
rect 1748 3217 1788 3223
rect 1796 3217 1900 3223
rect 3060 3217 3500 3223
rect 3572 3217 3772 3223
rect 3780 3217 4060 3223
rect 4068 3217 4396 3223
rect 4996 3217 5228 3223
rect 5268 3217 5996 3223
rect 6180 3217 6620 3223
rect 1410 3214 1470 3216
rect 1410 3206 1411 3214
rect 1420 3206 1421 3214
rect 1459 3206 1460 3214
rect 1469 3206 1470 3214
rect 1410 3204 1470 3206
rect 4418 3214 4478 3216
rect 4418 3206 4419 3214
rect 4428 3206 4429 3214
rect 4467 3206 4468 3214
rect 4477 3206 4478 3214
rect 4418 3204 4478 3206
rect 500 3197 508 3203
rect 1524 3197 1548 3203
rect 1556 3197 2156 3203
rect 2580 3197 2796 3203
rect 3444 3197 3468 3203
rect 3492 3197 3564 3203
rect 3652 3197 3852 3203
rect 4276 3197 4332 3203
rect 4500 3197 4956 3203
rect 4964 3197 5324 3203
rect 5332 3197 5468 3203
rect 5588 3197 5628 3203
rect 5684 3197 6156 3203
rect 6196 3197 7052 3203
rect 1204 3177 1500 3183
rect 1732 3177 1740 3183
rect 2132 3177 2300 3183
rect 2308 3177 2412 3183
rect 2420 3177 2588 3183
rect 2596 3177 2716 3183
rect 2772 3177 3148 3183
rect 3172 3177 3868 3183
rect 3956 3177 4156 3183
rect 4269 3183 4275 3196
rect 4164 3177 4275 3183
rect 4372 3177 4668 3183
rect 4868 3177 5068 3183
rect 5076 3177 5164 3183
rect 5620 3177 5820 3183
rect 5988 3177 6348 3183
rect 6356 3177 6396 3183
rect 6676 3177 7196 3183
rect 372 3157 556 3163
rect 628 3157 764 3163
rect 788 3157 908 3163
rect 1316 3157 1324 3163
rect 2164 3157 2332 3163
rect 3444 3157 3516 3163
rect 3540 3157 3660 3163
rect 3684 3157 3692 3163
rect 3700 3157 3964 3163
rect 3988 3157 4060 3163
rect 4116 3157 4604 3163
rect 4612 3157 4716 3163
rect 5005 3157 5827 3163
rect 548 3137 668 3143
rect 740 3137 748 3143
rect 820 3137 844 3143
rect 948 3137 1148 3143
rect 1172 3137 1212 3143
rect 1268 3137 1292 3143
rect 1332 3137 1356 3143
rect 1812 3137 2060 3143
rect 2100 3137 2156 3143
rect 2628 3137 2764 3143
rect 5005 3143 5011 3157
rect 2788 3137 5011 3143
rect 5028 3137 5036 3143
rect 5044 3137 5052 3143
rect 5156 3137 5260 3143
rect 5268 3137 5500 3143
rect 5524 3137 5724 3143
rect 5821 3143 5827 3157
rect 5844 3157 6108 3163
rect 6116 3157 6668 3163
rect 7156 3157 7180 3163
rect 5821 3137 6252 3143
rect 6285 3137 6332 3143
rect 388 3117 444 3123
rect 628 3117 636 3123
rect 708 3117 780 3123
rect 900 3117 1052 3123
rect 1060 3117 1276 3123
rect 1284 3117 1324 3123
rect 1812 3117 1932 3123
rect 1972 3117 1980 3123
rect 1988 3117 2092 3123
rect 2388 3117 2444 3123
rect 2836 3117 2924 3123
rect 2932 3117 3180 3123
rect 3284 3117 3740 3123
rect 3860 3117 3932 3123
rect 3940 3117 4044 3123
rect 4052 3117 4076 3123
rect 4116 3117 4220 3123
rect 4260 3117 4444 3123
rect 4452 3117 4636 3123
rect 4653 3117 4716 3123
rect 20 3097 124 3103
rect 164 3097 268 3103
rect 324 3097 396 3103
rect 484 3097 524 3103
rect 532 3097 652 3103
rect 692 3097 700 3103
rect 893 3103 899 3116
rect 740 3097 899 3103
rect 1348 3097 1388 3103
rect 1524 3097 1548 3103
rect 1620 3097 1820 3103
rect 1860 3097 2380 3103
rect 2516 3097 2524 3103
rect 2612 3097 2668 3103
rect 3220 3097 3260 3103
rect 3380 3097 3692 3103
rect 3732 3097 3772 3103
rect 3780 3097 3980 3103
rect 4068 3097 4172 3103
rect 4228 3097 4316 3103
rect 4340 3097 4515 3103
rect 84 3077 108 3083
rect 116 3077 332 3083
rect 340 3077 380 3083
rect 564 3077 572 3083
rect 1156 3077 1276 3083
rect 1588 3077 1708 3083
rect 1821 3083 1827 3096
rect 1821 3077 2348 3083
rect 2628 3077 2732 3083
rect 2804 3077 2892 3083
rect 2900 3077 2972 3083
rect 2996 3077 3068 3083
rect 3188 3077 3244 3083
rect 3252 3077 3596 3083
rect 3796 3077 4492 3083
rect 4509 3083 4515 3097
rect 4653 3103 4659 3117
rect 4756 3117 5228 3123
rect 5300 3117 5500 3123
rect 5572 3117 5612 3123
rect 5620 3117 6028 3123
rect 6285 3123 6291 3137
rect 6612 3137 6748 3143
rect 6756 3137 6908 3143
rect 7076 3137 7180 3143
rect 6036 3117 6291 3123
rect 6580 3117 6620 3123
rect 6628 3117 6844 3123
rect 6852 3117 6972 3123
rect 7172 3117 7292 3123
rect 4580 3097 4659 3103
rect 4708 3097 4844 3103
rect 4861 3097 4876 3103
rect 4509 3077 4732 3083
rect 4861 3083 4867 3097
rect 4884 3097 5580 3103
rect 5700 3097 5996 3103
rect 6292 3097 6444 3103
rect 6532 3097 6636 3103
rect 6660 3097 6812 3103
rect 6820 3097 7036 3103
rect 4804 3077 4867 3083
rect 4948 3077 5132 3083
rect 5380 3077 5452 3083
rect 5524 3077 5596 3083
rect 5940 3077 6060 3083
rect 6164 3077 6588 3083
rect 6708 3077 7116 3083
rect 7124 3077 7276 3083
rect 132 3057 156 3063
rect 164 3057 172 3063
rect 180 3057 316 3063
rect 372 3057 460 3063
rect 788 3057 908 3063
rect 1492 3057 1612 3063
rect 1796 3057 1836 3063
rect 1860 3057 1980 3063
rect 2084 3057 2140 3063
rect 2660 3057 2828 3063
rect 2836 3057 3196 3063
rect 3204 3057 3276 3063
rect 3284 3057 3420 3063
rect 3492 3057 3612 3063
rect 3764 3057 3804 3063
rect 3892 3057 4588 3063
rect 4596 3057 4684 3063
rect 4724 3057 5228 3063
rect 5332 3057 5596 3063
rect 5604 3057 5788 3063
rect 5796 3057 5852 3063
rect 5860 3057 5900 3063
rect 6260 3057 6300 3063
rect 6308 3057 6556 3063
rect 6772 3057 6828 3063
rect 6900 3057 6988 3063
rect 7108 3057 7164 3063
rect 164 3037 492 3043
rect 1572 3037 1612 3043
rect 1693 3037 1724 3043
rect 1693 3023 1699 3037
rect 2116 3037 2188 3043
rect 2196 3037 2396 3043
rect 2564 3037 2812 3043
rect 3140 3037 3260 3043
rect 3396 3037 3564 3043
rect 3588 3037 3628 3043
rect 3636 3037 3676 3043
rect 3844 3037 4380 3043
rect 4388 3037 4908 3043
rect 4916 3037 4940 3043
rect 4948 3037 5116 3043
rect 5140 3037 5244 3043
rect 5252 3037 5420 3043
rect 5460 3037 5932 3043
rect 6020 3037 6060 3043
rect 6068 3037 6220 3043
rect 6228 3037 6332 3043
rect 6676 3037 6844 3043
rect 6884 3037 6892 3043
rect 6900 3037 6956 3043
rect 7060 3037 7116 3043
rect 7140 3037 7164 3043
rect 1556 3017 1699 3023
rect 2068 3017 2204 3023
rect 2388 3017 2572 3023
rect 3524 3017 3820 3023
rect 3876 3017 3948 3023
rect 4884 3017 4892 3023
rect 4909 3017 5100 3023
rect 2914 3014 2974 3016
rect 2914 3006 2915 3014
rect 2924 3006 2925 3014
rect 2963 3006 2964 3014
rect 2973 3006 2974 3014
rect 2914 3004 2974 3006
rect 804 2997 1084 3003
rect 1092 2997 1148 3003
rect 1252 2997 1596 3003
rect 1684 2997 1740 3003
rect 1748 2997 1820 3003
rect 1940 2997 1964 3003
rect 2244 2997 2300 3003
rect 3796 2997 3884 3003
rect 4052 2997 4220 3003
rect 4525 3003 4531 3016
rect 4909 3003 4915 3017
rect 5108 3017 5836 3023
rect 6004 3017 6316 3023
rect 6580 3017 6716 3023
rect 6996 3017 7244 3023
rect 5922 3014 5982 3016
rect 5922 3006 5923 3014
rect 5932 3006 5933 3014
rect 5971 3006 5972 3014
rect 5981 3006 5982 3014
rect 5922 3004 5982 3006
rect 4525 2997 4915 3003
rect 4964 2997 4972 3003
rect 5012 2997 5260 3003
rect 6020 2997 6092 3003
rect 6276 2997 6492 3003
rect 6509 2997 6908 3003
rect 6509 2984 6515 2997
rect 6948 2997 7100 3003
rect 660 2977 684 2983
rect 692 2977 812 2983
rect 820 2977 1100 2983
rect 1236 2977 1260 2983
rect 2340 2977 2572 2983
rect 2740 2977 2828 2983
rect 3460 2977 3532 2983
rect 3540 2977 4284 2983
rect 4292 2977 4764 2983
rect 4772 2977 4812 2983
rect 4884 2977 6092 2983
rect 6164 2977 6348 2983
rect 6356 2977 6380 2983
rect 6452 2977 6508 2983
rect 6596 2977 6668 2983
rect 6964 2977 7052 2983
rect 7124 2977 7148 2983
rect 1060 2957 1084 2963
rect 1108 2957 1132 2963
rect 1140 2957 1180 2963
rect 1348 2957 1388 2963
rect 1412 2957 1516 2963
rect 1780 2957 1804 2963
rect 1844 2957 1932 2963
rect 2164 2957 2220 2963
rect 2292 2957 2460 2963
rect 3572 2957 3612 2963
rect 4212 2957 4236 2963
rect 4244 2957 4252 2963
rect 4516 2957 4700 2963
rect 4740 2957 4844 2963
rect 4852 2957 5004 2963
rect 5012 2957 5068 2963
rect 5444 2957 5628 2963
rect 5780 2957 5884 2963
rect 6324 2957 6460 2963
rect 6500 2957 6508 2963
rect 6516 2957 6860 2963
rect 7124 2957 7148 2963
rect 7156 2957 7276 2963
rect 7348 2957 7388 2963
rect 7396 2957 7443 2963
rect 84 2937 140 2943
rect 148 2937 220 2943
rect 436 2937 460 2943
rect 964 2937 988 2943
rect 996 2937 1212 2943
rect 1220 2937 1244 2943
rect 1252 2937 1324 2943
rect 1332 2937 1516 2943
rect 1556 2937 1580 2943
rect 1748 2937 1836 2943
rect 1892 2937 1948 2943
rect 2036 2937 2268 2943
rect 2292 2937 2460 2943
rect 2612 2937 2652 2943
rect 2660 2937 2780 2943
rect 3188 2937 3340 2943
rect 3508 2937 3580 2943
rect 4100 2937 4188 2943
rect 4196 2937 4348 2943
rect 4356 2937 4364 2943
rect 4372 2937 4556 2943
rect 4564 2937 4828 2943
rect 5060 2937 5372 2943
rect 5572 2937 5660 2943
rect 5732 2937 5772 2943
rect 5828 2937 6220 2943
rect 6228 2937 6620 2943
rect 7044 2937 7084 2943
rect 7092 2937 7276 2943
rect 36 2917 92 2923
rect 756 2917 988 2923
rect 1044 2917 1260 2923
rect 1268 2917 1292 2923
rect 1348 2917 1356 2923
rect 1524 2917 2092 2923
rect 2164 2917 2412 2923
rect 2420 2917 2508 2923
rect 2884 2917 3276 2923
rect 3284 2917 3388 2923
rect 3396 2917 3436 2923
rect 3444 2917 3516 2923
rect 3588 2917 3644 2923
rect 3780 2917 3788 2923
rect 3796 2917 3820 2923
rect 4004 2917 4492 2923
rect 4516 2917 4620 2923
rect 4852 2917 4988 2923
rect 5172 2917 5244 2923
rect 5364 2917 5404 2923
rect 5508 2917 5628 2923
rect 5645 2917 5996 2923
rect 244 2897 348 2903
rect 381 2897 604 2903
rect 381 2884 387 2897
rect 852 2897 908 2903
rect 1332 2897 2220 2903
rect 2260 2897 2316 2903
rect 2372 2897 2444 2903
rect 2452 2897 2460 2903
rect 3220 2897 3308 2903
rect 3476 2897 3548 2903
rect 3572 2897 3612 2903
rect 3668 2897 4332 2903
rect 4356 2897 4675 2903
rect 4973 2897 4988 2903
rect 308 2877 380 2883
rect 388 2877 412 2883
rect 532 2877 556 2883
rect 708 2877 796 2883
rect 884 2877 908 2883
rect 1076 2877 1244 2883
rect 1300 2877 1564 2883
rect 1668 2877 1708 2883
rect 1732 2877 1740 2883
rect 1748 2877 1964 2883
rect 2116 2877 2172 2883
rect 2221 2883 2227 2896
rect 2221 2877 2572 2883
rect 3236 2877 3292 2883
rect 4196 2877 4236 2883
rect 4340 2877 4540 2883
rect 4644 2877 4652 2883
rect 4669 2883 4675 2897
rect 4996 2897 5036 2903
rect 5076 2897 5420 2903
rect 5645 2903 5651 2917
rect 6036 2917 6108 2923
rect 6420 2917 6492 2923
rect 6564 2917 6636 2923
rect 6644 2917 6684 2923
rect 6788 2917 7116 2923
rect 7236 2917 7308 2923
rect 5428 2897 5651 2903
rect 5668 2897 5708 2903
rect 5844 2897 5996 2903
rect 6093 2897 6268 2903
rect 4669 2877 5180 2883
rect 5220 2877 5420 2883
rect 5524 2877 5532 2883
rect 5636 2877 5740 2883
rect 6093 2883 6099 2897
rect 6292 2897 6412 2903
rect 6436 2897 6476 2903
rect 6484 2897 6556 2903
rect 6644 2897 6748 2903
rect 6772 2897 6860 2903
rect 7229 2903 7235 2916
rect 6868 2897 7235 2903
rect 7412 2897 7443 2903
rect 5748 2877 6099 2883
rect 6116 2877 6476 2883
rect 6948 2877 7212 2883
rect 228 2857 540 2863
rect 548 2857 620 2863
rect 692 2857 716 2863
rect 820 2857 924 2863
rect 1012 2857 1132 2863
rect 1492 2857 1820 2863
rect 1844 2857 1964 2863
rect 2244 2857 2268 2863
rect 2356 2857 2396 2863
rect 3716 2857 3756 2863
rect 3764 2857 4300 2863
rect 4372 2857 5036 2863
rect 5140 2857 5980 2863
rect 6132 2857 6764 2863
rect 6932 2857 7052 2863
rect 388 2837 716 2843
rect 1076 2837 1100 2843
rect 1540 2837 1580 2843
rect 1636 2837 1772 2843
rect 1908 2837 1996 2843
rect 452 2817 940 2823
rect 948 2817 1212 2823
rect 1316 2817 1388 2823
rect 2285 2823 2291 2856
rect 3028 2837 6284 2843
rect 1508 2817 2291 2823
rect 2836 2817 3052 2823
rect 4244 2817 4268 2823
rect 4500 2817 5004 2823
rect 5060 2817 5132 2823
rect 5172 2817 5196 2823
rect 5284 2817 5292 2823
rect 5364 2817 6012 2823
rect 6244 2817 6300 2823
rect 6308 2817 7164 2823
rect 1410 2814 1470 2816
rect 1410 2806 1411 2814
rect 1420 2806 1421 2814
rect 1459 2806 1460 2814
rect 1469 2806 1470 2814
rect 1410 2804 1470 2806
rect 4418 2814 4478 2816
rect 4418 2806 4419 2814
rect 4428 2806 4429 2814
rect 4467 2806 4468 2814
rect 4477 2806 4478 2814
rect 4418 2804 4478 2806
rect 324 2797 588 2803
rect 596 2797 668 2803
rect 1028 2797 1068 2803
rect 1156 2797 1196 2803
rect 1204 2797 1324 2803
rect 1700 2797 1980 2803
rect 2292 2797 3564 2803
rect 4013 2797 4108 2803
rect 884 2777 1516 2783
rect 1572 2777 1795 2783
rect 260 2757 300 2763
rect 516 2757 668 2763
rect 916 2757 956 2763
rect 1012 2757 1036 2763
rect 1284 2757 1324 2763
rect 1620 2757 1660 2763
rect 1789 2763 1795 2777
rect 4013 2783 4019 2797
rect 4516 2797 4556 2803
rect 4660 2797 4908 2803
rect 4916 2797 5036 2803
rect 5124 2797 5148 2803
rect 5156 2797 5580 2803
rect 5588 2797 5788 2803
rect 6068 2797 6636 2803
rect 6644 2797 6972 2803
rect 6980 2797 7212 2803
rect 7220 2797 7324 2803
rect 1812 2777 4019 2783
rect 4036 2777 4092 2783
rect 4100 2777 4972 2783
rect 5012 2777 5836 2783
rect 6468 2777 6508 2783
rect 6516 2777 6828 2783
rect 1789 2757 2060 2763
rect 2068 2757 2380 2763
rect 2388 2757 2444 2763
rect 2596 2757 6508 2763
rect 6660 2757 6684 2763
rect 276 2737 300 2743
rect 404 2737 460 2743
rect 468 2737 508 2743
rect 532 2737 844 2743
rect 852 2737 1116 2743
rect 1156 2737 1372 2743
rect 1380 2737 1548 2743
rect 1556 2737 1612 2743
rect 1620 2737 1676 2743
rect 1908 2737 1932 2743
rect 2084 2737 2108 2743
rect 2116 2737 2172 2743
rect 2180 2737 2236 2743
rect 2820 2737 2828 2743
rect 2836 2737 2860 2743
rect 3316 2737 3356 2743
rect 3492 2737 3916 2743
rect 4148 2737 4316 2743
rect 4548 2737 4652 2743
rect 4868 2737 4940 2743
rect 5028 2737 5068 2743
rect 5092 2737 5100 2743
rect 5284 2737 5388 2743
rect 5540 2737 5772 2743
rect 5812 2737 7100 2743
rect 404 2717 572 2723
rect 628 2717 652 2723
rect 660 2717 828 2723
rect 964 2717 1036 2723
rect 1348 2717 1788 2723
rect 1828 2717 2019 2723
rect 2013 2704 2019 2717
rect 2212 2717 2348 2723
rect 2516 2717 2540 2723
rect 3124 2717 3164 2723
rect 3300 2717 3340 2723
rect 3348 2717 3420 2723
rect 3428 2717 3468 2723
rect 3636 2717 3724 2723
rect 3876 2717 4044 2723
rect 4132 2717 4156 2723
rect 4164 2717 4220 2723
rect 4260 2717 4515 2723
rect 68 2697 108 2703
rect 164 2697 172 2703
rect 340 2697 364 2703
rect 388 2697 460 2703
rect 468 2697 524 2703
rect 708 2697 732 2703
rect 804 2697 860 2703
rect 1012 2697 1036 2703
rect 1220 2697 1260 2703
rect 1380 2697 1484 2703
rect 1492 2697 1564 2703
rect 1572 2697 1628 2703
rect 1636 2697 1692 2703
rect 1748 2697 1788 2703
rect 1828 2697 1884 2703
rect 1892 2697 1900 2703
rect 1956 2697 1980 2703
rect 2020 2697 2124 2703
rect 2132 2697 2188 2703
rect 2196 2697 2252 2703
rect 2372 2697 2476 2703
rect 2532 2697 2556 2703
rect 2612 2697 3132 2703
rect 3396 2697 3468 2703
rect 3476 2697 3580 2703
rect 4004 2697 4412 2703
rect 4509 2703 4515 2717
rect 4532 2717 4675 2723
rect 4669 2704 4675 2717
rect 4788 2717 4844 2723
rect 4884 2717 4908 2723
rect 5044 2717 5084 2723
rect 5156 2717 5212 2723
rect 5437 2717 5468 2723
rect 4509 2697 4588 2703
rect 4612 2697 4636 2703
rect 4676 2697 4748 2703
rect 4804 2697 4940 2703
rect 4980 2697 5036 2703
rect 5437 2703 5443 2717
rect 5716 2717 5788 2723
rect 6340 2717 6460 2723
rect 6612 2717 6796 2723
rect 5076 2697 5443 2703
rect 5460 2697 5548 2703
rect 5796 2697 6668 2703
rect 6708 2697 6780 2703
rect 6868 2697 6876 2703
rect 356 2677 380 2683
rect 1124 2677 1724 2683
rect 1805 2677 1852 2683
rect 84 2657 108 2663
rect 596 2657 764 2663
rect 861 2657 972 2663
rect 861 2643 867 2657
rect 1524 2657 1580 2663
rect 1805 2663 1811 2677
rect 1876 2677 1916 2683
rect 1940 2677 2044 2683
rect 2724 2677 2732 2683
rect 2836 2677 2956 2683
rect 2996 2677 3020 2683
rect 3268 2677 3340 2683
rect 3389 2683 3395 2696
rect 3348 2677 3395 2683
rect 3732 2677 3772 2683
rect 3780 2677 3948 2683
rect 4180 2677 4268 2683
rect 4308 2677 5020 2683
rect 5092 2677 5164 2683
rect 5316 2677 5356 2683
rect 5412 2677 5516 2683
rect 5748 2677 5852 2683
rect 6276 2677 6332 2683
rect 6564 2677 6588 2683
rect 6644 2677 6668 2683
rect 6964 2677 7116 2683
rect 7124 2677 7292 2683
rect 1636 2657 1811 2663
rect 1828 2657 1836 2663
rect 1956 2657 2284 2663
rect 2500 2657 2556 2663
rect 2708 2657 3164 2663
rect 4308 2657 4332 2663
rect 4356 2657 4380 2663
rect 4628 2657 4764 2663
rect 4836 2657 4860 2663
rect 4884 2657 4908 2663
rect 4932 2657 4972 2663
rect 5060 2657 5212 2663
rect 6020 2657 6092 2663
rect 6100 2657 6316 2663
rect 6548 2657 6588 2663
rect 6724 2657 6908 2663
rect 292 2637 867 2643
rect 884 2637 908 2643
rect 932 2637 1804 2643
rect 1844 2637 2412 2643
rect 2484 2637 3004 2643
rect 3060 2637 3372 2643
rect 3796 2637 4092 2643
rect 4100 2637 4236 2643
rect 4244 2637 5308 2643
rect 5620 2637 5644 2643
rect 5780 2637 5836 2643
rect 5908 2637 6252 2643
rect 6276 2637 6348 2643
rect 6452 2637 6476 2643
rect 6660 2637 6716 2643
rect 6724 2637 6988 2643
rect 6996 2637 7068 2643
rect 68 2617 156 2623
rect 164 2617 188 2623
rect 196 2617 2700 2623
rect 3540 2617 4700 2623
rect 4740 2617 5084 2623
rect 5140 2617 5164 2623
rect 5188 2617 5516 2623
rect 6212 2617 6620 2623
rect 6932 2617 7100 2623
rect 2914 2614 2974 2616
rect 2914 2606 2915 2614
rect 2924 2606 2925 2614
rect 2963 2606 2964 2614
rect 2973 2606 2974 2614
rect 2914 2604 2974 2606
rect 5922 2614 5982 2616
rect 5922 2606 5923 2614
rect 5932 2606 5933 2614
rect 5971 2606 5972 2614
rect 5981 2606 5982 2614
rect 5922 2604 5982 2606
rect 1044 2597 2476 2603
rect 2516 2597 2684 2603
rect 3789 2597 4172 2603
rect 3789 2584 3795 2597
rect 4196 2597 4268 2603
rect 4740 2597 4828 2603
rect 4852 2597 4876 2603
rect 4916 2597 4940 2603
rect 5172 2597 5196 2603
rect 5268 2597 5436 2603
rect 5460 2597 5532 2603
rect 6516 2597 6556 2603
rect 6756 2597 6796 2603
rect 6820 2597 7084 2603
rect 7092 2597 7228 2603
rect 1300 2577 1724 2583
rect 1748 2577 1996 2583
rect 2004 2577 2044 2583
rect 2292 2577 2348 2583
rect 2436 2577 2476 2583
rect 2612 2577 2668 2583
rect 2724 2577 2780 2583
rect 2836 2577 2844 2583
rect 3284 2577 3324 2583
rect 3700 2577 3788 2583
rect 4532 2577 4652 2583
rect 4724 2577 4844 2583
rect 4996 2577 5148 2583
rect 5156 2577 5244 2583
rect 5268 2577 5292 2583
rect 5364 2577 6588 2583
rect 6596 2577 7020 2583
rect 7028 2577 7116 2583
rect 7188 2577 7276 2583
rect 84 2557 220 2563
rect 660 2557 764 2563
rect 964 2557 1020 2563
rect 1140 2557 1244 2563
rect 1508 2557 1612 2563
rect 1892 2557 1964 2563
rect 2260 2557 2332 2563
rect 2420 2557 2876 2563
rect 3140 2557 3372 2563
rect 3380 2557 3692 2563
rect 3876 2557 4060 2563
rect 4292 2557 4316 2563
rect 4324 2557 4412 2563
rect 4420 2557 4556 2563
rect 4564 2557 4940 2563
rect 4948 2557 5068 2563
rect 5076 2557 5452 2563
rect 5556 2557 5740 2563
rect 6116 2557 6124 2563
rect 6212 2557 6284 2563
rect 6292 2557 6684 2563
rect 6708 2557 7036 2563
rect 52 2537 131 2543
rect 125 2524 131 2537
rect 612 2537 684 2543
rect 1780 2537 1996 2543
rect 2324 2537 2540 2543
rect 2644 2537 2652 2543
rect 2660 2537 2668 2543
rect 2692 2537 2748 2543
rect 2868 2537 2876 2543
rect 2884 2537 2972 2543
rect 2996 2537 3132 2543
rect 3316 2537 3500 2543
rect 3508 2537 3660 2543
rect 4004 2537 4204 2543
rect 4212 2537 4300 2543
rect 4580 2537 4764 2543
rect 4820 2537 4828 2543
rect 4868 2537 4892 2543
rect 4957 2537 4988 2543
rect 20 2517 76 2523
rect 132 2517 156 2523
rect 276 2517 364 2523
rect 596 2517 620 2523
rect 676 2517 924 2523
rect 932 2517 1148 2523
rect 1220 2517 1308 2523
rect 1364 2517 1468 2523
rect 1508 2517 1548 2523
rect 1748 2517 1772 2523
rect 1988 2517 2028 2523
rect 2068 2517 2124 2523
rect 2196 2517 2220 2523
rect 2372 2517 2428 2523
rect 2436 2517 2588 2523
rect 2756 2517 2876 2523
rect 3076 2517 3228 2523
rect 3588 2517 3596 2523
rect 3684 2517 3756 2523
rect 4036 2517 4076 2523
rect 4180 2517 4252 2523
rect 4276 2517 4604 2523
rect 4676 2517 4876 2523
rect 4957 2523 4963 2537
rect 5044 2537 5100 2543
rect 5172 2537 5260 2543
rect 5332 2537 5356 2543
rect 5549 2543 5555 2556
rect 5444 2537 5555 2543
rect 5860 2537 5932 2543
rect 6244 2537 6284 2543
rect 6420 2537 6524 2543
rect 6612 2537 6812 2543
rect 6868 2537 6988 2543
rect 7012 2537 7180 2543
rect 7316 2537 7340 2543
rect 4900 2517 4963 2523
rect 4980 2517 5036 2523
rect 5044 2517 5356 2523
rect 5460 2517 5500 2523
rect 5540 2517 5548 2523
rect 5684 2517 5772 2523
rect 6004 2517 6140 2523
rect 6228 2517 6412 2523
rect 6452 2517 6659 2523
rect 100 2497 284 2503
rect 564 2497 1164 2503
rect 1172 2497 1180 2503
rect 1364 2497 1548 2503
rect 1876 2497 2268 2503
rect 2324 2497 2348 2503
rect 2388 2497 2524 2503
rect 2532 2497 3036 2503
rect 3156 2497 3676 2503
rect 4228 2497 4380 2503
rect 4388 2497 4780 2503
rect 4852 2497 5036 2503
rect 5124 2497 5180 2503
rect 5268 2497 5452 2503
rect 5492 2497 5548 2503
rect 5780 2497 5884 2503
rect 5892 2497 5996 2503
rect 6004 2497 6140 2503
rect 6148 2497 6188 2503
rect 6388 2497 6460 2503
rect 6612 2497 6636 2503
rect 6653 2503 6659 2517
rect 6676 2517 7164 2523
rect 7188 2517 7244 2523
rect 7332 2517 7388 2523
rect 6653 2497 6748 2503
rect 7028 2497 7084 2503
rect 7204 2497 7228 2503
rect 7364 2497 7404 2503
rect 7412 2497 7443 2503
rect 324 2477 492 2483
rect 1236 2477 1516 2483
rect 1796 2477 1836 2483
rect 1860 2477 1948 2483
rect 2228 2477 2348 2483
rect 2852 2477 2924 2483
rect 3044 2477 3116 2483
rect 3124 2477 3244 2483
rect 3604 2477 3980 2483
rect 4084 2477 4108 2483
rect 4116 2477 4652 2483
rect 4660 2477 5068 2483
rect 5076 2477 5372 2483
rect 5556 2477 5564 2483
rect 6212 2477 6620 2483
rect 6916 2477 7132 2483
rect 260 2457 300 2463
rect 468 2457 1708 2463
rect 1732 2457 2108 2463
rect 2196 2457 2300 2463
rect 3796 2457 4492 2463
rect 4532 2457 4588 2463
rect 4596 2457 4732 2463
rect 4740 2457 4796 2463
rect 4804 2457 4908 2463
rect 4916 2457 5196 2463
rect 5204 2457 5276 2463
rect 5348 2457 5404 2463
rect 5412 2457 5468 2463
rect 5748 2457 5884 2463
rect 5892 2457 6268 2463
rect 6365 2457 6476 2463
rect 356 2437 604 2443
rect 644 2437 956 2443
rect 964 2437 1116 2443
rect 1124 2437 1212 2443
rect 1300 2437 1692 2443
rect 2052 2437 3164 2443
rect 4196 2437 4716 2443
rect 4756 2437 4780 2443
rect 4884 2437 5027 2443
rect 212 2417 492 2423
rect 1748 2417 1868 2423
rect 1876 2417 1916 2423
rect 1956 2417 2236 2423
rect 2308 2417 3052 2423
rect 3092 2417 3148 2423
rect 4148 2417 4332 2423
rect 4564 2417 5004 2423
rect 5021 2423 5027 2437
rect 5044 2437 5324 2443
rect 5396 2437 5836 2443
rect 6020 2437 6124 2443
rect 6365 2443 6371 2457
rect 6292 2437 6371 2443
rect 5021 2417 5516 2423
rect 5764 2417 6476 2423
rect 6564 2417 6892 2423
rect 6900 2417 7260 2423
rect 1410 2414 1470 2416
rect 1410 2406 1411 2414
rect 1420 2406 1421 2414
rect 1459 2406 1460 2414
rect 1469 2406 1470 2414
rect 1410 2404 1470 2406
rect 4418 2414 4478 2416
rect 4418 2406 4419 2414
rect 4428 2406 4429 2414
rect 4467 2406 4468 2414
rect 4477 2406 4478 2414
rect 4418 2404 4478 2406
rect 1588 2397 1788 2403
rect 1860 2397 1900 2403
rect 2132 2397 2220 2403
rect 3028 2397 4403 2403
rect 244 2377 348 2383
rect 420 2377 636 2383
rect 740 2377 1116 2383
rect 1540 2377 1596 2383
rect 1668 2377 1676 2383
rect 1780 2377 2060 2383
rect 2068 2377 2284 2383
rect 2301 2377 2508 2383
rect 340 2357 540 2363
rect 564 2357 652 2363
rect 948 2357 1004 2363
rect 1012 2357 1628 2363
rect 1636 2357 1644 2363
rect 1652 2357 1804 2363
rect 2301 2363 2307 2377
rect 3140 2377 3324 2383
rect 3604 2377 4348 2383
rect 4397 2383 4403 2397
rect 4788 2397 4908 2403
rect 4916 2397 5084 2403
rect 5108 2397 5324 2403
rect 5364 2397 6028 2403
rect 6292 2397 6348 2403
rect 6404 2397 6492 2403
rect 6500 2397 6796 2403
rect 4397 2377 4460 2383
rect 4477 2377 4700 2383
rect 2084 2357 2307 2363
rect 2372 2357 2380 2363
rect 2708 2357 3244 2363
rect 3444 2357 4044 2363
rect 4068 2357 4172 2363
rect 4477 2363 4483 2377
rect 4724 2377 4972 2383
rect 5044 2377 5260 2383
rect 5300 2377 5516 2383
rect 5524 2377 6108 2383
rect 6132 2377 6524 2383
rect 4324 2357 4483 2363
rect 4500 2357 4796 2363
rect 4932 2357 5052 2363
rect 5316 2357 5388 2363
rect 5460 2357 5532 2363
rect 5597 2357 5660 2363
rect 308 2337 364 2343
rect 372 2337 412 2343
rect 564 2337 588 2343
rect 628 2337 684 2343
rect 788 2337 956 2343
rect 1108 2337 1180 2343
rect 1204 2337 1564 2343
rect 1620 2337 1756 2343
rect 1828 2337 1932 2343
rect 2020 2337 2172 2343
rect 2388 2337 2604 2343
rect 3060 2337 4572 2343
rect 4628 2337 5251 2343
rect 212 2317 524 2323
rect 788 2317 844 2323
rect 932 2317 956 2323
rect 1060 2317 1180 2323
rect 1188 2317 1292 2323
rect 1476 2317 2044 2323
rect 2077 2317 2156 2323
rect 2077 2304 2083 2317
rect 2276 2317 2300 2323
rect 2516 2317 2556 2323
rect 2596 2317 2988 2323
rect 3028 2317 3132 2323
rect 3380 2317 3420 2323
rect 3428 2317 3532 2323
rect 3540 2317 3564 2323
rect 3956 2317 4092 2323
rect 4132 2317 4364 2323
rect 4388 2317 4940 2323
rect 4964 2317 5132 2323
rect 5140 2317 5164 2323
rect 5172 2317 5228 2323
rect 5245 2323 5251 2337
rect 5597 2343 5603 2357
rect 5684 2357 5836 2363
rect 5844 2357 6092 2363
rect 6100 2357 6572 2363
rect 5268 2337 5603 2343
rect 5620 2337 5660 2343
rect 5700 2337 5788 2343
rect 5812 2337 6060 2343
rect 6340 2337 6428 2343
rect 6452 2337 6572 2343
rect 6580 2337 6684 2343
rect 7076 2337 7148 2343
rect 7156 2337 7260 2343
rect 7300 2337 7356 2343
rect 5245 2317 5772 2323
rect 5876 2317 6508 2323
rect 6612 2317 6652 2323
rect 7300 2317 7324 2323
rect 100 2297 124 2303
rect 132 2297 204 2303
rect 484 2297 604 2303
rect 740 2297 764 2303
rect 772 2297 1196 2303
rect 1220 2297 1388 2303
rect 1396 2297 1612 2303
rect 1828 2297 1884 2303
rect 1908 2297 1964 2303
rect 2020 2297 2076 2303
rect 2148 2297 2412 2303
rect 2548 2297 2668 2303
rect 2836 2297 2844 2303
rect 2900 2297 3148 2303
rect 3348 2297 3388 2303
rect 3444 2297 3452 2303
rect 3684 2297 3868 2303
rect 4100 2297 4108 2303
rect 4116 2297 4140 2303
rect 4260 2297 4300 2303
rect 4317 2297 4492 2303
rect 84 2277 108 2283
rect 148 2277 316 2283
rect 404 2277 476 2283
rect 900 2277 940 2283
rect 980 2277 1388 2283
rect 1428 2277 1644 2283
rect 2036 2277 2092 2283
rect 2100 2277 2332 2283
rect 2532 2277 2604 2283
rect 2660 2277 2780 2283
rect 2788 2277 2796 2283
rect 2836 2277 2860 2283
rect 3268 2277 3372 2283
rect 3469 2283 3475 2296
rect 3428 2277 3612 2283
rect 4317 2283 4323 2297
rect 4644 2297 4684 2303
rect 4692 2297 4748 2303
rect 4852 2297 5020 2303
rect 5124 2297 5164 2303
rect 5172 2297 5228 2303
rect 5364 2297 5436 2303
rect 5508 2297 5724 2303
rect 5732 2297 6124 2303
rect 6132 2297 6220 2303
rect 6260 2297 6748 2303
rect 3828 2277 4323 2283
rect 4372 2277 4428 2283
rect 4484 2277 4636 2283
rect 4660 2277 4684 2283
rect 4692 2277 4700 2283
rect 4916 2277 4972 2283
rect 5012 2277 5052 2283
rect 5140 2277 5580 2283
rect 5716 2277 5756 2283
rect 5780 2277 6028 2283
rect 6228 2277 6508 2283
rect 6516 2277 6636 2283
rect 6852 2277 6956 2283
rect 6964 2277 7132 2283
rect 7348 2277 7356 2283
rect 20 2257 92 2263
rect 164 2257 220 2263
rect 996 2257 1100 2263
rect 1140 2257 1164 2263
rect 1412 2257 1548 2263
rect 1572 2257 1820 2263
rect 1876 2257 1916 2263
rect 1924 2257 2012 2263
rect 2020 2257 2076 2263
rect 2212 2257 2348 2263
rect 2356 2257 2380 2263
rect 2484 2257 3036 2263
rect 3300 2257 3372 2263
rect 3396 2257 3468 2263
rect 3476 2257 3532 2263
rect 3652 2257 4380 2263
rect 4500 2257 4748 2263
rect 4829 2257 5475 2263
rect 180 2237 412 2243
rect 564 2237 588 2243
rect 852 2237 1052 2243
rect 1284 2237 1324 2243
rect 1620 2237 1628 2243
rect 1684 2237 1724 2243
rect 1748 2237 1820 2243
rect 1908 2237 1916 2243
rect 1924 2237 1948 2243
rect 2244 2237 2348 2243
rect 2548 2237 2652 2243
rect 4829 2243 4835 2257
rect 2980 2237 4835 2243
rect 4852 2237 4908 2243
rect 5092 2237 5244 2243
rect 5252 2237 5260 2243
rect 5332 2237 5372 2243
rect 5469 2243 5475 2257
rect 5492 2257 5500 2263
rect 5572 2257 5628 2263
rect 5636 2257 5692 2263
rect 5700 2257 5820 2263
rect 5828 2257 6220 2263
rect 6228 2257 6252 2263
rect 6269 2257 6332 2263
rect 5469 2237 5644 2243
rect 5901 2237 5932 2243
rect 868 2217 1052 2223
rect 1172 2217 1596 2223
rect 1757 2217 2307 2223
rect 756 2197 972 2203
rect 1156 2197 1372 2203
rect 1757 2203 1763 2217
rect 1588 2197 1763 2203
rect 1780 2197 1836 2203
rect 1844 2197 1884 2203
rect 2301 2203 2307 2217
rect 2324 2217 2860 2223
rect 3188 2217 5868 2223
rect 2914 2214 2974 2216
rect 2914 2206 2915 2214
rect 2924 2206 2925 2214
rect 2963 2206 2964 2214
rect 2973 2206 2974 2214
rect 2914 2204 2974 2206
rect 2301 2197 2444 2203
rect 2500 2197 2716 2203
rect 3300 2197 3516 2203
rect 3524 2197 3564 2203
rect 3956 2197 5084 2203
rect 5124 2197 5484 2203
rect 5604 2197 5660 2203
rect 5860 2197 5884 2203
rect 68 2177 124 2183
rect 132 2177 172 2183
rect 356 2177 595 2183
rect 589 2164 595 2177
rect 1204 2177 1228 2183
rect 1396 2177 1532 2183
rect 1556 2177 1612 2183
rect 1620 2177 1948 2183
rect 1972 2177 2044 2183
rect 2116 2177 2243 2183
rect 100 2157 140 2163
rect 372 2157 428 2163
rect 596 2157 620 2163
rect 628 2157 700 2163
rect 1124 2157 1148 2163
rect 1172 2157 1228 2163
rect 1268 2157 1420 2163
rect 1524 2157 1900 2163
rect 1924 2157 1964 2163
rect 1972 2157 2028 2163
rect 2068 2157 2172 2163
rect 2180 2157 2220 2163
rect 2237 2163 2243 2177
rect 2260 2177 2348 2183
rect 2397 2177 2787 2183
rect 2397 2163 2403 2177
rect 2237 2157 2403 2163
rect 2420 2157 2508 2163
rect 2781 2163 2787 2177
rect 2804 2177 3292 2183
rect 3444 2177 3484 2183
rect 3508 2177 3548 2183
rect 4308 2177 4332 2183
rect 4404 2177 4428 2183
rect 4500 2177 4908 2183
rect 4948 2177 5196 2183
rect 5220 2177 5260 2183
rect 5300 2177 5452 2183
rect 5476 2177 5676 2183
rect 5796 2177 5868 2183
rect 5901 2183 5907 2237
rect 6269 2243 6275 2257
rect 6356 2257 6444 2263
rect 6468 2257 6492 2263
rect 6644 2257 6796 2263
rect 6852 2257 7404 2263
rect 6068 2237 6275 2243
rect 6324 2237 6556 2243
rect 7012 2237 7244 2243
rect 6068 2217 6828 2223
rect 7204 2217 7260 2223
rect 7300 2217 7324 2223
rect 5922 2214 5982 2216
rect 5922 2206 5923 2214
rect 5932 2206 5933 2214
rect 5971 2206 5972 2214
rect 5981 2206 5982 2214
rect 5922 2204 5982 2206
rect 6068 2197 6460 2203
rect 6772 2197 6876 2203
rect 7284 2197 7292 2203
rect 5901 2177 5939 2183
rect 5933 2164 5939 2177
rect 6036 2177 6300 2183
rect 6324 2177 6764 2183
rect 7204 2177 7276 2183
rect 2781 2157 3020 2163
rect 3476 2157 3676 2163
rect 3796 2157 4044 2163
rect 4276 2157 4300 2163
rect 4532 2157 4940 2163
rect 5012 2157 5324 2163
rect 5428 2157 5788 2163
rect 5844 2157 5916 2163
rect 5940 2157 6076 2163
rect 6084 2157 6492 2163
rect 6500 2157 6572 2163
rect 6733 2157 7164 2163
rect 6733 2144 6739 2157
rect 7284 2157 7308 2163
rect 36 2137 156 2143
rect 164 2137 428 2143
rect 452 2137 508 2143
rect 964 2137 1260 2143
rect 1300 2137 1612 2143
rect 1796 2137 1980 2143
rect 2164 2137 2204 2143
rect 2292 2137 2300 2143
rect 2356 2137 2604 2143
rect 2644 2137 2780 2143
rect 2868 2137 3020 2143
rect 3108 2137 3196 2143
rect 3204 2137 3500 2143
rect 3780 2137 3932 2143
rect 3940 2137 4124 2143
rect 4276 2137 4300 2143
rect 4340 2137 4556 2143
rect 4564 2137 4652 2143
rect 4724 2137 4940 2143
rect 4964 2137 5100 2143
rect 5188 2137 5580 2143
rect 5620 2137 5948 2143
rect 5981 2137 6060 2143
rect 132 2117 172 2123
rect 404 2117 476 2123
rect 612 2117 700 2123
rect 708 2117 748 2123
rect 756 2117 828 2123
rect 836 2117 860 2123
rect 996 2117 1212 2123
rect 1396 2117 1548 2123
rect 1700 2117 1772 2123
rect 1860 2117 1916 2123
rect 2004 2117 2412 2123
rect 2420 2117 2572 2123
rect 3101 2123 3107 2136
rect 2900 2117 3107 2123
rect 3188 2117 3260 2123
rect 3604 2117 3724 2123
rect 3988 2117 4524 2123
rect 4532 2117 4540 2123
rect 4548 2117 4636 2123
rect 4772 2117 4860 2123
rect 4884 2117 4892 2123
rect 5108 2117 5132 2123
rect 5156 2117 5452 2123
rect 5524 2117 5532 2123
rect 5981 2123 5987 2137
rect 6260 2137 6332 2143
rect 6349 2137 6380 2143
rect 5549 2117 5987 2123
rect 244 2097 604 2103
rect 916 2097 940 2103
rect 948 2097 1052 2103
rect 1060 2097 1100 2103
rect 1108 2097 1372 2103
rect 1380 2097 1484 2103
rect 1492 2097 1852 2103
rect 2036 2097 2140 2103
rect 2164 2097 2284 2103
rect 2372 2097 2396 2103
rect 2404 2097 2444 2103
rect 2468 2097 2524 2103
rect 2548 2097 2572 2103
rect 2628 2097 2828 2103
rect 3012 2097 3020 2103
rect 3172 2097 3948 2103
rect 4004 2097 4332 2103
rect 4372 2097 4716 2103
rect 4740 2097 4828 2103
rect 4852 2097 4972 2103
rect 5076 2097 5244 2103
rect 5252 2097 5308 2103
rect 5396 2097 5427 2103
rect 372 2077 428 2083
rect 516 2077 556 2083
rect 692 2077 812 2083
rect 916 2077 956 2083
rect 1188 2077 1468 2083
rect 1508 2077 1644 2083
rect 1924 2077 2220 2083
rect 2804 2077 3971 2083
rect 388 2057 444 2063
rect 452 2057 1443 2063
rect 436 2037 572 2043
rect 1108 2037 1340 2043
rect 1348 2037 1420 2043
rect 1437 2043 1443 2057
rect 1716 2057 2092 2063
rect 2100 2057 2108 2063
rect 2196 2057 2428 2063
rect 3156 2057 3212 2063
rect 3556 2057 3580 2063
rect 3965 2063 3971 2077
rect 4020 2077 4060 2083
rect 4196 2077 4364 2083
rect 4404 2077 4524 2083
rect 4548 2077 5004 2083
rect 5044 2077 5052 2083
rect 5108 2077 5148 2083
rect 5204 2077 5228 2083
rect 5268 2077 5292 2083
rect 5348 2077 5372 2083
rect 5396 2077 5404 2083
rect 5421 2083 5427 2097
rect 5549 2103 5555 2117
rect 6349 2123 6355 2137
rect 6484 2137 6508 2143
rect 6516 2137 6732 2143
rect 6852 2137 6908 2143
rect 6932 2137 7068 2143
rect 6036 2117 6355 2123
rect 6372 2117 6508 2123
rect 6564 2117 6636 2123
rect 6660 2117 6796 2123
rect 6804 2117 6956 2123
rect 5476 2097 5555 2103
rect 5652 2097 5804 2103
rect 5956 2097 6060 2103
rect 6132 2097 6284 2103
rect 6324 2097 6620 2103
rect 6708 2097 6748 2103
rect 6772 2097 6876 2103
rect 6884 2097 6924 2103
rect 7348 2097 7404 2103
rect 5421 2077 6540 2083
rect 7044 2077 7372 2083
rect 3965 2057 5484 2063
rect 5524 2057 5564 2063
rect 5908 2057 6028 2063
rect 6036 2057 6364 2063
rect 6372 2057 6444 2063
rect 6452 2057 6716 2063
rect 1437 2037 2108 2043
rect 2644 2037 2796 2043
rect 3140 2037 3212 2043
rect 3220 2037 3308 2043
rect 3572 2037 3612 2043
rect 3828 2037 4012 2043
rect 4148 2037 6035 2043
rect 468 2017 892 2023
rect 1556 2017 1660 2023
rect 1764 2017 1868 2023
rect 2020 2017 2124 2023
rect 2452 2017 2643 2023
rect 1410 2014 1470 2016
rect 1410 2006 1411 2014
rect 1420 2006 1421 2014
rect 1459 2006 1460 2014
rect 1469 2006 1470 2014
rect 1410 2004 1470 2006
rect 564 1997 1020 2003
rect 1524 1997 2444 2003
rect 2637 2003 2643 2017
rect 2660 2017 2892 2023
rect 3044 2017 4396 2023
rect 4532 2017 4604 2023
rect 5172 2017 5340 2023
rect 5348 2017 5436 2023
rect 5460 2017 5596 2023
rect 5924 2017 6012 2023
rect 6029 2023 6035 2037
rect 6068 2037 6412 2043
rect 6029 2017 6764 2023
rect 7124 2017 7196 2023
rect 4418 2014 4478 2016
rect 4418 2006 4419 2014
rect 4428 2006 4429 2014
rect 4467 2006 4468 2014
rect 4477 2006 4478 2014
rect 4418 2004 4478 2006
rect 2637 1997 2876 2003
rect 3252 1997 3356 2003
rect 3892 1997 4067 2003
rect 532 1977 652 1983
rect 980 1977 1372 1983
rect 1380 1977 1692 1983
rect 1732 1977 2188 1983
rect 2676 1977 2780 1983
rect 2788 1977 2924 1983
rect 3044 1977 4028 1983
rect 4061 1983 4067 1997
rect 4580 1997 4908 2003
rect 5172 1997 5532 2003
rect 5549 1997 6076 2003
rect 4061 1977 4620 1983
rect 4756 1977 4860 1983
rect 4900 1977 5180 1983
rect 5220 1977 5324 1983
rect 5549 1983 5555 1997
rect 6212 1997 6700 2003
rect 5380 1977 5555 1983
rect 5565 1977 6140 1983
rect 484 1957 1516 1963
rect 1556 1957 1708 1963
rect 1741 1957 2780 1963
rect 372 1937 572 1943
rect 676 1937 716 1943
rect 724 1937 1036 1943
rect 1076 1937 1164 1943
rect 1412 1937 1580 1943
rect 1741 1943 1747 1957
rect 2804 1957 2988 1963
rect 2996 1957 3292 1963
rect 3300 1957 3692 1963
rect 3812 1957 4316 1963
rect 4356 1957 4492 1963
rect 4516 1957 4780 1963
rect 5565 1963 5571 1977
rect 6180 1977 6460 1983
rect 4916 1957 5571 1963
rect 6036 1957 6060 1963
rect 6084 1957 7004 1963
rect 1668 1937 1747 1943
rect 1764 1937 1836 1943
rect 1860 1937 2188 1943
rect 2308 1937 2348 1943
rect 2404 1937 2460 1943
rect 2916 1937 3132 1943
rect 3876 1937 4060 1943
rect 4148 1937 4236 1943
rect 4269 1937 4556 1943
rect 180 1917 300 1923
rect 532 1917 636 1923
rect 660 1917 860 1923
rect 1172 1917 1212 1923
rect 1524 1917 1596 1923
rect 1636 1917 1676 1923
rect 1700 1917 1788 1923
rect 1972 1917 2012 1923
rect 2164 1917 2300 1923
rect 2356 1917 2412 1923
rect 2420 1917 2764 1923
rect 2788 1917 3036 1923
rect 3124 1917 3164 1923
rect 3396 1917 3468 1923
rect 3668 1917 3900 1923
rect 4020 1917 4092 1923
rect 4269 1923 4275 1937
rect 4596 1937 4812 1943
rect 4884 1937 5452 1943
rect 5476 1937 5612 1943
rect 5796 1937 5932 1943
rect 6004 1937 6076 1943
rect 6084 1937 6140 1943
rect 6308 1937 6396 1943
rect 6404 1937 6796 1943
rect 7092 1937 7180 1943
rect 7188 1937 7196 1943
rect 4205 1917 4275 1923
rect 52 1897 67 1903
rect 20 1877 44 1883
rect 61 1883 67 1897
rect 116 1897 236 1903
rect 244 1897 556 1903
rect 596 1897 652 1903
rect 692 1897 796 1903
rect 1044 1897 1116 1903
rect 1172 1897 1212 1903
rect 1332 1897 1484 1903
rect 1620 1897 1660 1903
rect 1812 1897 1836 1903
rect 2052 1897 2076 1903
rect 2084 1897 2220 1903
rect 2228 1897 2316 1903
rect 2388 1897 2492 1903
rect 2532 1897 2556 1903
rect 2564 1897 2652 1903
rect 2756 1897 2796 1903
rect 2932 1897 3052 1903
rect 3060 1897 3100 1903
rect 3332 1897 3356 1903
rect 3460 1897 3500 1903
rect 3524 1897 3548 1903
rect 3556 1897 3628 1903
rect 3636 1897 3724 1903
rect 3732 1897 3788 1903
rect 3796 1897 3836 1903
rect 3924 1897 3964 1903
rect 4205 1903 4211 1917
rect 4292 1917 4348 1923
rect 4596 1917 4620 1923
rect 4644 1917 4716 1923
rect 4836 1917 5260 1923
rect 5364 1917 5452 1923
rect 5540 1917 6012 1923
rect 6036 1917 6092 1923
rect 6484 1917 6540 1923
rect 6548 1917 6620 1923
rect 6628 1917 6668 1923
rect 6724 1917 6764 1923
rect 7028 1917 7068 1923
rect 7076 1917 7443 1923
rect 4036 1897 4211 1903
rect 4228 1897 4508 1903
rect 4532 1897 4588 1903
rect 4596 1897 4652 1903
rect 4724 1897 4732 1903
rect 4772 1897 4844 1903
rect 4948 1897 5148 1903
rect 5412 1897 5596 1903
rect 5668 1897 5804 1903
rect 5908 1897 6172 1903
rect 6292 1897 6684 1903
rect 6772 1897 6908 1903
rect 7076 1897 7148 1903
rect 7188 1897 7308 1903
rect 7437 1897 7443 1917
rect 61 1877 140 1883
rect 148 1877 204 1883
rect 628 1877 716 1883
rect 788 1877 812 1883
rect 836 1877 876 1883
rect 1044 1877 1068 1883
rect 1220 1877 1276 1883
rect 1652 1877 1708 1883
rect 1716 1877 1868 1883
rect 1876 1877 2252 1883
rect 2260 1877 2268 1883
rect 2308 1877 2332 1883
rect 2452 1877 2460 1883
rect 2468 1877 2476 1883
rect 2548 1877 2588 1883
rect 2596 1877 2636 1883
rect 2708 1877 2716 1883
rect 2724 1877 2812 1883
rect 2820 1877 3084 1883
rect 3092 1877 3180 1883
rect 3348 1877 3388 1883
rect 3716 1877 3884 1883
rect 3892 1877 4028 1883
rect 4084 1877 4092 1883
rect 4164 1877 4268 1883
rect 4548 1877 4604 1883
rect 4612 1877 4668 1883
rect 4756 1877 5132 1883
rect 5140 1877 5516 1883
rect 5540 1877 5548 1883
rect 5844 1877 5916 1883
rect 5940 1877 6028 1883
rect 6084 1877 6412 1883
rect 6420 1877 6572 1883
rect 6580 1877 6844 1883
rect 6964 1877 6972 1883
rect 6980 1877 7004 1883
rect 7012 1877 7260 1883
rect 212 1857 268 1863
rect 420 1857 444 1863
rect 1188 1857 1276 1863
rect 1556 1857 1612 1863
rect 1620 1857 1772 1863
rect 1844 1857 1916 1863
rect 2004 1857 2060 1863
rect 2100 1857 2476 1863
rect 2500 1857 2732 1863
rect 2788 1857 2908 1863
rect 3060 1857 3084 1863
rect 3172 1857 3452 1863
rect 3588 1857 3724 1863
rect 3732 1857 3756 1863
rect 3764 1857 3820 1863
rect 4068 1857 4204 1863
rect 4244 1857 4572 1863
rect 4660 1857 4876 1863
rect 4916 1857 5468 1863
rect 5524 1857 5571 1863
rect 468 1837 524 1843
rect 1524 1837 2012 1843
rect 2148 1837 2284 1843
rect 2292 1837 2716 1843
rect 2884 1837 4092 1843
rect 4196 1837 4220 1843
rect 4228 1837 4252 1843
rect 4292 1837 4588 1843
rect 4628 1837 4716 1843
rect 4804 1837 5548 1843
rect 5565 1843 5571 1857
rect 5588 1857 6300 1863
rect 6308 1857 6316 1863
rect 6356 1857 6444 1863
rect 6452 1857 6588 1863
rect 6596 1857 6796 1863
rect 7124 1857 7260 1863
rect 5565 1837 5683 1843
rect 740 1817 940 1823
rect 1732 1817 1772 1823
rect 1972 1817 2204 1823
rect 2484 1817 2492 1823
rect 2500 1817 2572 1823
rect 2708 1817 2780 1823
rect 3380 1817 3420 1823
rect 3428 1817 3516 1823
rect 3524 1817 3564 1823
rect 3572 1817 4012 1823
rect 4020 1817 4300 1823
rect 4324 1817 4348 1823
rect 4356 1817 4396 1823
rect 4628 1817 5660 1823
rect 5677 1823 5683 1837
rect 5748 1837 6460 1843
rect 6500 1837 7180 1843
rect 7188 1837 7324 1843
rect 5677 1817 5900 1823
rect 6036 1817 6076 1823
rect 7124 1817 7180 1823
rect 2914 1814 2974 1816
rect 2914 1806 2915 1814
rect 2924 1806 2925 1814
rect 2963 1806 2964 1814
rect 2973 1806 2974 1814
rect 2914 1804 2974 1806
rect 5922 1814 5982 1816
rect 5922 1806 5923 1814
rect 5932 1806 5933 1814
rect 5971 1806 5972 1814
rect 5981 1806 5982 1814
rect 5922 1804 5982 1806
rect 1604 1797 1948 1803
rect 1956 1797 2012 1803
rect 2020 1797 2076 1803
rect 2212 1797 2316 1803
rect 3236 1797 3324 1803
rect 3332 1797 3436 1803
rect 3444 1797 3532 1803
rect 3764 1797 4076 1803
rect 4340 1797 4588 1803
rect 4605 1797 4828 1803
rect 1220 1777 1388 1783
rect 1652 1777 1868 1783
rect 2116 1777 2124 1783
rect 2132 1777 2476 1783
rect 2548 1777 2604 1783
rect 3076 1777 3244 1783
rect 3524 1777 3628 1783
rect 3636 1777 3772 1783
rect 3956 1777 3980 1783
rect 4212 1777 4316 1783
rect 4605 1783 4611 1797
rect 5012 1797 5276 1803
rect 5300 1797 5708 1803
rect 6020 1797 6044 1803
rect 6516 1797 6700 1803
rect 6708 1797 6780 1803
rect 4340 1777 4611 1783
rect 4644 1777 4700 1783
rect 4756 1777 5388 1783
rect 5444 1777 5708 1783
rect 5748 1777 5756 1783
rect 5764 1777 6044 1783
rect 6052 1777 6364 1783
rect 6372 1777 6620 1783
rect 7252 1777 7292 1783
rect 100 1757 140 1763
rect 148 1757 700 1763
rect 756 1757 796 1763
rect 852 1757 940 1763
rect 1028 1757 1564 1763
rect 1940 1757 2284 1763
rect 2340 1757 2508 1763
rect 2692 1757 2732 1763
rect 2884 1757 3004 1763
rect 3012 1757 3132 1763
rect 3140 1757 3212 1763
rect 3220 1757 3260 1763
rect 3277 1757 3740 1763
rect 84 1737 172 1743
rect 340 1737 428 1743
rect 468 1737 492 1743
rect 500 1737 604 1743
rect 772 1737 844 1743
rect 1076 1737 1340 1743
rect 1556 1737 1612 1743
rect 1620 1737 1692 1743
rect 1716 1737 1756 1743
rect 1764 1737 1836 1743
rect 2068 1737 2252 1743
rect 2372 1737 2396 1743
rect 2404 1737 2476 1743
rect 2564 1737 2732 1743
rect 3060 1737 3100 1743
rect 3277 1743 3283 1757
rect 3988 1757 4012 1763
rect 4228 1757 4524 1763
rect 4564 1757 4908 1763
rect 5092 1757 5148 1763
rect 5348 1757 5404 1763
rect 5428 1757 5708 1763
rect 5780 1757 6492 1763
rect 6660 1757 6908 1763
rect 7156 1757 7340 1763
rect 3188 1737 3283 1743
rect 3380 1737 3388 1743
rect 3604 1737 3692 1743
rect 3700 1737 4396 1743
rect 4660 1737 5123 1743
rect 196 1717 268 1723
rect 276 1717 348 1723
rect 356 1717 396 1723
rect 461 1723 467 1736
rect 420 1717 467 1723
rect 820 1717 972 1723
rect 1140 1717 1164 1723
rect 1172 1717 1484 1723
rect 1636 1717 1836 1723
rect 1844 1717 1916 1723
rect 2036 1717 2108 1723
rect 2244 1717 2268 1723
rect 2452 1717 2540 1723
rect 2772 1717 2812 1723
rect 3012 1717 3052 1723
rect 3268 1717 3276 1723
rect 3284 1717 3420 1723
rect 3476 1717 3596 1723
rect 3748 1717 3756 1723
rect 3764 1717 3788 1723
rect 4036 1717 4124 1723
rect 4132 1717 4204 1723
rect 4500 1717 4556 1723
rect 4628 1717 4668 1723
rect 4996 1717 5068 1723
rect 5117 1723 5123 1737
rect 5245 1737 5340 1743
rect 5245 1723 5251 1737
rect 5364 1737 5420 1743
rect 5492 1737 5740 1743
rect 5844 1737 5875 1743
rect 5117 1717 5251 1723
rect 5268 1717 5452 1723
rect 5460 1717 5548 1723
rect 5556 1717 5788 1723
rect 5796 1717 5852 1723
rect 5869 1723 5875 1737
rect 5908 1737 5996 1743
rect 6196 1737 6252 1743
rect 6580 1737 6588 1743
rect 7060 1737 7308 1743
rect 5869 1717 6316 1723
rect 6436 1717 6492 1723
rect 6548 1717 6652 1723
rect 7044 1717 7116 1723
rect 7236 1717 7260 1723
rect 7268 1717 7292 1723
rect 180 1697 204 1703
rect 388 1697 476 1703
rect 484 1697 588 1703
rect 596 1697 636 1703
rect 660 1697 748 1703
rect 756 1697 892 1703
rect 900 1697 1004 1703
rect 1124 1697 1228 1703
rect 1236 1697 1292 1703
rect 1636 1697 2092 1703
rect 2116 1697 2259 1703
rect 756 1677 780 1683
rect 836 1677 956 1683
rect 1700 1677 1756 1683
rect 1764 1677 1820 1683
rect 1908 1677 1932 1683
rect 1940 1677 1996 1683
rect 2004 1677 2060 1683
rect 2068 1677 2236 1683
rect 2253 1683 2259 1697
rect 2324 1697 2348 1703
rect 2388 1697 2508 1703
rect 2724 1697 2828 1703
rect 2852 1697 2988 1703
rect 2996 1697 3164 1703
rect 3204 1697 3868 1703
rect 3876 1697 4108 1703
rect 4308 1697 4540 1703
rect 4580 1697 4716 1703
rect 4724 1697 4748 1703
rect 4756 1697 4780 1703
rect 4788 1697 4892 1703
rect 4900 1697 5068 1703
rect 5076 1697 5372 1703
rect 5396 1697 5516 1703
rect 5588 1697 5644 1703
rect 5652 1697 5692 1703
rect 5716 1697 6252 1703
rect 7188 1697 7228 1703
rect 7412 1697 7443 1703
rect 2253 1677 2588 1683
rect 3636 1677 3660 1683
rect 3988 1677 4044 1683
rect 4100 1677 4636 1683
rect 4676 1677 4684 1683
rect 4708 1677 4764 1683
rect 4804 1677 4844 1683
rect 4932 1677 5132 1683
rect 5268 1677 5292 1683
rect 5533 1683 5539 1696
rect 5364 1677 5539 1683
rect 5604 1677 5820 1683
rect 5860 1677 6076 1683
rect 6116 1677 6556 1683
rect 6564 1677 7180 1683
rect 7204 1677 7276 1683
rect 52 1657 668 1663
rect 676 1657 1116 1663
rect 1300 1657 1340 1663
rect 2164 1657 2332 1663
rect 2356 1657 2396 1663
rect 2660 1657 3660 1663
rect 3684 1657 4323 1663
rect 660 1637 892 1643
rect 964 1637 1084 1643
rect 1140 1637 1148 1643
rect 1156 1637 1628 1643
rect 1716 1637 3052 1643
rect 3668 1637 3724 1643
rect 3972 1637 3996 1643
rect 4317 1643 4323 1657
rect 4564 1657 4588 1663
rect 5188 1657 5324 1663
rect 5332 1657 5452 1663
rect 5556 1657 5580 1663
rect 5636 1657 5980 1663
rect 6180 1657 6204 1663
rect 6292 1657 7404 1663
rect 4317 1637 5612 1643
rect 5693 1637 5884 1643
rect 900 1617 1276 1623
rect 1284 1617 1324 1623
rect 1748 1617 1804 1623
rect 1876 1617 2092 1623
rect 2132 1617 3772 1623
rect 3780 1617 4236 1623
rect 4500 1617 4716 1623
rect 4756 1617 4812 1623
rect 5693 1623 5699 1637
rect 5892 1637 6524 1643
rect 4980 1617 5699 1623
rect 5716 1617 6220 1623
rect 6308 1617 7164 1623
rect 7172 1617 7212 1623
rect 1410 1614 1470 1616
rect 1410 1606 1411 1614
rect 1420 1606 1421 1614
rect 1459 1606 1460 1614
rect 1469 1606 1470 1614
rect 1410 1604 1470 1606
rect 4418 1614 4478 1616
rect 4418 1606 4419 1614
rect 4428 1606 4429 1614
rect 4467 1606 4468 1614
rect 4477 1606 4478 1614
rect 4418 1604 4478 1606
rect 500 1597 540 1603
rect 788 1597 956 1603
rect 996 1597 1068 1603
rect 1524 1597 3676 1603
rect 3732 1597 3788 1603
rect 4164 1597 4364 1603
rect 4532 1597 4748 1603
rect 5060 1597 5212 1603
rect 5412 1597 5420 1603
rect 5460 1597 5628 1603
rect 5700 1597 6204 1603
rect 868 1577 876 1583
rect 932 1577 2915 1583
rect 628 1557 700 1563
rect 740 1557 796 1563
rect 804 1557 860 1563
rect 1076 1557 1212 1563
rect 1236 1557 1308 1563
rect 1572 1557 1740 1563
rect 1780 1557 1868 1563
rect 2004 1557 2204 1563
rect 2340 1557 2428 1563
rect 2909 1563 2915 1577
rect 3108 1577 3196 1583
rect 3204 1577 3980 1583
rect 4260 1577 4604 1583
rect 4660 1577 4684 1583
rect 5284 1577 5532 1583
rect 5540 1577 6124 1583
rect 2909 1557 3340 1563
rect 3348 1557 3644 1563
rect 4100 1557 4764 1563
rect 4884 1557 5292 1563
rect 5396 1557 5404 1563
rect 5732 1557 6268 1563
rect 6276 1557 6348 1563
rect 6468 1557 7180 1563
rect 7204 1557 7276 1563
rect 500 1537 748 1543
rect 756 1537 924 1543
rect 980 1537 1004 1543
rect 1021 1537 1068 1543
rect 676 1517 764 1523
rect 788 1517 828 1523
rect 884 1517 940 1523
rect 1021 1523 1027 1537
rect 1172 1537 1596 1543
rect 1604 1537 1852 1543
rect 2068 1537 2252 1543
rect 2276 1537 2380 1543
rect 2404 1537 3084 1543
rect 3732 1537 3804 1543
rect 4276 1537 4460 1543
rect 4820 1537 5036 1543
rect 5124 1537 5324 1543
rect 5332 1537 5420 1543
rect 5812 1537 6044 1543
rect 6356 1537 6364 1543
rect 6372 1537 7324 1543
rect 964 1517 1027 1523
rect 1044 1517 1052 1523
rect 1092 1517 1244 1523
rect 1540 1517 1724 1523
rect 1732 1517 1804 1523
rect 1860 1517 1980 1523
rect 2100 1517 2172 1523
rect 2228 1517 2364 1523
rect 2452 1517 2588 1523
rect 2612 1517 2828 1523
rect 2868 1517 2908 1523
rect 3012 1517 3020 1523
rect 3060 1517 3212 1523
rect 3668 1517 3916 1523
rect 4116 1517 4172 1523
rect 4388 1517 4412 1523
rect 4420 1517 4748 1523
rect 4948 1517 5004 1523
rect 5012 1517 5020 1523
rect 5092 1517 5596 1523
rect 5876 1517 5900 1523
rect 6004 1517 6172 1523
rect 6260 1517 6444 1523
rect 6516 1517 6524 1523
rect 6532 1517 6572 1523
rect 6996 1517 7036 1523
rect 7252 1517 7283 1523
rect 7277 1504 7283 1517
rect 52 1497 108 1503
rect 324 1497 700 1503
rect 724 1497 780 1503
rect 788 1497 844 1503
rect 957 1497 972 1503
rect 324 1477 380 1483
rect 388 1477 556 1483
rect 957 1483 963 1497
rect 1172 1497 1212 1503
rect 1284 1497 1404 1503
rect 1572 1497 1612 1503
rect 1620 1497 1676 1503
rect 1684 1497 1756 1503
rect 1844 1497 1884 1503
rect 2196 1497 2236 1503
rect 2292 1497 2764 1503
rect 2804 1497 3116 1503
rect 3156 1497 3180 1503
rect 3556 1497 3612 1503
rect 3636 1497 3708 1503
rect 3716 1497 3756 1503
rect 3764 1497 3836 1503
rect 3860 1497 4332 1503
rect 4372 1497 4524 1503
rect 4548 1497 4556 1503
rect 4596 1497 4604 1503
rect 4900 1497 5020 1503
rect 5140 1497 5308 1503
rect 5316 1497 5436 1503
rect 5668 1497 5788 1503
rect 5908 1497 6140 1503
rect 6580 1497 7004 1503
rect 4813 1484 4819 1496
rect 820 1477 963 1483
rect 980 1477 1036 1483
rect 1380 1477 1555 1483
rect 20 1457 44 1463
rect 68 1457 140 1463
rect 148 1457 204 1463
rect 212 1457 492 1463
rect 516 1457 652 1463
rect 884 1457 1132 1463
rect 1188 1457 1532 1463
rect 1549 1463 1555 1477
rect 1588 1477 1644 1483
rect 1716 1477 2060 1483
rect 2100 1477 2268 1483
rect 2292 1477 2460 1483
rect 2484 1477 2492 1483
rect 2500 1477 2604 1483
rect 2644 1477 2700 1483
rect 2740 1477 3388 1483
rect 3428 1477 3436 1483
rect 3828 1477 4076 1483
rect 4084 1477 4236 1483
rect 4372 1477 4508 1483
rect 4532 1477 4716 1483
rect 4724 1477 4796 1483
rect 5069 1483 5075 1496
rect 5012 1477 5043 1483
rect 5069 1477 5180 1483
rect 1549 1457 1596 1463
rect 1652 1457 1788 1463
rect 1940 1457 2076 1463
rect 2228 1457 2300 1463
rect 2324 1457 2652 1463
rect 2676 1457 2700 1463
rect 2708 1457 2796 1463
rect 2804 1457 2892 1463
rect 3140 1457 3260 1463
rect 3268 1457 3612 1463
rect 3908 1457 3980 1463
rect 4292 1457 4508 1463
rect 4564 1457 4700 1463
rect 4820 1457 5020 1463
rect 5037 1463 5043 1477
rect 5236 1477 5292 1483
rect 5332 1477 5372 1483
rect 5860 1477 5916 1483
rect 6228 1477 6540 1483
rect 6548 1477 7052 1483
rect 7060 1477 7212 1483
rect 7220 1477 7308 1483
rect 7316 1477 7356 1483
rect 5037 1457 5212 1463
rect 5556 1457 5564 1463
rect 5732 1457 5772 1463
rect 5780 1457 5820 1463
rect 5828 1457 5868 1463
rect 5876 1457 6060 1463
rect 6340 1457 6380 1463
rect 6388 1457 6476 1463
rect 6868 1457 7068 1463
rect 7252 1457 7292 1463
rect 212 1437 236 1443
rect 244 1437 332 1443
rect 340 1437 476 1443
rect 532 1437 588 1443
rect 660 1437 684 1443
rect 1140 1437 1260 1443
rect 1316 1437 1980 1443
rect 2020 1437 2124 1443
rect 2212 1437 2284 1443
rect 2308 1437 2460 1443
rect 2516 1437 2572 1443
rect 2580 1437 2636 1443
rect 2644 1437 2684 1443
rect 2692 1437 2796 1443
rect 2804 1437 2876 1443
rect 2884 1437 3068 1443
rect 3252 1437 3420 1443
rect 3604 1437 3724 1443
rect 3924 1437 4163 1443
rect 100 1417 156 1423
rect 164 1417 220 1423
rect 525 1423 531 1436
rect 228 1417 531 1423
rect 948 1417 988 1423
rect 1012 1417 1020 1423
rect 1076 1417 1180 1423
rect 1332 1417 1372 1423
rect 1396 1417 2348 1423
rect 2372 1417 2483 1423
rect 228 1397 268 1403
rect 276 1397 364 1403
rect 852 1397 908 1403
rect 1028 1397 2396 1403
rect 2477 1403 2483 1417
rect 2500 1417 2556 1423
rect 2564 1417 2668 1423
rect 3044 1417 3084 1423
rect 3156 1417 3484 1423
rect 3508 1417 4140 1423
rect 4157 1423 4163 1437
rect 4244 1437 4492 1443
rect 4628 1437 4652 1443
rect 4676 1437 4828 1443
rect 4884 1437 5084 1443
rect 5428 1437 6076 1443
rect 6148 1437 6396 1443
rect 6420 1437 6428 1443
rect 6772 1437 6972 1443
rect 6996 1437 7004 1443
rect 7012 1437 7052 1443
rect 7060 1437 7308 1443
rect 4157 1417 4428 1423
rect 4516 1417 4556 1423
rect 4580 1417 4892 1423
rect 4916 1417 5180 1423
rect 5204 1417 5308 1423
rect 6068 1417 6156 1423
rect 6164 1417 6220 1423
rect 6916 1417 6988 1423
rect 7284 1417 7372 1423
rect 2914 1414 2974 1416
rect 2914 1406 2915 1414
rect 2924 1406 2925 1414
rect 2963 1406 2964 1414
rect 2973 1406 2974 1414
rect 2914 1404 2974 1406
rect 5922 1414 5982 1416
rect 5922 1406 5923 1414
rect 5932 1406 5933 1414
rect 5971 1406 5972 1414
rect 5981 1406 5982 1414
rect 5922 1404 5982 1406
rect 2477 1397 2652 1403
rect 2669 1397 2860 1403
rect 164 1377 252 1383
rect 397 1377 972 1383
rect 397 1363 403 1377
rect 1108 1377 1260 1383
rect 1332 1377 1500 1383
rect 2036 1377 2044 1383
rect 2068 1377 2300 1383
rect 2404 1377 2428 1383
rect 2484 1377 2540 1383
rect 2580 1377 2604 1383
rect 2669 1383 2675 1397
rect 3124 1397 3276 1403
rect 3373 1397 3564 1403
rect 2660 1377 2675 1383
rect 2708 1377 2860 1383
rect 2884 1377 2908 1383
rect 3156 1377 3196 1383
rect 3373 1383 3379 1397
rect 3876 1397 4307 1403
rect 3300 1377 3379 1383
rect 3396 1377 3884 1383
rect 4301 1383 4307 1397
rect 4324 1397 4780 1403
rect 4788 1397 4844 1403
rect 4852 1397 5484 1403
rect 6164 1397 6188 1403
rect 6212 1397 6444 1403
rect 6532 1397 6668 1403
rect 6964 1397 7084 1403
rect 7092 1397 7164 1403
rect 7300 1397 7404 1403
rect 4301 1377 4652 1383
rect 4740 1377 4764 1383
rect 4788 1377 5011 1383
rect 276 1357 403 1363
rect 420 1357 524 1363
rect 612 1357 700 1363
rect 708 1357 812 1363
rect 1236 1357 1340 1363
rect 1428 1357 1548 1363
rect 1556 1357 1692 1363
rect 1940 1357 2092 1363
rect 2260 1357 2300 1363
rect 2340 1357 2588 1363
rect 2612 1357 2732 1363
rect 2772 1357 2819 1363
rect 2813 1344 2819 1357
rect 2836 1357 2860 1363
rect 2900 1357 2924 1363
rect 2948 1357 3404 1363
rect 3620 1357 3692 1363
rect 3780 1357 3996 1363
rect 4084 1357 4300 1363
rect 4404 1357 4940 1363
rect 5005 1363 5011 1377
rect 5028 1377 5052 1383
rect 5076 1377 5356 1383
rect 5492 1377 5516 1383
rect 5668 1377 5708 1383
rect 5716 1377 5820 1383
rect 5828 1377 5932 1383
rect 6020 1377 6540 1383
rect 6660 1377 6716 1383
rect 7188 1377 7308 1383
rect 5005 1357 5244 1363
rect 5268 1357 5468 1363
rect 5508 1357 7116 1363
rect 7316 1357 7340 1363
rect 516 1337 668 1343
rect 772 1337 1628 1343
rect 1684 1337 1708 1343
rect 1796 1337 1964 1343
rect 1988 1337 2060 1343
rect 2404 1337 2412 1343
rect 2452 1337 2524 1343
rect 2548 1337 2588 1343
rect 2644 1337 2684 1343
rect 2724 1337 2780 1343
rect 2820 1337 2924 1343
rect 2941 1337 3068 1343
rect 148 1317 188 1323
rect 196 1317 220 1323
rect 596 1317 620 1323
rect 852 1317 892 1323
rect 932 1317 1036 1323
rect 1076 1317 1100 1323
rect 1156 1317 1180 1323
rect 1620 1317 1660 1323
rect 1684 1317 1708 1323
rect 1908 1317 1964 1323
rect 1988 1317 1996 1323
rect 2004 1317 2044 1323
rect 2084 1317 2172 1323
rect 2228 1317 2268 1323
rect 2420 1317 2444 1323
rect 2468 1317 2604 1323
rect 2628 1317 2636 1323
rect 2676 1317 2732 1323
rect 2756 1317 2844 1323
rect 2941 1323 2947 1337
rect 3092 1337 3100 1343
rect 3268 1337 3356 1343
rect 3476 1337 3596 1343
rect 3652 1337 3836 1343
rect 3924 1337 3964 1343
rect 4125 1337 4572 1343
rect 2868 1317 2947 1323
rect 3044 1317 3324 1323
rect 3444 1317 3548 1323
rect 4125 1323 4131 1337
rect 4596 1337 4780 1343
rect 4964 1337 4988 1343
rect 4996 1337 5036 1343
rect 5044 1337 5084 1343
rect 5220 1337 5340 1343
rect 5348 1337 5388 1343
rect 5396 1337 5436 1343
rect 5444 1337 5484 1343
rect 5604 1337 5628 1343
rect 5636 1337 5868 1343
rect 5876 1337 6108 1343
rect 6116 1337 6172 1343
rect 6436 1337 6476 1343
rect 6596 1337 6732 1343
rect 6868 1337 6876 1343
rect 7156 1337 7356 1343
rect 3572 1317 4131 1323
rect 4148 1317 4556 1323
rect 4612 1317 4620 1323
rect 4740 1317 4956 1323
rect 4980 1317 5196 1323
rect 5252 1317 5459 1323
rect -35 1297 12 1303
rect 820 1297 1148 1303
rect 1156 1297 1164 1303
rect 1204 1297 1484 1303
rect 1748 1297 1756 1303
rect 1764 1297 1868 1303
rect 1876 1297 2076 1303
rect 2100 1297 2252 1303
rect 2276 1297 2284 1303
rect 2308 1297 2380 1303
rect 2420 1297 3036 1303
rect 3060 1297 3148 1303
rect 3236 1297 3276 1303
rect 3469 1297 4012 1303
rect 3469 1284 3475 1297
rect 4148 1297 4300 1303
rect 4452 1297 4492 1303
rect 4500 1297 4636 1303
rect 4644 1297 4796 1303
rect 4852 1297 4876 1303
rect 4900 1297 4988 1303
rect 4996 1297 5004 1303
rect 5188 1297 5228 1303
rect 5236 1297 5276 1303
rect 5453 1303 5459 1317
rect 5476 1317 5532 1323
rect 5588 1317 5692 1323
rect 6260 1317 6300 1323
rect 6388 1317 6412 1323
rect 6500 1317 6604 1323
rect 6612 1317 6796 1323
rect 6852 1317 6892 1323
rect 7028 1317 7068 1323
rect 7108 1317 7164 1323
rect 7284 1317 7340 1323
rect 7348 1317 7372 1323
rect 5453 1297 5916 1303
rect 6436 1297 6540 1303
rect 6548 1297 6684 1303
rect 6708 1297 6764 1303
rect 6772 1297 6876 1303
rect 6884 1297 7020 1303
rect 7124 1297 7260 1303
rect 372 1277 1084 1283
rect 1092 1277 3468 1283
rect 3556 1277 4716 1283
rect 4724 1277 5532 1283
rect 5860 1277 6204 1283
rect 6404 1277 6508 1283
rect 6596 1277 6924 1283
rect 740 1257 1267 1263
rect 1261 1244 1267 1257
rect 1764 1257 1772 1263
rect 1844 1257 3932 1263
rect 3940 1257 4076 1263
rect 4100 1257 4412 1263
rect 4676 1257 4828 1263
rect 4836 1257 5116 1263
rect 5156 1257 5420 1263
rect 6212 1257 6220 1263
rect 6404 1257 6412 1263
rect 6612 1257 6668 1263
rect 6740 1257 6908 1263
rect 116 1237 428 1243
rect 436 1237 1196 1243
rect 1268 1237 1404 1243
rect 1412 1237 1564 1243
rect 1572 1237 2364 1243
rect 2372 1237 3020 1243
rect 3044 1237 3628 1243
rect 3636 1237 3676 1243
rect 3940 1237 4268 1243
rect 4356 1237 4572 1243
rect 4596 1237 4844 1243
rect 4852 1237 5132 1243
rect 5204 1237 5308 1243
rect 5316 1237 5340 1243
rect 5716 1237 6028 1243
rect 6084 1237 6284 1243
rect 6733 1243 6739 1256
rect 6292 1237 6739 1243
rect 692 1217 1004 1223
rect 1012 1217 1292 1223
rect 1636 1217 1724 1223
rect 1748 1217 1772 1223
rect 1812 1217 1884 1223
rect 1988 1217 2012 1223
rect 2084 1217 2092 1223
rect 2260 1217 3644 1223
rect 3652 1217 3820 1223
rect 3997 1217 4172 1223
rect 1410 1214 1470 1216
rect 1410 1206 1411 1214
rect 1420 1206 1421 1214
rect 1459 1206 1460 1214
rect 1469 1206 1470 1214
rect 1410 1204 1470 1206
rect 868 1197 876 1203
rect 932 1197 1100 1203
rect 1140 1197 1388 1203
rect 1492 1197 2412 1203
rect 2436 1197 2444 1203
rect 2468 1197 2572 1203
rect 2596 1197 2668 1203
rect 2676 1197 2764 1203
rect 2804 1197 2812 1203
rect 2836 1197 2876 1203
rect 2900 1197 3100 1203
rect 3108 1197 3116 1203
rect 3188 1197 3372 1203
rect 3380 1197 3500 1203
rect 3540 1197 3564 1203
rect 3997 1203 4003 1217
rect 4564 1217 4764 1223
rect 4788 1217 4908 1223
rect 4932 1217 5260 1223
rect 5316 1217 6028 1223
rect 6484 1217 6860 1223
rect 4418 1214 4478 1216
rect 4418 1206 4419 1214
rect 4428 1206 4429 1214
rect 4467 1206 4468 1214
rect 4477 1206 4478 1214
rect 4418 1204 4478 1206
rect 3588 1197 4003 1203
rect 4020 1197 4172 1203
rect 4644 1197 4764 1203
rect 4948 1197 5052 1203
rect 5380 1197 6252 1203
rect 6612 1197 6620 1203
rect 356 1177 1580 1183
rect 1588 1177 2316 1183
rect 2324 1177 4204 1183
rect 4372 1177 4908 1183
rect 4916 1177 5084 1183
rect 5604 1177 5644 1183
rect 5700 1177 5836 1183
rect 6564 1177 6748 1183
rect 388 1157 1324 1163
rect 1348 1157 1500 1163
rect 1524 1157 1772 1163
rect 1780 1157 1996 1163
rect 2036 1157 2348 1163
rect 2356 1157 3340 1163
rect 3348 1157 4364 1163
rect 4644 1157 4684 1163
rect 4692 1157 4732 1163
rect 4756 1157 4972 1163
rect 5012 1157 5372 1163
rect 5469 1157 6156 1163
rect 772 1137 972 1143
rect 996 1137 1116 1143
rect 1140 1137 1212 1143
rect 1220 1137 1644 1143
rect 1652 1137 1852 1143
rect 1860 1137 1932 1143
rect 1972 1137 3372 1143
rect 3380 1137 3660 1143
rect 3668 1137 3788 1143
rect 4068 1137 4156 1143
rect 4164 1137 4236 1143
rect 4244 1137 4348 1143
rect 4388 1137 4428 1143
rect 4580 1137 4668 1143
rect 4676 1137 4716 1143
rect 5469 1143 5475 1157
rect 6548 1157 6604 1163
rect 6621 1157 6828 1163
rect 4948 1137 5475 1143
rect 5485 1137 5724 1143
rect 5485 1124 5491 1137
rect 6621 1143 6627 1157
rect 7188 1157 7308 1163
rect 6276 1137 6627 1143
rect 6644 1137 6780 1143
rect 228 1117 284 1123
rect 292 1117 348 1123
rect 484 1117 668 1123
rect 884 1117 940 1123
rect 964 1117 1004 1123
rect 1044 1117 1116 1123
rect 1140 1117 1148 1123
rect 1172 1117 1516 1123
rect 1540 1117 1692 1123
rect 1700 1117 2044 1123
rect 2068 1117 2188 1123
rect 2260 1117 2444 1123
rect 2484 1117 2492 1123
rect 2532 1117 2572 1123
rect 2580 1117 2636 1123
rect 2644 1117 2860 1123
rect 2868 1117 2972 1123
rect 2980 1117 3164 1123
rect 3236 1117 3308 1123
rect 3341 1117 3484 1123
rect 20 1097 300 1103
rect 308 1097 380 1103
rect 596 1097 700 1103
rect 708 1097 716 1103
rect 820 1097 892 1103
rect 916 1097 924 1103
rect 948 1097 1164 1103
rect 1236 1097 1292 1103
rect 1396 1097 1484 1103
rect 1492 1097 1564 1103
rect 1572 1097 1612 1103
rect 1716 1097 1804 1103
rect 1812 1097 1948 1103
rect 1956 1097 3132 1103
rect 3341 1103 3347 1117
rect 3620 1117 3628 1123
rect 3668 1117 3980 1123
rect 4004 1117 4028 1123
rect 4180 1117 4908 1123
rect 4916 1117 5468 1123
rect 5620 1117 5772 1123
rect 6244 1117 6300 1123
rect 6452 1117 6620 1123
rect 6628 1117 6892 1123
rect 7012 1117 7212 1123
rect 7332 1117 7356 1123
rect 3156 1097 3347 1103
rect 3380 1097 3404 1103
rect 3460 1097 3708 1103
rect 3764 1097 3884 1103
rect 3908 1097 3987 1103
rect 180 1077 236 1083
rect 292 1077 316 1083
rect 404 1077 508 1083
rect 516 1077 556 1083
rect 564 1077 636 1083
rect 724 1077 764 1083
rect 877 1077 1244 1083
rect 877 1064 883 1077
rect 1604 1077 1667 1083
rect 52 1057 108 1063
rect 276 1057 380 1063
rect 468 1057 652 1063
rect 660 1057 684 1063
rect 692 1057 876 1063
rect 996 1057 1036 1063
rect 1060 1057 1388 1063
rect 1540 1057 1612 1063
rect 1661 1063 1667 1077
rect 1684 1077 1836 1083
rect 1844 1077 1900 1083
rect 1940 1077 1996 1083
rect 2004 1077 2124 1083
rect 2132 1077 2940 1083
rect 2996 1077 3084 1083
rect 3092 1077 3436 1083
rect 3700 1077 3756 1083
rect 3764 1077 3964 1083
rect 3981 1083 3987 1097
rect 4052 1097 4140 1103
rect 4148 1097 4220 1103
rect 4340 1097 4412 1103
rect 4596 1097 4668 1103
rect 4676 1097 4684 1103
rect 4708 1097 4732 1103
rect 4980 1097 5100 1103
rect 5140 1097 5292 1103
rect 5405 1097 5436 1103
rect 3981 1077 4156 1083
rect 4221 1083 4227 1096
rect 4221 1077 4364 1083
rect 4372 1077 4588 1083
rect 4740 1077 4764 1083
rect 4772 1077 4972 1083
rect 5060 1077 5148 1083
rect 5156 1077 5196 1083
rect 5204 1077 5276 1083
rect 5405 1083 5411 1097
rect 5540 1097 5548 1103
rect 5588 1097 5756 1103
rect 5860 1097 6252 1103
rect 6308 1097 6940 1103
rect 6948 1097 7068 1103
rect 5364 1077 5411 1083
rect 5428 1077 5516 1083
rect 5524 1077 5564 1083
rect 5572 1077 5676 1083
rect 5684 1077 5820 1083
rect 5908 1077 6204 1083
rect 6228 1077 6428 1083
rect 6500 1077 6556 1083
rect 6596 1077 6636 1083
rect 6692 1077 6812 1083
rect 6884 1077 7020 1083
rect 1661 1057 1692 1063
rect 1748 1057 1756 1063
rect 1828 1057 1916 1063
rect 1940 1057 1948 1063
rect 1972 1057 1996 1063
rect 2052 1057 2252 1063
rect 2276 1057 2284 1063
rect 2308 1057 2412 1063
rect 2452 1057 2748 1063
rect 2772 1057 2812 1063
rect 2852 1057 3116 1063
rect 3204 1057 3228 1063
rect 3252 1057 3324 1063
rect 3348 1057 3388 1063
rect 3732 1057 4524 1063
rect 4548 1057 4620 1063
rect 4628 1057 4940 1063
rect 4964 1057 5116 1063
rect 5172 1057 5212 1063
rect 5476 1057 5580 1063
rect 5764 1057 6236 1063
rect 6484 1057 6524 1063
rect 6877 1063 6883 1076
rect 6532 1057 6883 1063
rect 7012 1057 7356 1063
rect 340 1037 492 1043
rect 548 1037 732 1043
rect 852 1037 1132 1043
rect 1204 1037 1340 1043
rect 1588 1037 2396 1043
rect 2404 1037 3580 1043
rect 3652 1037 3692 1043
rect 3748 1037 4332 1043
rect 4372 1037 6956 1043
rect 6964 1037 7276 1043
rect 493 1023 499 1036
rect 493 1017 588 1023
rect 596 1017 764 1023
rect 772 1017 1068 1023
rect 1076 1017 1292 1023
rect 1332 1017 2892 1023
rect 3028 1017 3052 1023
rect 3124 1017 3196 1023
rect 3204 1017 3276 1023
rect 3348 1017 3500 1023
rect 3892 1017 3900 1023
rect 4093 1017 4252 1023
rect 2914 1014 2974 1016
rect 2914 1006 2915 1014
rect 2924 1006 2925 1014
rect 2963 1006 2964 1014
rect 2973 1006 2974 1014
rect 2914 1004 2974 1006
rect 132 997 236 1003
rect 388 997 652 1003
rect 948 997 956 1003
rect 980 997 1260 1003
rect 1332 997 1548 1003
rect 1572 997 1900 1003
rect 1924 997 2044 1003
rect 2061 997 2300 1003
rect 420 977 556 983
rect 644 977 844 983
rect 1108 977 1132 983
rect 1380 977 1612 983
rect 2061 983 2067 997
rect 2324 997 2700 1003
rect 2717 997 2828 1003
rect 1748 977 2067 983
rect 2084 977 2092 983
rect 2228 977 2284 983
rect 2340 977 2476 983
rect 2500 977 2556 983
rect 2717 983 2723 997
rect 2852 997 2892 1003
rect 3028 997 3516 1003
rect 4093 1003 4099 1017
rect 4372 1017 4428 1023
rect 4532 1017 4748 1023
rect 5012 1017 5260 1023
rect 5380 1017 5532 1023
rect 5636 1017 5868 1023
rect 6100 1017 6236 1023
rect 6244 1017 6460 1023
rect 6612 1017 6716 1023
rect 6964 1017 6988 1023
rect 7044 1017 7084 1023
rect 5922 1014 5982 1016
rect 5922 1006 5923 1014
rect 5932 1006 5933 1014
rect 5971 1006 5972 1014
rect 5981 1006 5982 1014
rect 5922 1004 5982 1006
rect 3668 997 4099 1003
rect 4116 997 4172 1003
rect 4980 997 5260 1003
rect 5428 997 5452 1003
rect 5764 997 5884 1003
rect 5997 997 6876 1003
rect 2580 977 2723 983
rect 2740 977 2828 983
rect 2868 977 2924 983
rect 3236 977 3276 983
rect 3348 977 3548 983
rect 3812 977 3964 983
rect 4100 977 4124 983
rect 4148 977 4188 983
rect 4196 977 4284 983
rect 4500 977 4652 983
rect 4660 977 4668 983
rect 4852 977 5068 983
rect 5380 977 5468 983
rect 5492 977 5644 983
rect 5780 977 5804 983
rect 5812 977 5900 983
rect 5997 983 6003 997
rect 6980 997 7244 1003
rect 5924 977 6003 983
rect 6020 977 6220 983
rect 6388 977 6492 983
rect 6516 977 6988 983
rect 7204 977 7260 983
rect 132 957 332 963
rect 404 957 460 963
rect 468 957 508 963
rect 516 957 620 963
rect 628 957 716 963
rect 804 957 940 963
rect 948 957 1020 963
rect 1108 957 1164 963
rect 1172 957 1196 963
rect 1284 957 1500 963
rect 1556 957 1580 963
rect 1732 957 1900 963
rect 1940 957 2156 963
rect 2196 957 2252 963
rect 2276 957 2451 963
rect 116 937 204 943
rect 212 937 268 943
rect 724 937 796 943
rect 820 937 860 943
rect 1492 937 1564 943
rect 1572 937 1596 943
rect 1636 937 1971 943
rect 100 917 300 923
rect 388 917 428 923
rect 788 917 860 923
rect 1236 917 1292 923
rect 1316 917 1356 923
rect 1476 917 1820 923
rect 1860 917 1868 923
rect 1924 917 1948 923
rect 1965 923 1971 937
rect 1988 937 2108 943
rect 2164 937 2428 943
rect 2445 943 2451 957
rect 2468 957 2620 963
rect 2692 957 2716 963
rect 2724 957 2764 963
rect 2772 957 2860 963
rect 2900 957 3020 963
rect 3060 957 3260 963
rect 3268 957 3372 963
rect 3428 957 3532 963
rect 3636 957 3836 963
rect 3844 957 4028 963
rect 4036 957 4204 963
rect 4285 963 4291 976
rect 4285 957 4556 963
rect 4564 957 4572 963
rect 4948 957 5036 963
rect 5044 957 5100 963
rect 5268 957 5548 963
rect 5572 957 5932 963
rect 6132 957 6140 963
rect 6596 957 6604 963
rect 6612 957 6684 963
rect 7044 957 7164 963
rect 7252 957 7324 963
rect 2445 937 2892 943
rect 3012 937 3052 943
rect 3076 937 3148 943
rect 3364 937 3436 943
rect 3716 937 3756 943
rect 3780 937 3836 943
rect 3844 937 3900 943
rect 3908 937 4300 943
rect 4340 937 5324 943
rect 5364 937 5436 943
rect 5444 937 5500 943
rect 5588 937 5692 943
rect 5700 937 5772 943
rect 5828 937 5884 943
rect 5924 937 6076 943
rect 6164 937 6188 943
rect 6212 937 6252 943
rect 6260 937 6348 943
rect 6404 937 6652 943
rect 6660 937 6828 943
rect 6932 937 7036 943
rect 7060 937 7228 943
rect 7236 937 7340 943
rect 1965 917 2188 923
rect 2228 917 2380 923
rect 2420 917 2460 923
rect 2580 917 2588 923
rect 2612 917 2716 923
rect 2804 917 2844 923
rect 2868 917 3020 923
rect 3044 917 3084 923
rect 3156 917 3196 923
rect 3252 917 3708 923
rect 3764 917 3820 923
rect 3828 917 3884 923
rect 3892 917 4284 923
rect 4404 917 4524 923
rect 4900 917 4956 923
rect 5012 917 5068 923
rect 5092 917 5148 923
rect 5348 917 5452 923
rect 5476 917 5564 923
rect 5668 917 5724 923
rect 5780 917 5820 923
rect 5876 917 5900 923
rect 5908 917 6012 923
rect 6068 917 6092 923
rect 6180 917 6204 923
rect 6308 917 6380 923
rect 6436 917 6620 923
rect 6708 917 6764 923
rect 6948 917 7068 923
rect 7092 917 7148 923
rect 7220 917 7324 923
rect -35 897 12 903
rect 308 897 380 903
rect 1364 897 1532 903
rect 1796 897 1852 903
rect 1892 897 1900 903
rect 1908 897 1932 903
rect 2004 897 2300 903
rect 2324 897 2572 903
rect 2612 897 2636 903
rect 2708 897 2876 903
rect 2900 897 3324 903
rect 3348 897 3372 903
rect 3396 897 3596 903
rect 3764 897 3852 903
rect 3956 897 4124 903
rect 4148 897 4172 903
rect 4292 897 4748 903
rect 4772 897 4908 903
rect 4948 897 5020 903
rect 5140 897 5260 903
rect 5316 897 5404 903
rect 5748 897 5756 903
rect 6196 897 6268 903
rect 6532 897 6588 903
rect 6788 897 6844 903
rect 6884 897 6988 903
rect 7092 897 7228 903
rect 276 877 556 883
rect 820 877 1468 883
rect 1524 877 1868 883
rect 1876 877 2060 883
rect 2228 877 3180 883
rect 3412 877 3436 883
rect 3924 877 3996 883
rect 4621 877 4716 883
rect 532 857 1676 863
rect 1684 857 3244 863
rect 3357 857 3516 863
rect 756 837 1580 843
rect 1716 837 2124 843
rect 2212 837 2307 843
rect 820 817 1084 823
rect 1492 817 1740 823
rect 2301 823 2307 837
rect 2356 837 2620 843
rect 2660 837 2796 843
rect 2820 837 2860 843
rect 2900 837 2940 843
rect 3357 843 3363 857
rect 3524 857 3612 863
rect 4621 863 4627 877
rect 5748 877 6156 883
rect 6644 877 6764 883
rect 6788 877 6860 883
rect 6932 877 7196 883
rect 3828 857 4627 863
rect 4644 857 4860 863
rect 4996 857 5068 863
rect 5796 857 5820 863
rect 5860 857 6300 863
rect 6612 857 6668 863
rect 6676 857 6812 863
rect 6820 857 6876 863
rect 3012 837 3363 843
rect 3556 837 3724 843
rect 4004 837 4172 843
rect 4180 837 4236 843
rect 4637 843 4643 856
rect 4244 837 4643 843
rect 5172 837 5836 843
rect 5924 837 6044 843
rect 6148 837 6316 843
rect 6484 837 7308 843
rect 2301 817 3484 823
rect 3892 817 4364 823
rect 4500 817 4924 823
rect 5108 817 5228 823
rect 5236 817 5372 823
rect 5428 817 5468 823
rect 5812 817 5932 823
rect 5940 817 6172 823
rect 1410 814 1470 816
rect 1410 806 1411 814
rect 1420 806 1421 814
rect 1459 806 1460 814
rect 1469 806 1470 814
rect 1410 804 1470 806
rect 4418 814 4478 816
rect 4418 806 4419 814
rect 4428 806 4429 814
rect 4467 806 4468 814
rect 4477 806 4478 814
rect 4418 804 4478 806
rect 1012 797 1212 803
rect 1876 797 2316 803
rect 2452 797 2684 803
rect 2804 797 2908 803
rect 2916 797 3004 803
rect 3028 797 3036 803
rect 3204 797 3276 803
rect 3412 797 3644 803
rect 3892 797 4076 803
rect 4756 797 4876 803
rect 4900 797 5212 803
rect 5332 797 5388 803
rect 5396 797 5420 803
rect 5540 797 5916 803
rect 5940 797 6972 803
rect 1204 777 1804 783
rect 2084 777 2700 783
rect 2884 777 3427 783
rect 692 757 908 763
rect 1140 757 1180 763
rect 1245 757 2307 763
rect 132 737 204 743
rect 548 737 572 743
rect 580 737 748 743
rect 836 737 908 743
rect 916 737 924 743
rect 1245 743 1251 757
rect 1156 737 1251 743
rect 1268 737 1500 743
rect 1620 737 1852 743
rect 1860 737 1964 743
rect 2301 743 2307 757
rect 2324 757 2636 763
rect 2708 757 2828 763
rect 2836 757 3244 763
rect 3421 763 3427 777
rect 3444 777 5308 783
rect 5684 777 5996 783
rect 6004 777 6076 783
rect 6084 777 6124 783
rect 7076 777 7372 783
rect 3421 757 3452 763
rect 3700 757 4028 763
rect 4068 757 5452 763
rect 5588 757 5708 763
rect 5860 757 6364 763
rect 6724 757 6908 763
rect 6916 757 7100 763
rect 7108 757 7244 763
rect 2301 737 2412 743
rect 2436 737 2460 743
rect 2484 737 2620 743
rect 2644 737 2876 743
rect 2884 737 3020 743
rect 3028 737 3212 743
rect 3284 737 3644 743
rect 3652 737 3660 743
rect 4724 737 4812 743
rect 4932 737 5276 743
rect 5332 737 5564 743
rect 5652 737 6460 743
rect 7060 737 7132 743
rect 7236 737 7276 743
rect 68 717 268 723
rect 404 717 460 723
rect 500 717 636 723
rect 749 717 1164 723
rect 749 704 755 717
rect 1613 723 1619 736
rect 1220 717 1619 723
rect 1716 717 1980 723
rect 2180 717 2204 723
rect 2212 717 2252 723
rect 2260 717 2540 723
rect 2548 717 3052 723
rect 3108 717 3292 723
rect 3300 717 3356 723
rect 3396 717 3484 723
rect 3572 717 3692 723
rect 3924 717 3996 723
rect 4052 717 4508 723
rect 4612 717 4819 723
rect 52 697 124 703
rect 292 697 412 703
rect 628 697 668 703
rect 740 697 748 703
rect 900 697 908 703
rect 1028 697 1084 703
rect 1156 697 1196 703
rect 1204 697 1244 703
rect 1252 697 1308 703
rect 1428 697 1516 703
rect 1668 697 1756 703
rect 1764 697 1836 703
rect 1892 697 1900 703
rect 1908 697 1948 703
rect 2068 697 2140 703
rect 2292 697 2316 703
rect 2324 697 2396 703
rect 2420 697 2476 703
rect 2500 697 2572 703
rect 2612 697 2668 703
rect 2676 697 2844 703
rect 2852 697 3004 703
rect 3156 697 3196 703
rect 3300 697 3420 703
rect 3828 697 3916 703
rect 4180 697 4236 703
rect 4692 697 4700 703
rect 4708 697 4796 703
rect 4813 703 4819 717
rect 4852 717 4876 723
rect 4884 717 4988 723
rect 5044 717 5228 723
rect 5236 717 5340 723
rect 5492 717 5548 723
rect 5652 717 5756 723
rect 6020 717 6284 723
rect 6500 717 6540 723
rect 6580 717 6700 723
rect 6900 717 6956 723
rect 6964 717 7116 723
rect 7124 717 7132 723
rect 7140 717 7196 723
rect 4813 697 4844 703
rect 4964 697 5100 703
rect 5284 697 5404 703
rect 5444 697 5516 703
rect 5572 697 5612 703
rect 5620 697 5692 703
rect 5700 697 5804 703
rect 5812 697 5884 703
rect 6036 697 6204 703
rect 6452 697 6604 703
rect 6820 697 6828 703
rect 6836 697 6860 703
rect 7076 697 7084 703
rect 452 677 556 683
rect 1885 683 1891 696
rect 1044 677 1891 683
rect 2036 677 2204 683
rect 2436 677 2524 683
rect 2644 677 2684 683
rect 2724 677 2883 683
rect 116 657 188 663
rect 324 657 364 663
rect 388 657 444 663
rect 564 657 636 663
rect 852 657 892 663
rect 1076 657 1116 663
rect 1140 657 1180 663
rect 1364 657 1548 663
rect 1892 657 2012 663
rect 2068 657 2092 663
rect 2196 657 2236 663
rect 2244 657 2284 663
rect 2388 657 2444 663
rect 2452 657 2508 663
rect 2516 657 2604 663
rect 2685 663 2691 676
rect 2685 657 2796 663
rect 2877 663 2883 677
rect 2900 677 3084 683
rect 3108 677 3116 683
rect 3236 677 3276 683
rect 3284 677 3308 683
rect 3348 677 3372 683
rect 3412 677 3452 683
rect 3764 677 3932 683
rect 3972 677 4044 683
rect 4084 677 4124 683
rect 4132 677 4252 683
rect 4260 677 4284 683
rect 4548 677 5068 683
rect 5268 677 5292 683
rect 5604 677 5660 683
rect 5732 677 5868 683
rect 6340 677 6380 683
rect 6388 677 6508 683
rect 6516 677 6588 683
rect 7108 677 7324 683
rect 2877 657 2940 663
rect 3316 657 3452 663
rect 3460 657 3468 663
rect 3476 657 3587 663
rect 148 637 364 643
rect 436 637 620 643
rect 628 637 700 643
rect 788 637 1340 643
rect 1348 637 1436 643
rect 2100 637 3404 643
rect 3492 637 3564 643
rect 3581 643 3587 657
rect 3668 657 3676 663
rect 3860 657 3884 663
rect 3892 657 3964 663
rect 4708 657 4972 663
rect 5412 657 5500 663
rect 5556 657 5932 663
rect 6004 657 6124 663
rect 6132 657 6156 663
rect 6164 657 6268 663
rect 6276 657 6572 663
rect 6772 657 6780 663
rect 6788 657 6828 663
rect 6852 657 6924 663
rect 7012 657 7036 663
rect 7124 657 7148 663
rect 7156 657 7276 663
rect 3581 637 3676 643
rect 3828 637 3916 643
rect 3940 637 4188 643
rect 5316 637 5420 643
rect 5501 637 6748 643
rect 340 617 716 623
rect 1012 617 1324 623
rect 1572 617 2876 623
rect 3012 617 3116 623
rect 3268 617 3388 623
rect 4596 617 4620 623
rect 5501 623 5507 637
rect 6756 637 6876 643
rect 6884 637 6972 643
rect 7044 637 7196 643
rect 7300 637 7340 643
rect 5268 617 5507 623
rect 5620 617 5715 623
rect 2914 614 2974 616
rect 2914 606 2915 614
rect 2924 606 2925 614
rect 2963 606 2964 614
rect 2973 606 2974 614
rect 2914 604 2974 606
rect 1060 597 1132 603
rect 1348 597 1468 603
rect 1604 597 2659 603
rect 164 577 252 583
rect 260 577 300 583
rect 532 577 556 583
rect 740 577 780 583
rect 2100 577 2300 583
rect 2340 577 2572 583
rect 2653 583 2659 597
rect 2676 597 2732 603
rect 2861 597 2892 603
rect 2861 583 2867 597
rect 3069 597 3756 603
rect 2653 577 2867 583
rect 3069 583 3075 597
rect 3892 597 3916 603
rect 4804 597 4828 603
rect 5076 597 5468 603
rect 5508 597 5692 603
rect 5709 603 5715 617
rect 5796 617 5820 623
rect 5844 617 5900 623
rect 6500 617 6652 623
rect 5922 614 5982 616
rect 5922 606 5923 614
rect 5932 606 5933 614
rect 5971 606 5972 614
rect 5981 606 5982 614
rect 5922 604 5982 606
rect 5709 597 5836 603
rect 6004 597 6131 603
rect 2884 577 3075 583
rect 3092 577 3772 583
rect 3860 577 4076 583
rect 4612 577 4876 583
rect 5012 577 5276 583
rect 5284 577 5532 583
rect 5652 577 5804 583
rect 5828 577 6108 583
rect 6125 583 6131 597
rect 6420 597 6428 603
rect 6580 597 6684 603
rect 6692 597 6700 603
rect 6708 597 7052 603
rect 6125 577 6620 583
rect 6660 577 7004 583
rect 7044 577 7084 583
rect 7092 577 7260 583
rect 324 557 412 563
rect 420 557 524 563
rect 644 557 700 563
rect 708 557 924 563
rect 932 557 1100 563
rect 1300 557 1372 563
rect 1380 557 1612 563
rect 1620 557 1644 563
rect 1972 557 2044 563
rect 2148 557 2364 563
rect 2436 557 2508 563
rect 2532 557 2620 563
rect 2628 557 2684 563
rect 2692 557 2748 563
rect 2820 557 2876 563
rect 3092 557 3132 563
rect 3188 557 3276 563
rect 3284 557 3324 563
rect 3380 557 3436 563
rect 3444 557 3708 563
rect 3716 557 3868 563
rect 3876 557 4140 563
rect 4820 557 4844 563
rect 4852 557 4940 563
rect 5412 557 5660 563
rect 5668 557 5676 563
rect 5684 557 5772 563
rect 5828 557 5868 563
rect 5885 557 5996 563
rect 269 537 572 543
rect 52 517 172 523
rect 269 523 275 537
rect 772 537 892 543
rect 948 537 1004 543
rect 1140 537 1196 543
rect 1204 537 1340 543
rect 1444 537 1516 543
rect 1524 537 1628 543
rect 2292 537 2316 543
rect 2324 537 2444 543
rect 2516 537 2748 543
rect 2756 537 2844 543
rect 3012 537 3068 543
rect 3124 537 3196 543
rect 3284 537 3356 543
rect 3492 537 3580 543
rect 3796 537 3836 543
rect 4244 537 4300 543
rect 4324 537 4364 543
rect 4500 537 4572 543
rect 4676 537 4716 543
rect 5108 537 5196 543
rect 5204 537 5228 543
rect 5236 537 5308 543
rect 5316 537 5452 543
rect 5460 537 5596 543
rect 5885 543 5891 557
rect 6084 557 6140 563
rect 6196 557 6236 563
rect 6548 557 6716 563
rect 6772 557 6956 563
rect 5780 537 5891 543
rect 5956 537 6092 543
rect 6100 537 6204 543
rect 6276 537 6476 543
rect 6708 537 6860 543
rect 7092 537 7100 543
rect 7140 537 7180 543
rect 228 517 275 523
rect 292 517 332 523
rect 612 517 796 523
rect 916 517 940 523
rect 1092 517 1228 523
rect 1348 517 1372 523
rect 1508 517 1564 523
rect 1908 517 2076 523
rect 2132 517 2172 523
rect 2196 517 2220 523
rect 2356 517 2428 523
rect 2532 517 2588 523
rect 2612 517 2636 523
rect 2788 517 3276 523
rect 3316 517 3356 523
rect 3412 517 3548 523
rect 3556 517 3612 523
rect 3636 517 3740 523
rect 3812 517 3884 523
rect 4004 517 4204 523
rect 4292 517 4508 523
rect 4708 517 4748 523
rect 4772 517 4892 523
rect 5028 517 5292 523
rect 5380 517 5484 523
rect 5508 517 5532 523
rect 5684 517 5756 523
rect 5764 517 5900 523
rect 5908 517 6156 523
rect 6164 517 6380 523
rect 6660 517 6716 523
rect 6948 517 6988 523
rect 7060 517 7292 523
rect 196 497 380 503
rect 404 497 556 503
rect 1140 497 1244 503
rect 1252 497 1292 503
rect 1300 497 1548 503
rect 1556 497 1708 503
rect 1716 497 1740 503
rect 1748 497 1788 503
rect 1796 497 1852 503
rect 2308 497 2556 503
rect 2836 497 3052 503
rect 3140 497 3180 503
rect 3476 497 3516 503
rect 4628 497 4652 503
rect 4756 497 4780 503
rect 4820 497 4876 503
rect 5476 497 5500 503
rect 5524 497 5580 503
rect 5716 497 5772 503
rect 5812 497 5868 503
rect 5876 497 6060 503
rect 6100 497 6492 503
rect 6996 497 7084 503
rect 132 477 348 483
rect 356 477 428 483
rect 1044 477 1132 483
rect 1220 477 1484 483
rect 2868 477 3116 483
rect 3540 477 3644 483
rect 3652 477 3676 483
rect 4260 477 6780 483
rect 6996 477 7020 483
rect 7028 477 7068 483
rect 7108 477 7132 483
rect 596 457 1724 463
rect 2004 457 2300 463
rect 2612 457 2652 463
rect 2660 457 2796 463
rect 2804 457 2988 463
rect 2996 457 3164 463
rect 4308 457 5260 463
rect 5300 457 5628 463
rect 5652 457 6028 463
rect 6068 457 6956 463
rect 916 437 1004 443
rect 1204 437 1580 443
rect 2500 437 2540 443
rect 2548 437 3164 443
rect 3172 437 3180 443
rect 3540 437 3884 443
rect 4132 437 4348 443
rect 4564 437 5308 443
rect 5604 437 5772 443
rect 5821 437 6163 443
rect 1492 417 1612 423
rect 1620 417 1804 423
rect 1812 417 1836 423
rect 2100 417 3532 423
rect 4708 417 4716 423
rect 5172 417 5708 423
rect 5821 423 5827 437
rect 5748 417 5827 423
rect 5844 417 6060 423
rect 6157 423 6163 437
rect 6180 437 6492 443
rect 6740 437 6780 443
rect 7012 437 7180 443
rect 6157 417 6220 423
rect 6676 417 6748 423
rect 1410 414 1470 416
rect 1410 406 1411 414
rect 1420 406 1421 414
rect 1459 406 1460 414
rect 1469 406 1470 414
rect 1410 404 1470 406
rect 4418 414 4478 416
rect 4418 406 4419 414
rect 4428 406 4429 414
rect 4467 406 4468 414
rect 4477 406 4478 414
rect 4418 404 4478 406
rect 3700 397 3836 403
rect 3860 397 3916 403
rect 4068 397 4108 403
rect 4708 397 4732 403
rect 4740 397 5260 403
rect 5364 397 5644 403
rect 5812 397 7020 403
rect 788 377 908 383
rect 916 377 1260 383
rect 1268 377 1548 383
rect 1556 377 2028 383
rect 2036 377 2332 383
rect 3668 377 4156 383
rect 4756 377 4796 383
rect 4868 377 5020 383
rect 5028 377 5100 383
rect 5613 377 5820 383
rect 5613 364 5619 377
rect 5988 377 6140 383
rect 6164 377 6188 383
rect 6212 377 6316 383
rect 6372 377 6524 383
rect 6532 377 6876 383
rect 340 357 508 363
rect 996 357 1148 363
rect 1924 357 1980 363
rect 3588 357 3644 363
rect 3668 357 3900 363
rect 4244 357 4268 363
rect 4772 357 4972 363
rect 5492 357 5612 363
rect 5668 357 6012 363
rect 6020 357 6252 363
rect 6260 357 6284 363
rect 6292 357 6316 363
rect 6324 357 6412 363
rect 6500 357 6764 363
rect 1028 337 1084 343
rect 1444 337 1692 343
rect 1956 337 1964 343
rect 2084 337 2092 343
rect 2900 337 3036 343
rect 3044 337 3260 343
rect 3405 337 5116 343
rect 3405 324 3411 337
rect 5252 337 5388 343
rect 5476 337 5548 343
rect 5748 337 5859 343
rect 132 317 348 323
rect 388 317 508 323
rect 1012 317 1420 323
rect 1428 317 2156 323
rect 2164 317 2172 323
rect 2196 317 2284 323
rect 3220 317 3404 323
rect 3444 317 3468 323
rect 3524 317 3580 323
rect 3700 317 3820 323
rect 3828 317 3948 323
rect 3956 317 4348 323
rect 4372 317 4428 323
rect 4676 317 4828 323
rect 4836 317 4876 323
rect 5540 317 5548 323
rect 5732 317 5772 323
rect 5853 323 5859 337
rect 5876 337 6019 343
rect 5853 317 5996 323
rect 6013 323 6019 337
rect 6164 337 6220 343
rect 6228 337 6572 343
rect 6804 337 6860 343
rect 6996 337 7036 343
rect 6013 317 6028 323
rect 6052 317 6124 323
rect 6132 317 6172 323
rect 6484 317 6684 323
rect 6788 317 7276 323
rect 7284 317 7292 323
rect 84 297 92 303
rect 356 297 428 303
rect 484 297 684 303
rect 948 297 1052 303
rect 1060 297 1388 303
rect 1396 297 2220 303
rect 2820 297 2844 303
rect 2852 297 2876 303
rect 2884 297 3052 303
rect 3092 297 3180 303
rect 3268 297 3308 303
rect 3348 297 3452 303
rect 3668 297 5196 303
rect 5204 297 5324 303
rect 5588 297 5660 303
rect 5700 297 5836 303
rect 5844 297 6044 303
rect 6388 297 6508 303
rect 6836 297 6924 303
rect 6996 297 7164 303
rect 68 277 108 283
rect 116 277 172 283
rect 228 277 332 283
rect 340 277 396 283
rect 452 277 492 283
rect 532 277 604 283
rect 612 277 700 283
rect 836 277 860 283
rect 868 277 1068 283
rect 1300 277 1388 283
rect 1524 277 1996 283
rect 2052 277 2076 283
rect 2164 277 2204 283
rect 2788 277 2828 283
rect 2836 277 2892 283
rect 3188 277 3212 283
rect 3300 277 3500 283
rect 3636 277 3708 283
rect 3732 277 3900 283
rect 3956 277 3980 283
rect 3988 277 4172 283
rect 4180 277 4252 283
rect 4260 277 4268 283
rect 4308 277 4396 283
rect 4404 277 4476 283
rect 4564 277 4716 283
rect 4772 277 4796 283
rect 4996 277 5276 283
rect 5348 277 5388 283
rect 5748 277 5884 283
rect 5892 277 6092 283
rect 6132 277 6204 283
rect 6356 277 6396 283
rect 6404 277 6556 283
rect 6644 277 6876 283
rect 7012 277 7036 283
rect 7044 277 7068 283
rect 7092 277 7116 283
rect 7140 277 7180 283
rect 7188 277 7276 283
rect 212 257 444 263
rect 580 257 620 263
rect 628 257 796 263
rect 804 257 828 263
rect 884 257 956 263
rect 996 257 1036 263
rect 1076 257 1116 263
rect 1332 257 1676 263
rect 1828 257 1916 263
rect 1924 257 1980 263
rect 2020 257 2124 263
rect 2308 257 2572 263
rect 2676 257 3004 263
rect 3108 257 3132 263
rect 3140 257 3260 263
rect 3268 257 3372 263
rect 3588 257 3772 263
rect 3780 257 3852 263
rect 4212 257 4236 263
rect 4244 257 4284 263
rect 4372 257 4412 263
rect 4548 257 4636 263
rect 4660 257 4764 263
rect 4772 257 4844 263
rect 5341 263 5347 276
rect 5268 257 5468 263
rect 5492 257 5756 263
rect 5764 257 5804 263
rect 5812 257 5996 263
rect 6036 257 6156 263
rect 6196 257 6284 263
rect 6292 257 6380 263
rect 6468 257 6588 263
rect 6708 257 7228 263
rect 84 237 476 243
rect 500 237 604 243
rect 660 237 988 243
rect 1172 237 1548 243
rect 1940 237 2012 243
rect 2388 237 2460 243
rect 2468 237 2540 243
rect 2660 237 2700 243
rect 2868 237 3100 243
rect 4100 237 4204 243
rect 4244 237 4332 243
rect 4612 237 4668 243
rect 5044 237 5676 243
rect 5700 237 6108 243
rect 6116 237 6396 243
rect 6404 237 6620 243
rect 6628 237 6652 243
rect 6660 237 6700 243
rect 20 217 204 223
rect 324 217 444 223
rect 653 223 659 236
rect 564 217 659 223
rect 948 217 972 223
rect 2612 217 2716 223
rect 3460 217 4828 223
rect 4836 217 5596 223
rect 5668 217 5900 223
rect 6116 217 6188 223
rect 6436 217 6716 223
rect 6724 217 6748 223
rect 6756 217 6796 223
rect 2914 214 2974 216
rect 2914 206 2915 214
rect 2924 206 2925 214
rect 2963 206 2964 214
rect 2973 206 2974 214
rect 2914 204 2974 206
rect 5922 214 5982 216
rect 5922 206 5923 214
rect 5932 206 5933 214
rect 5971 206 5972 214
rect 5981 206 5982 214
rect 5922 204 5982 206
rect 93 197 284 203
rect 93 184 99 197
rect 404 197 748 203
rect 788 197 1027 203
rect 68 177 92 183
rect 276 177 492 183
rect 500 177 572 183
rect 708 177 892 183
rect 900 177 940 183
rect 1021 183 1027 197
rect 1044 197 2108 203
rect 2180 197 2627 203
rect 1021 177 1196 183
rect 1700 177 1868 183
rect 2100 177 2204 183
rect 2420 177 2508 183
rect 2564 177 2604 183
rect 2621 183 2627 197
rect 2804 197 2892 203
rect 4292 197 4364 203
rect 5204 197 5404 203
rect 5460 197 5612 203
rect 5748 197 5772 203
rect 6004 197 6124 203
rect 6141 197 6508 203
rect 2621 177 2924 183
rect 3188 177 3356 183
rect 3364 177 3660 183
rect 3876 177 4755 183
rect 4749 164 4755 177
rect 4932 177 5644 183
rect 5684 177 5868 183
rect 6141 183 6147 197
rect 6516 197 6972 203
rect 6980 197 7052 203
rect 5908 177 6147 183
rect 6180 177 6188 183
rect 6212 177 6691 183
rect 180 157 204 163
rect 324 157 364 163
rect 484 157 620 163
rect 644 157 764 163
rect 1236 157 1372 163
rect 1572 157 1644 163
rect 1764 157 2108 163
rect 2116 157 2396 163
rect 2436 157 2588 163
rect 2628 157 2652 163
rect 2724 157 2828 163
rect 2948 157 3244 163
rect 3268 157 3276 163
rect 3284 157 3340 163
rect 3348 157 3484 163
rect 3700 157 4076 163
rect 4756 157 5356 163
rect 5412 157 5484 163
rect 5508 157 5676 163
rect 5972 157 6300 163
rect 6548 157 6604 163
rect 6685 163 6691 177
rect 6772 177 6892 183
rect 6900 177 7020 183
rect 7076 177 7116 183
rect 6685 157 6732 163
rect 7172 157 7388 163
rect 68 137 268 143
rect 292 137 332 143
rect 436 137 524 143
rect 756 137 1052 143
rect 1108 137 1244 143
rect 1396 137 1532 143
rect 1636 137 1820 143
rect 2340 137 2476 143
rect 2596 137 2636 143
rect 2653 143 2659 156
rect 2653 137 2732 143
rect 3060 137 3132 143
rect 3316 137 3436 143
rect 3860 137 3884 143
rect 4116 137 4380 143
rect 4388 137 4572 143
rect 4804 137 4876 143
rect 4884 137 4940 143
rect 4948 137 5004 143
rect 5012 137 5164 143
rect 5284 137 5443 143
rect 628 117 668 123
rect 676 117 716 123
rect 1076 117 1132 123
rect 1140 117 1276 123
rect 1284 117 1516 123
rect 1668 117 1868 123
rect 1876 117 1964 123
rect 1972 117 2012 123
rect 2148 117 2268 123
rect 2292 117 2524 123
rect 2532 117 2620 123
rect 2628 117 2716 123
rect 2916 117 3020 123
rect 3028 117 3324 123
rect 3668 117 3756 123
rect 3844 117 3868 123
rect 3940 117 4140 123
rect 4196 117 4252 123
rect 4260 117 4348 123
rect 4980 117 5004 123
rect 5380 117 5420 123
rect 5437 123 5443 137
rect 5540 137 5596 143
rect 5620 137 6748 143
rect 6788 137 6988 143
rect 6996 137 7356 143
rect 5437 117 6412 123
rect 6484 117 6668 123
rect 6676 117 6844 123
rect 6884 117 6908 123
rect 7060 117 7084 123
rect 7108 117 7148 123
rect -35 97 12 103
rect 564 97 652 103
rect 692 97 1724 103
rect 2324 97 2348 103
rect 2372 97 2444 103
rect 2452 97 2476 103
rect 2564 97 2636 103
rect 2644 97 3068 103
rect 3140 97 3212 103
rect 3316 97 3356 103
rect 3860 97 3884 103
rect 4084 97 4156 103
rect 4820 97 4956 103
rect 5940 97 6012 103
rect 6084 97 6188 103
rect 6228 97 6268 103
rect 6644 97 6700 103
rect 6884 97 6956 103
rect 6964 97 7148 103
rect 7156 97 7260 103
rect 1780 77 2540 83
rect 5892 77 6172 83
rect 6212 77 6428 83
rect 6756 77 6908 83
rect 6932 77 7100 83
rect 3812 57 3836 63
rect 4068 37 4092 43
rect 4052 17 4060 23
rect 4244 17 4252 23
rect 4756 17 4780 23
rect 4996 17 5068 23
rect 1410 14 1470 16
rect 1410 6 1411 14
rect 1420 6 1421 14
rect 1459 6 1460 14
rect 1469 6 1470 14
rect 1410 4 1470 6
rect 4418 14 4478 16
rect 4418 6 4419 14
rect 4428 6 4429 14
rect 4467 6 4468 14
rect 4477 6 4478 14
rect 4418 4 4478 6
<< m4contact >>
rect 2916 5406 2923 5414
rect 2923 5406 2924 5414
rect 2928 5406 2933 5414
rect 2933 5406 2935 5414
rect 2935 5406 2936 5414
rect 2940 5406 2943 5414
rect 2943 5406 2945 5414
rect 2945 5406 2948 5414
rect 2952 5406 2953 5414
rect 2953 5406 2955 5414
rect 2955 5406 2960 5414
rect 2964 5406 2965 5414
rect 2965 5406 2972 5414
rect 5924 5406 5931 5414
rect 5931 5406 5932 5414
rect 5936 5406 5941 5414
rect 5941 5406 5943 5414
rect 5943 5406 5944 5414
rect 5948 5406 5951 5414
rect 5951 5406 5953 5414
rect 5953 5406 5956 5414
rect 5960 5406 5961 5414
rect 5961 5406 5963 5414
rect 5963 5406 5968 5414
rect 5972 5406 5973 5414
rect 5973 5406 5980 5414
rect 7340 5396 7348 5404
rect 6988 5376 6996 5384
rect 4108 5336 4116 5344
rect 7308 5336 7316 5344
rect 5132 5316 5140 5324
rect 6412 5316 6420 5324
rect 972 5296 980 5304
rect 1580 5296 1588 5304
rect 3980 5296 3988 5304
rect 5292 5296 5300 5304
rect 6604 5296 6612 5304
rect 7244 5276 7252 5284
rect 268 5256 276 5264
rect 4940 5256 4948 5264
rect 6124 5256 6132 5264
rect 6220 5256 6228 5264
rect 6444 5256 6452 5264
rect 1324 5216 1332 5224
rect 1412 5206 1419 5214
rect 1419 5206 1420 5214
rect 1424 5206 1429 5214
rect 1429 5206 1431 5214
rect 1431 5206 1432 5214
rect 1436 5206 1439 5214
rect 1439 5206 1441 5214
rect 1441 5206 1444 5214
rect 1448 5206 1449 5214
rect 1449 5206 1451 5214
rect 1451 5206 1456 5214
rect 1460 5206 1461 5214
rect 1461 5206 1468 5214
rect 4420 5206 4427 5214
rect 4427 5206 4428 5214
rect 4432 5206 4437 5214
rect 4437 5206 4439 5214
rect 4439 5206 4440 5214
rect 4444 5206 4447 5214
rect 4447 5206 4449 5214
rect 4449 5206 4452 5214
rect 4456 5206 4457 5214
rect 4457 5206 4459 5214
rect 4459 5206 4464 5214
rect 4468 5206 4469 5214
rect 4469 5206 4476 5214
rect 1580 5196 1588 5204
rect 4236 5196 4244 5204
rect 5772 5196 5780 5204
rect 6092 5196 6100 5204
rect 6124 5196 6132 5204
rect 6892 5196 6900 5204
rect 2060 5156 2068 5164
rect 3468 5156 3476 5164
rect 3756 5156 3764 5164
rect 6700 5156 6708 5164
rect 6732 5156 6740 5164
rect 1644 5136 1652 5144
rect 3948 5136 3956 5144
rect 764 5116 772 5124
rect 3468 5116 3476 5124
rect 3820 5116 3828 5124
rect 812 5096 820 5104
rect 1868 5096 1876 5104
rect 1964 5096 1972 5104
rect 3148 5096 3156 5104
rect 3372 5096 3380 5104
rect 3436 5096 3444 5104
rect 3724 5096 3732 5104
rect 4044 5096 4052 5104
rect 5420 5096 5428 5104
rect 6060 5096 6068 5104
rect 1804 5076 1812 5084
rect 1740 5056 1748 5064
rect 2028 5076 2036 5084
rect 268 5016 276 5024
rect 972 5016 980 5024
rect 1996 5036 2004 5044
rect 3660 5076 3668 5084
rect 4684 5076 4692 5084
rect 6188 5076 6196 5084
rect 6636 5076 6644 5084
rect 3500 5056 3508 5064
rect 4908 5056 4916 5064
rect 4716 5036 4724 5044
rect 1740 5016 1748 5024
rect 6828 5036 6836 5044
rect 2916 5006 2923 5014
rect 2923 5006 2924 5014
rect 2928 5006 2933 5014
rect 2933 5006 2935 5014
rect 2935 5006 2936 5014
rect 2940 5006 2943 5014
rect 2943 5006 2945 5014
rect 2945 5006 2948 5014
rect 2952 5006 2953 5014
rect 2953 5006 2955 5014
rect 2955 5006 2960 5014
rect 2964 5006 2965 5014
rect 2965 5006 2972 5014
rect 5924 5006 5931 5014
rect 5931 5006 5932 5014
rect 5936 5006 5941 5014
rect 5941 5006 5943 5014
rect 5943 5006 5944 5014
rect 5948 5006 5951 5014
rect 5951 5006 5953 5014
rect 5953 5006 5956 5014
rect 5960 5006 5961 5014
rect 5961 5006 5963 5014
rect 5963 5006 5968 5014
rect 5972 5006 5973 5014
rect 5973 5006 5980 5014
rect 3180 4996 3188 5004
rect 3820 4996 3828 5004
rect 4108 4996 4116 5004
rect 5132 4996 5140 5004
rect 6540 4996 6548 5004
rect 1036 4976 1044 4984
rect 1644 4976 1652 4984
rect 2508 4956 2516 4964
rect 3756 4956 3764 4964
rect 3948 4956 3956 4964
rect 3980 4956 3988 4964
rect 4716 4956 4724 4964
rect 1036 4936 1044 4944
rect 2316 4936 2324 4944
rect 2444 4936 2452 4944
rect 5100 4936 5108 4944
rect 6668 4976 6676 4984
rect 7052 4976 7060 4984
rect 6156 4956 6164 4964
rect 6540 4956 6548 4964
rect 3180 4916 3188 4924
rect 5004 4916 5012 4924
rect 5484 4916 5492 4924
rect 6060 4936 6068 4944
rect 6156 4916 6164 4924
rect 6540 4916 6548 4924
rect 1804 4896 1812 4904
rect 3372 4896 3380 4904
rect 1196 4876 1204 4884
rect 3660 4896 3668 4904
rect 5068 4896 5076 4904
rect 1996 4856 2004 4864
rect 5420 4856 5428 4864
rect 7180 4876 7188 4884
rect 3372 4836 3380 4844
rect 5004 4836 5012 4844
rect 5868 4836 5876 4844
rect 1412 4806 1419 4814
rect 1419 4806 1420 4814
rect 1424 4806 1429 4814
rect 1429 4806 1431 4814
rect 1431 4806 1432 4814
rect 1436 4806 1439 4814
rect 1439 4806 1441 4814
rect 1441 4806 1444 4814
rect 1448 4806 1449 4814
rect 1449 4806 1451 4814
rect 1451 4806 1456 4814
rect 1460 4806 1461 4814
rect 1461 4806 1468 4814
rect 4420 4806 4427 4814
rect 4427 4806 4428 4814
rect 4432 4806 4437 4814
rect 4437 4806 4439 4814
rect 4439 4806 4440 4814
rect 4444 4806 4447 4814
rect 4447 4806 4449 4814
rect 4449 4806 4452 4814
rect 4456 4806 4457 4814
rect 4457 4806 4459 4814
rect 4459 4806 4464 4814
rect 4468 4806 4469 4814
rect 4469 4806 4476 4814
rect 1964 4796 1972 4804
rect 2764 4796 2772 4804
rect 4044 4776 4052 4784
rect 4108 4776 4116 4784
rect 4908 4796 4916 4804
rect 6956 4796 6964 4804
rect 5132 4776 5140 4784
rect 6028 4776 6036 4784
rect 2764 4756 2772 4764
rect 1260 4736 1268 4744
rect 2028 4736 2036 4744
rect 2188 4736 2196 4744
rect 5004 4756 5012 4764
rect 7084 4756 7092 4764
rect 5324 4736 5332 4744
rect 7148 4736 7156 4744
rect 2156 4716 2164 4724
rect 300 4696 308 4704
rect 1996 4696 2004 4704
rect 5100 4696 5108 4704
rect 5836 4696 5844 4704
rect 6188 4716 6196 4724
rect 6572 4716 6580 4724
rect 7276 4716 7284 4724
rect 6252 4696 6260 4704
rect 6668 4696 6676 4704
rect 6764 4696 6772 4704
rect 7116 4696 7124 4704
rect 1612 4676 1620 4684
rect 2156 4676 2164 4684
rect 4076 4676 4084 4684
rect 4236 4676 4244 4684
rect 4748 4676 4756 4684
rect 4876 4676 4884 4684
rect 4908 4676 4916 4684
rect 1804 4636 1812 4644
rect 1996 4656 2004 4664
rect 5004 4656 5012 4664
rect 5196 4676 5204 4684
rect 5292 4676 5300 4684
rect 5324 4656 5332 4664
rect 6188 4656 6196 4664
rect 6220 4656 6228 4664
rect 6636 4656 6644 4664
rect 6700 4656 6708 4664
rect 588 4616 596 4624
rect 1868 4616 1876 4624
rect 6412 4616 6420 4624
rect 6988 4616 6996 4624
rect 7212 4616 7220 4624
rect 2916 4606 2923 4614
rect 2923 4606 2924 4614
rect 2928 4606 2933 4614
rect 2933 4606 2935 4614
rect 2935 4606 2936 4614
rect 2940 4606 2943 4614
rect 2943 4606 2945 4614
rect 2945 4606 2948 4614
rect 2952 4606 2953 4614
rect 2953 4606 2955 4614
rect 2955 4606 2960 4614
rect 2964 4606 2965 4614
rect 2965 4606 2972 4614
rect 5924 4606 5931 4614
rect 5931 4606 5932 4614
rect 5936 4606 5941 4614
rect 5941 4606 5943 4614
rect 5943 4606 5944 4614
rect 5948 4606 5951 4614
rect 5951 4606 5953 4614
rect 5953 4606 5956 4614
rect 5960 4606 5961 4614
rect 5961 4606 5963 4614
rect 5963 4606 5968 4614
rect 5972 4606 5973 4614
rect 5973 4606 5980 4614
rect 1004 4596 1012 4604
rect 4108 4596 4116 4604
rect 6188 4596 6196 4604
rect 6380 4596 6388 4604
rect 1580 4576 1588 4584
rect 6284 4576 6292 4584
rect 1292 4536 1300 4544
rect 1676 4536 1684 4544
rect 2508 4536 2516 4544
rect 4684 4536 4692 4544
rect 4908 4536 4916 4544
rect 6156 4556 6164 4564
rect 6700 4556 6708 4564
rect 7020 4556 7028 4564
rect 1196 4516 1204 4524
rect 1228 4516 1236 4524
rect 3948 4516 3956 4524
rect 4556 4516 4564 4524
rect 4940 4516 4948 4524
rect 1132 4496 1140 4504
rect 1548 4496 1556 4504
rect 3148 4496 3156 4504
rect 3532 4496 3540 4504
rect 2572 4476 2580 4484
rect 4556 4476 4564 4484
rect 6060 4496 6068 4504
rect 6636 4516 6644 4524
rect 7084 4516 7092 4524
rect 6476 4496 6484 4504
rect 6700 4496 6708 4504
rect 6540 4476 6548 4484
rect 6604 4476 6612 4484
rect 300 4456 308 4464
rect 556 4456 564 4464
rect 4716 4456 4724 4464
rect 460 4436 468 4444
rect 2156 4436 2164 4444
rect 3724 4416 3732 4424
rect 5484 4416 5492 4424
rect 6092 4436 6100 4444
rect 1412 4406 1419 4414
rect 1419 4406 1420 4414
rect 1424 4406 1429 4414
rect 1429 4406 1431 4414
rect 1431 4406 1432 4414
rect 1436 4406 1439 4414
rect 1439 4406 1441 4414
rect 1441 4406 1444 4414
rect 1448 4406 1449 4414
rect 1449 4406 1451 4414
rect 1451 4406 1456 4414
rect 1460 4406 1461 4414
rect 1461 4406 1468 4414
rect 4420 4406 4427 4414
rect 4427 4406 4428 4414
rect 4432 4406 4437 4414
rect 4437 4406 4439 4414
rect 4439 4406 4440 4414
rect 4444 4406 4447 4414
rect 4447 4406 4449 4414
rect 4449 4406 4452 4414
rect 4456 4406 4457 4414
rect 4457 4406 4459 4414
rect 4459 4406 4464 4414
rect 4468 4406 4469 4414
rect 4469 4406 4476 4414
rect 4876 4396 4884 4404
rect 6668 4396 6676 4404
rect 6796 4396 6804 4404
rect 7148 4396 7156 4404
rect 1868 4376 1876 4384
rect 3692 4376 3700 4384
rect 5484 4376 5492 4384
rect 6572 4376 6580 4384
rect 6092 4356 6100 4364
rect 6124 4356 6132 4364
rect 428 4336 436 4344
rect 2188 4336 2196 4344
rect 5036 4336 5044 4344
rect 5804 4336 5812 4344
rect 6668 4336 6676 4344
rect 7116 4336 7124 4344
rect 7148 4336 7156 4344
rect 108 4316 116 4324
rect 3596 4296 3604 4304
rect 4684 4316 4692 4324
rect 6060 4316 6068 4324
rect 6572 4316 6580 4324
rect 5036 4296 5044 4304
rect 5004 4276 5012 4284
rect 588 4256 596 4264
rect 1196 4256 1204 4264
rect 2316 4256 2324 4264
rect 4972 4256 4980 4264
rect 1100 4236 1108 4244
rect 4108 4236 4116 4244
rect 4140 4236 4148 4244
rect 5292 4256 5300 4264
rect 5612 4256 5620 4264
rect 6092 4256 6100 4264
rect 7116 4256 7124 4264
rect 5100 4236 5108 4244
rect 5164 4236 5172 4244
rect 3308 4216 3316 4224
rect 2916 4206 2923 4214
rect 2923 4206 2924 4214
rect 2928 4206 2933 4214
rect 2933 4206 2935 4214
rect 2935 4206 2936 4214
rect 2940 4206 2943 4214
rect 2943 4206 2945 4214
rect 2945 4206 2948 4214
rect 2952 4206 2953 4214
rect 2953 4206 2955 4214
rect 2955 4206 2960 4214
rect 2964 4206 2965 4214
rect 2965 4206 2972 4214
rect 748 4176 756 4184
rect 1132 4176 1140 4184
rect 6028 4236 6036 4244
rect 6380 4236 6388 4244
rect 6412 4236 6420 4244
rect 7180 4236 7188 4244
rect 6316 4216 6324 4224
rect 7244 4216 7252 4224
rect 5924 4206 5931 4214
rect 5931 4206 5932 4214
rect 5936 4206 5941 4214
rect 5941 4206 5943 4214
rect 5943 4206 5944 4214
rect 5948 4206 5951 4214
rect 5951 4206 5953 4214
rect 5953 4206 5956 4214
rect 5960 4206 5961 4214
rect 5961 4206 5963 4214
rect 5963 4206 5968 4214
rect 5972 4206 5973 4214
rect 5973 4206 5980 4214
rect 6124 4196 6132 4204
rect 5132 4176 5140 4184
rect 5324 4176 5332 4184
rect 5516 4176 5524 4184
rect 108 4156 116 4164
rect 2540 4156 2548 4164
rect 5772 4156 5780 4164
rect 5804 4156 5812 4164
rect 6284 4196 6292 4204
rect 7212 4176 7220 4184
rect 6892 4156 6900 4164
rect 1548 4136 1556 4144
rect 1676 4136 1684 4144
rect 5164 4136 5172 4144
rect 5484 4136 5492 4144
rect 5868 4136 5876 4144
rect 6028 4136 6036 4144
rect 6252 4136 6260 4144
rect 6668 4136 6676 4144
rect 7308 4136 7316 4144
rect 2636 4116 2644 4124
rect 3916 4116 3924 4124
rect 4044 4116 4052 4124
rect 4268 4116 4276 4124
rect 5804 4116 5812 4124
rect 6060 4116 6068 4124
rect 7244 4116 7252 4124
rect 7372 4116 7380 4124
rect 748 4096 756 4104
rect 1932 4096 1940 4104
rect 4940 4096 4948 4104
rect 6540 4096 6548 4104
rect 7084 4096 7092 4104
rect 1068 4076 1076 4084
rect 1324 4076 1332 4084
rect 1836 4076 1844 4084
rect 1964 4076 1972 4084
rect 3532 4076 3540 4084
rect 4076 4076 4084 4084
rect 4716 4076 4724 4084
rect 1548 4056 1556 4064
rect 2444 4056 2452 4064
rect 460 4036 468 4044
rect 4140 4036 4148 4044
rect 5196 4056 5204 4064
rect 6156 4076 6164 4084
rect 7276 4076 7284 4084
rect 7308 4076 7316 4084
rect 6316 4056 6324 4064
rect 6924 4036 6932 4044
rect 4204 4016 4212 4024
rect 4556 4016 4564 4024
rect 6444 4016 6452 4024
rect 1412 4006 1419 4014
rect 1419 4006 1420 4014
rect 1424 4006 1429 4014
rect 1429 4006 1431 4014
rect 1431 4006 1432 4014
rect 1436 4006 1439 4014
rect 1439 4006 1441 4014
rect 1441 4006 1444 4014
rect 1448 4006 1449 4014
rect 1449 4006 1451 4014
rect 1451 4006 1456 4014
rect 1460 4006 1461 4014
rect 1461 4006 1468 4014
rect 4420 4006 4427 4014
rect 4427 4006 4428 4014
rect 4432 4006 4437 4014
rect 4437 4006 4439 4014
rect 4439 4006 4440 4014
rect 4444 4006 4447 4014
rect 4447 4006 4449 4014
rect 4449 4006 4452 4014
rect 4456 4006 4457 4014
rect 4457 4006 4459 4014
rect 4459 4006 4464 4014
rect 4468 4006 4469 4014
rect 4469 4006 4476 4014
rect 2092 3996 2100 4004
rect 4844 3996 4852 4004
rect 5260 3996 5268 4004
rect 6220 3996 6228 4004
rect 812 3976 820 3984
rect 1996 3976 2004 3984
rect 2700 3976 2708 3984
rect 3372 3976 3380 3984
rect 6732 3976 6740 3984
rect 4684 3956 4692 3964
rect 4780 3956 4788 3964
rect 5196 3956 5204 3964
rect 172 3936 180 3944
rect 1100 3936 1108 3944
rect 4812 3936 4820 3944
rect 5164 3936 5172 3944
rect 2060 3916 2068 3924
rect 2348 3916 2356 3924
rect 2764 3916 2772 3924
rect 684 3896 692 3904
rect 876 3896 884 3904
rect 3692 3896 3700 3904
rect 3724 3896 3732 3904
rect 4044 3896 4052 3904
rect 4076 3896 4084 3904
rect 140 3876 148 3884
rect 428 3876 436 3884
rect 2508 3876 2516 3884
rect 2828 3856 2836 3864
rect 4716 3876 4724 3884
rect 4812 3876 4820 3884
rect 4876 3896 4884 3904
rect 4972 3896 4980 3904
rect 5804 3896 5812 3904
rect 6412 3896 6420 3904
rect 6476 3916 6484 3924
rect 7180 3916 7188 3924
rect 5580 3876 5588 3884
rect 684 3836 692 3844
rect 3948 3836 3956 3844
rect 4204 3836 4212 3844
rect 5100 3836 5108 3844
rect 1196 3816 1204 3824
rect 2916 3806 2923 3814
rect 2923 3806 2924 3814
rect 2928 3806 2933 3814
rect 2933 3806 2935 3814
rect 2935 3806 2936 3814
rect 2940 3806 2943 3814
rect 2943 3806 2945 3814
rect 2945 3806 2948 3814
rect 2952 3806 2953 3814
rect 2953 3806 2955 3814
rect 2955 3806 2960 3814
rect 2964 3806 2965 3814
rect 2965 3806 2972 3814
rect 620 3796 628 3804
rect 4364 3796 4372 3804
rect 4908 3816 4916 3824
rect 4940 3816 4948 3824
rect 6412 3836 6420 3844
rect 5924 3806 5931 3814
rect 5931 3806 5932 3814
rect 5936 3806 5941 3814
rect 5941 3806 5943 3814
rect 5943 3806 5944 3814
rect 5948 3806 5951 3814
rect 5951 3806 5953 3814
rect 5953 3806 5956 3814
rect 5960 3806 5961 3814
rect 5961 3806 5963 3814
rect 5963 3806 5968 3814
rect 5972 3806 5973 3814
rect 5973 3806 5980 3814
rect 5164 3796 5172 3804
rect 5324 3796 5332 3804
rect 204 3776 212 3784
rect 684 3776 692 3784
rect 1292 3776 1300 3784
rect 3692 3776 3700 3784
rect 172 3756 180 3764
rect 876 3756 884 3764
rect 5868 3776 5876 3784
rect 6764 3796 6772 3804
rect 972 3756 980 3764
rect 1868 3756 1876 3764
rect 2316 3756 2324 3764
rect 4972 3756 4980 3764
rect 5260 3756 5268 3764
rect 6348 3756 6356 3764
rect 460 3736 468 3744
rect 588 3736 596 3744
rect 1612 3736 1620 3744
rect 2540 3736 2548 3744
rect 2604 3736 2612 3744
rect 3948 3736 3956 3744
rect 4076 3736 4084 3744
rect 4844 3736 4852 3744
rect 5228 3736 5236 3744
rect 1836 3716 1844 3724
rect 2156 3716 2164 3724
rect 4652 3716 4660 3724
rect 4748 3716 4756 3724
rect 4940 3716 4948 3724
rect 5516 3716 5524 3724
rect 5612 3716 5620 3724
rect 5836 3716 5844 3724
rect 1004 3696 1012 3704
rect 940 3676 948 3684
rect 972 3676 980 3684
rect 3820 3696 3828 3704
rect 4108 3696 4116 3704
rect 4716 3696 4724 3704
rect 3980 3676 3988 3684
rect 4908 3676 4916 3684
rect 5100 3676 5108 3684
rect 5132 3676 5140 3684
rect 1292 3636 1300 3644
rect 1324 3636 1332 3644
rect 3660 3636 3668 3644
rect 5612 3656 5620 3664
rect 7116 3656 7124 3664
rect 4716 3636 4724 3644
rect 5548 3636 5556 3644
rect 6636 3636 6644 3644
rect 6860 3636 6868 3644
rect 7148 3636 7156 3644
rect 3692 3616 3700 3624
rect 4524 3616 4532 3624
rect 5164 3616 5172 3624
rect 5292 3616 5300 3624
rect 1412 3606 1419 3614
rect 1419 3606 1420 3614
rect 1424 3606 1429 3614
rect 1429 3606 1431 3614
rect 1431 3606 1432 3614
rect 1436 3606 1439 3614
rect 1439 3606 1441 3614
rect 1441 3606 1444 3614
rect 1448 3606 1449 3614
rect 1449 3606 1451 3614
rect 1451 3606 1456 3614
rect 1460 3606 1461 3614
rect 1461 3606 1468 3614
rect 4420 3606 4427 3614
rect 4427 3606 4428 3614
rect 4432 3606 4437 3614
rect 4437 3606 4439 3614
rect 4439 3606 4440 3614
rect 4444 3606 4447 3614
rect 4447 3606 4449 3614
rect 4449 3606 4452 3614
rect 4456 3606 4457 3614
rect 4457 3606 4459 3614
rect 4459 3606 4464 3614
rect 4468 3606 4469 3614
rect 4469 3606 4476 3614
rect 3916 3596 3924 3604
rect 4012 3596 4020 3604
rect 972 3576 980 3584
rect 2636 3576 2644 3584
rect 3020 3576 3028 3584
rect 6892 3596 6900 3604
rect 5612 3576 5620 3584
rect 5676 3576 5684 3584
rect 5868 3576 5876 3584
rect 6220 3576 6228 3584
rect 6956 3576 6964 3584
rect 2476 3556 2484 3564
rect 2572 3556 2580 3564
rect 4236 3556 4244 3564
rect 6796 3556 6804 3564
rect 6988 3556 6996 3564
rect 4780 3536 4788 3544
rect 5836 3536 5844 3544
rect 6476 3536 6484 3544
rect 7212 3536 7220 3544
rect 2348 3516 2356 3524
rect 4108 3516 4116 3524
rect 4844 3516 4852 3524
rect 5772 3516 5780 3524
rect 5804 3516 5812 3524
rect 6828 3516 6836 3524
rect 1516 3496 1524 3504
rect 2156 3496 2164 3504
rect 2380 3496 2388 3504
rect 3692 3496 3700 3504
rect 5036 3496 5044 3504
rect 5068 3496 5076 3504
rect 5644 3496 5652 3504
rect 7020 3496 7028 3504
rect 7052 3496 7060 3504
rect 7276 3496 7284 3504
rect 492 3476 500 3484
rect 876 3476 884 3484
rect 2700 3476 2708 3484
rect 4108 3476 4116 3484
rect 4588 3476 4596 3484
rect 5468 3476 5476 3484
rect 6444 3476 6452 3484
rect 6476 3476 6484 3484
rect 6604 3476 6612 3484
rect 1644 3456 1652 3464
rect 3628 3456 3636 3464
rect 4524 3456 4532 3464
rect 3820 3436 3828 3444
rect 4812 3436 4820 3444
rect 556 3416 564 3424
rect 1612 3416 1620 3424
rect 5324 3436 5332 3444
rect 5452 3436 5460 3444
rect 2916 3406 2923 3414
rect 2923 3406 2924 3414
rect 2928 3406 2933 3414
rect 2933 3406 2935 3414
rect 2935 3406 2936 3414
rect 2940 3406 2943 3414
rect 2943 3406 2945 3414
rect 2945 3406 2948 3414
rect 2952 3406 2953 3414
rect 2953 3406 2955 3414
rect 2955 3406 2960 3414
rect 2964 3406 2965 3414
rect 2965 3406 2972 3414
rect 3980 3396 3988 3404
rect 4268 3396 4276 3404
rect 5164 3396 5172 3404
rect 6508 3416 6516 3424
rect 6540 3416 6548 3424
rect 5924 3406 5931 3414
rect 5931 3406 5932 3414
rect 5936 3406 5941 3414
rect 5941 3406 5943 3414
rect 5943 3406 5944 3414
rect 5948 3406 5951 3414
rect 5951 3406 5953 3414
rect 5953 3406 5956 3414
rect 5960 3406 5961 3414
rect 5961 3406 5963 3414
rect 5963 3406 5968 3414
rect 5972 3406 5973 3414
rect 5973 3406 5980 3414
rect 5260 3396 5268 3404
rect 6348 3396 6356 3404
rect 2764 3376 2772 3384
rect 3660 3376 3668 3384
rect 3948 3376 3956 3384
rect 4364 3376 4372 3384
rect 4524 3376 4532 3384
rect 812 3336 820 3344
rect 1004 3336 1012 3344
rect 1292 3336 1300 3344
rect 1644 3336 1652 3344
rect 2476 3356 2484 3364
rect 4044 3356 4052 3364
rect 4748 3356 4756 3364
rect 2732 3336 2740 3344
rect 108 3316 116 3324
rect 876 3316 884 3324
rect 4716 3316 4724 3324
rect 4780 3336 4788 3344
rect 5100 3356 5108 3364
rect 4588 3296 4596 3304
rect 5068 3336 5076 3344
rect 4812 3316 4820 3324
rect 5836 3316 5844 3324
rect 6220 3316 6228 3324
rect 6700 3316 6708 3324
rect 5612 3296 5620 3304
rect 6604 3296 6612 3304
rect 1868 3276 1876 3284
rect 1964 3256 1972 3264
rect 1996 3256 2004 3264
rect 3404 3256 3412 3264
rect 5036 3276 5044 3284
rect 7148 3296 7156 3304
rect 7180 3296 7188 3304
rect 4780 3256 4788 3264
rect 5420 3256 5428 3264
rect 2508 3236 2516 3244
rect 5740 3236 5748 3244
rect 5260 3216 5268 3224
rect 1412 3206 1419 3214
rect 1419 3206 1420 3214
rect 1424 3206 1429 3214
rect 1429 3206 1431 3214
rect 1431 3206 1432 3214
rect 1436 3206 1439 3214
rect 1439 3206 1441 3214
rect 1441 3206 1444 3214
rect 1448 3206 1449 3214
rect 1449 3206 1451 3214
rect 1451 3206 1456 3214
rect 1460 3206 1461 3214
rect 1461 3206 1468 3214
rect 4420 3206 4427 3214
rect 4427 3206 4428 3214
rect 4432 3206 4437 3214
rect 4437 3206 4439 3214
rect 4439 3206 4440 3214
rect 4444 3206 4447 3214
rect 4447 3206 4449 3214
rect 4449 3206 4452 3214
rect 4456 3206 4457 3214
rect 4457 3206 4459 3214
rect 4459 3206 4464 3214
rect 4468 3206 4469 3214
rect 4469 3206 4476 3214
rect 492 3196 500 3204
rect 1516 3196 1524 3204
rect 2156 3196 2164 3204
rect 4332 3196 4340 3204
rect 5324 3196 5332 3204
rect 5644 3196 5652 3204
rect 5676 3196 5684 3204
rect 1740 3176 1748 3184
rect 3148 3176 3156 3184
rect 5484 3176 5492 3184
rect 908 3156 916 3164
rect 1324 3156 1332 3164
rect 3436 3156 3444 3164
rect 3692 3156 3700 3164
rect 3980 3156 3988 3164
rect 4108 3156 4116 3164
rect 748 3136 756 3144
rect 844 3136 852 3144
rect 1260 3136 1268 3144
rect 1292 3136 1300 3144
rect 1356 3136 1364 3144
rect 2092 3136 2100 3144
rect 5836 3156 5844 3164
rect 7148 3156 7156 3164
rect 7180 3156 7188 3164
rect 6252 3136 6260 3144
rect 620 3116 628 3124
rect 1772 3116 1780 3124
rect 1804 3116 1812 3124
rect 1964 3116 1972 3124
rect 2220 3116 2228 3124
rect 2668 3116 2676 3124
rect 3180 3116 3188 3124
rect 4108 3116 4116 3124
rect 684 3096 692 3104
rect 972 3096 980 3104
rect 1260 3096 1268 3104
rect 1548 3096 1556 3104
rect 1612 3096 1620 3104
rect 2380 3096 2388 3104
rect 2508 3096 2516 3104
rect 3980 3096 3988 3104
rect 4012 3096 4020 3104
rect 4332 3096 4340 3104
rect 556 3076 564 3084
rect 2348 3076 2356 3084
rect 5228 3116 5236 3124
rect 5612 3116 5620 3124
rect 4844 3096 4852 3104
rect 4876 3096 4884 3104
rect 5580 3096 5588 3104
rect 7244 3096 7252 3104
rect 4940 3076 4948 3084
rect 5132 3076 5140 3084
rect 6700 3076 6708 3084
rect 1612 3056 1620 3064
rect 1772 3056 1780 3064
rect 3564 3036 3572 3044
rect 3628 3036 3636 3044
rect 6668 3036 6676 3044
rect 2572 3016 2580 3024
rect 4140 3016 4148 3024
rect 4524 3016 4532 3024
rect 4876 3016 4884 3024
rect 2916 3006 2923 3014
rect 2923 3006 2924 3014
rect 2928 3006 2933 3014
rect 2933 3006 2935 3014
rect 2935 3006 2936 3014
rect 2940 3006 2943 3014
rect 2943 3006 2945 3014
rect 2945 3006 2948 3014
rect 2952 3006 2953 3014
rect 2953 3006 2955 3014
rect 2955 3006 2960 3014
rect 2964 3006 2965 3014
rect 2965 3006 2972 3014
rect 1740 2996 1748 3004
rect 5924 3006 5931 3014
rect 5931 3006 5932 3014
rect 5936 3006 5941 3014
rect 5941 3006 5943 3014
rect 5943 3006 5944 3014
rect 5948 3006 5951 3014
rect 5951 3006 5953 3014
rect 5953 3006 5956 3014
rect 5960 3006 5961 3014
rect 5961 3006 5963 3014
rect 5963 3006 5968 3014
rect 5972 3006 5973 3014
rect 5973 3006 5980 3014
rect 4972 2996 4980 3004
rect 7212 2996 7220 3004
rect 4812 2976 4820 2984
rect 6444 2976 6452 2984
rect 7116 2976 7124 2984
rect 1804 2956 1812 2964
rect 1836 2956 1844 2964
rect 2284 2956 2292 2964
rect 4236 2956 4244 2964
rect 5068 2956 5076 2964
rect 6508 2956 6516 2964
rect 7340 2956 7348 2964
rect 1324 2936 1332 2944
rect 1580 2936 1588 2944
rect 2604 2936 2612 2944
rect 3404 2936 3412 2944
rect 4364 2936 4372 2944
rect 6220 2936 6228 2944
rect 1036 2916 1044 2924
rect 1260 2916 1268 2924
rect 1356 2916 1364 2924
rect 2156 2916 2164 2924
rect 2412 2916 2420 2924
rect 3788 2916 3796 2924
rect 3820 2916 3828 2924
rect 4652 2916 4660 2924
rect 4716 2916 4724 2924
rect 5100 2916 5108 2924
rect 844 2896 852 2904
rect 2220 2896 2228 2904
rect 2444 2896 2452 2904
rect 3564 2896 3572 2904
rect 556 2876 564 2884
rect 1708 2876 1716 2884
rect 1740 2876 1748 2884
rect 1964 2876 1972 2884
rect 4332 2876 4340 2884
rect 4652 2876 4660 2884
rect 5068 2896 5076 2904
rect 5420 2896 5428 2904
rect 6412 2916 6420 2924
rect 5516 2876 5524 2884
rect 1004 2856 1012 2864
rect 4300 2856 4308 2864
rect 5036 2856 5044 2864
rect 5132 2856 5140 2864
rect 6924 2856 6932 2864
rect 1068 2836 1076 2844
rect 1100 2836 1108 2844
rect 3020 2836 3028 2844
rect 6284 2836 6292 2844
rect 3052 2816 3060 2824
rect 5004 2816 5012 2824
rect 5164 2816 5172 2824
rect 5196 2816 5204 2824
rect 5292 2816 5300 2824
rect 5356 2816 5364 2824
rect 1412 2806 1419 2814
rect 1419 2806 1420 2814
rect 1424 2806 1429 2814
rect 1429 2806 1431 2814
rect 1431 2806 1432 2814
rect 1436 2806 1439 2814
rect 1439 2806 1441 2814
rect 1441 2806 1444 2814
rect 1448 2806 1449 2814
rect 1449 2806 1451 2814
rect 1451 2806 1456 2814
rect 1460 2806 1461 2814
rect 1461 2806 1468 2814
rect 4420 2806 4427 2814
rect 4427 2806 4428 2814
rect 4432 2806 4437 2814
rect 4437 2806 4439 2814
rect 4439 2806 4440 2814
rect 4444 2806 4447 2814
rect 4447 2806 4449 2814
rect 4449 2806 4452 2814
rect 4456 2806 4457 2814
rect 4457 2806 4459 2814
rect 4459 2806 4464 2814
rect 4468 2806 4469 2814
rect 4469 2806 4476 2814
rect 3628 2796 3636 2804
rect 5004 2776 5012 2784
rect 5836 2776 5844 2784
rect 2380 2756 2388 2764
rect 6508 2756 6516 2764
rect 1836 2736 1844 2744
rect 2828 2736 2836 2744
rect 2860 2736 2868 2744
rect 3308 2736 3316 2744
rect 4940 2736 4948 2744
rect 5068 2736 5076 2744
rect 5100 2736 5108 2744
rect 5772 2736 5780 2744
rect 5804 2736 5812 2744
rect 652 2716 660 2724
rect 1036 2716 1044 2724
rect 2508 2716 2516 2724
rect 172 2696 180 2704
rect 1900 2696 1908 2704
rect 5068 2696 5076 2704
rect 6668 2696 6676 2704
rect 6860 2696 6868 2704
rect 108 2656 116 2664
rect 2732 2676 2740 2684
rect 4300 2676 4308 2684
rect 5196 2676 5204 2684
rect 6220 2676 6228 2684
rect 6636 2676 6644 2684
rect 1836 2656 1844 2664
rect 4876 2656 4884 2664
rect 4908 2656 4916 2664
rect 6668 2656 6676 2664
rect 7020 2656 7028 2664
rect 2476 2636 2484 2644
rect 3372 2636 3380 2644
rect 5612 2636 5620 2644
rect 6476 2636 6484 2644
rect 2916 2606 2923 2614
rect 2923 2606 2924 2614
rect 2928 2606 2933 2614
rect 2933 2606 2935 2614
rect 2935 2606 2936 2614
rect 2940 2606 2943 2614
rect 2943 2606 2945 2614
rect 2945 2606 2948 2614
rect 2952 2606 2953 2614
rect 2953 2606 2955 2614
rect 2955 2606 2960 2614
rect 2964 2606 2965 2614
rect 2965 2606 2972 2614
rect 5924 2606 5931 2614
rect 5931 2606 5932 2614
rect 5936 2606 5941 2614
rect 5941 2606 5943 2614
rect 5943 2606 5944 2614
rect 5948 2606 5951 2614
rect 5951 2606 5953 2614
rect 5953 2606 5956 2614
rect 5960 2606 5961 2614
rect 5961 2606 5963 2614
rect 5963 2606 5968 2614
rect 5972 2606 5973 2614
rect 5973 2606 5980 2614
rect 2476 2596 2484 2604
rect 4268 2596 4276 2604
rect 4940 2596 4948 2604
rect 5164 2596 5172 2604
rect 5452 2596 5460 2604
rect 2284 2576 2292 2584
rect 2828 2576 2836 2584
rect 4716 2576 4724 2584
rect 5292 2576 5300 2584
rect 6124 2556 6132 2564
rect 2316 2536 2324 2544
rect 2668 2536 2676 2544
rect 2860 2536 2868 2544
rect 4812 2536 4820 2544
rect 3596 2516 3604 2524
rect 4876 2516 4884 2524
rect 5260 2536 5268 2544
rect 5324 2536 5332 2544
rect 5356 2536 5364 2544
rect 7308 2536 7316 2544
rect 7340 2536 7348 2544
rect 5036 2516 5044 2524
rect 5548 2516 5556 2524
rect 6412 2516 6420 2524
rect 1868 2496 1876 2504
rect 3148 2496 3156 2504
rect 4204 2496 4212 2504
rect 4844 2496 4852 2504
rect 5260 2496 5268 2504
rect 7404 2496 7412 2504
rect 748 2476 756 2484
rect 2220 2476 2228 2484
rect 3980 2476 3988 2484
rect 4652 2476 4660 2484
rect 5548 2476 5556 2484
rect 1708 2456 1716 2464
rect 2188 2456 2196 2464
rect 3788 2456 3796 2464
rect 5196 2456 5204 2464
rect 1292 2436 1300 2444
rect 3340 2436 3348 2444
rect 4716 2436 4724 2444
rect 4780 2436 4788 2444
rect 492 2416 500 2424
rect 1740 2416 1748 2424
rect 4140 2416 4148 2424
rect 4556 2416 4564 2424
rect 5516 2416 5524 2424
rect 6892 2416 6900 2424
rect 1412 2406 1419 2414
rect 1419 2406 1420 2414
rect 1424 2406 1429 2414
rect 1429 2406 1431 2414
rect 1431 2406 1432 2414
rect 1436 2406 1439 2414
rect 1439 2406 1441 2414
rect 1441 2406 1444 2414
rect 1448 2406 1449 2414
rect 1449 2406 1451 2414
rect 1451 2406 1456 2414
rect 1460 2406 1461 2414
rect 1461 2406 1468 2414
rect 4420 2406 4427 2414
rect 4427 2406 4428 2414
rect 4432 2406 4437 2414
rect 4437 2406 4439 2414
rect 4439 2406 4440 2414
rect 4444 2406 4447 2414
rect 4447 2406 4449 2414
rect 4449 2406 4452 2414
rect 4456 2406 4457 2414
rect 4457 2406 4459 2414
rect 4459 2406 4464 2414
rect 4468 2406 4469 2414
rect 4469 2406 4476 2414
rect 1900 2396 1908 2404
rect 1676 2376 1684 2384
rect 2284 2376 2292 2384
rect 1644 2356 1652 2364
rect 5324 2396 5332 2404
rect 6284 2396 6292 2404
rect 6348 2396 6356 2404
rect 2380 2356 2388 2364
rect 3244 2356 3252 2364
rect 4044 2356 4052 2364
rect 7212 2376 7220 2384
rect 588 2336 596 2344
rect 1612 2336 1620 2344
rect 204 2316 212 2324
rect 3628 2316 3636 2324
rect 6060 2336 6068 2344
rect 5772 2316 5780 2324
rect 44 2296 52 2304
rect 1900 2296 1908 2304
rect 2412 2296 2420 2304
rect 2444 2296 2452 2304
rect 2828 2296 2836 2304
rect 3436 2296 3444 2304
rect 4108 2296 4116 2304
rect 4300 2296 4308 2304
rect 2796 2276 2804 2284
rect 2860 2276 2868 2284
rect 4748 2296 4756 2304
rect 5164 2296 5172 2304
rect 5228 2296 5236 2304
rect 6124 2296 6132 2304
rect 4364 2276 4372 2284
rect 4652 2276 4660 2284
rect 4684 2276 4692 2284
rect 4844 2276 4852 2284
rect 5580 2276 5588 2284
rect 5612 2276 5620 2284
rect 5772 2276 5780 2284
rect 6028 2276 6036 2284
rect 6636 2276 6644 2284
rect 7340 2276 7348 2284
rect 1164 2256 1172 2264
rect 2380 2256 2388 2264
rect 2476 2256 2484 2264
rect 4748 2256 4756 2264
rect 172 2236 180 2244
rect 588 2236 596 2244
rect 1324 2236 1332 2244
rect 1612 2236 1620 2244
rect 4908 2236 4916 2244
rect 4972 2236 4980 2244
rect 5484 2256 5492 2264
rect 6220 2256 6228 2264
rect 5644 2236 5652 2244
rect 1772 2196 1780 2204
rect 3180 2216 3188 2224
rect 5868 2216 5876 2224
rect 2916 2206 2923 2214
rect 2923 2206 2924 2214
rect 2928 2206 2933 2214
rect 2933 2206 2935 2214
rect 2935 2206 2936 2214
rect 2940 2206 2943 2214
rect 2943 2206 2945 2214
rect 2945 2206 2948 2214
rect 2952 2206 2953 2214
rect 2953 2206 2955 2214
rect 2955 2206 2960 2214
rect 2964 2206 2965 2214
rect 2965 2206 2972 2214
rect 1196 2176 1204 2184
rect 1228 2176 1236 2184
rect 1164 2156 1172 2164
rect 1900 2156 1908 2164
rect 1964 2156 1972 2164
rect 4300 2176 4308 2184
rect 4332 2176 4340 2184
rect 4940 2176 4948 2184
rect 5196 2176 5204 2184
rect 5292 2176 5300 2184
rect 5452 2176 5460 2184
rect 7404 2256 7412 2264
rect 5924 2206 5931 2214
rect 5931 2206 5932 2214
rect 5936 2206 5941 2214
rect 5941 2206 5943 2214
rect 5943 2206 5944 2214
rect 5948 2206 5951 2214
rect 5951 2206 5953 2214
rect 5953 2206 5956 2214
rect 5960 2206 5961 2214
rect 5961 2206 5963 2214
rect 5963 2206 5968 2214
rect 5972 2206 5973 2214
rect 5973 2206 5980 2214
rect 6060 2196 6068 2204
rect 7276 2196 7284 2204
rect 3788 2156 3796 2164
rect 5004 2156 5012 2164
rect 5836 2156 5844 2164
rect 6572 2156 6580 2164
rect 1612 2136 1620 2144
rect 2284 2136 2292 2144
rect 2348 2136 2356 2144
rect 2860 2136 2868 2144
rect 4300 2136 4308 2144
rect 4332 2136 4340 2144
rect 4940 2136 4948 2144
rect 5612 2136 5620 2144
rect 1548 2116 1556 2124
rect 1772 2116 1780 2124
rect 2412 2116 2420 2124
rect 2572 2116 2580 2124
rect 4876 2116 4884 2124
rect 5100 2116 5108 2124
rect 5516 2116 5524 2124
rect 2156 2096 2164 2104
rect 2444 2096 2452 2104
rect 3020 2096 3028 2104
rect 4332 2096 4340 2104
rect 4844 2096 4852 2104
rect 908 2076 916 2084
rect 2796 2076 2804 2084
rect 428 2036 436 2044
rect 1708 2056 1716 2064
rect 4012 2076 4020 2084
rect 4524 2076 4532 2084
rect 5004 2076 5012 2084
rect 5036 2076 5044 2084
rect 5196 2076 5204 2084
rect 5260 2076 5268 2084
rect 5292 2076 5300 2084
rect 5388 2076 5396 2084
rect 6028 2116 6036 2124
rect 7340 2116 7348 2124
rect 6060 2096 6068 2104
rect 6316 2096 6324 2104
rect 5484 2056 5492 2064
rect 3212 2036 3220 2044
rect 3564 2036 3572 2044
rect 3820 2036 3828 2044
rect 1708 2016 1716 2024
rect 1868 2016 1876 2024
rect 2124 2016 2132 2024
rect 1412 2006 1419 2014
rect 1419 2006 1420 2014
rect 1424 2006 1429 2014
rect 1429 2006 1431 2014
rect 1431 2006 1432 2014
rect 1436 2006 1439 2014
rect 1439 2006 1441 2014
rect 1441 2006 1444 2014
rect 1448 2006 1449 2014
rect 1449 2006 1451 2014
rect 1451 2006 1456 2014
rect 1460 2006 1461 2014
rect 1461 2006 1468 2014
rect 1516 1996 1524 2004
rect 4524 2016 4532 2024
rect 4812 2016 4820 2024
rect 5452 2016 5460 2024
rect 6060 2036 6068 2044
rect 4420 2006 4427 2014
rect 4427 2006 4428 2014
rect 4432 2006 4437 2014
rect 4437 2006 4439 2014
rect 4439 2006 4440 2014
rect 4444 2006 4447 2014
rect 4447 2006 4449 2014
rect 4449 2006 4452 2014
rect 4456 2006 4457 2014
rect 4457 2006 4459 2014
rect 4459 2006 4464 2014
rect 4468 2006 4469 2014
rect 4469 2006 4476 2014
rect 3244 1996 3252 2004
rect 652 1976 660 1984
rect 2188 1976 2196 1984
rect 4044 1976 4052 1984
rect 4908 1996 4916 2004
rect 5164 1996 5172 2004
rect 6700 1996 6708 2004
rect 1516 1956 1524 1964
rect 716 1936 724 1944
rect 2348 1936 2356 1944
rect 1164 1916 1172 1924
rect 3084 1916 3092 1924
rect 4588 1936 4596 1944
rect 5452 1936 5460 1944
rect 2220 1896 2228 1904
rect 5260 1916 5268 1924
rect 6028 1916 6036 1924
rect 4716 1896 4724 1904
rect 1708 1876 1716 1884
rect 2252 1876 2260 1884
rect 2700 1876 2708 1884
rect 4076 1876 4084 1884
rect 4748 1876 4756 1884
rect 5132 1876 5140 1884
rect 5548 1876 5556 1884
rect 6028 1876 6036 1884
rect 6412 1876 6420 1884
rect 6956 1876 6964 1884
rect 1612 1856 1620 1864
rect 2092 1856 2100 1864
rect 2476 1856 2484 1864
rect 3052 1856 3060 1864
rect 4652 1856 4660 1864
rect 4908 1856 4916 1864
rect 1516 1836 1524 1844
rect 4588 1836 4596 1844
rect 5580 1856 5588 1864
rect 6316 1856 6324 1864
rect 7116 1856 7124 1864
rect 1772 1816 1780 1824
rect 5740 1836 5748 1844
rect 6028 1816 6036 1824
rect 6188 1816 6196 1824
rect 2916 1806 2923 1814
rect 2923 1806 2924 1814
rect 2928 1806 2933 1814
rect 2933 1806 2935 1814
rect 2935 1806 2936 1814
rect 2940 1806 2943 1814
rect 2943 1806 2945 1814
rect 2945 1806 2948 1814
rect 2952 1806 2953 1814
rect 2953 1806 2955 1814
rect 2955 1806 2960 1814
rect 2964 1806 2965 1814
rect 2965 1806 2972 1814
rect 5924 1806 5931 1814
rect 5931 1806 5932 1814
rect 5936 1806 5941 1814
rect 5941 1806 5943 1814
rect 5943 1806 5944 1814
rect 5948 1806 5951 1814
rect 5951 1806 5953 1814
rect 5953 1806 5956 1814
rect 5960 1806 5961 1814
rect 5961 1806 5963 1814
rect 5963 1806 5968 1814
rect 5972 1806 5973 1814
rect 5973 1806 5980 1814
rect 4076 1796 4084 1804
rect 1644 1776 1652 1784
rect 4748 1776 4756 1784
rect 5708 1776 5716 1784
rect 2476 1736 2484 1744
rect 4012 1756 4020 1764
rect 4524 1756 4532 1764
rect 5420 1756 5428 1764
rect 7148 1756 7156 1764
rect 3372 1736 3380 1744
rect 1836 1716 1844 1724
rect 2156 1716 2164 1724
rect 2220 1716 2228 1724
rect 2444 1716 2452 1724
rect 3756 1716 3764 1724
rect 4620 1716 4628 1724
rect 5068 1716 5076 1724
rect 5132 1736 5140 1744
rect 5836 1736 5844 1744
rect 5548 1716 5556 1724
rect 6572 1736 6580 1744
rect 7116 1716 7124 1724
rect 652 1696 660 1704
rect 1228 1696 1236 1704
rect 2092 1696 2100 1704
rect 2348 1696 2356 1704
rect 2380 1696 2388 1704
rect 4300 1696 4308 1704
rect 4716 1696 4724 1704
rect 5708 1696 5716 1704
rect 7180 1696 7188 1704
rect 7404 1696 7412 1704
rect 3628 1676 3636 1684
rect 3980 1676 3988 1684
rect 4684 1676 4692 1684
rect 5260 1676 5268 1684
rect 44 1656 52 1664
rect 2156 1656 2164 1664
rect 3660 1656 3668 1664
rect 1132 1636 1140 1644
rect 1708 1636 1716 1644
rect 7404 1656 7412 1664
rect 1324 1616 1332 1624
rect 1868 1616 1876 1624
rect 2092 1616 2100 1624
rect 2124 1616 2132 1624
rect 1412 1606 1419 1614
rect 1419 1606 1420 1614
rect 1424 1606 1429 1614
rect 1429 1606 1431 1614
rect 1431 1606 1432 1614
rect 1436 1606 1439 1614
rect 1439 1606 1441 1614
rect 1441 1606 1444 1614
rect 1448 1606 1449 1614
rect 1449 1606 1451 1614
rect 1451 1606 1456 1614
rect 1460 1606 1461 1614
rect 1461 1606 1468 1614
rect 4420 1606 4427 1614
rect 4427 1606 4428 1614
rect 4432 1606 4437 1614
rect 4437 1606 4439 1614
rect 4439 1606 4440 1614
rect 4444 1606 4447 1614
rect 4447 1606 4449 1614
rect 4449 1606 4452 1614
rect 4456 1606 4457 1614
rect 4457 1606 4459 1614
rect 4459 1606 4464 1614
rect 4468 1606 4469 1614
rect 4469 1606 4476 1614
rect 4524 1596 4532 1604
rect 4748 1596 4756 1604
rect 5420 1596 5428 1604
rect 876 1576 884 1584
rect 1068 1556 1076 1564
rect 1740 1556 1748 1564
rect 1996 1556 2004 1564
rect 3340 1556 3348 1564
rect 5388 1556 5396 1564
rect 492 1536 500 1544
rect 748 1536 756 1544
rect 1164 1536 1172 1544
rect 2060 1536 2068 1544
rect 3308 1536 3316 1544
rect 4268 1536 4276 1544
rect 6348 1536 6356 1544
rect 1036 1516 1044 1524
rect 1804 1516 1812 1524
rect 2604 1516 2612 1524
rect 2860 1516 2868 1524
rect 3020 1516 3028 1524
rect 3660 1516 3668 1524
rect 5004 1516 5012 1524
rect 5740 1516 5748 1524
rect 5868 1516 5876 1524
rect 6252 1516 6260 1524
rect 6508 1516 6516 1524
rect 716 1496 724 1504
rect 1612 1496 1620 1504
rect 1996 1496 2004 1504
rect 3244 1496 3252 1504
rect 4556 1496 4564 1504
rect 4588 1496 4596 1504
rect 4812 1496 4820 1504
rect 7020 1496 7028 1504
rect 1068 1476 1076 1484
rect 876 1456 884 1464
rect 2092 1476 2100 1484
rect 2284 1476 2292 1484
rect 2476 1476 2484 1484
rect 2636 1476 2644 1484
rect 2700 1476 2708 1484
rect 2732 1476 2740 1484
rect 3436 1476 3444 1484
rect 4364 1476 4372 1484
rect 1932 1456 1940 1464
rect 4556 1456 4564 1464
rect 4812 1456 4820 1464
rect 6220 1476 6228 1484
rect 7308 1476 7316 1484
rect 5548 1456 5556 1464
rect 2796 1436 2804 1444
rect 3244 1436 3252 1444
rect 940 1416 948 1424
rect 1004 1416 1012 1424
rect 1324 1416 1332 1424
rect 908 1396 916 1404
rect 3084 1416 3092 1424
rect 4140 1416 4148 1424
rect 4172 1436 4180 1444
rect 4876 1436 4884 1444
rect 6412 1436 6420 1444
rect 6988 1436 6996 1444
rect 4908 1416 4916 1424
rect 7372 1416 7380 1424
rect 2916 1406 2923 1414
rect 2923 1406 2924 1414
rect 2928 1406 2933 1414
rect 2933 1406 2935 1414
rect 2935 1406 2936 1414
rect 2940 1406 2943 1414
rect 2943 1406 2945 1414
rect 2945 1406 2948 1414
rect 2952 1406 2953 1414
rect 2953 1406 2955 1414
rect 2955 1406 2960 1414
rect 2964 1406 2965 1414
rect 2965 1406 2972 1414
rect 5924 1406 5931 1414
rect 5931 1406 5932 1414
rect 5936 1406 5941 1414
rect 5941 1406 5943 1414
rect 5943 1406 5944 1414
rect 5948 1406 5951 1414
rect 5951 1406 5953 1414
rect 5953 1406 5956 1414
rect 5960 1406 5961 1414
rect 5961 1406 5963 1414
rect 5963 1406 5968 1414
rect 5972 1406 5973 1414
rect 5973 1406 5980 1414
rect 1100 1376 1108 1384
rect 2028 1376 2036 1384
rect 2572 1376 2580 1384
rect 2604 1376 2612 1384
rect 3308 1396 3316 1404
rect 2860 1376 2868 1384
rect 3148 1376 3156 1384
rect 3564 1396 3572 1404
rect 4780 1396 4788 1404
rect 6188 1396 6196 1404
rect 7404 1396 7412 1404
rect 812 1356 820 1364
rect 1228 1356 1236 1364
rect 1708 1356 1716 1364
rect 2092 1356 2100 1364
rect 5068 1376 5076 1384
rect 7116 1356 7124 1364
rect 2220 1336 2228 1344
rect 2412 1336 2420 1344
rect 44 1316 52 1324
rect 844 1316 852 1324
rect 1676 1316 1684 1324
rect 1708 1316 1716 1324
rect 1996 1316 2004 1324
rect 2060 1316 2068 1324
rect 2460 1316 2468 1324
rect 2636 1316 2644 1324
rect 2732 1316 2740 1324
rect 3084 1336 3092 1344
rect 3436 1316 3444 1324
rect 6860 1336 6868 1344
rect 7148 1336 7156 1344
rect 4140 1316 4148 1324
rect 4556 1316 4564 1324
rect 4620 1316 4628 1324
rect 1164 1296 1172 1304
rect 1740 1296 1748 1304
rect 2284 1296 2292 1304
rect 2380 1296 2388 1304
rect 2412 1296 2420 1304
rect 4300 1296 4308 1304
rect 4844 1296 4852 1304
rect 7276 1316 7284 1324
rect 7116 1296 7124 1304
rect 1772 1256 1780 1264
rect 1836 1256 1844 1264
rect 6220 1256 6228 1264
rect 6412 1256 6420 1264
rect 4588 1236 4596 1244
rect 1772 1216 1780 1224
rect 1804 1216 1812 1224
rect 2092 1216 2100 1224
rect 2156 1216 2164 1224
rect 2252 1216 2260 1224
rect 3820 1216 3828 1224
rect 1412 1206 1419 1214
rect 1419 1206 1420 1214
rect 1424 1206 1429 1214
rect 1429 1206 1431 1214
rect 1431 1206 1432 1214
rect 1436 1206 1439 1214
rect 1439 1206 1441 1214
rect 1441 1206 1444 1214
rect 1448 1206 1449 1214
rect 1449 1206 1451 1214
rect 1451 1206 1456 1214
rect 1460 1206 1461 1214
rect 1461 1206 1468 1214
rect 876 1196 884 1204
rect 2412 1196 2420 1204
rect 2444 1196 2452 1204
rect 2572 1196 2580 1204
rect 2796 1196 2804 1204
rect 3116 1196 3124 1204
rect 3148 1196 3156 1204
rect 4172 1216 4180 1224
rect 4908 1216 4916 1224
rect 6028 1216 6036 1224
rect 6860 1216 6868 1224
rect 4420 1206 4427 1214
rect 4427 1206 4428 1214
rect 4432 1206 4437 1214
rect 4437 1206 4439 1214
rect 4439 1206 4440 1214
rect 4444 1206 4447 1214
rect 4447 1206 4449 1214
rect 4449 1206 4452 1214
rect 4456 1206 4457 1214
rect 4457 1206 4459 1214
rect 4459 1206 4464 1214
rect 4468 1206 4469 1214
rect 4469 1206 4476 1214
rect 4940 1196 4948 1204
rect 6604 1196 6612 1204
rect 4908 1176 4916 1184
rect 1324 1156 1332 1164
rect 1996 1156 2004 1164
rect 2028 1156 2036 1164
rect 4972 1156 4980 1164
rect 1932 1136 1940 1144
rect 1964 1136 1972 1144
rect 3372 1136 3380 1144
rect 3788 1136 3796 1144
rect 4716 1136 4724 1144
rect 7180 1156 7188 1164
rect 940 1116 948 1124
rect 1036 1116 1044 1124
rect 1132 1116 1140 1124
rect 2060 1116 2068 1124
rect 2252 1116 2260 1124
rect 2444 1116 2452 1124
rect 2476 1116 2484 1124
rect 2508 1116 2516 1124
rect 812 1096 820 1104
rect 908 1096 916 1104
rect 3148 1096 3156 1104
rect 3628 1116 3636 1124
rect 3660 1116 3668 1124
rect 5484 1116 5492 1124
rect 5868 1116 5876 1124
rect 7212 1116 7220 1124
rect 844 1076 852 1084
rect 3436 1076 3444 1084
rect 4044 1096 4052 1104
rect 4684 1096 4692 1104
rect 4780 1096 4788 1104
rect 4972 1096 4980 1104
rect 5356 1096 5364 1104
rect 5548 1096 5556 1104
rect 5580 1096 5588 1104
rect 7340 1096 7348 1104
rect 7308 1076 7316 1084
rect 1740 1056 1748 1064
rect 1932 1056 1940 1064
rect 2252 1056 2260 1064
rect 2284 1056 2292 1064
rect 2444 1056 2452 1064
rect 4524 1056 4532 1064
rect 4940 1056 4948 1064
rect 5580 1056 5588 1064
rect 5740 1056 5748 1064
rect 1580 1036 1588 1044
rect 4332 1036 4340 1044
rect 4364 1036 4372 1044
rect 1324 1016 1332 1024
rect 3020 1016 3028 1024
rect 3884 1016 3892 1024
rect 2916 1006 2923 1014
rect 2923 1006 2924 1014
rect 2928 1006 2933 1014
rect 2933 1006 2935 1014
rect 2935 1006 2936 1014
rect 2940 1006 2943 1014
rect 2943 1006 2945 1014
rect 2945 1006 2948 1014
rect 2952 1006 2953 1014
rect 2953 1006 2955 1014
rect 2955 1006 2960 1014
rect 2964 1006 2965 1014
rect 2965 1006 2972 1014
rect 940 996 948 1004
rect 1900 996 1908 1004
rect 1132 976 1140 984
rect 1740 976 1748 984
rect 2300 996 2308 1004
rect 2700 996 2708 1004
rect 2092 976 2100 984
rect 2828 996 2836 1004
rect 4524 1016 4532 1024
rect 5868 1016 5876 1024
rect 5924 1006 5931 1014
rect 5931 1006 5932 1014
rect 5936 1006 5941 1014
rect 5941 1006 5943 1014
rect 5943 1006 5944 1014
rect 5948 1006 5951 1014
rect 5951 1006 5953 1014
rect 5953 1006 5956 1014
rect 5960 1006 5961 1014
rect 5961 1006 5963 1014
rect 5963 1006 5968 1014
rect 5972 1006 5973 1014
rect 5973 1006 5980 1014
rect 4812 996 4820 1004
rect 5260 996 5268 1004
rect 5420 996 5428 1004
rect 2860 976 2868 984
rect 3276 976 3284 984
rect 4652 976 4660 984
rect 1932 956 1940 964
rect 1868 916 1876 924
rect 3052 956 3060 964
rect 6124 956 6132 964
rect 6604 956 6612 964
rect 3436 936 3444 944
rect 3756 936 3764 944
rect 4332 936 4340 944
rect 6188 936 6196 944
rect 2572 916 2580 924
rect 5004 916 5012 924
rect 7212 916 7220 924
rect 1772 896 1780 904
rect 1900 896 1908 904
rect 2316 896 2324 904
rect 2604 896 2612 904
rect 2700 896 2708 904
rect 3756 896 3764 904
rect 3916 896 3924 904
rect 5740 896 5748 904
rect 6764 896 6772 904
rect 2220 876 2228 884
rect 3244 856 3252 864
rect 1580 836 1588 844
rect 1708 836 1716 844
rect 5324 876 5332 884
rect 5068 856 5076 864
rect 6476 836 6484 844
rect 5228 816 5236 824
rect 5420 816 5428 824
rect 5804 816 5812 824
rect 1412 806 1419 814
rect 1419 806 1420 814
rect 1424 806 1429 814
rect 1429 806 1431 814
rect 1431 806 1432 814
rect 1436 806 1439 814
rect 1439 806 1441 814
rect 1441 806 1444 814
rect 1448 806 1449 814
rect 1449 806 1451 814
rect 1451 806 1456 814
rect 1460 806 1461 814
rect 1461 806 1468 814
rect 4420 806 4427 814
rect 4427 806 4428 814
rect 4432 806 4437 814
rect 4437 806 4439 814
rect 4439 806 4440 814
rect 4444 806 4447 814
rect 4447 806 4449 814
rect 4449 806 4452 814
rect 4456 806 4457 814
rect 4457 806 4459 814
rect 4459 806 4464 814
rect 4468 806 4469 814
rect 4469 806 4476 814
rect 1868 796 1876 804
rect 2316 796 2324 804
rect 3020 796 3028 804
rect 3404 796 3412 804
rect 4748 796 4756 804
rect 4876 796 4884 804
rect 1196 776 1204 784
rect 204 736 212 744
rect 1612 736 1620 744
rect 3436 776 3444 784
rect 5356 776 5364 784
rect 5676 776 5684 784
rect 2412 736 2420 744
rect 3660 736 3668 744
rect 4716 736 4724 744
rect 268 716 276 724
rect 4044 716 4052 724
rect 748 696 756 704
rect 908 696 916 704
rect 1900 696 1908 704
rect 2412 696 2420 704
rect 4684 696 4692 704
rect 4876 716 4884 724
rect 5644 716 5652 724
rect 5772 716 5780 724
rect 7212 716 7220 724
rect 6028 696 6036 704
rect 7084 696 7092 704
rect 3116 676 3124 684
rect 140 636 148 644
rect 3404 636 3412 644
rect 3660 656 3668 664
rect 3884 656 3892 664
rect 6124 656 6132 664
rect 6156 656 6164 664
rect 6764 656 6772 664
rect 3916 636 3924 644
rect 1004 616 1012 624
rect 3532 616 3540 624
rect 4908 616 4916 624
rect 5260 616 5268 624
rect 2916 606 2923 614
rect 2923 606 2924 614
rect 2928 606 2933 614
rect 2933 606 2935 614
rect 2935 606 2936 614
rect 2940 606 2943 614
rect 2943 606 2945 614
rect 2945 606 2948 614
rect 2952 606 2953 614
rect 2953 606 2955 614
rect 2955 606 2960 614
rect 2964 606 2965 614
rect 2965 606 2972 614
rect 76 576 84 584
rect 2572 576 2580 584
rect 3756 596 3764 604
rect 3884 596 3892 604
rect 5924 606 5931 614
rect 5931 606 5932 614
rect 5936 606 5941 614
rect 5941 606 5943 614
rect 5943 606 5944 614
rect 5948 606 5951 614
rect 5951 606 5953 614
rect 5953 606 5956 614
rect 5960 606 5961 614
rect 5961 606 5963 614
rect 5963 606 5968 614
rect 5972 606 5973 614
rect 5973 606 5980 614
rect 5836 596 5844 604
rect 5804 576 5812 584
rect 6412 596 6420 604
rect 6700 596 6708 604
rect 3372 556 3380 564
rect 4812 556 4820 564
rect 5228 556 5236 564
rect 5676 556 5684 564
rect 4364 536 4372 544
rect 5740 536 5748 544
rect 7084 536 7092 544
rect 908 516 916 524
rect 2604 516 2612 524
rect 3884 516 3892 524
rect 5484 516 5492 524
rect 1132 496 1140 504
rect 4748 496 4756 504
rect 4780 496 4788 504
rect 5516 496 5524 504
rect 7084 496 7092 504
rect 428 476 436 484
rect 6988 476 6996 484
rect 588 456 596 464
rect 1996 456 2004 464
rect 5260 456 5268 464
rect 6028 456 6036 464
rect 3180 436 3188 444
rect 4556 436 4564 444
rect 5772 436 5780 444
rect 3532 416 3540 424
rect 4716 416 4724 424
rect 5836 416 5844 424
rect 1412 406 1419 414
rect 1419 406 1420 414
rect 1424 406 1429 414
rect 1429 406 1431 414
rect 1431 406 1432 414
rect 1436 406 1439 414
rect 1439 406 1441 414
rect 1441 406 1444 414
rect 1448 406 1449 414
rect 1449 406 1451 414
rect 1451 406 1456 414
rect 1460 406 1461 414
rect 1461 406 1468 414
rect 4420 406 4427 414
rect 4427 406 4428 414
rect 4432 406 4437 414
rect 4437 406 4439 414
rect 4439 406 4440 414
rect 4444 406 4447 414
rect 4447 406 4449 414
rect 4449 406 4452 414
rect 4456 406 4457 414
rect 4457 406 4459 414
rect 4459 406 4464 414
rect 4468 406 4469 414
rect 4469 406 4476 414
rect 1548 376 1556 384
rect 2028 376 2036 384
rect 4236 356 4244 364
rect 1964 336 1972 344
rect 2092 336 2100 344
rect 4364 316 4372 324
rect 4876 316 4884 324
rect 5548 316 5556 324
rect 5868 336 5876 344
rect 7276 316 7284 324
rect 76 296 84 304
rect 3052 296 3060 304
rect 3660 296 3668 304
rect 5324 296 5332 304
rect 1068 276 1076 284
rect 1516 276 1524 284
rect 1996 276 2004 284
rect 2028 276 2036 284
rect 5740 276 5748 284
rect 7180 276 7188 284
rect 5484 256 5492 264
rect 6156 256 6164 264
rect 6700 256 6708 264
rect 6188 216 6196 224
rect 2916 206 2923 214
rect 2923 206 2924 214
rect 2928 206 2933 214
rect 2933 206 2935 214
rect 2935 206 2936 214
rect 2940 206 2943 214
rect 2943 206 2945 214
rect 2945 206 2948 214
rect 2952 206 2953 214
rect 2953 206 2955 214
rect 2955 206 2960 214
rect 2964 206 2965 214
rect 2965 206 2972 214
rect 5924 206 5931 214
rect 5931 206 5932 214
rect 5936 206 5941 214
rect 5941 206 5943 214
rect 5943 206 5944 214
rect 5948 206 5951 214
rect 5951 206 5953 214
rect 5953 206 5956 214
rect 5960 206 5961 214
rect 5961 206 5963 214
rect 5963 206 5968 214
rect 5972 206 5973 214
rect 5973 206 5980 214
rect 748 196 756 204
rect 4364 196 4372 204
rect 5612 196 5620 204
rect 3660 176 3668 184
rect 6156 176 6164 184
rect 6188 176 6196 184
rect 204 156 212 164
rect 3276 156 3284 164
rect 5484 156 5492 164
rect 6700 176 6708 184
rect 268 136 276 144
rect 748 136 756 144
rect 1068 116 1076 124
rect 1516 116 1524 124
rect 1964 116 1972 124
rect 5612 136 5620 144
rect 6988 136 6996 144
rect 6220 96 6228 104
rect 7148 96 7156 104
rect 4716 76 4724 84
rect 4044 16 4052 24
rect 4236 16 4244 24
rect 4780 16 4788 24
rect 5068 16 5076 24
rect 6412 16 6420 24
rect 1412 6 1419 14
rect 1419 6 1420 14
rect 1424 6 1429 14
rect 1429 6 1431 14
rect 1431 6 1432 14
rect 1436 6 1439 14
rect 1439 6 1441 14
rect 1441 6 1444 14
rect 1448 6 1449 14
rect 1449 6 1451 14
rect 1451 6 1456 14
rect 1460 6 1461 14
rect 1461 6 1468 14
rect 4420 6 4427 14
rect 4427 6 4428 14
rect 4432 6 4437 14
rect 4437 6 4439 14
rect 4439 6 4440 14
rect 4444 6 4447 14
rect 4447 6 4449 14
rect 4449 6 4452 14
rect 4456 6 4457 14
rect 4457 6 4459 14
rect 4459 6 4464 14
rect 4468 6 4469 14
rect 4469 6 4476 14
<< metal4 >>
rect 970 5304 982 5306
rect 970 5296 972 5304
rect 980 5296 982 5304
rect 266 5264 278 5266
rect 266 5256 268 5264
rect 276 5256 278 5264
rect 266 5024 278 5256
rect 762 5124 822 5126
rect 762 5116 764 5124
rect 772 5116 822 5124
rect 762 5114 822 5116
rect 810 5104 822 5114
rect 810 5096 812 5104
rect 820 5096 822 5104
rect 810 5094 822 5096
rect 266 5016 268 5024
rect 276 5016 278 5024
rect 266 5014 278 5016
rect 970 5024 982 5296
rect 970 5016 972 5024
rect 980 5016 982 5024
rect 970 5014 982 5016
rect 1322 5224 1334 5226
rect 1322 5216 1324 5224
rect 1332 5216 1334 5224
rect 1034 4984 1046 4986
rect 1034 4976 1036 4984
rect 1044 4976 1046 4984
rect 1034 4944 1046 4976
rect 1034 4936 1036 4944
rect 1044 4936 1046 4944
rect 1034 4934 1046 4936
rect 1194 4884 1206 4886
rect 1194 4876 1196 4884
rect 1204 4876 1206 4884
rect 298 4704 310 4706
rect 298 4696 300 4704
rect 308 4696 310 4704
rect 298 4464 310 4696
rect 586 4624 598 4626
rect 586 4616 588 4624
rect 596 4616 598 4624
rect 298 4456 300 4464
rect 308 4456 310 4464
rect 298 4454 310 4456
rect 554 4464 566 4466
rect 554 4456 556 4464
rect 564 4456 566 4464
rect 458 4444 470 4446
rect 458 4436 460 4444
rect 468 4436 470 4444
rect 426 4344 438 4346
rect 426 4336 428 4344
rect 436 4336 438 4344
rect 106 4324 118 4326
rect 106 4316 108 4324
rect 116 4316 118 4324
rect 106 4164 118 4316
rect 106 4156 108 4164
rect 116 4156 118 4164
rect 106 4154 118 4156
rect 170 3944 182 3946
rect 170 3936 172 3944
rect 180 3936 182 3944
rect 138 3884 150 3886
rect 138 3876 140 3884
rect 148 3876 150 3884
rect 106 3324 118 3326
rect 106 3316 108 3324
rect 116 3316 118 3324
rect 106 2664 118 3316
rect 106 2656 108 2664
rect 116 2656 118 2664
rect 106 2654 118 2656
rect 42 2304 54 2306
rect 42 2296 44 2304
rect 52 2296 54 2304
rect 42 1664 54 2296
rect 42 1656 44 1664
rect 52 1656 54 1664
rect 42 1324 54 1656
rect 42 1316 44 1324
rect 52 1316 54 1324
rect 42 1314 54 1316
rect 138 644 150 3876
rect 170 3764 182 3936
rect 426 3884 438 4336
rect 426 3876 428 3884
rect 436 3876 438 3884
rect 426 3874 438 3876
rect 458 4044 470 4436
rect 458 4036 460 4044
rect 468 4036 470 4044
rect 170 3756 172 3764
rect 180 3756 182 3764
rect 170 3754 182 3756
rect 202 3784 214 3786
rect 202 3776 204 3784
rect 212 3776 214 3784
rect 170 2704 182 2706
rect 170 2696 172 2704
rect 180 2696 182 2704
rect 170 2244 182 2696
rect 202 2324 214 3776
rect 458 3744 470 4036
rect 458 3736 460 3744
rect 468 3736 470 3744
rect 458 3734 470 3736
rect 490 3484 502 3486
rect 490 3476 492 3484
rect 500 3476 502 3484
rect 490 3204 502 3476
rect 554 3424 566 4456
rect 586 4264 598 4616
rect 586 4256 588 4264
rect 596 4256 598 4264
rect 586 4254 598 4256
rect 1002 4604 1014 4606
rect 1002 4596 1004 4604
rect 1012 4596 1014 4604
rect 746 4184 758 4186
rect 746 4176 748 4184
rect 756 4176 758 4184
rect 746 4104 758 4176
rect 746 4096 748 4104
rect 756 4096 758 4104
rect 746 4094 758 4096
rect 810 3984 822 3986
rect 810 3976 812 3984
rect 820 3976 822 3984
rect 682 3904 694 3906
rect 682 3896 684 3904
rect 692 3896 694 3904
rect 682 3844 694 3896
rect 682 3836 684 3844
rect 692 3836 694 3844
rect 682 3834 694 3836
rect 618 3804 630 3806
rect 618 3796 620 3804
rect 628 3796 630 3804
rect 554 3416 556 3424
rect 564 3416 566 3424
rect 554 3414 566 3416
rect 586 3744 598 3746
rect 586 3736 588 3744
rect 596 3736 598 3744
rect 490 3196 492 3204
rect 500 3196 502 3204
rect 490 3194 502 3196
rect 554 3084 566 3086
rect 554 3076 556 3084
rect 564 3076 566 3084
rect 554 2884 566 3076
rect 554 2876 556 2884
rect 564 2876 566 2884
rect 554 2874 566 2876
rect 202 2316 204 2324
rect 212 2316 214 2324
rect 202 2314 214 2316
rect 490 2424 502 2426
rect 490 2416 492 2424
rect 500 2416 502 2424
rect 170 2236 172 2244
rect 180 2236 182 2244
rect 170 2234 182 2236
rect 426 2044 438 2046
rect 426 2036 428 2044
rect 436 2036 438 2044
rect 138 636 140 644
rect 148 636 150 644
rect 138 634 150 636
rect 202 744 214 746
rect 202 736 204 744
rect 212 736 214 744
rect 74 584 86 586
rect 74 576 76 584
rect 84 576 86 584
rect 74 304 86 576
rect 74 296 76 304
rect 84 296 86 304
rect 74 294 86 296
rect 202 164 214 736
rect 202 156 204 164
rect 212 156 214 164
rect 202 154 214 156
rect 266 724 278 726
rect 266 716 268 724
rect 276 716 278 724
rect 266 144 278 716
rect 426 484 438 2036
rect 490 1544 502 2416
rect 586 2344 598 3736
rect 618 3124 630 3796
rect 618 3116 620 3124
rect 628 3116 630 3124
rect 618 3114 630 3116
rect 682 3784 694 3786
rect 682 3776 684 3784
rect 692 3776 694 3784
rect 682 3104 694 3776
rect 810 3344 822 3976
rect 874 3904 886 3906
rect 874 3896 876 3904
rect 884 3896 886 3904
rect 874 3764 886 3896
rect 874 3756 876 3764
rect 884 3756 886 3764
rect 874 3754 886 3756
rect 970 3764 982 3766
rect 970 3756 972 3764
rect 980 3756 982 3764
rect 938 3684 950 3686
rect 938 3676 940 3684
rect 948 3676 950 3684
rect 810 3336 812 3344
rect 820 3336 822 3344
rect 810 3334 822 3336
rect 874 3484 886 3486
rect 874 3476 876 3484
rect 884 3476 886 3484
rect 874 3324 886 3476
rect 874 3316 876 3324
rect 884 3316 886 3324
rect 874 3314 886 3316
rect 906 3164 918 3166
rect 906 3156 908 3164
rect 916 3156 918 3164
rect 682 3096 684 3104
rect 692 3096 694 3104
rect 682 3094 694 3096
rect 746 3144 758 3146
rect 746 3136 748 3144
rect 756 3136 758 3144
rect 586 2336 588 2344
rect 596 2336 598 2344
rect 586 2334 598 2336
rect 650 2724 662 2726
rect 650 2716 652 2724
rect 660 2716 662 2724
rect 490 1536 492 1544
rect 500 1536 502 1544
rect 490 1534 502 1536
rect 586 2244 598 2246
rect 586 2236 588 2244
rect 596 2236 598 2244
rect 426 476 428 484
rect 436 476 438 484
rect 426 474 438 476
rect 586 464 598 2236
rect 650 1984 662 2716
rect 746 2484 758 3136
rect 842 3144 854 3146
rect 842 3136 844 3144
rect 852 3136 854 3144
rect 842 2904 854 3136
rect 842 2896 844 2904
rect 852 2896 854 2904
rect 842 2894 854 2896
rect 746 2476 748 2484
rect 756 2476 758 2484
rect 746 2474 758 2476
rect 650 1976 652 1984
rect 660 1976 662 1984
rect 650 1704 662 1976
rect 906 2084 918 3156
rect 906 2076 908 2084
rect 916 2076 918 2084
rect 650 1696 652 1704
rect 660 1696 662 1704
rect 650 1694 662 1696
rect 714 1944 726 1946
rect 714 1936 716 1944
rect 724 1936 726 1944
rect 714 1504 726 1936
rect 874 1584 886 1586
rect 874 1576 876 1584
rect 884 1576 886 1584
rect 714 1496 716 1504
rect 724 1496 726 1504
rect 714 1494 726 1496
rect 746 1544 758 1546
rect 746 1536 748 1544
rect 756 1536 758 1544
rect 746 704 758 1536
rect 874 1464 886 1576
rect 874 1456 876 1464
rect 884 1456 886 1464
rect 874 1454 886 1456
rect 906 1404 918 2076
rect 938 1424 950 3676
rect 970 3684 982 3756
rect 1002 3704 1014 4596
rect 1194 4524 1206 4876
rect 1258 4744 1270 4746
rect 1258 4736 1260 4744
rect 1268 4736 1270 4744
rect 1194 4516 1196 4524
rect 1204 4516 1206 4524
rect 1194 4514 1206 4516
rect 1226 4524 1238 4526
rect 1226 4516 1228 4524
rect 1236 4516 1238 4524
rect 1130 4504 1142 4506
rect 1130 4496 1132 4504
rect 1140 4496 1142 4504
rect 1098 4244 1110 4246
rect 1098 4236 1100 4244
rect 1108 4236 1110 4244
rect 1002 3696 1004 3704
rect 1012 3696 1014 3704
rect 1002 3694 1014 3696
rect 1066 4084 1078 4086
rect 1066 4076 1068 4084
rect 1076 4076 1078 4084
rect 970 3676 972 3684
rect 980 3676 982 3684
rect 970 3674 982 3676
rect 970 3584 982 3586
rect 970 3576 972 3584
rect 980 3576 982 3584
rect 970 3104 982 3576
rect 970 3096 972 3104
rect 980 3096 982 3104
rect 970 3094 982 3096
rect 1002 3344 1014 3346
rect 1002 3336 1004 3344
rect 1012 3336 1014 3344
rect 1002 2864 1014 3336
rect 1002 2856 1004 2864
rect 1012 2856 1014 2864
rect 1002 2854 1014 2856
rect 1034 2924 1046 2926
rect 1034 2916 1036 2924
rect 1044 2916 1046 2924
rect 1034 2724 1046 2916
rect 1066 2844 1078 4076
rect 1098 3944 1110 4236
rect 1130 4184 1142 4496
rect 1130 4176 1132 4184
rect 1140 4176 1142 4184
rect 1130 4174 1142 4176
rect 1194 4264 1206 4266
rect 1194 4256 1196 4264
rect 1204 4256 1206 4264
rect 1098 3936 1100 3944
rect 1108 3936 1110 3944
rect 1098 3934 1110 3936
rect 1194 3824 1206 4256
rect 1194 3816 1196 3824
rect 1204 3816 1206 3824
rect 1194 3814 1206 3816
rect 1066 2836 1068 2844
rect 1076 2836 1078 2844
rect 1066 2834 1078 2836
rect 1098 2844 1110 2846
rect 1098 2836 1100 2844
rect 1108 2836 1110 2844
rect 1034 2716 1036 2724
rect 1044 2716 1046 2724
rect 1034 2714 1046 2716
rect 1066 1564 1078 1566
rect 1066 1556 1068 1564
rect 1076 1556 1078 1564
rect 1034 1524 1046 1526
rect 1034 1516 1036 1524
rect 1044 1516 1046 1524
rect 938 1416 940 1424
rect 948 1416 950 1424
rect 938 1414 950 1416
rect 1002 1424 1014 1426
rect 1002 1416 1004 1424
rect 1012 1416 1014 1424
rect 906 1396 908 1404
rect 916 1396 918 1404
rect 906 1394 918 1396
rect 810 1364 822 1366
rect 810 1356 812 1364
rect 820 1356 822 1364
rect 810 1104 822 1356
rect 810 1096 812 1104
rect 820 1096 822 1104
rect 810 1094 822 1096
rect 842 1324 854 1326
rect 842 1316 844 1324
rect 852 1316 854 1324
rect 842 1084 854 1316
rect 874 1204 886 1206
rect 874 1196 876 1204
rect 884 1196 886 1204
rect 874 1126 886 1196
rect 874 1114 918 1126
rect 906 1104 918 1114
rect 906 1096 908 1104
rect 916 1096 918 1104
rect 906 1094 918 1096
rect 938 1124 950 1126
rect 938 1116 940 1124
rect 948 1116 950 1124
rect 842 1076 844 1084
rect 852 1076 854 1084
rect 842 1074 854 1076
rect 938 1004 950 1116
rect 938 996 940 1004
rect 948 996 950 1004
rect 938 994 950 996
rect 746 696 748 704
rect 756 696 758 704
rect 746 694 758 696
rect 906 704 918 706
rect 906 696 908 704
rect 916 696 918 704
rect 906 524 918 696
rect 1002 624 1014 1416
rect 1034 1124 1046 1516
rect 1066 1484 1078 1556
rect 1066 1476 1068 1484
rect 1076 1476 1078 1484
rect 1066 1474 1078 1476
rect 1098 1384 1110 2836
rect 1162 2264 1174 2266
rect 1162 2256 1164 2264
rect 1172 2256 1174 2264
rect 1162 2164 1174 2256
rect 1162 2156 1164 2164
rect 1172 2156 1174 2164
rect 1162 2154 1174 2156
rect 1194 2184 1206 2186
rect 1194 2176 1196 2184
rect 1204 2176 1206 2184
rect 1162 1924 1174 1926
rect 1162 1916 1164 1924
rect 1172 1916 1174 1924
rect 1098 1376 1100 1384
rect 1108 1376 1110 1384
rect 1098 1374 1110 1376
rect 1130 1644 1142 1646
rect 1130 1636 1132 1644
rect 1140 1636 1142 1644
rect 1034 1116 1036 1124
rect 1044 1116 1046 1124
rect 1034 1114 1046 1116
rect 1130 1124 1142 1636
rect 1162 1544 1174 1916
rect 1162 1536 1164 1544
rect 1172 1536 1174 1544
rect 1162 1304 1174 1536
rect 1162 1296 1164 1304
rect 1172 1296 1174 1304
rect 1162 1294 1174 1296
rect 1130 1116 1132 1124
rect 1140 1116 1142 1124
rect 1130 1114 1142 1116
rect 1002 616 1004 624
rect 1012 616 1014 624
rect 1002 614 1014 616
rect 1130 984 1142 986
rect 1130 976 1132 984
rect 1140 976 1142 984
rect 906 516 908 524
rect 916 516 918 524
rect 906 514 918 516
rect 1130 504 1142 976
rect 1194 784 1206 2176
rect 1226 2184 1238 4516
rect 1258 3144 1270 4736
rect 1290 4544 1302 4546
rect 1290 4536 1292 4544
rect 1300 4536 1302 4544
rect 1290 3784 1302 4536
rect 1322 4084 1334 5216
rect 1322 4076 1324 4084
rect 1332 4076 1334 4084
rect 1322 4074 1334 4076
rect 1408 5214 1472 5416
rect 2912 5414 2976 5416
rect 2912 5406 2916 5414
rect 2924 5406 2928 5414
rect 2936 5406 2940 5414
rect 2948 5406 2952 5414
rect 2960 5406 2964 5414
rect 2972 5406 2976 5414
rect 1408 5206 1412 5214
rect 1420 5206 1424 5214
rect 1432 5206 1436 5214
rect 1444 5206 1448 5214
rect 1456 5206 1460 5214
rect 1468 5206 1472 5214
rect 1408 4814 1472 5206
rect 1578 5304 1590 5306
rect 1578 5296 1580 5304
rect 1588 5296 1590 5304
rect 1578 5204 1590 5296
rect 1578 5196 1580 5204
rect 1588 5196 1590 5204
rect 1578 5194 1590 5196
rect 2058 5164 2070 5166
rect 2058 5156 2060 5164
rect 2068 5156 2070 5164
rect 1642 5144 1654 5146
rect 1642 5136 1644 5144
rect 1652 5136 1654 5144
rect 1642 4984 1654 5136
rect 1866 5104 1878 5106
rect 1866 5096 1868 5104
rect 1876 5096 1878 5104
rect 1802 5084 1814 5086
rect 1802 5076 1804 5084
rect 1812 5076 1814 5084
rect 1738 5064 1750 5066
rect 1738 5056 1740 5064
rect 1748 5056 1750 5064
rect 1738 5024 1750 5056
rect 1738 5016 1740 5024
rect 1748 5016 1750 5024
rect 1738 5014 1750 5016
rect 1642 4976 1644 4984
rect 1652 4976 1654 4984
rect 1642 4974 1654 4976
rect 1408 4806 1412 4814
rect 1420 4806 1424 4814
rect 1432 4806 1436 4814
rect 1444 4806 1448 4814
rect 1456 4806 1460 4814
rect 1468 4806 1472 4814
rect 1408 4414 1472 4806
rect 1802 4904 1814 5076
rect 1802 4896 1804 4904
rect 1812 4896 1814 4904
rect 1610 4684 1622 4686
rect 1610 4676 1612 4684
rect 1620 4676 1622 4684
rect 1578 4584 1590 4586
rect 1578 4576 1580 4584
rect 1588 4576 1590 4584
rect 1408 4406 1412 4414
rect 1420 4406 1424 4414
rect 1432 4406 1436 4414
rect 1444 4406 1448 4414
rect 1456 4406 1460 4414
rect 1468 4406 1472 4414
rect 1290 3776 1292 3784
rect 1300 3776 1302 3784
rect 1290 3774 1302 3776
rect 1408 4014 1472 4406
rect 1546 4504 1558 4506
rect 1546 4496 1548 4504
rect 1556 4496 1558 4504
rect 1546 4144 1558 4496
rect 1546 4136 1548 4144
rect 1556 4136 1558 4144
rect 1546 4064 1558 4136
rect 1546 4056 1548 4064
rect 1556 4056 1558 4064
rect 1546 4054 1558 4056
rect 1408 4006 1412 4014
rect 1420 4006 1424 4014
rect 1432 4006 1436 4014
rect 1444 4006 1448 4014
rect 1456 4006 1460 4014
rect 1468 4006 1472 4014
rect 1290 3644 1302 3646
rect 1290 3636 1292 3644
rect 1300 3636 1302 3644
rect 1290 3344 1302 3636
rect 1290 3336 1292 3344
rect 1300 3336 1302 3344
rect 1290 3334 1302 3336
rect 1322 3644 1334 3646
rect 1322 3636 1324 3644
rect 1332 3636 1334 3644
rect 1322 3164 1334 3636
rect 1322 3156 1324 3164
rect 1332 3156 1334 3164
rect 1322 3154 1334 3156
rect 1408 3614 1472 4006
rect 1408 3606 1412 3614
rect 1420 3606 1424 3614
rect 1432 3606 1436 3614
rect 1444 3606 1448 3614
rect 1456 3606 1460 3614
rect 1468 3606 1472 3614
rect 1408 3214 1472 3606
rect 1408 3206 1412 3214
rect 1420 3206 1424 3214
rect 1432 3206 1436 3214
rect 1444 3206 1448 3214
rect 1456 3206 1460 3214
rect 1468 3206 1472 3214
rect 1258 3136 1260 3144
rect 1268 3136 1270 3144
rect 1258 3134 1270 3136
rect 1290 3144 1302 3146
rect 1290 3136 1292 3144
rect 1300 3136 1302 3144
rect 1258 3104 1270 3106
rect 1258 3096 1260 3104
rect 1268 3096 1270 3104
rect 1258 2924 1270 3096
rect 1258 2916 1260 2924
rect 1268 2916 1270 2924
rect 1258 2914 1270 2916
rect 1290 2444 1302 3136
rect 1354 3144 1366 3146
rect 1354 3136 1356 3144
rect 1364 3136 1366 3144
rect 1290 2436 1292 2444
rect 1300 2436 1302 2444
rect 1290 2434 1302 2436
rect 1322 2944 1334 2946
rect 1322 2936 1324 2944
rect 1332 2936 1334 2944
rect 1322 2244 1334 2936
rect 1354 2924 1366 3136
rect 1354 2916 1356 2924
rect 1364 2916 1366 2924
rect 1354 2914 1366 2916
rect 1322 2236 1324 2244
rect 1332 2236 1334 2244
rect 1322 2234 1334 2236
rect 1408 2814 1472 3206
rect 1514 3504 1526 3506
rect 1514 3496 1516 3504
rect 1524 3496 1526 3504
rect 1514 3204 1526 3496
rect 1514 3196 1516 3204
rect 1524 3196 1526 3204
rect 1514 3194 1526 3196
rect 1408 2806 1412 2814
rect 1420 2806 1424 2814
rect 1432 2806 1436 2814
rect 1444 2806 1448 2814
rect 1456 2806 1460 2814
rect 1468 2806 1472 2814
rect 1408 2414 1472 2806
rect 1408 2406 1412 2414
rect 1420 2406 1424 2414
rect 1432 2406 1436 2414
rect 1444 2406 1448 2414
rect 1456 2406 1460 2414
rect 1468 2406 1472 2414
rect 1226 2176 1228 2184
rect 1236 2176 1238 2184
rect 1226 2174 1238 2176
rect 1408 2014 1472 2406
rect 1408 2006 1412 2014
rect 1420 2006 1424 2014
rect 1432 2006 1436 2014
rect 1444 2006 1448 2014
rect 1456 2006 1460 2014
rect 1468 2006 1472 2014
rect 1546 3104 1558 3106
rect 1546 3096 1548 3104
rect 1556 3096 1558 3104
rect 1546 2124 1558 3096
rect 1578 2944 1590 4576
rect 1610 3744 1622 4676
rect 1802 4644 1814 4896
rect 1802 4636 1804 4644
rect 1812 4636 1814 4644
rect 1802 4634 1814 4636
rect 1866 4624 1878 5096
rect 1962 5104 1974 5106
rect 1962 5096 1964 5104
rect 1972 5096 1974 5104
rect 1962 4804 1974 5096
rect 2026 5084 2038 5086
rect 2026 5076 2028 5084
rect 2036 5076 2038 5084
rect 1994 5044 2006 5046
rect 1994 5036 1996 5044
rect 2004 5036 2006 5044
rect 1994 4864 2006 5036
rect 1994 4856 1996 4864
rect 2004 4856 2006 4864
rect 1994 4854 2006 4856
rect 1962 4796 1964 4804
rect 1972 4796 1974 4804
rect 1962 4794 1974 4796
rect 2026 4744 2038 5076
rect 2026 4736 2028 4744
rect 2036 4736 2038 4744
rect 2026 4734 2038 4736
rect 1866 4616 1868 4624
rect 1876 4616 1878 4624
rect 1866 4614 1878 4616
rect 1994 4704 2006 4706
rect 1994 4696 1996 4704
rect 2004 4696 2006 4704
rect 1994 4664 2006 4696
rect 1994 4656 1996 4664
rect 2004 4656 2006 4664
rect 1674 4544 1686 4546
rect 1674 4536 1676 4544
rect 1684 4536 1686 4544
rect 1674 4144 1686 4536
rect 1674 4136 1676 4144
rect 1684 4136 1686 4144
rect 1674 4134 1686 4136
rect 1866 4384 1878 4386
rect 1866 4376 1868 4384
rect 1876 4376 1878 4384
rect 1610 3736 1612 3744
rect 1620 3736 1622 3744
rect 1610 3734 1622 3736
rect 1834 4084 1846 4086
rect 1834 4076 1836 4084
rect 1844 4076 1846 4084
rect 1834 3724 1846 4076
rect 1866 3764 1878 4376
rect 1866 3756 1868 3764
rect 1876 3756 1878 3764
rect 1866 3754 1878 3756
rect 1930 4104 1942 4106
rect 1930 4096 1932 4104
rect 1940 4096 1942 4104
rect 1834 3716 1836 3724
rect 1844 3716 1846 3724
rect 1834 3714 1846 3716
rect 1642 3464 1654 3466
rect 1642 3456 1644 3464
rect 1652 3456 1654 3464
rect 1610 3424 1622 3426
rect 1610 3416 1612 3424
rect 1620 3416 1622 3424
rect 1610 3104 1622 3416
rect 1642 3344 1654 3456
rect 1642 3336 1644 3344
rect 1652 3336 1654 3344
rect 1642 3334 1654 3336
rect 1866 3284 1878 3286
rect 1866 3276 1868 3284
rect 1876 3276 1878 3284
rect 1610 3096 1612 3104
rect 1620 3096 1622 3104
rect 1610 3094 1622 3096
rect 1738 3184 1750 3186
rect 1738 3176 1740 3184
rect 1748 3176 1750 3184
rect 1578 2936 1580 2944
rect 1588 2936 1590 2944
rect 1578 2934 1590 2936
rect 1610 3064 1622 3066
rect 1610 3056 1612 3064
rect 1620 3056 1622 3064
rect 1610 2344 1622 3056
rect 1738 3004 1750 3176
rect 1770 3124 1782 3126
rect 1770 3116 1772 3124
rect 1780 3116 1782 3124
rect 1770 3064 1782 3116
rect 1770 3056 1772 3064
rect 1780 3056 1782 3064
rect 1770 3054 1782 3056
rect 1802 3124 1814 3126
rect 1802 3116 1804 3124
rect 1812 3116 1814 3124
rect 1738 2996 1740 3004
rect 1748 2996 1750 3004
rect 1738 2994 1750 2996
rect 1802 2964 1814 3116
rect 1802 2956 1804 2964
rect 1812 2956 1814 2964
rect 1802 2954 1814 2956
rect 1834 2964 1846 2966
rect 1834 2956 1836 2964
rect 1844 2956 1846 2964
rect 1834 2926 1846 2956
rect 1706 2914 1846 2926
rect 1706 2884 1718 2914
rect 1706 2876 1708 2884
rect 1716 2876 1718 2884
rect 1706 2874 1718 2876
rect 1738 2884 1750 2886
rect 1738 2876 1740 2884
rect 1748 2876 1750 2884
rect 1706 2464 1718 2466
rect 1706 2456 1708 2464
rect 1716 2456 1718 2464
rect 1674 2384 1686 2386
rect 1674 2376 1676 2384
rect 1684 2376 1686 2384
rect 1610 2336 1612 2344
rect 1620 2336 1622 2344
rect 1610 2334 1622 2336
rect 1642 2364 1654 2366
rect 1642 2356 1644 2364
rect 1652 2356 1654 2364
rect 1546 2116 1548 2124
rect 1556 2116 1558 2124
rect 1226 1704 1238 1706
rect 1226 1696 1228 1704
rect 1236 1696 1238 1704
rect 1226 1364 1238 1696
rect 1322 1624 1334 1626
rect 1322 1616 1324 1624
rect 1332 1616 1334 1624
rect 1322 1424 1334 1616
rect 1322 1416 1324 1424
rect 1332 1416 1334 1424
rect 1322 1414 1334 1416
rect 1408 1614 1472 2006
rect 1514 2004 1526 2006
rect 1514 1996 1516 2004
rect 1524 1996 1526 2004
rect 1514 1964 1526 1996
rect 1514 1956 1516 1964
rect 1524 1956 1526 1964
rect 1514 1954 1526 1956
rect 1408 1606 1412 1614
rect 1420 1606 1424 1614
rect 1432 1606 1436 1614
rect 1444 1606 1448 1614
rect 1456 1606 1460 1614
rect 1468 1606 1472 1614
rect 1226 1356 1228 1364
rect 1236 1356 1238 1364
rect 1226 1354 1238 1356
rect 1408 1214 1472 1606
rect 1408 1206 1412 1214
rect 1420 1206 1424 1214
rect 1432 1206 1436 1214
rect 1444 1206 1448 1214
rect 1456 1206 1460 1214
rect 1468 1206 1472 1214
rect 1322 1164 1334 1166
rect 1322 1156 1324 1164
rect 1332 1156 1334 1164
rect 1322 1024 1334 1156
rect 1322 1016 1324 1024
rect 1332 1016 1334 1024
rect 1322 1014 1334 1016
rect 1194 776 1196 784
rect 1204 776 1206 784
rect 1194 774 1206 776
rect 1408 814 1472 1206
rect 1408 806 1412 814
rect 1420 806 1424 814
rect 1432 806 1436 814
rect 1444 806 1448 814
rect 1456 806 1460 814
rect 1468 806 1472 814
rect 1130 496 1132 504
rect 1140 496 1142 504
rect 1130 494 1142 496
rect 586 456 588 464
rect 596 456 598 464
rect 586 454 598 456
rect 1408 414 1472 806
rect 1408 406 1412 414
rect 1420 406 1424 414
rect 1432 406 1436 414
rect 1444 406 1448 414
rect 1456 406 1460 414
rect 1468 406 1472 414
rect 1066 284 1078 286
rect 1066 276 1068 284
rect 1076 276 1078 284
rect 266 136 268 144
rect 276 136 278 144
rect 266 134 278 136
rect 746 204 758 206
rect 746 196 748 204
rect 756 196 758 204
rect 746 144 758 196
rect 746 136 748 144
rect 756 136 758 144
rect 746 134 758 136
rect 1066 124 1078 276
rect 1066 116 1068 124
rect 1076 116 1078 124
rect 1066 114 1078 116
rect 1408 14 1472 406
rect 1514 1844 1526 1846
rect 1514 1836 1516 1844
rect 1524 1836 1526 1844
rect 1514 284 1526 1836
rect 1546 384 1558 2116
rect 1610 2244 1622 2246
rect 1610 2236 1612 2244
rect 1620 2236 1622 2244
rect 1610 2144 1622 2236
rect 1610 2136 1612 2144
rect 1620 2136 1622 2144
rect 1610 1864 1622 2136
rect 1610 1856 1612 1864
rect 1620 1856 1622 1864
rect 1610 1854 1622 1856
rect 1642 1784 1654 2356
rect 1642 1776 1644 1784
rect 1652 1776 1654 1784
rect 1642 1774 1654 1776
rect 1610 1504 1622 1506
rect 1610 1496 1612 1504
rect 1620 1496 1622 1504
rect 1578 1044 1590 1046
rect 1578 1036 1580 1044
rect 1588 1036 1590 1044
rect 1578 844 1590 1036
rect 1578 836 1580 844
rect 1588 836 1590 844
rect 1578 834 1590 836
rect 1610 744 1622 1496
rect 1674 1324 1686 2376
rect 1706 2064 1718 2456
rect 1706 2056 1708 2064
rect 1716 2056 1718 2064
rect 1706 2054 1718 2056
rect 1738 2424 1750 2876
rect 1834 2744 1846 2746
rect 1834 2736 1836 2744
rect 1844 2736 1846 2744
rect 1834 2664 1846 2736
rect 1834 2656 1836 2664
rect 1844 2656 1846 2664
rect 1834 2654 1846 2656
rect 1866 2504 1878 3276
rect 1866 2496 1868 2504
rect 1876 2496 1878 2504
rect 1866 2494 1878 2496
rect 1898 2704 1910 2706
rect 1898 2696 1900 2704
rect 1908 2696 1910 2704
rect 1738 2416 1740 2424
rect 1748 2416 1750 2424
rect 1706 2024 1718 2026
rect 1706 2016 1708 2024
rect 1716 2016 1718 2024
rect 1706 1884 1718 2016
rect 1706 1876 1708 1884
rect 1716 1876 1718 1884
rect 1706 1874 1718 1876
rect 1706 1644 1718 1646
rect 1706 1636 1708 1644
rect 1716 1636 1718 1644
rect 1706 1364 1718 1636
rect 1706 1356 1708 1364
rect 1716 1356 1718 1364
rect 1706 1354 1718 1356
rect 1738 1564 1750 2416
rect 1898 2404 1910 2696
rect 1898 2396 1900 2404
rect 1908 2396 1910 2404
rect 1898 2394 1910 2396
rect 1898 2304 1910 2306
rect 1898 2296 1900 2304
rect 1908 2296 1910 2304
rect 1770 2204 1782 2206
rect 1770 2196 1772 2204
rect 1780 2196 1782 2204
rect 1770 2124 1782 2196
rect 1898 2164 1910 2296
rect 1898 2156 1900 2164
rect 1908 2156 1910 2164
rect 1898 2154 1910 2156
rect 1770 2116 1772 2124
rect 1780 2116 1782 2124
rect 1770 2114 1782 2116
rect 1866 2024 1878 2026
rect 1866 2016 1868 2024
rect 1876 2016 1878 2024
rect 1738 1556 1740 1564
rect 1748 1556 1750 1564
rect 1674 1316 1676 1324
rect 1684 1316 1686 1324
rect 1674 1314 1686 1316
rect 1706 1324 1718 1326
rect 1706 1316 1708 1324
rect 1716 1316 1718 1324
rect 1706 844 1718 1316
rect 1738 1304 1750 1556
rect 1738 1296 1740 1304
rect 1748 1296 1750 1304
rect 1738 1294 1750 1296
rect 1770 1824 1782 1826
rect 1770 1816 1772 1824
rect 1780 1816 1782 1824
rect 1770 1264 1782 1816
rect 1834 1724 1846 1726
rect 1834 1716 1836 1724
rect 1844 1716 1846 1724
rect 1770 1256 1772 1264
rect 1780 1256 1782 1264
rect 1770 1254 1782 1256
rect 1802 1524 1814 1526
rect 1802 1516 1804 1524
rect 1812 1516 1814 1524
rect 1770 1224 1782 1226
rect 1770 1216 1772 1224
rect 1780 1216 1782 1224
rect 1738 1064 1750 1066
rect 1738 1056 1740 1064
rect 1748 1056 1750 1064
rect 1738 984 1750 1056
rect 1738 976 1740 984
rect 1748 976 1750 984
rect 1738 974 1750 976
rect 1770 904 1782 1216
rect 1802 1224 1814 1516
rect 1834 1264 1846 1716
rect 1866 1624 1878 2016
rect 1866 1616 1868 1624
rect 1876 1616 1878 1624
rect 1866 1614 1878 1616
rect 1930 1464 1942 4096
rect 1962 4084 1974 4086
rect 1962 4076 1964 4084
rect 1972 4076 1974 4084
rect 1962 3264 1974 4076
rect 1994 3984 2006 4656
rect 1994 3976 1996 3984
rect 2004 3976 2006 3984
rect 1994 3974 2006 3976
rect 2058 3924 2070 5156
rect 2912 5014 2976 5406
rect 4106 5344 4118 5346
rect 4106 5336 4108 5344
rect 4116 5336 4118 5344
rect 3978 5304 3990 5306
rect 3978 5296 3980 5304
rect 3988 5296 3990 5304
rect 3466 5164 3478 5166
rect 3466 5156 3468 5164
rect 3476 5156 3478 5164
rect 3466 5124 3478 5156
rect 3466 5116 3468 5124
rect 3476 5116 3478 5124
rect 3466 5114 3478 5116
rect 3754 5164 3766 5166
rect 3754 5156 3756 5164
rect 3764 5156 3766 5164
rect 2912 5006 2916 5014
rect 2924 5006 2928 5014
rect 2936 5006 2940 5014
rect 2948 5006 2952 5014
rect 2960 5006 2964 5014
rect 2972 5006 2976 5014
rect 2506 4964 2518 4966
rect 2506 4956 2508 4964
rect 2516 4956 2518 4964
rect 2314 4944 2326 4946
rect 2314 4936 2316 4944
rect 2324 4936 2326 4944
rect 2186 4744 2198 4746
rect 2186 4736 2188 4744
rect 2196 4736 2198 4744
rect 2154 4724 2166 4726
rect 2154 4716 2156 4724
rect 2164 4716 2166 4724
rect 2154 4684 2166 4716
rect 2154 4676 2156 4684
rect 2164 4676 2166 4684
rect 2154 4674 2166 4676
rect 2154 4444 2166 4446
rect 2154 4436 2156 4444
rect 2164 4436 2166 4444
rect 2058 3916 2060 3924
rect 2068 3916 2070 3924
rect 2058 3914 2070 3916
rect 2090 4004 2102 4006
rect 2090 3996 2092 4004
rect 2100 3996 2102 4004
rect 1962 3256 1964 3264
rect 1972 3256 1974 3264
rect 1962 3254 1974 3256
rect 1994 3264 2006 3266
rect 1994 3256 1996 3264
rect 2004 3256 2006 3264
rect 1962 3124 1974 3126
rect 1962 3116 1964 3124
rect 1972 3116 1974 3124
rect 1962 2884 1974 3116
rect 1962 2876 1964 2884
rect 1972 2876 1974 2884
rect 1962 2874 1974 2876
rect 1930 1456 1932 1464
rect 1940 1456 1942 1464
rect 1930 1454 1942 1456
rect 1962 2164 1974 2166
rect 1962 2156 1964 2164
rect 1972 2156 1974 2164
rect 1834 1256 1836 1264
rect 1844 1256 1846 1264
rect 1834 1254 1846 1256
rect 1802 1216 1804 1224
rect 1812 1216 1814 1224
rect 1802 1214 1814 1216
rect 1930 1144 1942 1146
rect 1930 1136 1932 1144
rect 1940 1136 1942 1144
rect 1930 1064 1942 1136
rect 1962 1144 1974 2156
rect 1994 1564 2006 3256
rect 2090 3144 2102 3996
rect 2154 3724 2166 4436
rect 2186 4344 2198 4736
rect 2186 4336 2188 4344
rect 2196 4336 2198 4344
rect 2186 4334 2198 4336
rect 2314 4264 2326 4936
rect 2314 4256 2316 4264
rect 2324 4256 2326 4264
rect 2314 4254 2326 4256
rect 2442 4944 2454 4946
rect 2442 4936 2444 4944
rect 2452 4936 2454 4944
rect 2442 4064 2454 4936
rect 2442 4056 2444 4064
rect 2452 4056 2454 4064
rect 2442 4054 2454 4056
rect 2506 4544 2518 4956
rect 2762 4804 2774 4806
rect 2762 4796 2764 4804
rect 2772 4796 2774 4804
rect 2762 4764 2774 4796
rect 2762 4756 2764 4764
rect 2772 4756 2774 4764
rect 2762 4754 2774 4756
rect 2506 4536 2508 4544
rect 2516 4536 2518 4544
rect 2346 3924 2358 3926
rect 2346 3916 2348 3924
rect 2356 3916 2358 3924
rect 2154 3716 2156 3724
rect 2164 3716 2166 3724
rect 2154 3714 2166 3716
rect 2314 3764 2326 3766
rect 2314 3756 2316 3764
rect 2324 3756 2326 3764
rect 2090 3136 2092 3144
rect 2100 3136 2102 3144
rect 2090 3134 2102 3136
rect 2154 3504 2166 3506
rect 2154 3496 2156 3504
rect 2164 3496 2166 3504
rect 2154 3204 2166 3496
rect 2154 3196 2156 3204
rect 2164 3196 2166 3204
rect 2154 2924 2166 3196
rect 2154 2916 2156 2924
rect 2164 2916 2166 2924
rect 2154 2914 2166 2916
rect 2218 3124 2230 3126
rect 2218 3116 2220 3124
rect 2228 3116 2230 3124
rect 2218 2904 2230 3116
rect 2218 2896 2220 2904
rect 2228 2896 2230 2904
rect 2218 2484 2230 2896
rect 2282 2964 2294 2966
rect 2282 2956 2284 2964
rect 2292 2956 2294 2964
rect 2282 2584 2294 2956
rect 2282 2576 2284 2584
rect 2292 2576 2294 2584
rect 2282 2574 2294 2576
rect 2314 2544 2326 3756
rect 2346 3524 2358 3916
rect 2506 3884 2518 4536
rect 2912 4614 2976 5006
rect 2912 4606 2916 4614
rect 2924 4606 2928 4614
rect 2936 4606 2940 4614
rect 2948 4606 2952 4614
rect 2960 4606 2964 4614
rect 2972 4606 2976 4614
rect 2570 4484 2582 4486
rect 2570 4476 2572 4484
rect 2580 4476 2582 4484
rect 2506 3876 2508 3884
rect 2516 3876 2518 3884
rect 2346 3516 2348 3524
rect 2356 3516 2358 3524
rect 2346 3514 2358 3516
rect 2474 3564 2486 3566
rect 2474 3556 2476 3564
rect 2484 3556 2486 3564
rect 2378 3504 2390 3506
rect 2378 3496 2380 3504
rect 2388 3496 2390 3504
rect 2378 3104 2390 3496
rect 2474 3364 2486 3556
rect 2474 3356 2476 3364
rect 2484 3356 2486 3364
rect 2474 3354 2486 3356
rect 2506 3244 2518 3876
rect 2538 4164 2550 4166
rect 2538 4156 2540 4164
rect 2548 4156 2550 4164
rect 2538 3744 2550 4156
rect 2538 3736 2540 3744
rect 2548 3736 2550 3744
rect 2538 3734 2550 3736
rect 2570 3564 2582 4476
rect 2912 4214 2976 4606
rect 3146 5104 3158 5106
rect 3146 5096 3148 5104
rect 3156 5096 3158 5104
rect 3146 4504 3158 5096
rect 3370 5104 3382 5106
rect 3370 5096 3372 5104
rect 3380 5096 3382 5104
rect 3178 5004 3190 5006
rect 3178 4996 3180 5004
rect 3188 4996 3190 5004
rect 3178 4924 3190 4996
rect 3178 4916 3180 4924
rect 3188 4916 3190 4924
rect 3178 4914 3190 4916
rect 3370 4904 3382 5096
rect 3434 5104 3446 5106
rect 3434 5096 3436 5104
rect 3444 5096 3446 5104
rect 3434 5086 3446 5096
rect 3722 5104 3734 5106
rect 3722 5096 3724 5104
rect 3732 5096 3734 5104
rect 3434 5074 3510 5086
rect 3498 5064 3510 5074
rect 3498 5056 3500 5064
rect 3508 5056 3510 5064
rect 3498 5054 3510 5056
rect 3658 5084 3670 5086
rect 3658 5076 3660 5084
rect 3668 5076 3670 5084
rect 3370 4896 3372 4904
rect 3380 4896 3382 4904
rect 3370 4894 3382 4896
rect 3658 4904 3670 5076
rect 3658 4896 3660 4904
rect 3668 4896 3670 4904
rect 3658 4894 3670 4896
rect 3146 4496 3148 4504
rect 3156 4496 3158 4504
rect 3146 4494 3158 4496
rect 3370 4844 3382 4846
rect 3370 4836 3372 4844
rect 3380 4836 3382 4844
rect 2912 4206 2916 4214
rect 2924 4206 2928 4214
rect 2936 4206 2940 4214
rect 2948 4206 2952 4214
rect 2960 4206 2964 4214
rect 2972 4206 2976 4214
rect 2634 4124 2646 4126
rect 2634 4116 2636 4124
rect 2644 4116 2646 4124
rect 2570 3556 2572 3564
rect 2580 3556 2582 3564
rect 2570 3554 2582 3556
rect 2602 3744 2614 3746
rect 2602 3736 2604 3744
rect 2612 3736 2614 3744
rect 2506 3236 2508 3244
rect 2516 3236 2518 3244
rect 2506 3234 2518 3236
rect 2378 3096 2380 3104
rect 2388 3096 2390 3104
rect 2378 3094 2390 3096
rect 2506 3104 2518 3106
rect 2506 3096 2508 3104
rect 2516 3096 2518 3104
rect 2314 2536 2316 2544
rect 2324 2536 2326 2544
rect 2314 2534 2326 2536
rect 2346 3084 2358 3086
rect 2346 3076 2348 3084
rect 2356 3076 2358 3084
rect 2218 2476 2220 2484
rect 2228 2476 2230 2484
rect 2218 2474 2230 2476
rect 2186 2464 2198 2466
rect 2186 2456 2188 2464
rect 2196 2456 2198 2464
rect 2154 2104 2166 2106
rect 2154 2096 2156 2104
rect 2164 2096 2166 2104
rect 2122 2024 2134 2026
rect 2122 2016 2124 2024
rect 2132 2016 2134 2024
rect 2090 1864 2102 1866
rect 2090 1856 2092 1864
rect 2100 1856 2102 1864
rect 2090 1704 2102 1856
rect 2090 1696 2092 1704
rect 2100 1696 2102 1704
rect 2090 1694 2102 1696
rect 1994 1556 1996 1564
rect 2004 1556 2006 1564
rect 1994 1554 2006 1556
rect 2090 1624 2102 1626
rect 2090 1616 2092 1624
rect 2100 1616 2102 1624
rect 2058 1544 2070 1546
rect 2058 1536 2060 1544
rect 2068 1536 2070 1544
rect 1994 1504 2006 1506
rect 1994 1496 1996 1504
rect 2004 1496 2006 1504
rect 1994 1324 2006 1496
rect 1994 1316 1996 1324
rect 2004 1316 2006 1324
rect 1994 1314 2006 1316
rect 2026 1384 2038 1386
rect 2026 1376 2028 1384
rect 2036 1376 2038 1384
rect 1962 1136 1964 1144
rect 1972 1136 1974 1144
rect 1962 1134 1974 1136
rect 1994 1164 2006 1166
rect 1994 1156 1996 1164
rect 2004 1156 2006 1164
rect 1994 1126 2006 1156
rect 2026 1164 2038 1376
rect 2058 1324 2070 1536
rect 2090 1484 2102 1616
rect 2122 1624 2134 2016
rect 2154 1724 2166 2096
rect 2186 1984 2198 2456
rect 2282 2384 2294 2386
rect 2282 2376 2284 2384
rect 2292 2376 2294 2384
rect 2282 2144 2294 2376
rect 2282 2136 2284 2144
rect 2292 2136 2294 2144
rect 2282 2134 2294 2136
rect 2346 2144 2358 3076
rect 2410 2924 2422 2926
rect 2410 2916 2412 2924
rect 2420 2916 2422 2924
rect 2378 2764 2390 2766
rect 2378 2756 2380 2764
rect 2388 2756 2390 2764
rect 2378 2364 2390 2756
rect 2378 2356 2380 2364
rect 2388 2356 2390 2364
rect 2378 2354 2390 2356
rect 2410 2304 2422 2916
rect 2410 2296 2412 2304
rect 2420 2296 2422 2304
rect 2410 2294 2422 2296
rect 2442 2904 2454 2906
rect 2442 2896 2444 2904
rect 2452 2896 2454 2904
rect 2442 2304 2454 2896
rect 2506 2724 2518 3096
rect 2506 2716 2508 2724
rect 2516 2716 2518 2724
rect 2506 2714 2518 2716
rect 2570 3024 2582 3026
rect 2570 3016 2572 3024
rect 2580 3016 2582 3024
rect 2474 2644 2486 2646
rect 2474 2636 2476 2644
rect 2484 2636 2486 2644
rect 2474 2604 2486 2636
rect 2474 2596 2476 2604
rect 2484 2596 2486 2604
rect 2474 2594 2486 2596
rect 2442 2296 2444 2304
rect 2452 2296 2454 2304
rect 2442 2294 2454 2296
rect 2346 2136 2348 2144
rect 2356 2136 2358 2144
rect 2346 2134 2358 2136
rect 2378 2264 2390 2266
rect 2378 2256 2380 2264
rect 2388 2256 2390 2264
rect 2186 1976 2188 1984
rect 2196 1976 2198 1984
rect 2186 1974 2198 1976
rect 2346 1944 2358 1946
rect 2346 1936 2348 1944
rect 2356 1936 2358 1944
rect 2154 1716 2156 1724
rect 2164 1716 2166 1724
rect 2154 1714 2166 1716
rect 2218 1904 2230 1906
rect 2218 1896 2220 1904
rect 2228 1896 2230 1904
rect 2218 1724 2230 1896
rect 2218 1716 2220 1724
rect 2228 1716 2230 1724
rect 2218 1714 2230 1716
rect 2250 1884 2262 1886
rect 2250 1876 2252 1884
rect 2260 1876 2262 1884
rect 2122 1616 2124 1624
rect 2132 1616 2134 1624
rect 2122 1614 2134 1616
rect 2154 1664 2166 1666
rect 2154 1656 2156 1664
rect 2164 1656 2166 1664
rect 2090 1476 2092 1484
rect 2100 1476 2102 1484
rect 2090 1474 2102 1476
rect 2058 1316 2060 1324
rect 2068 1316 2070 1324
rect 2058 1314 2070 1316
rect 2090 1364 2102 1366
rect 2090 1356 2092 1364
rect 2100 1356 2102 1364
rect 2090 1224 2102 1356
rect 2090 1216 2092 1224
rect 2100 1216 2102 1224
rect 2090 1214 2102 1216
rect 2154 1224 2166 1656
rect 2154 1216 2156 1224
rect 2164 1216 2166 1224
rect 2154 1214 2166 1216
rect 2218 1344 2230 1346
rect 2218 1336 2220 1344
rect 2228 1336 2230 1344
rect 2026 1156 2028 1164
rect 2036 1156 2038 1164
rect 2026 1154 2038 1156
rect 1994 1124 2070 1126
rect 1994 1116 2060 1124
rect 2068 1116 2070 1124
rect 1994 1114 2070 1116
rect 1930 1056 1932 1064
rect 1940 1056 1942 1064
rect 1930 1054 1942 1056
rect 1898 1004 1910 1006
rect 1898 996 1900 1004
rect 1908 996 1910 1004
rect 1898 966 1910 996
rect 2090 984 2102 986
rect 2090 976 2092 984
rect 2100 976 2102 984
rect 1898 964 1942 966
rect 1898 956 1932 964
rect 1940 956 1942 964
rect 1898 954 1942 956
rect 1770 896 1772 904
rect 1780 896 1782 904
rect 1770 894 1782 896
rect 1866 924 1878 926
rect 1866 916 1868 924
rect 1876 916 1878 924
rect 1706 836 1708 844
rect 1716 836 1718 844
rect 1706 834 1718 836
rect 1866 804 1878 916
rect 1866 796 1868 804
rect 1876 796 1878 804
rect 1866 794 1878 796
rect 1898 904 1910 906
rect 1898 896 1900 904
rect 1908 896 1910 904
rect 1610 736 1612 744
rect 1620 736 1622 744
rect 1610 734 1622 736
rect 1898 704 1910 896
rect 1898 696 1900 704
rect 1908 696 1910 704
rect 1898 694 1910 696
rect 1546 376 1548 384
rect 1556 376 1558 384
rect 1546 374 1558 376
rect 1994 464 2006 466
rect 1994 456 1996 464
rect 2004 456 2006 464
rect 1514 276 1516 284
rect 1524 276 1526 284
rect 1514 124 1526 276
rect 1514 116 1516 124
rect 1524 116 1526 124
rect 1514 114 1526 116
rect 1962 344 1974 346
rect 1962 336 1964 344
rect 1972 336 1974 344
rect 1962 124 1974 336
rect 1994 284 2006 456
rect 1994 276 1996 284
rect 2004 276 2006 284
rect 1994 274 2006 276
rect 2026 384 2038 386
rect 2026 376 2028 384
rect 2036 376 2038 384
rect 2026 284 2038 376
rect 2090 344 2102 976
rect 2218 884 2230 1336
rect 2250 1224 2262 1876
rect 2346 1704 2358 1936
rect 2346 1696 2348 1704
rect 2356 1696 2358 1704
rect 2346 1694 2358 1696
rect 2378 1704 2390 2256
rect 2474 2264 2486 2266
rect 2474 2256 2476 2264
rect 2484 2256 2486 2264
rect 2378 1696 2380 1704
rect 2388 1696 2390 1704
rect 2282 1484 2294 1486
rect 2282 1476 2284 1484
rect 2292 1476 2294 1484
rect 2282 1304 2294 1476
rect 2282 1296 2284 1304
rect 2292 1296 2294 1304
rect 2282 1294 2294 1296
rect 2378 1304 2390 1696
rect 2410 2124 2422 2126
rect 2410 2116 2412 2124
rect 2420 2116 2422 2124
rect 2410 1344 2422 2116
rect 2442 2104 2454 2106
rect 2442 2096 2444 2104
rect 2452 2096 2454 2104
rect 2442 1724 2454 2096
rect 2474 1864 2486 2256
rect 2570 2124 2582 3016
rect 2602 2944 2614 3736
rect 2634 3584 2646 4116
rect 2634 3576 2636 3584
rect 2644 3576 2646 3584
rect 2634 3574 2646 3576
rect 2698 3984 2710 3986
rect 2698 3976 2700 3984
rect 2708 3976 2710 3984
rect 2698 3484 2710 3976
rect 2698 3476 2700 3484
rect 2708 3476 2710 3484
rect 2698 3474 2710 3476
rect 2762 3924 2774 3926
rect 2762 3916 2764 3924
rect 2772 3916 2774 3924
rect 2762 3384 2774 3916
rect 2762 3376 2764 3384
rect 2772 3376 2774 3384
rect 2762 3374 2774 3376
rect 2826 3864 2838 3866
rect 2826 3856 2828 3864
rect 2836 3856 2838 3864
rect 2730 3344 2742 3346
rect 2730 3336 2732 3344
rect 2740 3336 2742 3344
rect 2602 2936 2604 2944
rect 2612 2936 2614 2944
rect 2602 2934 2614 2936
rect 2666 3124 2678 3126
rect 2666 3116 2668 3124
rect 2676 3116 2678 3124
rect 2666 2544 2678 3116
rect 2730 2684 2742 3336
rect 2826 2744 2838 3856
rect 2912 3814 2976 4206
rect 2912 3806 2916 3814
rect 2924 3806 2928 3814
rect 2936 3806 2940 3814
rect 2948 3806 2952 3814
rect 2960 3806 2964 3814
rect 2972 3806 2976 3814
rect 2912 3414 2976 3806
rect 3306 4224 3318 4226
rect 3306 4216 3308 4224
rect 3316 4216 3318 4224
rect 2912 3406 2916 3414
rect 2924 3406 2928 3414
rect 2936 3406 2940 3414
rect 2948 3406 2952 3414
rect 2960 3406 2964 3414
rect 2972 3406 2976 3414
rect 2912 3014 2976 3406
rect 2912 3006 2916 3014
rect 2924 3006 2928 3014
rect 2936 3006 2940 3014
rect 2948 3006 2952 3014
rect 2960 3006 2964 3014
rect 2972 3006 2976 3014
rect 2826 2736 2828 2744
rect 2836 2736 2838 2744
rect 2826 2734 2838 2736
rect 2858 2744 2870 2746
rect 2858 2736 2860 2744
rect 2868 2736 2870 2744
rect 2730 2676 2732 2684
rect 2740 2676 2742 2684
rect 2730 2674 2742 2676
rect 2666 2536 2668 2544
rect 2676 2536 2678 2544
rect 2666 2534 2678 2536
rect 2826 2584 2838 2586
rect 2826 2576 2828 2584
rect 2836 2576 2838 2584
rect 2826 2304 2838 2576
rect 2858 2544 2870 2736
rect 2858 2536 2860 2544
rect 2868 2536 2870 2544
rect 2858 2534 2870 2536
rect 2912 2614 2976 3006
rect 3018 3584 3030 3586
rect 3018 3576 3020 3584
rect 3028 3576 3030 3584
rect 3018 2844 3030 3576
rect 3018 2836 3020 2844
rect 3028 2836 3030 2844
rect 3018 2834 3030 2836
rect 3146 3184 3158 3186
rect 3146 3176 3148 3184
rect 3156 3176 3158 3184
rect 2912 2606 2916 2614
rect 2924 2606 2928 2614
rect 2936 2606 2940 2614
rect 2948 2606 2952 2614
rect 2960 2606 2964 2614
rect 2972 2606 2976 2614
rect 2826 2296 2828 2304
rect 2836 2296 2838 2304
rect 2826 2294 2838 2296
rect 2570 2116 2572 2124
rect 2580 2116 2582 2124
rect 2570 2114 2582 2116
rect 2794 2284 2806 2286
rect 2794 2276 2796 2284
rect 2804 2276 2806 2284
rect 2794 2084 2806 2276
rect 2858 2284 2870 2286
rect 2858 2276 2860 2284
rect 2868 2276 2870 2284
rect 2858 2144 2870 2276
rect 2858 2136 2860 2144
rect 2868 2136 2870 2144
rect 2858 2134 2870 2136
rect 2912 2214 2976 2606
rect 2912 2206 2916 2214
rect 2924 2206 2928 2214
rect 2936 2206 2940 2214
rect 2948 2206 2952 2214
rect 2960 2206 2964 2214
rect 2972 2206 2976 2214
rect 2794 2076 2796 2084
rect 2804 2076 2806 2084
rect 2794 2074 2806 2076
rect 2474 1856 2476 1864
rect 2484 1856 2486 1864
rect 2474 1854 2486 1856
rect 2698 1884 2710 1886
rect 2698 1876 2700 1884
rect 2708 1876 2710 1884
rect 2442 1716 2444 1724
rect 2452 1716 2454 1724
rect 2442 1714 2454 1716
rect 2474 1744 2486 1746
rect 2474 1736 2476 1744
rect 2484 1736 2486 1744
rect 2474 1484 2486 1736
rect 2474 1476 2476 1484
rect 2484 1476 2486 1484
rect 2474 1474 2486 1476
rect 2602 1524 2614 1526
rect 2602 1516 2604 1524
rect 2612 1516 2614 1524
rect 2410 1336 2412 1344
rect 2420 1336 2422 1344
rect 2410 1334 2422 1336
rect 2570 1384 2582 1386
rect 2570 1376 2572 1384
rect 2580 1376 2582 1384
rect 2442 1324 2470 1326
rect 2442 1316 2460 1324
rect 2468 1316 2470 1324
rect 2442 1314 2470 1316
rect 2378 1296 2380 1304
rect 2388 1296 2390 1304
rect 2378 1294 2390 1296
rect 2410 1304 2422 1306
rect 2410 1296 2412 1304
rect 2420 1296 2422 1304
rect 2250 1216 2252 1224
rect 2260 1216 2262 1224
rect 2250 1214 2262 1216
rect 2410 1204 2422 1296
rect 2410 1196 2412 1204
rect 2420 1196 2422 1204
rect 2410 1194 2422 1196
rect 2442 1204 2454 1314
rect 2442 1196 2444 1204
rect 2452 1196 2454 1204
rect 2442 1194 2454 1196
rect 2570 1204 2582 1376
rect 2602 1384 2614 1516
rect 2602 1376 2604 1384
rect 2612 1376 2614 1384
rect 2602 1374 2614 1376
rect 2634 1484 2646 1486
rect 2634 1476 2636 1484
rect 2644 1476 2646 1484
rect 2634 1324 2646 1476
rect 2698 1484 2710 1876
rect 2912 1814 2976 2206
rect 3050 2824 3062 2826
rect 3050 2816 3052 2824
rect 3060 2816 3062 2824
rect 2912 1806 2916 1814
rect 2924 1806 2928 1814
rect 2936 1806 2940 1814
rect 2948 1806 2952 1814
rect 2960 1806 2964 1814
rect 2972 1806 2976 1814
rect 2858 1524 2870 1526
rect 2858 1516 2860 1524
rect 2868 1516 2870 1524
rect 2698 1476 2700 1484
rect 2708 1476 2710 1484
rect 2698 1474 2710 1476
rect 2730 1484 2742 1486
rect 2730 1476 2732 1484
rect 2740 1476 2742 1484
rect 2634 1316 2636 1324
rect 2644 1316 2646 1324
rect 2634 1314 2646 1316
rect 2730 1324 2742 1476
rect 2730 1316 2732 1324
rect 2740 1316 2742 1324
rect 2730 1314 2742 1316
rect 2794 1444 2806 1446
rect 2794 1436 2796 1444
rect 2804 1436 2806 1444
rect 2570 1196 2572 1204
rect 2580 1196 2582 1204
rect 2570 1194 2582 1196
rect 2794 1204 2806 1436
rect 2858 1384 2870 1516
rect 2858 1376 2860 1384
rect 2868 1376 2870 1384
rect 2858 1374 2870 1376
rect 2912 1414 2976 1806
rect 3018 2104 3030 2106
rect 3018 2096 3020 2104
rect 3028 2096 3030 2104
rect 3018 1524 3030 2096
rect 3050 1864 3062 2816
rect 3146 2504 3158 3176
rect 3146 2496 3148 2504
rect 3156 2496 3158 2504
rect 3146 2494 3158 2496
rect 3178 3124 3190 3126
rect 3178 3116 3180 3124
rect 3188 3116 3190 3124
rect 3178 2224 3190 3116
rect 3306 2744 3318 4216
rect 3370 3984 3382 4836
rect 3530 4504 3542 4506
rect 3530 4496 3532 4504
rect 3540 4496 3542 4504
rect 3530 4084 3542 4496
rect 3722 4424 3734 5096
rect 3754 4964 3766 5156
rect 3946 5144 3958 5146
rect 3946 5136 3948 5144
rect 3956 5136 3958 5144
rect 3818 5124 3830 5126
rect 3818 5116 3820 5124
rect 3828 5116 3830 5124
rect 3818 5004 3830 5116
rect 3818 4996 3820 5004
rect 3828 4996 3830 5004
rect 3818 4994 3830 4996
rect 3754 4956 3756 4964
rect 3764 4956 3766 4964
rect 3754 4954 3766 4956
rect 3946 4964 3958 5136
rect 3946 4956 3948 4964
rect 3956 4956 3958 4964
rect 3946 4954 3958 4956
rect 3978 4964 3990 5296
rect 3978 4956 3980 4964
rect 3988 4956 3990 4964
rect 3978 4954 3990 4956
rect 4042 5104 4054 5106
rect 4042 5096 4044 5104
rect 4052 5096 4054 5104
rect 4042 4784 4054 5096
rect 4106 5004 4118 5336
rect 4416 5214 4480 5416
rect 5920 5414 5984 5416
rect 5920 5406 5924 5414
rect 5932 5406 5936 5414
rect 5944 5406 5948 5414
rect 5956 5406 5960 5414
rect 5968 5406 5972 5414
rect 5980 5406 5984 5414
rect 5130 5324 5142 5326
rect 5130 5316 5132 5324
rect 5140 5316 5142 5324
rect 4416 5206 4420 5214
rect 4428 5206 4432 5214
rect 4440 5206 4444 5214
rect 4452 5206 4456 5214
rect 4464 5206 4468 5214
rect 4476 5206 4480 5214
rect 4106 4996 4108 5004
rect 4116 4996 4118 5004
rect 4106 4994 4118 4996
rect 4234 5204 4246 5206
rect 4234 5196 4236 5204
rect 4244 5196 4246 5204
rect 4042 4776 4044 4784
rect 4052 4776 4054 4784
rect 4042 4774 4054 4776
rect 4106 4784 4118 4786
rect 4106 4776 4108 4784
rect 4116 4776 4118 4784
rect 4074 4684 4086 4686
rect 4074 4676 4076 4684
rect 4084 4676 4086 4684
rect 3722 4416 3724 4424
rect 3732 4416 3734 4424
rect 3690 4384 3702 4386
rect 3690 4376 3692 4384
rect 3700 4376 3702 4384
rect 3530 4076 3532 4084
rect 3540 4076 3542 4084
rect 3530 4074 3542 4076
rect 3594 4304 3606 4306
rect 3594 4296 3596 4304
rect 3604 4296 3606 4304
rect 3370 3976 3372 3984
rect 3380 3976 3382 3984
rect 3370 3974 3382 3976
rect 3402 3264 3414 3266
rect 3402 3256 3404 3264
rect 3412 3256 3414 3264
rect 3402 2944 3414 3256
rect 3402 2936 3404 2944
rect 3412 2936 3414 2944
rect 3402 2934 3414 2936
rect 3434 3164 3446 3166
rect 3434 3156 3436 3164
rect 3444 3156 3446 3164
rect 3306 2736 3308 2744
rect 3316 2736 3318 2744
rect 3306 2734 3318 2736
rect 3370 2644 3382 2646
rect 3370 2636 3372 2644
rect 3380 2636 3382 2644
rect 3338 2444 3350 2446
rect 3338 2436 3340 2444
rect 3348 2436 3350 2444
rect 3178 2216 3180 2224
rect 3188 2216 3190 2224
rect 3178 2214 3190 2216
rect 3242 2364 3254 2366
rect 3242 2356 3244 2364
rect 3252 2356 3254 2364
rect 3210 2044 3222 2046
rect 3210 2036 3212 2044
rect 3220 2036 3222 2044
rect 3050 1856 3052 1864
rect 3060 1856 3062 1864
rect 3050 1854 3062 1856
rect 3082 1924 3094 1926
rect 3082 1916 3084 1924
rect 3092 1916 3094 1924
rect 3018 1516 3020 1524
rect 3028 1516 3030 1524
rect 3018 1514 3030 1516
rect 3082 1424 3094 1916
rect 3082 1416 3084 1424
rect 3092 1416 3094 1424
rect 3082 1414 3094 1416
rect 2912 1406 2916 1414
rect 2924 1406 2928 1414
rect 2936 1406 2940 1414
rect 2948 1406 2952 1414
rect 2960 1406 2964 1414
rect 2972 1406 2976 1414
rect 2794 1196 2796 1204
rect 2804 1196 2806 1204
rect 2794 1194 2806 1196
rect 2410 1154 2486 1166
rect 2250 1124 2262 1126
rect 2250 1116 2252 1124
rect 2260 1116 2262 1124
rect 2250 1064 2262 1116
rect 2410 1086 2422 1154
rect 2250 1056 2252 1064
rect 2260 1056 2262 1064
rect 2250 1054 2262 1056
rect 2282 1074 2422 1086
rect 2442 1124 2454 1126
rect 2442 1116 2444 1124
rect 2452 1116 2454 1124
rect 2282 1064 2294 1074
rect 2282 1056 2284 1064
rect 2292 1056 2294 1064
rect 2282 1054 2294 1056
rect 2442 1064 2454 1116
rect 2474 1124 2486 1154
rect 2474 1116 2476 1124
rect 2484 1116 2486 1124
rect 2474 1114 2486 1116
rect 2506 1124 2518 1126
rect 2506 1116 2508 1124
rect 2516 1116 2518 1124
rect 2442 1056 2444 1064
rect 2452 1056 2454 1064
rect 2442 1054 2454 1056
rect 2506 1046 2518 1116
rect 2474 1034 2518 1046
rect 2474 1006 2486 1034
rect 2912 1014 2976 1406
rect 3146 1384 3158 1386
rect 3146 1376 3148 1384
rect 3156 1376 3158 1384
rect 3082 1344 3094 1346
rect 3082 1336 3084 1344
rect 3092 1336 3094 1344
rect 3082 1086 3094 1336
rect 3114 1204 3126 1206
rect 3114 1196 3116 1204
rect 3124 1196 3126 1204
rect 3114 1126 3126 1196
rect 3146 1204 3158 1376
rect 3146 1196 3148 1204
rect 3156 1196 3158 1204
rect 3146 1194 3158 1196
rect 3114 1114 3158 1126
rect 3146 1104 3158 1114
rect 3146 1096 3148 1104
rect 3156 1096 3158 1104
rect 3146 1094 3158 1096
rect 3082 1074 3126 1086
rect 2912 1006 2916 1014
rect 2924 1006 2928 1014
rect 2936 1006 2940 1014
rect 2948 1006 2952 1014
rect 2960 1006 2964 1014
rect 2972 1006 2976 1014
rect 2298 1004 2486 1006
rect 2298 996 2300 1004
rect 2308 996 2486 1004
rect 2298 994 2486 996
rect 2698 1004 2710 1006
rect 2698 996 2700 1004
rect 2708 996 2710 1004
rect 2570 924 2582 926
rect 2570 916 2572 924
rect 2580 916 2582 924
rect 2218 876 2220 884
rect 2228 876 2230 884
rect 2218 874 2230 876
rect 2314 904 2326 906
rect 2314 896 2316 904
rect 2324 896 2326 904
rect 2314 804 2326 896
rect 2314 796 2316 804
rect 2324 796 2326 804
rect 2314 794 2326 796
rect 2410 744 2422 746
rect 2410 736 2412 744
rect 2420 736 2422 744
rect 2410 704 2422 736
rect 2410 696 2412 704
rect 2420 696 2422 704
rect 2410 694 2422 696
rect 2570 584 2582 916
rect 2570 576 2572 584
rect 2580 576 2582 584
rect 2570 574 2582 576
rect 2602 904 2614 906
rect 2602 896 2604 904
rect 2612 896 2614 904
rect 2602 524 2614 896
rect 2698 904 2710 996
rect 2826 1004 2870 1006
rect 2826 996 2828 1004
rect 2836 996 2870 1004
rect 2826 994 2870 996
rect 2858 984 2870 994
rect 2858 976 2860 984
rect 2868 976 2870 984
rect 2858 974 2870 976
rect 2698 896 2700 904
rect 2708 896 2710 904
rect 2698 894 2710 896
rect 2602 516 2604 524
rect 2612 516 2614 524
rect 2602 514 2614 516
rect 2912 614 2976 1006
rect 3018 1024 3030 1026
rect 3018 1016 3020 1024
rect 3028 1016 3030 1024
rect 3018 804 3030 1016
rect 3018 796 3020 804
rect 3028 796 3030 804
rect 3018 794 3030 796
rect 3050 964 3062 966
rect 3050 956 3052 964
rect 3060 956 3062 964
rect 2912 606 2916 614
rect 2924 606 2928 614
rect 2936 606 2940 614
rect 2948 606 2952 614
rect 2960 606 2964 614
rect 2972 606 2976 614
rect 2090 336 2092 344
rect 2100 336 2102 344
rect 2090 334 2102 336
rect 2026 276 2028 284
rect 2036 276 2038 284
rect 2026 274 2038 276
rect 1962 116 1964 124
rect 1972 116 1974 124
rect 1962 114 1974 116
rect 2912 214 2976 606
rect 3050 304 3062 956
rect 3114 684 3126 1074
rect 3210 1046 3222 2036
rect 3242 2004 3254 2356
rect 3242 1996 3244 2004
rect 3252 1996 3254 2004
rect 3242 1994 3254 1996
rect 3338 1564 3350 2436
rect 3370 1744 3382 2636
rect 3434 2304 3446 3156
rect 3562 3044 3574 3046
rect 3562 3036 3564 3044
rect 3572 3036 3574 3044
rect 3562 2904 3574 3036
rect 3562 2896 3564 2904
rect 3572 2896 3574 2904
rect 3562 2894 3574 2896
rect 3594 2524 3606 4296
rect 3690 3904 3702 4376
rect 3690 3896 3692 3904
rect 3700 3896 3702 3904
rect 3690 3894 3702 3896
rect 3722 3904 3734 4416
rect 3946 4524 3958 4526
rect 3946 4516 3948 4524
rect 3956 4516 3958 4524
rect 3722 3896 3724 3904
rect 3732 3896 3734 3904
rect 3722 3894 3734 3896
rect 3914 4124 3926 4126
rect 3914 4116 3916 4124
rect 3924 4116 3926 4124
rect 3690 3784 3702 3786
rect 3690 3776 3692 3784
rect 3700 3776 3702 3784
rect 3658 3644 3670 3646
rect 3658 3636 3660 3644
rect 3668 3636 3670 3644
rect 3626 3464 3638 3466
rect 3626 3456 3628 3464
rect 3636 3456 3638 3464
rect 3626 3044 3638 3456
rect 3658 3384 3670 3636
rect 3690 3624 3702 3776
rect 3690 3616 3692 3624
rect 3700 3616 3702 3624
rect 3690 3614 3702 3616
rect 3818 3704 3830 3706
rect 3818 3696 3820 3704
rect 3828 3696 3830 3704
rect 3658 3376 3660 3384
rect 3668 3376 3670 3384
rect 3658 3374 3670 3376
rect 3690 3504 3702 3506
rect 3690 3496 3692 3504
rect 3700 3496 3702 3504
rect 3690 3164 3702 3496
rect 3690 3156 3692 3164
rect 3700 3156 3702 3164
rect 3690 3154 3702 3156
rect 3818 3444 3830 3696
rect 3914 3604 3926 4116
rect 3946 3844 3958 4516
rect 4042 4124 4054 4126
rect 4042 4116 4044 4124
rect 4052 4116 4054 4124
rect 4042 3904 4054 4116
rect 4074 4084 4086 4676
rect 4106 4604 4118 4776
rect 4234 4684 4246 5196
rect 4234 4676 4236 4684
rect 4244 4676 4246 4684
rect 4234 4674 4246 4676
rect 4416 4814 4480 5206
rect 4938 5264 4950 5266
rect 4938 5256 4940 5264
rect 4948 5256 4950 5264
rect 4416 4806 4420 4814
rect 4428 4806 4432 4814
rect 4440 4806 4444 4814
rect 4452 4806 4456 4814
rect 4464 4806 4468 4814
rect 4476 4806 4480 4814
rect 4106 4596 4108 4604
rect 4116 4596 4118 4604
rect 4106 4594 4118 4596
rect 4416 4414 4480 4806
rect 4682 5084 4694 5086
rect 4682 5076 4684 5084
rect 4692 5076 4694 5084
rect 4682 4544 4694 5076
rect 4906 5064 4918 5066
rect 4906 5056 4908 5064
rect 4916 5056 4918 5064
rect 4714 5044 4726 5046
rect 4714 5036 4716 5044
rect 4724 5036 4726 5044
rect 4714 4964 4726 5036
rect 4714 4956 4716 4964
rect 4724 4956 4726 4964
rect 4714 4954 4726 4956
rect 4906 4804 4918 5056
rect 4906 4796 4908 4804
rect 4916 4796 4918 4804
rect 4906 4794 4918 4796
rect 4682 4536 4684 4544
rect 4692 4536 4694 4544
rect 4682 4534 4694 4536
rect 4746 4684 4758 4686
rect 4746 4676 4748 4684
rect 4756 4676 4758 4684
rect 4416 4406 4420 4414
rect 4428 4406 4432 4414
rect 4440 4406 4444 4414
rect 4452 4406 4456 4414
rect 4464 4406 4468 4414
rect 4476 4406 4480 4414
rect 4074 4076 4076 4084
rect 4084 4076 4086 4084
rect 4074 4074 4086 4076
rect 4106 4244 4118 4246
rect 4106 4236 4108 4244
rect 4116 4236 4118 4244
rect 4042 3896 4044 3904
rect 4052 3896 4054 3904
rect 4042 3894 4054 3896
rect 4074 3904 4086 3906
rect 4074 3896 4076 3904
rect 4084 3896 4086 3904
rect 3946 3836 3948 3844
rect 3956 3836 3958 3844
rect 3946 3834 3958 3836
rect 3914 3596 3916 3604
rect 3924 3596 3926 3604
rect 3914 3594 3926 3596
rect 3946 3744 3958 3746
rect 3946 3736 3948 3744
rect 3956 3736 3958 3744
rect 3818 3436 3820 3444
rect 3828 3436 3830 3444
rect 3626 3036 3628 3044
rect 3636 3036 3638 3044
rect 3626 3034 3638 3036
rect 3786 2924 3798 2926
rect 3786 2916 3788 2924
rect 3796 2916 3798 2924
rect 3594 2516 3596 2524
rect 3604 2516 3606 2524
rect 3594 2514 3606 2516
rect 3626 2804 3638 2806
rect 3626 2796 3628 2804
rect 3636 2796 3638 2804
rect 3626 2324 3638 2796
rect 3786 2464 3798 2916
rect 3818 2924 3830 3436
rect 3946 3384 3958 3736
rect 4074 3744 4086 3896
rect 4074 3736 4076 3744
rect 4084 3736 4086 3744
rect 4074 3734 4086 3736
rect 4106 3704 4118 4236
rect 4138 4244 4150 4246
rect 4138 4236 4140 4244
rect 4148 4236 4150 4244
rect 4138 4044 4150 4236
rect 4138 4036 4140 4044
rect 4148 4036 4150 4044
rect 4138 4034 4150 4036
rect 4266 4124 4278 4126
rect 4266 4116 4268 4124
rect 4276 4116 4278 4124
rect 4106 3696 4108 3704
rect 4116 3696 4118 3704
rect 3978 3684 3990 3686
rect 3978 3676 3980 3684
rect 3988 3676 3990 3684
rect 3978 3404 3990 3676
rect 3978 3396 3980 3404
rect 3988 3396 3990 3404
rect 3978 3394 3990 3396
rect 4010 3604 4022 3606
rect 4010 3596 4012 3604
rect 4020 3596 4022 3604
rect 3946 3376 3948 3384
rect 3956 3376 3958 3384
rect 3946 3374 3958 3376
rect 3978 3164 3990 3166
rect 3978 3156 3980 3164
rect 3988 3156 3990 3164
rect 3978 3104 3990 3156
rect 3978 3096 3980 3104
rect 3988 3096 3990 3104
rect 3978 3094 3990 3096
rect 4010 3104 4022 3596
rect 4106 3524 4118 3696
rect 4106 3516 4108 3524
rect 4116 3516 4118 3524
rect 4106 3514 4118 3516
rect 4202 4024 4214 4026
rect 4202 4016 4204 4024
rect 4212 4016 4214 4024
rect 4202 3844 4214 4016
rect 4202 3836 4204 3844
rect 4212 3836 4214 3844
rect 4106 3484 4118 3486
rect 4106 3476 4108 3484
rect 4116 3476 4118 3484
rect 4010 3096 4012 3104
rect 4020 3096 4022 3104
rect 4010 3094 4022 3096
rect 4042 3364 4054 3366
rect 4042 3356 4044 3364
rect 4052 3356 4054 3364
rect 3818 2916 3820 2924
rect 3828 2916 3830 2924
rect 3818 2914 3830 2916
rect 3786 2456 3788 2464
rect 3796 2456 3798 2464
rect 3786 2454 3798 2456
rect 3978 2484 3990 2486
rect 3978 2476 3980 2484
rect 3988 2476 3990 2484
rect 3626 2316 3628 2324
rect 3636 2316 3638 2324
rect 3626 2314 3638 2316
rect 3434 2296 3436 2304
rect 3444 2296 3446 2304
rect 3434 2294 3446 2296
rect 3786 2164 3798 2166
rect 3786 2156 3788 2164
rect 3796 2156 3798 2164
rect 3370 1736 3372 1744
rect 3380 1736 3382 1744
rect 3370 1734 3382 1736
rect 3562 2044 3574 2046
rect 3562 2036 3564 2044
rect 3572 2036 3574 2044
rect 3338 1556 3340 1564
rect 3348 1556 3350 1564
rect 3338 1554 3350 1556
rect 3306 1544 3318 1546
rect 3306 1536 3308 1544
rect 3316 1536 3318 1544
rect 3114 676 3116 684
rect 3124 676 3126 684
rect 3114 674 3126 676
rect 3178 1034 3222 1046
rect 3242 1504 3254 1506
rect 3242 1496 3244 1504
rect 3252 1496 3254 1504
rect 3242 1444 3254 1496
rect 3242 1436 3244 1444
rect 3252 1436 3254 1444
rect 3178 444 3190 1034
rect 3242 864 3254 1436
rect 3306 1404 3318 1536
rect 3306 1396 3308 1404
rect 3316 1396 3318 1404
rect 3306 1394 3318 1396
rect 3434 1484 3446 1486
rect 3434 1476 3436 1484
rect 3444 1476 3446 1484
rect 3434 1324 3446 1476
rect 3562 1404 3574 2036
rect 3754 1724 3766 1726
rect 3754 1716 3756 1724
rect 3764 1716 3766 1724
rect 3562 1396 3564 1404
rect 3572 1396 3574 1404
rect 3562 1394 3574 1396
rect 3626 1684 3638 1686
rect 3626 1676 3628 1684
rect 3636 1676 3638 1684
rect 3434 1316 3436 1324
rect 3444 1316 3446 1324
rect 3434 1314 3446 1316
rect 3370 1144 3382 1146
rect 3370 1136 3372 1144
rect 3380 1136 3382 1144
rect 3242 856 3244 864
rect 3252 856 3254 864
rect 3242 854 3254 856
rect 3274 984 3286 986
rect 3274 976 3276 984
rect 3284 976 3286 984
rect 3178 436 3180 444
rect 3188 436 3190 444
rect 3178 434 3190 436
rect 3050 296 3052 304
rect 3060 296 3062 304
rect 3050 294 3062 296
rect 2912 206 2916 214
rect 2924 206 2928 214
rect 2936 206 2940 214
rect 2948 206 2952 214
rect 2960 206 2964 214
rect 2972 206 2976 214
rect 1408 6 1412 14
rect 1420 6 1424 14
rect 1432 6 1436 14
rect 1444 6 1448 14
rect 1456 6 1460 14
rect 1468 6 1472 14
rect 1408 -10 1472 6
rect 2912 -10 2976 206
rect 3274 164 3286 976
rect 3370 564 3382 1136
rect 3626 1124 3638 1676
rect 3658 1664 3670 1666
rect 3658 1656 3660 1664
rect 3668 1656 3670 1664
rect 3658 1524 3670 1656
rect 3658 1516 3660 1524
rect 3668 1516 3670 1524
rect 3658 1514 3670 1516
rect 3626 1116 3628 1124
rect 3636 1116 3638 1124
rect 3626 1114 3638 1116
rect 3658 1124 3670 1126
rect 3658 1116 3660 1124
rect 3668 1116 3670 1124
rect 3434 1084 3446 1086
rect 3434 1076 3436 1084
rect 3444 1076 3446 1084
rect 3434 944 3446 1076
rect 3434 936 3436 944
rect 3444 936 3446 944
rect 3402 804 3414 806
rect 3402 796 3404 804
rect 3412 796 3414 804
rect 3402 644 3414 796
rect 3434 784 3446 936
rect 3434 776 3436 784
rect 3444 776 3446 784
rect 3434 774 3446 776
rect 3658 744 3670 1116
rect 3754 944 3766 1716
rect 3786 1144 3798 2156
rect 3818 2044 3830 2046
rect 3818 2036 3820 2044
rect 3828 2036 3830 2044
rect 3818 1224 3830 2036
rect 3978 1684 3990 2476
rect 4042 2364 4054 3356
rect 4106 3164 4118 3476
rect 4106 3156 4108 3164
rect 4116 3156 4118 3164
rect 4106 3154 4118 3156
rect 4042 2356 4044 2364
rect 4052 2356 4054 2364
rect 4042 2354 4054 2356
rect 4106 3124 4118 3126
rect 4106 3116 4108 3124
rect 4116 3116 4118 3124
rect 4106 2304 4118 3116
rect 4138 3024 4150 3026
rect 4138 3016 4140 3024
rect 4148 3016 4150 3024
rect 4138 2424 4150 3016
rect 4202 2504 4214 3836
rect 4234 3564 4246 3566
rect 4234 3556 4236 3564
rect 4244 3556 4246 3564
rect 4234 2964 4246 3556
rect 4266 3404 4278 4116
rect 4416 4014 4480 4406
rect 4554 4524 4566 4526
rect 4554 4516 4556 4524
rect 4564 4516 4566 4524
rect 4554 4484 4566 4516
rect 4554 4476 4556 4484
rect 4564 4476 4566 4484
rect 4554 4024 4566 4476
rect 4714 4464 4726 4466
rect 4714 4456 4716 4464
rect 4724 4456 4726 4464
rect 4554 4016 4556 4024
rect 4564 4016 4566 4024
rect 4554 4014 4566 4016
rect 4682 4324 4694 4326
rect 4682 4316 4684 4324
rect 4692 4316 4694 4324
rect 4416 4006 4420 4014
rect 4428 4006 4432 4014
rect 4440 4006 4444 4014
rect 4452 4006 4456 4014
rect 4464 4006 4468 4014
rect 4476 4006 4480 4014
rect 4266 3396 4268 3404
rect 4276 3396 4278 3404
rect 4266 3394 4278 3396
rect 4362 3804 4374 3806
rect 4362 3796 4364 3804
rect 4372 3796 4374 3804
rect 4362 3384 4374 3796
rect 4362 3376 4364 3384
rect 4372 3376 4374 3384
rect 4362 3374 4374 3376
rect 4416 3614 4480 4006
rect 4682 3964 4694 4316
rect 4714 4084 4726 4456
rect 4714 4076 4716 4084
rect 4724 4076 4726 4084
rect 4714 4074 4726 4076
rect 4682 3956 4684 3964
rect 4692 3956 4694 3964
rect 4682 3954 4694 3956
rect 4714 3884 4726 3886
rect 4714 3876 4716 3884
rect 4724 3876 4726 3884
rect 4650 3724 4662 3726
rect 4650 3716 4652 3724
rect 4660 3716 4662 3724
rect 4416 3606 4420 3614
rect 4428 3606 4432 3614
rect 4440 3606 4444 3614
rect 4452 3606 4456 3614
rect 4464 3606 4468 3614
rect 4476 3606 4480 3614
rect 4416 3214 4480 3606
rect 4522 3624 4534 3626
rect 4522 3616 4524 3624
rect 4532 3616 4534 3624
rect 4522 3464 4534 3616
rect 4522 3456 4524 3464
rect 4532 3456 4534 3464
rect 4522 3454 4534 3456
rect 4586 3484 4598 3486
rect 4586 3476 4588 3484
rect 4596 3476 4598 3484
rect 4416 3206 4420 3214
rect 4428 3206 4432 3214
rect 4440 3206 4444 3214
rect 4452 3206 4456 3214
rect 4464 3206 4468 3214
rect 4476 3206 4480 3214
rect 4330 3204 4342 3206
rect 4330 3196 4332 3204
rect 4340 3196 4342 3204
rect 4330 3104 4342 3196
rect 4330 3096 4332 3104
rect 4340 3096 4342 3104
rect 4330 3094 4342 3096
rect 4234 2956 4236 2964
rect 4244 2956 4246 2964
rect 4234 2954 4246 2956
rect 4362 2944 4374 2946
rect 4362 2936 4364 2944
rect 4372 2936 4374 2944
rect 4330 2884 4342 2886
rect 4330 2876 4332 2884
rect 4340 2876 4342 2884
rect 4298 2864 4310 2866
rect 4298 2856 4300 2864
rect 4308 2856 4310 2864
rect 4298 2684 4310 2856
rect 4298 2676 4300 2684
rect 4308 2676 4310 2684
rect 4202 2496 4204 2504
rect 4212 2496 4214 2504
rect 4202 2494 4214 2496
rect 4266 2604 4278 2606
rect 4266 2596 4268 2604
rect 4276 2596 4278 2604
rect 4138 2416 4140 2424
rect 4148 2416 4150 2424
rect 4138 2414 4150 2416
rect 4106 2296 4108 2304
rect 4116 2296 4118 2304
rect 4106 2294 4118 2296
rect 4010 2084 4022 2086
rect 4010 2076 4012 2084
rect 4020 2076 4022 2084
rect 4010 1764 4022 2076
rect 4010 1756 4012 1764
rect 4020 1756 4022 1764
rect 4010 1754 4022 1756
rect 4042 1984 4054 1986
rect 4042 1976 4044 1984
rect 4052 1976 4054 1984
rect 3978 1676 3980 1684
rect 3988 1676 3990 1684
rect 3978 1674 3990 1676
rect 3818 1216 3820 1224
rect 3828 1216 3830 1224
rect 3818 1214 3830 1216
rect 3786 1136 3788 1144
rect 3796 1136 3798 1144
rect 3786 1134 3798 1136
rect 4042 1104 4054 1976
rect 4074 1884 4086 1886
rect 4074 1876 4076 1884
rect 4084 1876 4086 1884
rect 4074 1804 4086 1876
rect 4074 1796 4076 1804
rect 4084 1796 4086 1804
rect 4074 1794 4086 1796
rect 4266 1544 4278 2596
rect 4298 2304 4310 2676
rect 4298 2296 4300 2304
rect 4308 2296 4310 2304
rect 4298 2294 4310 2296
rect 4298 2184 4310 2186
rect 4298 2176 4300 2184
rect 4308 2176 4310 2184
rect 4298 2144 4310 2176
rect 4330 2184 4342 2876
rect 4362 2284 4374 2936
rect 4362 2276 4364 2284
rect 4372 2276 4374 2284
rect 4362 2274 4374 2276
rect 4416 2814 4480 3206
rect 4522 3384 4534 3386
rect 4522 3376 4524 3384
rect 4532 3376 4534 3384
rect 4522 3024 4534 3376
rect 4586 3304 4598 3476
rect 4586 3296 4588 3304
rect 4596 3296 4598 3304
rect 4586 3294 4598 3296
rect 4522 3016 4524 3024
rect 4532 3016 4534 3024
rect 4522 3014 4534 3016
rect 4650 2924 4662 3716
rect 4714 3704 4726 3876
rect 4746 3724 4758 4676
rect 4874 4684 4886 4686
rect 4874 4676 4876 4684
rect 4884 4676 4886 4684
rect 4874 4404 4886 4676
rect 4906 4684 4918 4686
rect 4906 4676 4908 4684
rect 4916 4676 4918 4684
rect 4906 4544 4918 4676
rect 4906 4536 4908 4544
rect 4916 4536 4918 4544
rect 4906 4534 4918 4536
rect 4938 4524 4950 5256
rect 5130 5004 5142 5316
rect 5130 4996 5132 5004
rect 5140 4996 5142 5004
rect 5002 4954 5078 4966
rect 5002 4924 5014 4954
rect 5002 4916 5004 4924
rect 5012 4916 5014 4924
rect 5002 4914 5014 4916
rect 5066 4904 5078 4954
rect 5066 4896 5068 4904
rect 5076 4896 5078 4904
rect 5066 4894 5078 4896
rect 5098 4944 5110 4946
rect 5098 4936 5100 4944
rect 5108 4936 5110 4944
rect 5002 4844 5014 4846
rect 5002 4836 5004 4844
rect 5012 4836 5014 4844
rect 5002 4764 5014 4836
rect 5002 4756 5004 4764
rect 5012 4756 5014 4764
rect 5002 4754 5014 4756
rect 5098 4704 5110 4936
rect 5130 4784 5142 4996
rect 5130 4776 5132 4784
rect 5140 4776 5142 4784
rect 5130 4774 5142 4776
rect 5290 5304 5302 5306
rect 5290 5296 5292 5304
rect 5300 5296 5302 5304
rect 5098 4696 5100 4704
rect 5108 4696 5110 4704
rect 5098 4694 5110 4696
rect 5194 4684 5206 4686
rect 5194 4676 5196 4684
rect 5204 4676 5206 4684
rect 4938 4516 4940 4524
rect 4948 4516 4950 4524
rect 4938 4514 4950 4516
rect 5002 4664 5014 4666
rect 5002 4656 5004 4664
rect 5012 4656 5014 4664
rect 4874 4396 4876 4404
rect 4884 4396 4886 4404
rect 4842 4004 4854 4006
rect 4842 3996 4844 4004
rect 4852 3996 4854 4004
rect 4746 3716 4748 3724
rect 4756 3716 4758 3724
rect 4746 3714 4758 3716
rect 4778 3964 4790 3966
rect 4778 3956 4780 3964
rect 4788 3956 4790 3964
rect 4714 3696 4716 3704
rect 4724 3696 4726 3704
rect 4714 3644 4726 3696
rect 4714 3636 4716 3644
rect 4724 3636 4726 3644
rect 4714 3634 4726 3636
rect 4778 3544 4790 3956
rect 4810 3944 4822 3946
rect 4810 3936 4812 3944
rect 4820 3936 4822 3944
rect 4810 3884 4822 3936
rect 4810 3876 4812 3884
rect 4820 3876 4822 3884
rect 4810 3874 4822 3876
rect 4778 3536 4780 3544
rect 4788 3536 4790 3544
rect 4746 3364 4758 3366
rect 4746 3356 4748 3364
rect 4756 3356 4758 3364
rect 4650 2916 4652 2924
rect 4660 2916 4662 2924
rect 4650 2914 4662 2916
rect 4714 3324 4726 3326
rect 4714 3316 4716 3324
rect 4724 3316 4726 3324
rect 4714 2924 4726 3316
rect 4714 2916 4716 2924
rect 4724 2916 4726 2924
rect 4714 2914 4726 2916
rect 4416 2806 4420 2814
rect 4428 2806 4432 2814
rect 4440 2806 4444 2814
rect 4452 2806 4456 2814
rect 4464 2806 4468 2814
rect 4476 2806 4480 2814
rect 4416 2414 4480 2806
rect 4650 2884 4662 2886
rect 4650 2876 4652 2884
rect 4660 2876 4662 2884
rect 4650 2484 4662 2876
rect 4650 2476 4652 2484
rect 4660 2476 4662 2484
rect 4416 2406 4420 2414
rect 4428 2406 4432 2414
rect 4440 2406 4444 2414
rect 4452 2406 4456 2414
rect 4464 2406 4468 2414
rect 4476 2406 4480 2414
rect 4330 2176 4332 2184
rect 4340 2176 4342 2184
rect 4330 2174 4342 2176
rect 4298 2136 4300 2144
rect 4308 2136 4310 2144
rect 4298 2134 4310 2136
rect 4330 2144 4342 2146
rect 4330 2136 4332 2144
rect 4340 2136 4342 2144
rect 4330 2104 4342 2136
rect 4330 2096 4332 2104
rect 4340 2096 4342 2104
rect 4330 2094 4342 2096
rect 4416 2014 4480 2406
rect 4554 2424 4566 2426
rect 4554 2416 4556 2424
rect 4564 2416 4566 2424
rect 4522 2084 4534 2086
rect 4522 2076 4524 2084
rect 4532 2076 4534 2084
rect 4522 2024 4534 2076
rect 4522 2016 4524 2024
rect 4532 2016 4534 2024
rect 4522 2014 4534 2016
rect 4416 2006 4420 2014
rect 4428 2006 4432 2014
rect 4440 2006 4444 2014
rect 4452 2006 4456 2014
rect 4464 2006 4468 2014
rect 4476 2006 4480 2014
rect 4266 1536 4268 1544
rect 4276 1536 4278 1544
rect 4266 1534 4278 1536
rect 4298 1704 4310 1706
rect 4298 1696 4300 1704
rect 4308 1696 4310 1704
rect 4170 1444 4182 1446
rect 4170 1436 4172 1444
rect 4180 1436 4182 1444
rect 4138 1424 4150 1426
rect 4138 1416 4140 1424
rect 4148 1416 4150 1424
rect 4138 1324 4150 1416
rect 4138 1316 4140 1324
rect 4148 1316 4150 1324
rect 4138 1314 4150 1316
rect 4170 1224 4182 1436
rect 4298 1304 4310 1696
rect 4416 1614 4480 2006
rect 4416 1606 4420 1614
rect 4428 1606 4432 1614
rect 4440 1606 4444 1614
rect 4452 1606 4456 1614
rect 4464 1606 4468 1614
rect 4476 1606 4480 1614
rect 4298 1296 4300 1304
rect 4308 1296 4310 1304
rect 4298 1294 4310 1296
rect 4362 1484 4374 1486
rect 4362 1476 4364 1484
rect 4372 1476 4374 1484
rect 4170 1216 4172 1224
rect 4180 1216 4182 1224
rect 4170 1214 4182 1216
rect 4042 1096 4044 1104
rect 4052 1096 4054 1104
rect 4042 1094 4054 1096
rect 4330 1044 4342 1046
rect 4330 1036 4332 1044
rect 4340 1036 4342 1044
rect 3754 936 3756 944
rect 3764 936 3766 944
rect 3754 934 3766 936
rect 3882 1024 3894 1026
rect 3882 1016 3884 1024
rect 3892 1016 3894 1024
rect 3658 736 3660 744
rect 3668 736 3670 744
rect 3658 734 3670 736
rect 3754 904 3766 906
rect 3754 896 3756 904
rect 3764 896 3766 904
rect 3402 636 3404 644
rect 3412 636 3414 644
rect 3402 634 3414 636
rect 3658 664 3670 666
rect 3658 656 3660 664
rect 3668 656 3670 664
rect 3370 556 3372 564
rect 3380 556 3382 564
rect 3370 554 3382 556
rect 3530 624 3542 626
rect 3530 616 3532 624
rect 3540 616 3542 624
rect 3530 424 3542 616
rect 3530 416 3532 424
rect 3540 416 3542 424
rect 3530 414 3542 416
rect 3658 304 3670 656
rect 3754 604 3766 896
rect 3882 664 3894 1016
rect 4330 944 4342 1036
rect 4330 936 4332 944
rect 4340 936 4342 944
rect 4330 934 4342 936
rect 4362 1044 4374 1476
rect 4362 1036 4364 1044
rect 4372 1036 4374 1044
rect 3882 656 3884 664
rect 3892 656 3894 664
rect 3882 654 3894 656
rect 3914 904 3926 906
rect 3914 896 3916 904
rect 3924 896 3926 904
rect 3914 644 3926 896
rect 3914 636 3916 644
rect 3924 636 3926 644
rect 3914 634 3926 636
rect 4042 724 4054 726
rect 4042 716 4044 724
rect 4052 716 4054 724
rect 3754 596 3756 604
rect 3764 596 3766 604
rect 3754 594 3766 596
rect 3882 604 3894 606
rect 3882 596 3884 604
rect 3892 596 3894 604
rect 3882 524 3894 596
rect 3882 516 3884 524
rect 3892 516 3894 524
rect 3882 514 3894 516
rect 3658 296 3660 304
rect 3668 296 3670 304
rect 3658 184 3670 296
rect 3658 176 3660 184
rect 3668 176 3670 184
rect 3658 174 3670 176
rect 3274 156 3276 164
rect 3284 156 3286 164
rect 3274 154 3286 156
rect 4042 24 4054 716
rect 4362 544 4374 1036
rect 4362 536 4364 544
rect 4372 536 4374 544
rect 4042 16 4044 24
rect 4052 16 4054 24
rect 4042 14 4054 16
rect 4234 364 4246 366
rect 4234 356 4236 364
rect 4244 356 4246 364
rect 4234 24 4246 356
rect 4362 324 4374 536
rect 4362 316 4364 324
rect 4372 316 4374 324
rect 4362 204 4374 316
rect 4362 196 4364 204
rect 4372 196 4374 204
rect 4362 194 4374 196
rect 4416 1214 4480 1606
rect 4522 1764 4534 1766
rect 4522 1756 4524 1764
rect 4532 1756 4534 1764
rect 4522 1604 4534 1756
rect 4522 1596 4524 1604
rect 4532 1596 4534 1604
rect 4522 1594 4534 1596
rect 4554 1504 4566 2416
rect 4650 2284 4662 2476
rect 4714 2584 4726 2586
rect 4714 2576 4716 2584
rect 4724 2576 4726 2584
rect 4714 2444 4726 2576
rect 4714 2436 4716 2444
rect 4724 2436 4726 2444
rect 4714 2434 4726 2436
rect 4746 2304 4758 3356
rect 4778 3344 4790 3536
rect 4842 3744 4854 3996
rect 4842 3736 4844 3744
rect 4852 3736 4854 3744
rect 4842 3524 4854 3736
rect 4842 3516 4844 3524
rect 4852 3516 4854 3524
rect 4778 3336 4780 3344
rect 4788 3336 4790 3344
rect 4778 3334 4790 3336
rect 4810 3444 4822 3446
rect 4810 3436 4812 3444
rect 4820 3436 4822 3444
rect 4810 3324 4822 3436
rect 4810 3316 4812 3324
rect 4820 3316 4822 3324
rect 4810 3314 4822 3316
rect 4778 3264 4790 3266
rect 4778 3256 4780 3264
rect 4788 3256 4790 3264
rect 4778 2444 4790 3256
rect 4842 3104 4854 3516
rect 4842 3096 4844 3104
rect 4852 3096 4854 3104
rect 4842 3094 4854 3096
rect 4874 3904 4886 4396
rect 5002 4284 5014 4656
rect 5034 4344 5046 4346
rect 5034 4336 5036 4344
rect 5044 4336 5046 4344
rect 5034 4304 5046 4336
rect 5034 4296 5036 4304
rect 5044 4296 5046 4304
rect 5034 4294 5046 4296
rect 5002 4276 5004 4284
rect 5012 4276 5014 4284
rect 5002 4274 5014 4276
rect 4970 4264 4982 4266
rect 4970 4256 4972 4264
rect 4980 4256 4982 4264
rect 4874 3896 4876 3904
rect 4884 3896 4886 3904
rect 4874 3104 4886 3896
rect 4938 4104 4950 4106
rect 4938 4096 4940 4104
rect 4948 4096 4950 4104
rect 4906 3824 4918 3826
rect 4906 3816 4908 3824
rect 4916 3816 4918 3824
rect 4906 3684 4918 3816
rect 4938 3824 4950 4096
rect 4938 3816 4940 3824
rect 4948 3816 4950 3824
rect 4938 3814 4950 3816
rect 4970 3904 4982 4256
rect 4970 3896 4972 3904
rect 4980 3896 4982 3904
rect 4970 3764 4982 3896
rect 5098 4244 5110 4246
rect 5098 4236 5100 4244
rect 5108 4236 5110 4244
rect 5098 3844 5110 4236
rect 5162 4244 5174 4246
rect 5162 4236 5164 4244
rect 5172 4236 5174 4244
rect 5098 3836 5100 3844
rect 5108 3836 5110 3844
rect 5098 3834 5110 3836
rect 5130 4184 5142 4186
rect 5130 4176 5132 4184
rect 5140 4176 5142 4184
rect 4970 3756 4972 3764
rect 4980 3756 4982 3764
rect 4970 3754 4982 3756
rect 4906 3676 4908 3684
rect 4916 3676 4918 3684
rect 4906 3674 4918 3676
rect 4938 3724 4950 3726
rect 4938 3716 4940 3724
rect 4948 3716 4950 3724
rect 4874 3096 4876 3104
rect 4884 3096 4886 3104
rect 4874 3094 4886 3096
rect 4938 3084 4950 3716
rect 5098 3684 5110 3686
rect 5098 3676 5100 3684
rect 5108 3676 5110 3684
rect 5034 3504 5046 3506
rect 5034 3496 5036 3504
rect 5044 3496 5046 3504
rect 5034 3284 5046 3496
rect 5066 3504 5078 3506
rect 5066 3496 5068 3504
rect 5076 3496 5078 3504
rect 5066 3344 5078 3496
rect 5066 3336 5068 3344
rect 5076 3336 5078 3344
rect 5066 3334 5078 3336
rect 5098 3364 5110 3676
rect 5130 3684 5142 4176
rect 5162 4144 5174 4236
rect 5162 4136 5164 4144
rect 5172 4136 5174 4144
rect 5162 4134 5174 4136
rect 5194 4064 5206 4676
rect 5290 4684 5302 5296
rect 5770 5204 5782 5206
rect 5770 5196 5772 5204
rect 5780 5196 5782 5204
rect 5418 5104 5430 5106
rect 5418 5096 5420 5104
rect 5428 5096 5430 5104
rect 5418 4864 5430 5096
rect 5418 4856 5420 4864
rect 5428 4856 5430 4864
rect 5418 4854 5430 4856
rect 5482 4924 5494 4926
rect 5482 4916 5484 4924
rect 5492 4916 5494 4924
rect 5290 4676 5292 4684
rect 5300 4676 5302 4684
rect 5290 4674 5302 4676
rect 5322 4744 5334 4746
rect 5322 4736 5324 4744
rect 5332 4736 5334 4744
rect 5322 4664 5334 4736
rect 5322 4656 5324 4664
rect 5332 4656 5334 4664
rect 5322 4654 5334 4656
rect 5482 4424 5494 4916
rect 5482 4416 5484 4424
rect 5492 4416 5494 4424
rect 5482 4414 5494 4416
rect 5482 4384 5494 4386
rect 5482 4376 5484 4384
rect 5492 4376 5494 4384
rect 5194 4056 5196 4064
rect 5204 4056 5206 4064
rect 5194 4054 5206 4056
rect 5290 4264 5302 4266
rect 5290 4256 5292 4264
rect 5300 4256 5302 4264
rect 5258 4004 5270 4006
rect 5258 3996 5260 4004
rect 5268 3996 5270 4004
rect 5194 3964 5206 3966
rect 5194 3956 5196 3964
rect 5204 3956 5206 3964
rect 5162 3944 5174 3946
rect 5162 3936 5164 3944
rect 5172 3936 5174 3944
rect 5162 3804 5174 3936
rect 5162 3796 5164 3804
rect 5172 3796 5174 3804
rect 5162 3794 5174 3796
rect 5130 3676 5132 3684
rect 5140 3676 5142 3684
rect 5130 3674 5142 3676
rect 5162 3624 5174 3626
rect 5162 3616 5164 3624
rect 5172 3616 5174 3624
rect 5162 3404 5174 3616
rect 5162 3396 5164 3404
rect 5172 3396 5174 3404
rect 5162 3394 5174 3396
rect 5098 3356 5100 3364
rect 5108 3356 5110 3364
rect 5034 3276 5036 3284
rect 5044 3276 5046 3284
rect 5034 3274 5046 3276
rect 4938 3076 4940 3084
rect 4948 3076 4950 3084
rect 4938 3074 4950 3076
rect 4874 3024 4886 3026
rect 4874 3016 4876 3024
rect 4884 3016 4886 3024
rect 4810 2984 4822 2986
rect 4810 2976 4812 2984
rect 4820 2976 4822 2984
rect 4810 2544 4822 2976
rect 4874 2664 4886 3016
rect 4970 3004 4982 3006
rect 4970 2996 4972 3004
rect 4980 2996 4982 3004
rect 4938 2744 4950 2746
rect 4938 2736 4940 2744
rect 4948 2736 4950 2744
rect 4874 2656 4876 2664
rect 4884 2656 4886 2664
rect 4874 2654 4886 2656
rect 4906 2664 4918 2666
rect 4906 2656 4908 2664
rect 4916 2656 4918 2664
rect 4810 2536 4812 2544
rect 4820 2536 4822 2544
rect 4810 2534 4822 2536
rect 4874 2524 4886 2526
rect 4874 2516 4876 2524
rect 4884 2516 4886 2524
rect 4778 2436 4780 2444
rect 4788 2436 4790 2444
rect 4778 2434 4790 2436
rect 4842 2504 4854 2506
rect 4842 2496 4844 2504
rect 4852 2496 4854 2504
rect 4746 2296 4748 2304
rect 4756 2296 4758 2304
rect 4746 2294 4758 2296
rect 4650 2276 4652 2284
rect 4660 2276 4662 2284
rect 4650 2274 4662 2276
rect 4682 2284 4694 2286
rect 4682 2276 4684 2284
rect 4692 2276 4694 2284
rect 4586 1944 4598 1946
rect 4586 1936 4588 1944
rect 4596 1936 4598 1944
rect 4586 1844 4598 1936
rect 4586 1836 4588 1844
rect 4596 1836 4598 1844
rect 4586 1834 4598 1836
rect 4650 1864 4662 1866
rect 4650 1856 4652 1864
rect 4660 1856 4662 1864
rect 4618 1724 4630 1726
rect 4618 1716 4620 1724
rect 4628 1716 4630 1724
rect 4554 1496 4556 1504
rect 4564 1496 4566 1504
rect 4554 1494 4566 1496
rect 4586 1504 4598 1506
rect 4586 1496 4588 1504
rect 4596 1496 4598 1504
rect 4416 1206 4420 1214
rect 4428 1206 4432 1214
rect 4440 1206 4444 1214
rect 4452 1206 4456 1214
rect 4464 1206 4468 1214
rect 4476 1206 4480 1214
rect 4416 814 4480 1206
rect 4554 1464 4566 1466
rect 4554 1456 4556 1464
rect 4564 1456 4566 1464
rect 4554 1324 4566 1456
rect 4554 1316 4556 1324
rect 4564 1316 4566 1324
rect 4522 1064 4534 1066
rect 4522 1056 4524 1064
rect 4532 1056 4534 1064
rect 4522 1024 4534 1056
rect 4522 1016 4524 1024
rect 4532 1016 4534 1024
rect 4522 1014 4534 1016
rect 4416 806 4420 814
rect 4428 806 4432 814
rect 4440 806 4444 814
rect 4452 806 4456 814
rect 4464 806 4468 814
rect 4476 806 4480 814
rect 4416 414 4480 806
rect 4554 444 4566 1316
rect 4586 1244 4598 1496
rect 4618 1324 4630 1716
rect 4618 1316 4620 1324
rect 4628 1316 4630 1324
rect 4618 1314 4630 1316
rect 4586 1236 4588 1244
rect 4596 1236 4598 1244
rect 4586 1234 4598 1236
rect 4650 984 4662 1856
rect 4682 1684 4694 2276
rect 4842 2284 4854 2496
rect 4842 2276 4844 2284
rect 4852 2276 4854 2284
rect 4842 2274 4854 2276
rect 4746 2264 4758 2266
rect 4746 2256 4748 2264
rect 4756 2256 4758 2264
rect 4714 1904 4726 1906
rect 4714 1896 4716 1904
rect 4724 1896 4726 1904
rect 4714 1704 4726 1896
rect 4746 1884 4758 2256
rect 4874 2124 4886 2516
rect 4906 2244 4918 2656
rect 4938 2604 4950 2736
rect 4938 2596 4940 2604
rect 4948 2596 4950 2604
rect 4938 2594 4950 2596
rect 4906 2236 4908 2244
rect 4916 2236 4918 2244
rect 4906 2234 4918 2236
rect 4970 2244 4982 2996
rect 5066 2964 5078 2966
rect 5066 2956 5068 2964
rect 5076 2956 5078 2964
rect 5066 2904 5078 2956
rect 5098 2924 5110 3356
rect 5098 2916 5100 2924
rect 5108 2916 5110 2924
rect 5098 2914 5110 2916
rect 5130 3084 5142 3086
rect 5130 3076 5132 3084
rect 5140 3076 5142 3084
rect 5066 2896 5068 2904
rect 5076 2896 5078 2904
rect 5066 2894 5078 2896
rect 5034 2864 5046 2866
rect 5034 2856 5036 2864
rect 5044 2856 5046 2864
rect 5002 2824 5014 2826
rect 5002 2816 5004 2824
rect 5012 2816 5014 2824
rect 5002 2784 5014 2816
rect 5002 2776 5004 2784
rect 5012 2776 5014 2784
rect 5002 2774 5014 2776
rect 4970 2236 4972 2244
rect 4980 2236 4982 2244
rect 4970 2234 4982 2236
rect 5034 2524 5046 2856
rect 5130 2864 5142 3076
rect 5130 2856 5132 2864
rect 5140 2856 5142 2864
rect 5066 2744 5078 2746
rect 5066 2736 5068 2744
rect 5076 2736 5078 2744
rect 5066 2704 5078 2736
rect 5066 2696 5068 2704
rect 5076 2696 5078 2704
rect 5066 2694 5078 2696
rect 5098 2744 5110 2746
rect 5098 2736 5100 2744
rect 5108 2736 5110 2744
rect 5034 2516 5036 2524
rect 5044 2516 5046 2524
rect 4938 2184 4950 2186
rect 4938 2176 4940 2184
rect 4948 2176 4950 2184
rect 4938 2144 4950 2176
rect 4938 2136 4940 2144
rect 4948 2136 4950 2144
rect 4938 2134 4950 2136
rect 5002 2164 5014 2166
rect 5002 2156 5004 2164
rect 5012 2156 5014 2164
rect 4874 2116 4876 2124
rect 4884 2116 4886 2124
rect 4874 2114 4886 2116
rect 4842 2104 4854 2106
rect 4842 2096 4844 2104
rect 4852 2096 4854 2104
rect 4746 1876 4748 1884
rect 4756 1876 4758 1884
rect 4746 1874 4758 1876
rect 4810 2024 4822 2026
rect 4810 2016 4812 2024
rect 4820 2016 4822 2024
rect 4714 1696 4716 1704
rect 4724 1696 4726 1704
rect 4714 1694 4726 1696
rect 4746 1784 4758 1786
rect 4746 1776 4748 1784
rect 4756 1776 4758 1784
rect 4682 1676 4684 1684
rect 4692 1676 4694 1684
rect 4682 1674 4694 1676
rect 4746 1604 4758 1776
rect 4746 1596 4748 1604
rect 4756 1596 4758 1604
rect 4746 1594 4758 1596
rect 4810 1504 4822 2016
rect 4810 1496 4812 1504
rect 4820 1496 4822 1504
rect 4810 1494 4822 1496
rect 4810 1464 4822 1466
rect 4810 1456 4812 1464
rect 4820 1456 4822 1464
rect 4778 1404 4790 1406
rect 4778 1396 4780 1404
rect 4788 1396 4790 1404
rect 4714 1144 4726 1146
rect 4714 1136 4716 1144
rect 4724 1136 4726 1144
rect 4650 976 4652 984
rect 4660 976 4662 984
rect 4650 974 4662 976
rect 4682 1104 4694 1106
rect 4682 1096 4684 1104
rect 4692 1096 4694 1104
rect 4682 704 4694 1096
rect 4714 744 4726 1136
rect 4778 1104 4790 1396
rect 4778 1096 4780 1104
rect 4788 1096 4790 1104
rect 4778 1094 4790 1096
rect 4810 1004 4822 1456
rect 4842 1304 4854 2096
rect 5002 2084 5014 2156
rect 5002 2076 5004 2084
rect 5012 2076 5014 2084
rect 5002 2074 5014 2076
rect 5034 2084 5046 2516
rect 5098 2124 5110 2736
rect 5098 2116 5100 2124
rect 5108 2116 5110 2124
rect 5098 2114 5110 2116
rect 5034 2076 5036 2084
rect 5044 2076 5046 2084
rect 5034 2074 5046 2076
rect 4906 2004 4918 2006
rect 4906 1996 4908 2004
rect 4916 1996 4918 2004
rect 4906 1864 4918 1996
rect 4906 1856 4908 1864
rect 4916 1856 4918 1864
rect 4906 1854 4918 1856
rect 5130 1884 5142 2856
rect 5162 2824 5174 2826
rect 5162 2816 5164 2824
rect 5172 2816 5174 2824
rect 5162 2604 5174 2816
rect 5194 2824 5206 3956
rect 5258 3764 5270 3996
rect 5258 3756 5260 3764
rect 5268 3756 5270 3764
rect 5258 3754 5270 3756
rect 5194 2816 5196 2824
rect 5204 2816 5206 2824
rect 5194 2814 5206 2816
rect 5226 3744 5238 3746
rect 5226 3736 5228 3744
rect 5236 3736 5238 3744
rect 5226 3124 5238 3736
rect 5290 3624 5302 4256
rect 5322 4184 5334 4186
rect 5322 4176 5324 4184
rect 5332 4176 5334 4184
rect 5322 3804 5334 4176
rect 5482 4144 5494 4376
rect 5610 4264 5622 4266
rect 5610 4256 5612 4264
rect 5620 4256 5622 4264
rect 5482 4136 5484 4144
rect 5492 4136 5494 4144
rect 5482 4134 5494 4136
rect 5514 4184 5526 4186
rect 5514 4176 5516 4184
rect 5524 4176 5526 4184
rect 5322 3796 5324 3804
rect 5332 3796 5334 3804
rect 5322 3794 5334 3796
rect 5514 3724 5526 4176
rect 5514 3716 5516 3724
rect 5524 3716 5526 3724
rect 5514 3714 5526 3716
rect 5578 3884 5590 3886
rect 5578 3876 5580 3884
rect 5588 3876 5590 3884
rect 5290 3616 5292 3624
rect 5300 3616 5302 3624
rect 5290 3614 5302 3616
rect 5546 3644 5558 3646
rect 5546 3636 5548 3644
rect 5556 3636 5558 3644
rect 5450 3484 5478 3486
rect 5450 3476 5468 3484
rect 5476 3476 5478 3484
rect 5450 3474 5478 3476
rect 5322 3444 5334 3446
rect 5322 3436 5324 3444
rect 5332 3436 5334 3444
rect 5258 3404 5270 3406
rect 5258 3396 5260 3404
rect 5268 3396 5270 3404
rect 5258 3224 5270 3396
rect 5258 3216 5260 3224
rect 5268 3216 5270 3224
rect 5258 3214 5270 3216
rect 5322 3204 5334 3436
rect 5450 3444 5462 3474
rect 5450 3436 5452 3444
rect 5460 3436 5462 3444
rect 5450 3434 5462 3436
rect 5322 3196 5324 3204
rect 5332 3196 5334 3204
rect 5322 3194 5334 3196
rect 5418 3264 5430 3266
rect 5418 3256 5420 3264
rect 5428 3256 5430 3264
rect 5226 3116 5228 3124
rect 5236 3116 5238 3124
rect 5162 2596 5164 2604
rect 5172 2596 5174 2604
rect 5162 2594 5174 2596
rect 5194 2684 5206 2686
rect 5194 2676 5196 2684
rect 5204 2676 5206 2684
rect 5194 2464 5206 2676
rect 5194 2456 5196 2464
rect 5204 2456 5206 2464
rect 5194 2454 5206 2456
rect 5162 2304 5174 2306
rect 5162 2296 5164 2304
rect 5172 2296 5174 2304
rect 5162 2004 5174 2296
rect 5226 2304 5238 3116
rect 5418 2904 5430 3256
rect 5418 2896 5420 2904
rect 5428 2896 5430 2904
rect 5418 2894 5430 2896
rect 5482 3184 5494 3186
rect 5482 3176 5484 3184
rect 5492 3176 5494 3184
rect 5290 2824 5302 2826
rect 5290 2816 5292 2824
rect 5300 2816 5302 2824
rect 5290 2584 5302 2816
rect 5290 2576 5292 2584
rect 5300 2576 5302 2584
rect 5290 2574 5302 2576
rect 5354 2824 5366 2826
rect 5354 2816 5356 2824
rect 5364 2816 5366 2824
rect 5258 2544 5270 2546
rect 5258 2536 5260 2544
rect 5268 2536 5270 2544
rect 5258 2504 5270 2536
rect 5258 2496 5260 2504
rect 5268 2496 5270 2504
rect 5258 2494 5270 2496
rect 5322 2544 5334 2546
rect 5322 2536 5324 2544
rect 5332 2536 5334 2544
rect 5322 2404 5334 2536
rect 5354 2544 5366 2816
rect 5354 2536 5356 2544
rect 5364 2536 5366 2544
rect 5354 2534 5366 2536
rect 5450 2604 5462 2606
rect 5450 2596 5452 2604
rect 5460 2596 5462 2604
rect 5322 2396 5324 2404
rect 5332 2396 5334 2404
rect 5322 2394 5334 2396
rect 5226 2296 5228 2304
rect 5236 2296 5238 2304
rect 5226 2294 5238 2296
rect 5194 2184 5206 2186
rect 5194 2176 5196 2184
rect 5204 2176 5206 2184
rect 5194 2084 5206 2176
rect 5290 2184 5302 2186
rect 5290 2176 5292 2184
rect 5300 2176 5302 2184
rect 5194 2076 5196 2084
rect 5204 2076 5206 2084
rect 5194 2074 5206 2076
rect 5258 2084 5270 2086
rect 5258 2076 5260 2084
rect 5268 2076 5270 2084
rect 5162 1996 5164 2004
rect 5172 1996 5174 2004
rect 5162 1994 5174 1996
rect 5258 1924 5270 2076
rect 5290 2084 5302 2176
rect 5450 2184 5462 2596
rect 5482 2264 5494 3176
rect 5482 2256 5484 2264
rect 5492 2256 5494 2264
rect 5482 2254 5494 2256
rect 5514 2884 5526 2886
rect 5514 2876 5516 2884
rect 5524 2876 5526 2884
rect 5514 2424 5526 2876
rect 5546 2524 5558 3636
rect 5546 2516 5548 2524
rect 5556 2516 5558 2524
rect 5546 2514 5558 2516
rect 5578 3104 5590 3876
rect 5610 3724 5622 4256
rect 5770 4164 5782 5196
rect 5920 5014 5984 5406
rect 7338 5404 7350 5406
rect 7338 5396 7340 5404
rect 7348 5396 7350 5404
rect 6986 5384 6998 5386
rect 6986 5376 6988 5384
rect 6996 5376 6998 5384
rect 6410 5324 6422 5326
rect 6410 5316 6412 5324
rect 6420 5316 6422 5324
rect 6122 5264 6134 5266
rect 6122 5256 6124 5264
rect 6132 5256 6134 5264
rect 6090 5204 6102 5206
rect 6090 5196 6092 5204
rect 6100 5196 6102 5204
rect 5920 5006 5924 5014
rect 5932 5006 5936 5014
rect 5944 5006 5948 5014
rect 5956 5006 5960 5014
rect 5968 5006 5972 5014
rect 5980 5006 5984 5014
rect 5866 4844 5878 4846
rect 5866 4836 5868 4844
rect 5876 4836 5878 4844
rect 5834 4704 5846 4706
rect 5834 4696 5836 4704
rect 5844 4696 5846 4704
rect 5770 4156 5772 4164
rect 5780 4156 5782 4164
rect 5770 4154 5782 4156
rect 5802 4344 5814 4346
rect 5802 4336 5804 4344
rect 5812 4336 5814 4344
rect 5802 4164 5814 4336
rect 5802 4156 5804 4164
rect 5812 4156 5814 4164
rect 5802 4154 5814 4156
rect 5802 4124 5814 4126
rect 5802 4116 5804 4124
rect 5812 4116 5814 4124
rect 5802 3904 5814 4116
rect 5802 3896 5804 3904
rect 5812 3896 5814 3904
rect 5802 3894 5814 3896
rect 5610 3716 5612 3724
rect 5620 3716 5622 3724
rect 5610 3664 5622 3716
rect 5834 3724 5846 4696
rect 5866 4144 5878 4836
rect 5866 4136 5868 4144
rect 5876 4136 5878 4144
rect 5866 4134 5878 4136
rect 5920 4614 5984 5006
rect 6058 5104 6070 5106
rect 6058 5096 6060 5104
rect 6068 5096 6070 5104
rect 6058 4944 6070 5096
rect 6058 4936 6060 4944
rect 6068 4936 6070 4944
rect 5920 4606 5924 4614
rect 5932 4606 5936 4614
rect 5944 4606 5948 4614
rect 5956 4606 5960 4614
rect 5968 4606 5972 4614
rect 5980 4606 5984 4614
rect 5920 4214 5984 4606
rect 5920 4206 5924 4214
rect 5932 4206 5936 4214
rect 5944 4206 5948 4214
rect 5956 4206 5960 4214
rect 5968 4206 5972 4214
rect 5980 4206 5984 4214
rect 5920 3814 5984 4206
rect 6026 4784 6038 4786
rect 6026 4776 6028 4784
rect 6036 4776 6038 4784
rect 6026 4244 6038 4776
rect 6026 4236 6028 4244
rect 6036 4236 6038 4244
rect 6026 4144 6038 4236
rect 6026 4136 6028 4144
rect 6036 4136 6038 4144
rect 6026 4134 6038 4136
rect 6058 4504 6070 4936
rect 6058 4496 6060 4504
rect 6068 4496 6070 4504
rect 6058 4324 6070 4496
rect 6090 4444 6102 5196
rect 6122 5204 6134 5256
rect 6122 5196 6124 5204
rect 6132 5196 6134 5204
rect 6122 5194 6134 5196
rect 6218 5264 6230 5266
rect 6218 5256 6220 5264
rect 6228 5256 6230 5264
rect 6186 5084 6198 5086
rect 6186 5076 6188 5084
rect 6196 5076 6198 5084
rect 6154 4964 6166 4966
rect 6154 4956 6156 4964
rect 6164 4956 6166 4964
rect 6154 4924 6166 4956
rect 6154 4916 6156 4924
rect 6164 4916 6166 4924
rect 6154 4914 6166 4916
rect 6186 4724 6198 5076
rect 6186 4716 6188 4724
rect 6196 4716 6198 4724
rect 6186 4714 6198 4716
rect 6186 4664 6198 4666
rect 6186 4656 6188 4664
rect 6196 4656 6198 4664
rect 6186 4604 6198 4656
rect 6218 4664 6230 5256
rect 6218 4656 6220 4664
rect 6228 4656 6230 4664
rect 6218 4654 6230 4656
rect 6250 4704 6262 4706
rect 6250 4696 6252 4704
rect 6260 4696 6262 4704
rect 6186 4596 6188 4604
rect 6196 4596 6198 4604
rect 6186 4594 6198 4596
rect 6090 4436 6092 4444
rect 6100 4436 6102 4444
rect 6090 4434 6102 4436
rect 6154 4564 6166 4566
rect 6154 4556 6156 4564
rect 6164 4556 6166 4564
rect 6058 4316 6060 4324
rect 6068 4316 6070 4324
rect 6058 4124 6070 4316
rect 6090 4364 6102 4366
rect 6090 4356 6092 4364
rect 6100 4356 6102 4364
rect 6090 4264 6102 4356
rect 6090 4256 6092 4264
rect 6100 4256 6102 4264
rect 6090 4254 6102 4256
rect 6122 4364 6134 4366
rect 6122 4356 6124 4364
rect 6132 4356 6134 4364
rect 6122 4204 6134 4356
rect 6122 4196 6124 4204
rect 6132 4196 6134 4204
rect 6122 4194 6134 4196
rect 6058 4116 6060 4124
rect 6068 4116 6070 4124
rect 6058 4114 6070 4116
rect 6154 4084 6166 4556
rect 6250 4144 6262 4696
rect 6410 4624 6422 5316
rect 6602 5304 6614 5306
rect 6602 5296 6604 5304
rect 6612 5296 6614 5304
rect 6410 4616 6412 4624
rect 6420 4616 6422 4624
rect 6410 4614 6422 4616
rect 6442 5264 6454 5266
rect 6442 5256 6444 5264
rect 6452 5256 6454 5264
rect 6378 4604 6390 4606
rect 6378 4596 6380 4604
rect 6388 4596 6390 4604
rect 6282 4584 6294 4586
rect 6282 4576 6284 4584
rect 6292 4576 6294 4584
rect 6282 4204 6294 4576
rect 6378 4244 6390 4596
rect 6378 4236 6380 4244
rect 6388 4236 6390 4244
rect 6378 4234 6390 4236
rect 6410 4244 6422 4246
rect 6410 4236 6412 4244
rect 6420 4236 6422 4244
rect 6282 4196 6284 4204
rect 6292 4196 6294 4204
rect 6282 4194 6294 4196
rect 6314 4224 6326 4226
rect 6314 4216 6316 4224
rect 6324 4216 6326 4224
rect 6250 4136 6252 4144
rect 6260 4136 6262 4144
rect 6250 4134 6262 4136
rect 6154 4076 6156 4084
rect 6164 4076 6166 4084
rect 6154 4074 6166 4076
rect 6314 4064 6326 4216
rect 6314 4056 6316 4064
rect 6324 4056 6326 4064
rect 6314 4054 6326 4056
rect 5920 3806 5924 3814
rect 5932 3806 5936 3814
rect 5944 3806 5948 3814
rect 5956 3806 5960 3814
rect 5968 3806 5972 3814
rect 5980 3806 5984 3814
rect 5834 3716 5836 3724
rect 5844 3716 5846 3724
rect 5834 3714 5846 3716
rect 5866 3784 5878 3786
rect 5866 3776 5868 3784
rect 5876 3776 5878 3784
rect 5610 3656 5612 3664
rect 5620 3656 5622 3664
rect 5610 3654 5622 3656
rect 5610 3584 5622 3586
rect 5610 3576 5612 3584
rect 5620 3576 5622 3584
rect 5610 3304 5622 3576
rect 5674 3584 5686 3586
rect 5674 3576 5676 3584
rect 5684 3576 5686 3584
rect 5610 3296 5612 3304
rect 5620 3296 5622 3304
rect 5610 3294 5622 3296
rect 5642 3504 5654 3506
rect 5642 3496 5644 3504
rect 5652 3496 5654 3504
rect 5642 3204 5654 3496
rect 5642 3196 5644 3204
rect 5652 3196 5654 3204
rect 5642 3194 5654 3196
rect 5674 3204 5686 3576
rect 5866 3584 5878 3776
rect 5866 3576 5868 3584
rect 5876 3576 5878 3584
rect 5866 3574 5878 3576
rect 5834 3544 5846 3546
rect 5834 3536 5836 3544
rect 5844 3536 5846 3544
rect 5770 3524 5782 3526
rect 5770 3516 5772 3524
rect 5780 3516 5782 3524
rect 5674 3196 5676 3204
rect 5684 3196 5686 3204
rect 5674 3194 5686 3196
rect 5738 3244 5750 3246
rect 5738 3236 5740 3244
rect 5748 3236 5750 3244
rect 5578 3096 5580 3104
rect 5588 3096 5590 3104
rect 5514 2416 5516 2424
rect 5524 2416 5526 2424
rect 5450 2176 5452 2184
rect 5460 2176 5462 2184
rect 5450 2174 5462 2176
rect 5514 2124 5526 2416
rect 5514 2116 5516 2124
rect 5524 2116 5526 2124
rect 5514 2114 5526 2116
rect 5546 2484 5558 2486
rect 5546 2476 5548 2484
rect 5556 2476 5558 2484
rect 5290 2076 5292 2084
rect 5300 2076 5302 2084
rect 5290 2074 5302 2076
rect 5386 2084 5398 2086
rect 5386 2076 5388 2084
rect 5396 2076 5398 2084
rect 5258 1916 5260 1924
rect 5268 1916 5270 1924
rect 5258 1914 5270 1916
rect 5130 1876 5132 1884
rect 5140 1876 5142 1884
rect 5130 1744 5142 1876
rect 5130 1736 5132 1744
rect 5140 1736 5142 1744
rect 5130 1734 5142 1736
rect 5066 1724 5078 1726
rect 5066 1716 5068 1724
rect 5076 1716 5078 1724
rect 5002 1524 5014 1526
rect 5002 1516 5004 1524
rect 5012 1516 5014 1524
rect 4842 1296 4844 1304
rect 4852 1296 4854 1304
rect 4842 1294 4854 1296
rect 4874 1444 4886 1446
rect 4874 1436 4876 1444
rect 4884 1436 4886 1444
rect 4810 996 4812 1004
rect 4820 996 4822 1004
rect 4714 736 4716 744
rect 4724 736 4726 744
rect 4714 734 4726 736
rect 4746 804 4758 806
rect 4746 796 4748 804
rect 4756 796 4758 804
rect 4682 696 4684 704
rect 4692 696 4694 704
rect 4682 694 4694 696
rect 4746 504 4758 796
rect 4810 564 4822 996
rect 4874 804 4886 1436
rect 4906 1424 4918 1426
rect 4906 1416 4908 1424
rect 4916 1416 4918 1424
rect 4906 1224 4918 1416
rect 4906 1216 4908 1224
rect 4916 1216 4918 1224
rect 4906 1214 4918 1216
rect 4938 1204 4950 1206
rect 4938 1196 4940 1204
rect 4948 1196 4950 1204
rect 4874 796 4876 804
rect 4884 796 4886 804
rect 4874 794 4886 796
rect 4906 1184 4918 1186
rect 4906 1176 4908 1184
rect 4916 1176 4918 1184
rect 4810 556 4812 564
rect 4820 556 4822 564
rect 4810 554 4822 556
rect 4874 724 4886 726
rect 4874 716 4876 724
rect 4884 716 4886 724
rect 4746 496 4748 504
rect 4756 496 4758 504
rect 4746 494 4758 496
rect 4778 504 4790 506
rect 4778 496 4780 504
rect 4788 496 4790 504
rect 4554 436 4556 444
rect 4564 436 4566 444
rect 4554 434 4566 436
rect 4416 406 4420 414
rect 4428 406 4432 414
rect 4440 406 4444 414
rect 4452 406 4456 414
rect 4464 406 4468 414
rect 4476 406 4480 414
rect 4234 16 4236 24
rect 4244 16 4246 24
rect 4234 14 4246 16
rect 4416 14 4480 406
rect 4714 424 4726 426
rect 4714 416 4716 424
rect 4724 416 4726 424
rect 4714 84 4726 416
rect 4714 76 4716 84
rect 4724 76 4726 84
rect 4714 74 4726 76
rect 4778 24 4790 496
rect 4874 324 4886 716
rect 4906 624 4918 1176
rect 4938 1064 4950 1196
rect 4970 1164 4982 1166
rect 4970 1156 4972 1164
rect 4980 1156 4982 1164
rect 4970 1104 4982 1156
rect 4970 1096 4972 1104
rect 4980 1096 4982 1104
rect 4970 1094 4982 1096
rect 4938 1056 4940 1064
rect 4948 1056 4950 1064
rect 4938 1054 4950 1056
rect 5002 924 5014 1516
rect 5066 1384 5078 1716
rect 5066 1376 5068 1384
rect 5076 1376 5078 1384
rect 5066 1374 5078 1376
rect 5258 1684 5270 1686
rect 5258 1676 5260 1684
rect 5268 1676 5270 1684
rect 5258 1004 5270 1676
rect 5386 1564 5398 2076
rect 5482 2064 5494 2066
rect 5482 2056 5484 2064
rect 5492 2056 5494 2064
rect 5450 2024 5462 2026
rect 5450 2016 5452 2024
rect 5460 2016 5462 2024
rect 5450 1944 5462 2016
rect 5450 1936 5452 1944
rect 5460 1936 5462 1944
rect 5450 1934 5462 1936
rect 5418 1764 5430 1766
rect 5418 1756 5420 1764
rect 5428 1756 5430 1764
rect 5418 1604 5430 1756
rect 5418 1596 5420 1604
rect 5428 1596 5430 1604
rect 5418 1594 5430 1596
rect 5386 1556 5388 1564
rect 5396 1556 5398 1564
rect 5386 1554 5398 1556
rect 5482 1124 5494 2056
rect 5546 1884 5558 2476
rect 5546 1876 5548 1884
rect 5556 1876 5558 1884
rect 5546 1874 5558 1876
rect 5578 2284 5590 3096
rect 5610 3124 5622 3126
rect 5610 3116 5612 3124
rect 5620 3116 5622 3124
rect 5610 2644 5622 3116
rect 5610 2636 5612 2644
rect 5620 2636 5622 2644
rect 5610 2634 5622 2636
rect 5578 2276 5580 2284
rect 5588 2276 5590 2284
rect 5578 1864 5590 2276
rect 5610 2284 5622 2286
rect 5610 2276 5612 2284
rect 5620 2276 5622 2284
rect 5610 2144 5622 2276
rect 5610 2136 5612 2144
rect 5620 2136 5622 2144
rect 5610 2134 5622 2136
rect 5642 2244 5654 2246
rect 5642 2236 5644 2244
rect 5652 2236 5654 2244
rect 5578 1856 5580 1864
rect 5588 1856 5590 1864
rect 5578 1854 5590 1856
rect 5546 1724 5558 1726
rect 5546 1716 5548 1724
rect 5556 1716 5558 1724
rect 5546 1464 5558 1716
rect 5546 1456 5548 1464
rect 5556 1456 5558 1464
rect 5546 1454 5558 1456
rect 5482 1116 5484 1124
rect 5492 1116 5494 1124
rect 5482 1114 5494 1116
rect 5258 996 5260 1004
rect 5268 996 5270 1004
rect 5258 994 5270 996
rect 5354 1104 5366 1106
rect 5354 1096 5356 1104
rect 5364 1096 5366 1104
rect 5002 916 5004 924
rect 5012 916 5014 924
rect 5002 914 5014 916
rect 5322 884 5334 886
rect 5322 876 5324 884
rect 5332 876 5334 884
rect 4906 616 4908 624
rect 4916 616 4918 624
rect 4906 614 4918 616
rect 5066 864 5078 866
rect 5066 856 5068 864
rect 5076 856 5078 864
rect 4874 316 4876 324
rect 4884 316 4886 324
rect 4874 314 4886 316
rect 4778 16 4780 24
rect 4788 16 4790 24
rect 4778 14 4790 16
rect 5066 24 5078 856
rect 5226 824 5238 826
rect 5226 816 5228 824
rect 5236 816 5238 824
rect 5226 564 5238 816
rect 5226 556 5228 564
rect 5236 556 5238 564
rect 5226 554 5238 556
rect 5258 624 5270 626
rect 5258 616 5260 624
rect 5268 616 5270 624
rect 5258 464 5270 616
rect 5258 456 5260 464
rect 5268 456 5270 464
rect 5258 454 5270 456
rect 5322 304 5334 876
rect 5354 784 5366 1096
rect 5546 1104 5558 1106
rect 5546 1096 5548 1104
rect 5556 1096 5558 1104
rect 5418 1004 5430 1006
rect 5418 996 5420 1004
rect 5428 996 5430 1004
rect 5418 824 5430 996
rect 5418 816 5420 824
rect 5428 816 5430 824
rect 5418 814 5430 816
rect 5354 776 5356 784
rect 5364 776 5366 784
rect 5354 774 5366 776
rect 5482 524 5526 526
rect 5482 516 5484 524
rect 5492 516 5526 524
rect 5482 514 5526 516
rect 5514 504 5526 514
rect 5514 496 5516 504
rect 5524 496 5526 504
rect 5514 494 5526 496
rect 5546 324 5558 1096
rect 5578 1104 5590 1106
rect 5578 1096 5580 1104
rect 5588 1096 5590 1104
rect 5578 1064 5590 1096
rect 5578 1056 5580 1064
rect 5588 1056 5590 1064
rect 5578 1054 5590 1056
rect 5642 724 5654 2236
rect 5738 1844 5750 3236
rect 5770 2744 5782 3516
rect 5770 2736 5772 2744
rect 5780 2736 5782 2744
rect 5770 2734 5782 2736
rect 5802 3524 5814 3526
rect 5802 3516 5804 3524
rect 5812 3516 5814 3524
rect 5802 2744 5814 3516
rect 5834 3324 5846 3536
rect 5834 3316 5836 3324
rect 5844 3316 5846 3324
rect 5834 3314 5846 3316
rect 5920 3414 5984 3806
rect 6218 4004 6230 4006
rect 6218 3996 6220 4004
rect 6228 3996 6230 4004
rect 6218 3584 6230 3996
rect 6410 3904 6422 4236
rect 6442 4024 6454 5256
rect 6538 5004 6550 5006
rect 6538 4996 6540 5004
rect 6548 4996 6550 5004
rect 6538 4964 6550 4996
rect 6538 4956 6540 4964
rect 6548 4956 6550 4964
rect 6538 4954 6550 4956
rect 6538 4924 6550 4926
rect 6538 4916 6540 4924
rect 6548 4916 6550 4924
rect 6442 4016 6444 4024
rect 6452 4016 6454 4024
rect 6442 4014 6454 4016
rect 6474 4504 6486 4506
rect 6474 4496 6476 4504
rect 6484 4496 6486 4504
rect 6410 3896 6412 3904
rect 6420 3896 6422 3904
rect 6410 3894 6422 3896
rect 6474 3924 6486 4496
rect 6538 4484 6550 4916
rect 6538 4476 6540 4484
rect 6548 4476 6550 4484
rect 6538 4474 6550 4476
rect 6570 4724 6582 4726
rect 6570 4716 6572 4724
rect 6580 4716 6582 4724
rect 6570 4384 6582 4716
rect 6602 4484 6614 5296
rect 6890 5204 6902 5206
rect 6890 5196 6892 5204
rect 6900 5196 6902 5204
rect 6698 5164 6710 5166
rect 6698 5156 6700 5164
rect 6708 5156 6710 5164
rect 6634 5084 6646 5086
rect 6634 5076 6636 5084
rect 6644 5076 6646 5084
rect 6634 4664 6646 5076
rect 6666 4984 6678 4986
rect 6666 4976 6668 4984
rect 6676 4976 6678 4984
rect 6666 4704 6678 4976
rect 6666 4696 6668 4704
rect 6676 4696 6678 4704
rect 6666 4694 6678 4696
rect 6634 4656 6636 4664
rect 6644 4656 6646 4664
rect 6634 4654 6646 4656
rect 6698 4664 6710 5156
rect 6698 4656 6700 4664
rect 6708 4656 6710 4664
rect 6698 4654 6710 4656
rect 6730 5164 6742 5166
rect 6730 5156 6732 5164
rect 6740 5156 6742 5164
rect 6698 4564 6710 4566
rect 6698 4556 6700 4564
rect 6708 4556 6710 4564
rect 6602 4476 6604 4484
rect 6612 4476 6614 4484
rect 6602 4474 6614 4476
rect 6634 4524 6646 4526
rect 6634 4516 6636 4524
rect 6644 4516 6646 4524
rect 6570 4376 6572 4384
rect 6580 4376 6582 4384
rect 6570 4324 6582 4376
rect 6570 4316 6572 4324
rect 6580 4316 6582 4324
rect 6570 4314 6582 4316
rect 6474 3916 6476 3924
rect 6484 3916 6486 3924
rect 6410 3844 6422 3846
rect 6410 3836 6412 3844
rect 6420 3836 6422 3844
rect 6218 3576 6220 3584
rect 6228 3576 6230 3584
rect 6218 3574 6230 3576
rect 6346 3764 6358 3766
rect 6346 3756 6348 3764
rect 6356 3756 6358 3764
rect 5920 3406 5924 3414
rect 5932 3406 5936 3414
rect 5944 3406 5948 3414
rect 5956 3406 5960 3414
rect 5968 3406 5972 3414
rect 5980 3406 5984 3414
rect 5834 3164 5846 3166
rect 5834 3156 5836 3164
rect 5844 3156 5846 3164
rect 5834 2784 5846 3156
rect 5834 2776 5836 2784
rect 5844 2776 5846 2784
rect 5834 2774 5846 2776
rect 5920 3014 5984 3406
rect 6346 3404 6358 3756
rect 6346 3396 6348 3404
rect 6356 3396 6358 3404
rect 6346 3394 6358 3396
rect 5920 3006 5924 3014
rect 5932 3006 5936 3014
rect 5944 3006 5948 3014
rect 5956 3006 5960 3014
rect 5968 3006 5972 3014
rect 5980 3006 5984 3014
rect 5802 2736 5804 2744
rect 5812 2736 5814 2744
rect 5802 2734 5814 2736
rect 5920 2614 5984 3006
rect 6218 3324 6230 3326
rect 6218 3316 6220 3324
rect 6228 3316 6230 3324
rect 6218 2944 6230 3316
rect 6218 2936 6220 2944
rect 6228 2936 6230 2944
rect 6218 2934 6230 2936
rect 6250 3144 6262 3146
rect 6250 3136 6252 3144
rect 6260 3136 6262 3144
rect 5920 2606 5924 2614
rect 5932 2606 5936 2614
rect 5944 2606 5948 2614
rect 5956 2606 5960 2614
rect 5968 2606 5972 2614
rect 5980 2606 5984 2614
rect 5770 2324 5782 2326
rect 5770 2316 5772 2324
rect 5780 2316 5782 2324
rect 5770 2284 5782 2316
rect 5770 2276 5772 2284
rect 5780 2276 5782 2284
rect 5770 2274 5782 2276
rect 5866 2224 5878 2226
rect 5866 2216 5868 2224
rect 5876 2216 5878 2224
rect 5738 1836 5740 1844
rect 5748 1836 5750 1844
rect 5706 1784 5718 1786
rect 5706 1776 5708 1784
rect 5716 1776 5718 1784
rect 5706 1704 5718 1776
rect 5706 1696 5708 1704
rect 5716 1696 5718 1704
rect 5706 1694 5718 1696
rect 5738 1524 5750 1836
rect 5834 2164 5846 2166
rect 5834 2156 5836 2164
rect 5844 2156 5846 2164
rect 5834 1744 5846 2156
rect 5834 1736 5836 1744
rect 5844 1736 5846 1744
rect 5834 1734 5846 1736
rect 5738 1516 5740 1524
rect 5748 1516 5750 1524
rect 5738 1514 5750 1516
rect 5866 1524 5878 2216
rect 5866 1516 5868 1524
rect 5876 1516 5878 1524
rect 5866 1124 5878 1516
rect 5866 1116 5868 1124
rect 5876 1116 5878 1124
rect 5866 1114 5878 1116
rect 5920 2214 5984 2606
rect 6218 2684 6230 2686
rect 6218 2676 6220 2684
rect 6228 2676 6230 2684
rect 6122 2564 6134 2566
rect 6122 2556 6124 2564
rect 6132 2556 6134 2564
rect 6058 2344 6070 2346
rect 6058 2336 6060 2344
rect 6068 2336 6070 2344
rect 5920 2206 5924 2214
rect 5932 2206 5936 2214
rect 5944 2206 5948 2214
rect 5956 2206 5960 2214
rect 5968 2206 5972 2214
rect 5980 2206 5984 2214
rect 5920 1814 5984 2206
rect 6026 2284 6038 2286
rect 6026 2276 6028 2284
rect 6036 2276 6038 2284
rect 6026 2124 6038 2276
rect 6058 2204 6070 2336
rect 6122 2304 6134 2556
rect 6122 2296 6124 2304
rect 6132 2296 6134 2304
rect 6122 2294 6134 2296
rect 6218 2264 6230 2676
rect 6218 2256 6220 2264
rect 6228 2256 6230 2264
rect 6218 2254 6230 2256
rect 6058 2196 6060 2204
rect 6068 2196 6070 2204
rect 6058 2194 6070 2196
rect 6026 2116 6028 2124
rect 6036 2116 6038 2124
rect 6026 2114 6038 2116
rect 6058 2104 6070 2106
rect 6058 2096 6060 2104
rect 6068 2096 6070 2104
rect 6058 2044 6070 2096
rect 6058 2036 6060 2044
rect 6068 2036 6070 2044
rect 6058 2034 6070 2036
rect 6026 1924 6038 1926
rect 6026 1916 6028 1924
rect 6036 1916 6038 1924
rect 6026 1884 6038 1916
rect 6026 1876 6028 1884
rect 6036 1876 6038 1884
rect 6026 1874 6038 1876
rect 5920 1806 5924 1814
rect 5932 1806 5936 1814
rect 5944 1806 5948 1814
rect 5956 1806 5960 1814
rect 5968 1806 5972 1814
rect 5980 1806 5984 1814
rect 5920 1414 5984 1806
rect 5920 1406 5924 1414
rect 5932 1406 5936 1414
rect 5944 1406 5948 1414
rect 5956 1406 5960 1414
rect 5968 1406 5972 1414
rect 5980 1406 5984 1414
rect 5738 1064 5750 1066
rect 5738 1056 5740 1064
rect 5748 1056 5750 1064
rect 5738 904 5750 1056
rect 5738 896 5740 904
rect 5748 896 5750 904
rect 5738 894 5750 896
rect 5866 1024 5878 1026
rect 5866 1016 5868 1024
rect 5876 1016 5878 1024
rect 5802 824 5814 826
rect 5802 816 5804 824
rect 5812 816 5814 824
rect 5642 716 5644 724
rect 5652 716 5654 724
rect 5642 714 5654 716
rect 5674 784 5686 786
rect 5674 776 5676 784
rect 5684 776 5686 784
rect 5674 564 5686 776
rect 5674 556 5676 564
rect 5684 556 5686 564
rect 5674 554 5686 556
rect 5770 724 5782 726
rect 5770 716 5772 724
rect 5780 716 5782 724
rect 5546 316 5548 324
rect 5556 316 5558 324
rect 5546 314 5558 316
rect 5738 544 5750 546
rect 5738 536 5740 544
rect 5748 536 5750 544
rect 5322 296 5324 304
rect 5332 296 5334 304
rect 5322 294 5334 296
rect 5738 284 5750 536
rect 5770 444 5782 716
rect 5802 584 5814 816
rect 5802 576 5804 584
rect 5812 576 5814 584
rect 5802 574 5814 576
rect 5834 604 5846 606
rect 5834 596 5836 604
rect 5844 596 5846 604
rect 5770 436 5772 444
rect 5780 436 5782 444
rect 5770 434 5782 436
rect 5834 424 5846 596
rect 5834 416 5836 424
rect 5844 416 5846 424
rect 5834 414 5846 416
rect 5866 344 5878 1016
rect 5866 336 5868 344
rect 5876 336 5878 344
rect 5866 334 5878 336
rect 5920 1014 5984 1406
rect 6026 1824 6038 1826
rect 6026 1816 6028 1824
rect 6036 1816 6038 1824
rect 6026 1224 6038 1816
rect 6186 1824 6198 1826
rect 6186 1816 6188 1824
rect 6196 1816 6198 1824
rect 6186 1404 6198 1816
rect 6250 1524 6262 3136
rect 6410 2924 6422 3836
rect 6474 3544 6486 3916
rect 6474 3536 6476 3544
rect 6484 3536 6486 3544
rect 6442 3484 6454 3486
rect 6442 3476 6444 3484
rect 6452 3476 6454 3484
rect 6442 2984 6454 3476
rect 6474 3484 6486 3536
rect 6474 3476 6476 3484
rect 6484 3476 6486 3484
rect 6474 3474 6486 3476
rect 6538 4104 6550 4106
rect 6538 4096 6540 4104
rect 6548 4096 6550 4104
rect 6442 2976 6444 2984
rect 6452 2976 6454 2984
rect 6442 2974 6454 2976
rect 6506 3424 6518 3426
rect 6506 3416 6508 3424
rect 6516 3416 6518 3424
rect 6506 2964 6518 3416
rect 6538 3424 6550 4096
rect 6634 3644 6646 4516
rect 6698 4504 6710 4556
rect 6698 4496 6700 4504
rect 6708 4496 6710 4504
rect 6666 4404 6678 4406
rect 6666 4396 6668 4404
rect 6676 4396 6678 4404
rect 6666 4344 6678 4396
rect 6666 4336 6668 4344
rect 6676 4336 6678 4344
rect 6666 4334 6678 4336
rect 6634 3636 6636 3644
rect 6644 3636 6646 3644
rect 6634 3634 6646 3636
rect 6666 4144 6678 4146
rect 6666 4136 6668 4144
rect 6676 4136 6678 4144
rect 6538 3416 6540 3424
rect 6548 3416 6550 3424
rect 6538 3414 6550 3416
rect 6602 3484 6614 3486
rect 6602 3476 6604 3484
rect 6612 3476 6614 3484
rect 6602 3304 6614 3476
rect 6602 3296 6604 3304
rect 6612 3296 6614 3304
rect 6602 3294 6614 3296
rect 6506 2956 6508 2964
rect 6516 2956 6518 2964
rect 6506 2954 6518 2956
rect 6666 3044 6678 4136
rect 6666 3036 6668 3044
rect 6676 3036 6678 3044
rect 6410 2916 6412 2924
rect 6420 2916 6422 2924
rect 6282 2844 6294 2846
rect 6282 2836 6284 2844
rect 6292 2836 6294 2844
rect 6282 2404 6294 2836
rect 6410 2524 6422 2916
rect 6506 2764 6518 2766
rect 6506 2756 6508 2764
rect 6516 2756 6518 2764
rect 6410 2516 6412 2524
rect 6420 2516 6422 2524
rect 6282 2396 6284 2404
rect 6292 2396 6294 2404
rect 6282 2394 6294 2396
rect 6346 2404 6358 2406
rect 6346 2396 6348 2404
rect 6356 2396 6358 2404
rect 6314 2104 6326 2106
rect 6314 2096 6316 2104
rect 6324 2096 6326 2104
rect 6314 1864 6326 2096
rect 6314 1856 6316 1864
rect 6324 1856 6326 1864
rect 6314 1854 6326 1856
rect 6346 1544 6358 2396
rect 6410 1884 6422 2516
rect 6410 1876 6412 1884
rect 6420 1876 6422 1884
rect 6410 1874 6422 1876
rect 6474 2644 6486 2646
rect 6474 2636 6476 2644
rect 6484 2636 6486 2644
rect 6346 1536 6348 1544
rect 6356 1536 6358 1544
rect 6346 1534 6358 1536
rect 6250 1516 6252 1524
rect 6260 1516 6262 1524
rect 6250 1514 6262 1516
rect 6186 1396 6188 1404
rect 6196 1396 6198 1404
rect 6186 1394 6198 1396
rect 6218 1484 6230 1486
rect 6218 1476 6220 1484
rect 6228 1476 6230 1484
rect 6218 1264 6230 1476
rect 6218 1256 6220 1264
rect 6228 1256 6230 1264
rect 6218 1254 6230 1256
rect 6410 1444 6422 1446
rect 6410 1436 6412 1444
rect 6420 1436 6422 1444
rect 6410 1264 6422 1436
rect 6410 1256 6412 1264
rect 6420 1256 6422 1264
rect 6410 1254 6422 1256
rect 6026 1216 6028 1224
rect 6036 1216 6038 1224
rect 6026 1214 6038 1216
rect 5920 1006 5924 1014
rect 5932 1006 5936 1014
rect 5944 1006 5948 1014
rect 5956 1006 5960 1014
rect 5968 1006 5972 1014
rect 5980 1006 5984 1014
rect 5920 614 5984 1006
rect 6122 964 6134 966
rect 6122 956 6124 964
rect 6132 956 6134 964
rect 5920 606 5924 614
rect 5932 606 5936 614
rect 5944 606 5948 614
rect 5956 606 5960 614
rect 5968 606 5972 614
rect 5980 606 5984 614
rect 5738 276 5740 284
rect 5748 276 5750 284
rect 5738 274 5750 276
rect 5482 264 5494 266
rect 5482 256 5484 264
rect 5492 256 5494 264
rect 5482 164 5494 256
rect 5920 214 5984 606
rect 6026 704 6038 706
rect 6026 696 6028 704
rect 6036 696 6038 704
rect 6026 464 6038 696
rect 6122 664 6134 956
rect 6186 944 6198 946
rect 6186 936 6188 944
rect 6196 936 6198 944
rect 6122 656 6124 664
rect 6132 656 6134 664
rect 6122 654 6134 656
rect 6154 664 6166 666
rect 6154 656 6156 664
rect 6164 656 6166 664
rect 6026 456 6028 464
rect 6036 456 6038 464
rect 6026 454 6038 456
rect 5920 206 5924 214
rect 5932 206 5936 214
rect 5944 206 5948 214
rect 5956 206 5960 214
rect 5968 206 5972 214
rect 5980 206 5984 214
rect 5482 156 5484 164
rect 5492 156 5494 164
rect 5482 154 5494 156
rect 5610 204 5622 206
rect 5610 196 5612 204
rect 5620 196 5622 204
rect 5610 144 5622 196
rect 5610 136 5612 144
rect 5620 136 5622 144
rect 5610 134 5622 136
rect 5066 16 5068 24
rect 5076 16 5078 24
rect 5066 14 5078 16
rect 4416 6 4420 14
rect 4428 6 4432 14
rect 4440 6 4444 14
rect 4452 6 4456 14
rect 4464 6 4468 14
rect 4476 6 4480 14
rect 4416 -10 4480 6
rect 5920 -10 5984 206
rect 6154 264 6166 656
rect 6154 256 6156 264
rect 6164 256 6166 264
rect 6154 184 6166 256
rect 6186 224 6198 936
rect 6474 844 6486 2636
rect 6506 1524 6518 2756
rect 6666 2704 6678 3036
rect 6666 2696 6668 2704
rect 6676 2696 6678 2704
rect 6634 2684 6646 2686
rect 6634 2676 6636 2684
rect 6644 2676 6646 2684
rect 6634 2284 6646 2676
rect 6666 2664 6678 2696
rect 6666 2656 6668 2664
rect 6676 2656 6678 2664
rect 6666 2654 6678 2656
rect 6698 3324 6710 4496
rect 6730 3984 6742 5156
rect 6826 5044 6838 5046
rect 6826 5036 6828 5044
rect 6836 5036 6838 5044
rect 6730 3976 6732 3984
rect 6740 3976 6742 3984
rect 6730 3974 6742 3976
rect 6762 4704 6774 4706
rect 6762 4696 6764 4704
rect 6772 4696 6774 4704
rect 6762 3804 6774 4696
rect 6762 3796 6764 3804
rect 6772 3796 6774 3804
rect 6762 3794 6774 3796
rect 6794 4404 6806 4406
rect 6794 4396 6796 4404
rect 6804 4396 6806 4404
rect 6794 3564 6806 4396
rect 6794 3556 6796 3564
rect 6804 3556 6806 3564
rect 6794 3554 6806 3556
rect 6826 3524 6838 5036
rect 6890 4164 6902 5196
rect 6890 4156 6892 4164
rect 6900 4156 6902 4164
rect 6890 4154 6902 4156
rect 6954 4804 6966 4806
rect 6954 4796 6956 4804
rect 6964 4796 6966 4804
rect 6922 4044 6934 4046
rect 6922 4036 6924 4044
rect 6932 4036 6934 4044
rect 6826 3516 6828 3524
rect 6836 3516 6838 3524
rect 6826 3514 6838 3516
rect 6858 3644 6870 3646
rect 6858 3636 6860 3644
rect 6868 3636 6870 3644
rect 6698 3316 6700 3324
rect 6708 3316 6710 3324
rect 6698 3084 6710 3316
rect 6698 3076 6700 3084
rect 6708 3076 6710 3084
rect 6634 2276 6636 2284
rect 6644 2276 6646 2284
rect 6634 2274 6646 2276
rect 6570 2164 6582 2166
rect 6570 2156 6572 2164
rect 6580 2156 6582 2164
rect 6570 1744 6582 2156
rect 6698 2004 6710 3076
rect 6858 2704 6870 3636
rect 6858 2696 6860 2704
rect 6868 2696 6870 2704
rect 6858 2694 6870 2696
rect 6890 3604 6902 3606
rect 6890 3596 6892 3604
rect 6900 3596 6902 3604
rect 6890 2424 6902 3596
rect 6922 2864 6934 4036
rect 6922 2856 6924 2864
rect 6932 2856 6934 2864
rect 6922 2854 6934 2856
rect 6954 3584 6966 4796
rect 6986 4624 6998 5376
rect 7306 5344 7318 5346
rect 7306 5336 7308 5344
rect 7316 5336 7318 5344
rect 7242 5284 7254 5286
rect 7242 5276 7244 5284
rect 7252 5276 7254 5284
rect 6986 4616 6988 4624
rect 6996 4616 6998 4624
rect 6986 4614 6998 4616
rect 7050 4984 7062 4986
rect 7050 4976 7052 4984
rect 7060 4976 7062 4984
rect 6954 3576 6956 3584
rect 6964 3576 6966 3584
rect 6890 2416 6892 2424
rect 6900 2416 6902 2424
rect 6890 2414 6902 2416
rect 6698 1996 6700 2004
rect 6708 1996 6710 2004
rect 6698 1994 6710 1996
rect 6954 1884 6966 3576
rect 7018 4564 7030 4566
rect 7018 4556 7020 4564
rect 7028 4556 7030 4564
rect 6954 1876 6956 1884
rect 6964 1876 6966 1884
rect 6954 1874 6966 1876
rect 6986 3564 6998 3566
rect 6986 3556 6988 3564
rect 6996 3556 6998 3564
rect 6570 1736 6572 1744
rect 6580 1736 6582 1744
rect 6570 1734 6582 1736
rect 6506 1516 6508 1524
rect 6516 1516 6518 1524
rect 6506 1514 6518 1516
rect 6986 1444 6998 3556
rect 7018 3504 7030 4556
rect 7018 3496 7020 3504
rect 7028 3496 7030 3504
rect 7018 3494 7030 3496
rect 7050 3504 7062 4976
rect 7178 4884 7190 4886
rect 7178 4876 7180 4884
rect 7188 4876 7190 4884
rect 7082 4764 7094 4766
rect 7082 4756 7084 4764
rect 7092 4756 7094 4764
rect 7082 4524 7094 4756
rect 7146 4744 7158 4746
rect 7146 4736 7148 4744
rect 7156 4736 7158 4744
rect 7082 4516 7084 4524
rect 7092 4516 7094 4524
rect 7082 4514 7094 4516
rect 7114 4704 7126 4706
rect 7114 4696 7116 4704
rect 7124 4696 7126 4704
rect 7114 4344 7126 4696
rect 7146 4404 7158 4736
rect 7146 4396 7148 4404
rect 7156 4396 7158 4404
rect 7146 4394 7158 4396
rect 7114 4336 7116 4344
rect 7124 4336 7126 4344
rect 7114 4334 7126 4336
rect 7146 4344 7158 4346
rect 7146 4336 7148 4344
rect 7156 4336 7158 4344
rect 7114 4264 7126 4266
rect 7114 4256 7116 4264
rect 7124 4256 7126 4264
rect 7050 3496 7052 3504
rect 7060 3496 7062 3504
rect 7050 3494 7062 3496
rect 7082 4104 7094 4106
rect 7082 4096 7084 4104
rect 7092 4096 7094 4104
rect 7018 2664 7030 2666
rect 7018 2656 7020 2664
rect 7028 2656 7030 2664
rect 7018 1504 7030 2656
rect 7018 1496 7020 1504
rect 7028 1496 7030 1504
rect 7018 1494 7030 1496
rect 6986 1436 6988 1444
rect 6996 1436 6998 1444
rect 6986 1434 6998 1436
rect 6858 1344 6870 1346
rect 6858 1336 6860 1344
rect 6868 1336 6870 1344
rect 6858 1224 6870 1336
rect 6858 1216 6860 1224
rect 6868 1216 6870 1224
rect 6858 1214 6870 1216
rect 6602 1204 6614 1206
rect 6602 1196 6604 1204
rect 6612 1196 6614 1204
rect 6602 964 6614 1196
rect 6602 956 6604 964
rect 6612 956 6614 964
rect 6602 954 6614 956
rect 6474 836 6476 844
rect 6484 836 6486 844
rect 6474 834 6486 836
rect 6762 904 6774 906
rect 6762 896 6764 904
rect 6772 896 6774 904
rect 6762 664 6774 896
rect 7082 704 7094 4096
rect 7114 3664 7126 4256
rect 7114 3656 7116 3664
rect 7124 3656 7126 3664
rect 7114 3654 7126 3656
rect 7146 3644 7158 4336
rect 7178 4244 7190 4876
rect 7178 4236 7180 4244
rect 7188 4236 7190 4244
rect 7178 4234 7190 4236
rect 7210 4624 7222 4626
rect 7210 4616 7212 4624
rect 7220 4616 7222 4624
rect 7210 4184 7222 4616
rect 7242 4224 7254 5276
rect 7242 4216 7244 4224
rect 7252 4216 7254 4224
rect 7242 4214 7254 4216
rect 7274 4724 7286 4726
rect 7274 4716 7276 4724
rect 7284 4716 7286 4724
rect 7210 4176 7212 4184
rect 7220 4176 7222 4184
rect 7210 4174 7222 4176
rect 7242 4124 7254 4126
rect 7242 4116 7244 4124
rect 7252 4116 7254 4124
rect 7146 3636 7148 3644
rect 7156 3636 7158 3644
rect 7146 3634 7158 3636
rect 7178 3924 7190 3926
rect 7178 3916 7180 3924
rect 7188 3916 7190 3924
rect 7146 3304 7158 3306
rect 7146 3296 7148 3304
rect 7156 3296 7158 3304
rect 7146 3164 7158 3296
rect 7178 3304 7190 3916
rect 7178 3296 7180 3304
rect 7188 3296 7190 3304
rect 7178 3294 7190 3296
rect 7210 3544 7222 3546
rect 7210 3536 7212 3544
rect 7220 3536 7222 3544
rect 7146 3156 7148 3164
rect 7156 3156 7158 3164
rect 7146 3154 7158 3156
rect 7178 3164 7190 3166
rect 7178 3156 7180 3164
rect 7188 3156 7190 3164
rect 7114 2984 7126 2986
rect 7114 2976 7116 2984
rect 7124 2976 7126 2984
rect 7114 1864 7126 2976
rect 7114 1856 7116 1864
rect 7124 1856 7126 1864
rect 7114 1854 7126 1856
rect 7146 1764 7158 1766
rect 7146 1756 7148 1764
rect 7156 1756 7158 1764
rect 7114 1724 7126 1726
rect 7114 1716 7116 1724
rect 7124 1716 7126 1724
rect 7114 1364 7126 1716
rect 7114 1356 7116 1364
rect 7124 1356 7126 1364
rect 7114 1304 7126 1356
rect 7114 1296 7116 1304
rect 7124 1296 7126 1304
rect 7114 1294 7126 1296
rect 7146 1344 7158 1756
rect 7178 1704 7190 3156
rect 7210 3004 7222 3536
rect 7242 3104 7254 4116
rect 7274 4084 7286 4716
rect 7306 4144 7318 5336
rect 7306 4136 7308 4144
rect 7316 4136 7318 4144
rect 7306 4134 7318 4136
rect 7274 4076 7276 4084
rect 7284 4076 7286 4084
rect 7274 4074 7286 4076
rect 7306 4084 7318 4086
rect 7306 4076 7308 4084
rect 7316 4076 7318 4084
rect 7242 3096 7244 3104
rect 7252 3096 7254 3104
rect 7242 3094 7254 3096
rect 7274 3504 7286 3506
rect 7274 3496 7276 3504
rect 7284 3496 7286 3504
rect 7210 2996 7212 3004
rect 7220 2996 7222 3004
rect 7210 2994 7222 2996
rect 7178 1696 7180 1704
rect 7188 1696 7190 1704
rect 7178 1694 7190 1696
rect 7210 2384 7222 2386
rect 7210 2376 7212 2384
rect 7220 2376 7222 2384
rect 7146 1336 7148 1344
rect 7156 1336 7158 1344
rect 7082 696 7084 704
rect 7092 696 7094 704
rect 7082 694 7094 696
rect 6762 656 6764 664
rect 6772 656 6774 664
rect 6762 654 6774 656
rect 6186 216 6188 224
rect 6196 216 6198 224
rect 6186 214 6198 216
rect 6410 604 6422 606
rect 6410 596 6412 604
rect 6420 596 6422 604
rect 6154 176 6156 184
rect 6164 176 6166 184
rect 6154 174 6166 176
rect 6186 184 6198 186
rect 6186 176 6188 184
rect 6196 176 6198 184
rect 6186 126 6198 176
rect 6186 114 6230 126
rect 6218 104 6230 114
rect 6218 96 6220 104
rect 6228 96 6230 104
rect 6218 94 6230 96
rect 6410 24 6422 596
rect 6698 604 6710 606
rect 6698 596 6700 604
rect 6708 596 6710 604
rect 6698 264 6710 596
rect 7082 544 7094 546
rect 7082 536 7084 544
rect 7092 536 7094 544
rect 7082 504 7094 536
rect 7082 496 7084 504
rect 7092 496 7094 504
rect 7082 494 7094 496
rect 6698 256 6700 264
rect 6708 256 6710 264
rect 6698 184 6710 256
rect 6698 176 6700 184
rect 6708 176 6710 184
rect 6698 174 6710 176
rect 6986 484 6998 486
rect 6986 476 6988 484
rect 6996 476 6998 484
rect 6986 144 6998 476
rect 6986 136 6988 144
rect 6996 136 6998 144
rect 6986 134 6998 136
rect 7146 104 7158 1336
rect 7178 1164 7190 1166
rect 7178 1156 7180 1164
rect 7188 1156 7190 1164
rect 7178 284 7190 1156
rect 7210 1124 7222 2376
rect 7274 2204 7286 3496
rect 7306 2544 7318 4076
rect 7338 2964 7350 5396
rect 7338 2956 7340 2964
rect 7348 2956 7350 2964
rect 7338 2954 7350 2956
rect 7370 4124 7382 4126
rect 7370 4116 7372 4124
rect 7380 4116 7382 4124
rect 7306 2536 7308 2544
rect 7316 2536 7318 2544
rect 7306 2534 7318 2536
rect 7338 2544 7350 2546
rect 7338 2536 7340 2544
rect 7348 2536 7350 2544
rect 7338 2284 7350 2536
rect 7338 2276 7340 2284
rect 7348 2276 7350 2284
rect 7338 2274 7350 2276
rect 7274 2196 7276 2204
rect 7284 2196 7286 2204
rect 7274 2194 7286 2196
rect 7338 2124 7350 2126
rect 7338 2116 7340 2124
rect 7348 2116 7350 2124
rect 7306 1484 7318 1486
rect 7306 1476 7308 1484
rect 7316 1476 7318 1484
rect 7210 1116 7212 1124
rect 7220 1116 7222 1124
rect 7210 924 7222 1116
rect 7210 916 7212 924
rect 7220 916 7222 924
rect 7210 724 7222 916
rect 7210 716 7212 724
rect 7220 716 7222 724
rect 7210 714 7222 716
rect 7274 1324 7286 1326
rect 7274 1316 7276 1324
rect 7284 1316 7286 1324
rect 7274 324 7286 1316
rect 7306 1084 7318 1476
rect 7338 1104 7350 2116
rect 7370 1424 7382 4116
rect 7402 2504 7414 2506
rect 7402 2496 7404 2504
rect 7412 2496 7414 2504
rect 7402 2264 7414 2496
rect 7402 2256 7404 2264
rect 7412 2256 7414 2264
rect 7402 2254 7414 2256
rect 7370 1416 7372 1424
rect 7380 1416 7382 1424
rect 7370 1414 7382 1416
rect 7402 1704 7414 1706
rect 7402 1696 7404 1704
rect 7412 1696 7414 1704
rect 7402 1664 7414 1696
rect 7402 1656 7404 1664
rect 7412 1656 7414 1664
rect 7402 1404 7414 1656
rect 7402 1396 7404 1404
rect 7412 1396 7414 1404
rect 7402 1394 7414 1396
rect 7338 1096 7340 1104
rect 7348 1096 7350 1104
rect 7338 1094 7350 1096
rect 7306 1076 7308 1084
rect 7316 1076 7318 1084
rect 7306 1074 7318 1076
rect 7274 316 7276 324
rect 7284 316 7286 324
rect 7274 314 7286 316
rect 7178 276 7180 284
rect 7188 276 7190 284
rect 7178 274 7190 276
rect 7146 96 7148 104
rect 7156 96 7158 104
rect 7146 94 7158 96
rect 6410 16 6412 24
rect 6420 16 6422 24
rect 6410 14 6422 16
use BUFX2  _2110_
timestamp 1596991774
transform -1 0 56 0 -1 210
box -4 -6 52 206
use XOR2X1  _2481_
timestamp 1596991774
transform -1 0 168 0 -1 210
box -4 -6 116 206
use XNOR2X1  _2477_
timestamp 1596991774
transform 1 0 168 0 -1 210
box -4 -6 116 206
use NAND2X1  _2488_
timestamp 1596991774
transform 1 0 8 0 1 210
box -4 -6 52 206
use NOR2X1  _2539_
timestamp 1596991774
transform 1 0 56 0 1 210
box -4 -6 52 206
use OAI21X1  _2494_
timestamp 1596991774
transform 1 0 104 0 1 210
box -4 -6 68 206
use NOR2X1  _2489_
timestamp 1596991774
transform -1 0 216 0 1 210
box -4 -6 52 206
use NOR2X1  _2482_
timestamp 1596991774
transform 1 0 280 0 -1 210
box -4 -6 52 206
use XNOR2X1  _2478_
timestamp 1596991774
transform -1 0 440 0 -1 210
box -4 -6 116 206
use INVX1  _2468_
timestamp 1596991774
transform 1 0 216 0 1 210
box -4 -6 36 206
use NAND2X1  _2469_
timestamp 1596991774
transform -1 0 296 0 1 210
box -4 -6 52 206
use INVX1  _2470_
timestamp 1596991774
transform 1 0 296 0 1 210
box -4 -6 36 206
use OAI21X1  _2490_
timestamp 1596991774
transform 1 0 328 0 1 210
box -4 -6 68 206
use NAND2X1  _2471_
timestamp 1596991774
transform 1 0 392 0 1 210
box -4 -6 52 206
use BUFX2  _2109_
timestamp 1596991774
transform 1 0 440 0 -1 210
box -4 -6 52 206
use AOI22X1  _2476_
timestamp 1596991774
transform 1 0 488 0 -1 210
box -4 -6 84 206
use NAND2X1  _2472_
timestamp 1596991774
transform 1 0 568 0 -1 210
box -4 -6 52 206
use NAND2X1  _2487_
timestamp 1596991774
transform -1 0 488 0 1 210
box -4 -6 52 206
use OAI21X1  _2474_
timestamp 1596991774
transform -1 0 552 0 1 210
box -4 -6 68 206
use INVX1  _2464_
timestamp 1596991774
transform -1 0 584 0 1 210
box -4 -6 36 206
use OAI21X1  _2467_
timestamp 1596991774
transform 1 0 584 0 1 210
box -4 -6 68 206
use NAND2X1  _2540_
timestamp 1596991774
transform 1 0 616 0 -1 210
box -4 -6 52 206
use NOR2X1  _2475_
timestamp 1596991774
transform -1 0 712 0 -1 210
box -4 -6 52 206
use XNOR2X1  _2473_
timestamp 1596991774
transform -1 0 824 0 -1 210
box -4 -6 116 206
use NAND2X1  _2466_
timestamp 1596991774
transform -1 0 696 0 1 210
box -4 -6 52 206
use XNOR2X1  _2465_
timestamp 1596991774
transform -1 0 808 0 1 210
box -4 -6 116 206
use INVX1  _3075_
timestamp 1596991774
transform 1 0 808 0 1 210
box -4 -6 36 206
use XOR2X1  _2462_
timestamp 1596991774
transform 1 0 824 0 -1 210
box -4 -6 116 206
use XNOR2X1  _2463_
timestamp 1596991774
transform -1 0 1048 0 -1 210
box -4 -6 116 206
use OAI22X1  _3076_
timestamp 1596991774
transform -1 0 920 0 1 210
box -4 -6 84 206
use INVX1  _3074_
timestamp 1596991774
transform -1 0 952 0 1 210
box -4 -6 36 206
use NOR2X1  _3077_
timestamp 1596991774
transform 1 0 952 0 1 210
box -4 -6 52 206
use OAI22X1  _3073_
timestamp 1596991774
transform 1 0 1000 0 1 210
box -4 -6 84 206
use INVX1  _3126_
timestamp 1596991774
transform 1 0 1048 0 -1 210
box -4 -6 36 206
use OAI22X1  _3128_
timestamp 1596991774
transform 1 0 1080 0 -1 210
box -4 -6 84 206
use INVX1  _3127_
timestamp 1596991774
transform -1 0 1192 0 -1 210
box -4 -6 36 206
use INVX1  _3100_
timestamp 1596991774
transform 1 0 1192 0 -1 210
box -4 -6 36 206
use INVX1  _3071_
timestamp 1596991774
transform -1 0 1112 0 1 210
box -4 -6 36 206
use INVX1  _3072_
timestamp 1596991774
transform -1 0 1144 0 1 210
box -4 -6 36 206
use NAND3X1  _3096_
timestamp 1596991774
transform 1 0 1144 0 1 210
box -4 -6 68 206
use NAND2X1  _3082_
timestamp 1596991774
transform 1 0 1208 0 1 210
box -4 -6 52 206
use OAI22X1  _3102_
timestamp 1596991774
transform 1 0 1224 0 -1 210
box -4 -6 84 206
use INVX1  _3101_
timestamp 1596991774
transform -1 0 1336 0 -1 210
box -4 -6 36 206
use INVX1  _3098_
timestamp 1596991774
transform 1 0 1336 0 -1 210
box -4 -6 36 206
use OAI21X1  _3083_
timestamp 1596991774
transform -1 0 1432 0 -1 210
box -4 -6 68 206
use NOR2X1  _3103_
timestamp 1596991774
transform 1 0 1256 0 1 210
box -4 -6 52 206
use NAND3X1  _3122_
timestamp 1596991774
transform 1 0 1304 0 1 210
box -4 -6 68 206
use OAI22X1  _3099_
timestamp 1596991774
transform -1 0 1448 0 1 210
box -4 -6 84 206
use FILL  SFILL14960x2100
timestamp 1596991774
transform 1 0 1496 0 1 210
box -4 -6 20 206
use FILL  SFILL14800x2100
timestamp 1596991774
transform 1 0 1480 0 1 210
box -4 -6 20 206
use FILL  SFILL14640x2100
timestamp 1596991774
transform 1 0 1464 0 1 210
box -4 -6 20 206
use FILL  SFILL14480x2100
timestamp 1596991774
transform 1 0 1448 0 1 210
box -4 -6 20 206
use FILL  SFILL14800x100
timestamp 1596991774
transform -1 0 1496 0 -1 210
box -4 -6 20 206
use FILL  SFILL14640x100
timestamp 1596991774
transform -1 0 1480 0 -1 210
box -4 -6 20 206
use FILL  SFILL14480x100
timestamp 1596991774
transform -1 0 1464 0 -1 210
box -4 -6 20 206
use FILL  SFILL14320x100
timestamp 1596991774
transform -1 0 1448 0 -1 210
box -4 -6 20 206
use INVX1  _3081_
timestamp 1596991774
transform -1 0 1528 0 -1 210
box -4 -6 36 206
use OAI21X1  _3109_
timestamp 1596991774
transform -1 0 1624 0 1 210
box -4 -6 68 206
use NAND2X1  _3108_
timestamp 1596991774
transform 1 0 1512 0 1 210
box -4 -6 52 206
use INVX1  _3078_
timestamp 1596991774
transform 1 0 1576 0 -1 210
box -4 -6 36 206
use NOR2X1  _3084_
timestamp 1596991774
transform -1 0 1576 0 -1 210
box -4 -6 52 206
use OAI22X1  _3080_
timestamp 1596991774
transform 1 0 1608 0 -1 210
box -4 -6 84 206
use INVX1  _3079_
timestamp 1596991774
transform -1 0 1720 0 -1 210
box -4 -6 36 206
use AOI21X1  _2541_
timestamp 1596991774
transform -1 0 1784 0 -1 210
box -4 -6 68 206
use INVX1  _3104_
timestamp 1596991774
transform -1 0 1816 0 -1 210
box -4 -6 36 206
use INVX1  _3107_
timestamp 1596991774
transform -1 0 1656 0 1 210
box -4 -6 36 206
use NOR2X1  _3110_
timestamp 1596991774
transform -1 0 1704 0 1 210
box -4 -6 52 206
use NAND2X1  _3030_
timestamp 1596991774
transform 1 0 1704 0 1 210
box -4 -6 52 206
use OAI21X1  _3031_
timestamp 1596991774
transform -1 0 1816 0 1 210
box -4 -6 68 206
use OAI22X1  _3106_
timestamp 1596991774
transform 1 0 1816 0 -1 210
box -4 -6 84 206
use INVX1  _3105_
timestamp 1596991774
transform -1 0 1928 0 -1 210
box -4 -6 36 206
use INVX1  _3026_
timestamp 1596991774
transform 1 0 1928 0 -1 210
box -4 -6 36 206
use OAI22X1  _3028_
timestamp 1596991774
transform 1 0 1960 0 -1 210
box -4 -6 84 206
use INVX1  _3029_
timestamp 1596991774
transform -1 0 1848 0 1 210
box -4 -6 36 206
use NAND2X1  _3056_
timestamp 1596991774
transform -1 0 1896 0 1 210
box -4 -6 52 206
use NOR2X1  _3032_
timestamp 1596991774
transform -1 0 1944 0 1 210
box -4 -6 52 206
use INVX1  _3023_
timestamp 1596991774
transform 1 0 1944 0 1 210
box -4 -6 36 206
use OAI22X1  _3024_
timestamp 1596991774
transform -1 0 2056 0 1 210
box -4 -6 84 206
use INVX1  _3027_
timestamp 1596991774
transform 1 0 2040 0 -1 210
box -4 -6 36 206
use INVX1  _3022_
timestamp 1596991774
transform -1 0 2104 0 -1 210
box -4 -6 36 206
use OAI21X1  _2461_
timestamp 1596991774
transform -1 0 2168 0 -1 210
box -4 -6 68 206
use XNOR2X1  _2447_
timestamp 1596991774
transform 1 0 2168 0 -1 210
box -4 -6 116 206
use NAND3X1  _3044_
timestamp 1596991774
transform -1 0 2120 0 1 210
box -4 -6 68 206
use NOR2X1  _3025_
timestamp 1596991774
transform 1 0 2120 0 1 210
box -4 -6 52 206
use OAI22X1  _3021_
timestamp 1596991774
transform 1 0 2168 0 1 210
box -4 -6 84 206
use NAND2X1  _2456_
timestamp 1596991774
transform 1 0 2280 0 -1 210
box -4 -6 52 206
use NOR2X1  _2459_
timestamp 1596991774
transform 1 0 2328 0 -1 210
box -4 -6 52 206
use AOI21X1  _2460_
timestamp 1596991774
transform -1 0 2440 0 -1 210
box -4 -6 68 206
use INVX1  _3020_
timestamp 1596991774
transform 1 0 2248 0 1 210
box -4 -6 36 206
use INVX1  _3019_
timestamp 1596991774
transform -1 0 2312 0 1 210
box -4 -6 36 206
use XNOR2X1  _2454_
timestamp 1596991774
transform -1 0 2424 0 1 210
box -4 -6 116 206
use NAND2X1  _2458_
timestamp 1596991774
transform -1 0 2488 0 -1 210
box -4 -6 52 206
use INVX1  _2457_
timestamp 1596991774
transform -1 0 2520 0 -1 210
box -4 -6 36 206
use NAND3X1  _2537_
timestamp 1596991774
transform 1 0 2520 0 -1 210
box -4 -6 68 206
use AOI21X1  _2453_
timestamp 1596991774
transform -1 0 2648 0 -1 210
box -4 -6 68 206
use INVX1  _3048_
timestamp 1596991774
transform -1 0 2456 0 1 210
box -4 -6 36 206
use XNOR2X1  _2455_
timestamp 1596991774
transform -1 0 2568 0 1 210
box -4 -6 116 206
use OR2X2  _2343_
timestamp 1596991774
transform -1 0 2632 0 1 210
box -4 -6 68 206
use NOR2X1  _2452_
timestamp 1596991774
transform 1 0 2648 0 -1 210
box -4 -6 52 206
use INVX1  _2451_
timestamp 1596991774
transform -1 0 2728 0 -1 210
box -4 -6 36 206
use XNOR2X1  _2446_
timestamp 1596991774
transform -1 0 2840 0 -1 210
box -4 -6 116 206
use INVX1  _2996_
timestamp 1596991774
transform -1 0 2664 0 1 210
box -4 -6 36 206
use XNOR2X1  _2443_
timestamp 1596991774
transform 1 0 2664 0 1 210
box -4 -6 116 206
use NAND2X1  _2437_
timestamp 1596991774
transform -1 0 2824 0 1 210
box -4 -6 52 206
use AND2X2  _2448_
timestamp 1596991774
transform 1 0 2824 0 1 210
box -4 -6 68 206
use BUFX2  _2098_
timestamp 1596991774
transform -1 0 2888 0 -1 210
box -4 -6 52 206
use FILL  SFILL29520x2100
timestamp 1596991774
transform 1 0 2952 0 1 210
box -4 -6 20 206
use FILL  SFILL29360x2100
timestamp 1596991774
transform 1 0 2936 0 1 210
box -4 -6 20 206
use FILL  SFILL29200x2100
timestamp 1596991774
transform 1 0 2920 0 1 210
box -4 -6 20 206
use FILL  SFILL29520x100
timestamp 1596991774
transform -1 0 2968 0 -1 210
box -4 -6 20 206
use INVX1  _2436_
timestamp 1596991774
transform -1 0 2920 0 1 210
box -4 -6 36 206
use AOI21X1  _2445_
timestamp 1596991774
transform 1 0 2888 0 -1 210
box -4 -6 68 206
use FILL  SFILL29680x2100
timestamp 1596991774
transform 1 0 2968 0 1 210
box -4 -6 20 206
use FILL  SFILL30000x100
timestamp 1596991774
transform -1 0 3016 0 -1 210
box -4 -6 20 206
use FILL  SFILL29840x100
timestamp 1596991774
transform -1 0 3000 0 -1 210
box -4 -6 20 206
use FILL  SFILL29680x100
timestamp 1596991774
transform -1 0 2984 0 -1 210
box -4 -6 20 206
use INVX1  _2898_
timestamp 1596991774
transform 1 0 2984 0 1 210
box -4 -6 36 206
use NAND2X1  _2442_
timestamp 1596991774
transform -1 0 3064 0 -1 210
box -4 -6 52 206
use OAI21X1  _2450_
timestamp 1596991774
transform -1 0 3128 0 -1 210
box -4 -6 68 206
use NAND2X1  _2439_
timestamp 1596991774
transform -1 0 3176 0 -1 210
box -4 -6 52 206
use NOR2X1  _2449_
timestamp 1596991774
transform 1 0 3176 0 -1 210
box -4 -6 52 206
use AOI22X1  _2899_
timestamp 1596991774
transform -1 0 3096 0 1 210
box -4 -6 84 206
use INVX1  _2900_
timestamp 1596991774
transform 1 0 3096 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_insert260
timestamp 1596991774
transform -1 0 3176 0 1 210
box -4 -6 52 206
use INVX1  _2897_
timestamp 1596991774
transform 1 0 3176 0 1 210
box -4 -6 36 206
use INVX1  _2611_
timestamp 1596991774
transform 1 0 3208 0 1 210
box -4 -6 36 206
use INVX1  _2438_
timestamp 1596991774
transform -1 0 3256 0 -1 210
box -4 -6 36 206
use NOR2X1  _2444_
timestamp 1596991774
transform 1 0 3256 0 -1 210
box -4 -6 52 206
use NAND2X1  _2441_
timestamp 1596991774
transform -1 0 3352 0 -1 210
box -4 -6 52 206
use INVX1  _2440_
timestamp 1596991774
transform 1 0 3352 0 -1 210
box -4 -6 36 206
use BUFX2  _2107_
timestamp 1596991774
transform 1 0 3384 0 -1 210
box -4 -6 52 206
use AOI22X1  _2613_
timestamp 1596991774
transform 1 0 3240 0 1 210
box -4 -6 84 206
use INVX1  _2612_
timestamp 1596991774
transform -1 0 3352 0 1 210
box -4 -6 36 206
use INVX1  _2614_
timestamp 1596991774
transform -1 0 3384 0 1 210
box -4 -6 36 206
use AOI22X1  _2616_
timestamp 1596991774
transform 1 0 3384 0 1 210
box -4 -6 84 206
use BUFX2  _2106_
timestamp 1596991774
transform 1 0 3432 0 -1 210
box -4 -6 52 206
use BUFX2  _2099_
timestamp 1596991774
transform 1 0 3480 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3638_
timestamp 1596991774
transform -1 0 3720 0 -1 210
box -4 -6 196 206
use NAND2X1  _2617_
timestamp 1596991774
transform -1 0 3512 0 1 210
box -4 -6 52 206
use INVX1  _3384_
timestamp 1596991774
transform -1 0 3544 0 1 210
box -4 -6 36 206
use NAND2X1  _3391_
timestamp 1596991774
transform 1 0 3544 0 1 210
box -4 -6 52 206
use NOR2X1  _3399_
timestamp 1596991774
transform 1 0 3592 0 1 210
box -4 -6 52 206
use BUFX2  _2115_
timestamp 1596991774
transform -1 0 3768 0 -1 210
box -4 -6 52 206
use INVX1  _3410_
timestamp 1596991774
transform -1 0 3800 0 -1 210
box -4 -6 36 206
use BUFX2  _2114_
timestamp 1596991774
transform -1 0 3848 0 -1 210
box -4 -6 52 206
use OAI21X1  _3400_
timestamp 1596991774
transform 1 0 3640 0 1 210
box -4 -6 68 206
use INVX1  _3390_
timestamp 1596991774
transform -1 0 3736 0 1 210
box -4 -6 36 206
use NOR2X1  _3392_
timestamp 1596991774
transform -1 0 3784 0 1 210
box -4 -6 52 206
use NAND2X1  _3393_
timestamp 1596991774
transform -1 0 3832 0 1 210
box -4 -6 52 206
use OAI21X1  _3389_
timestamp 1596991774
transform 1 0 3848 0 -1 210
box -4 -6 68 206
use INVX1  _3383_
timestamp 1596991774
transform 1 0 3912 0 -1 210
box -4 -6 36 206
use DFFPOSX1  _3420_
timestamp 1596991774
transform -1 0 4136 0 -1 210
box -4 -6 196 206
use AOI21X1  _3411_
timestamp 1596991774
transform 1 0 3832 0 1 210
box -4 -6 68 206
use OAI21X1  _3388_
timestamp 1596991774
transform -1 0 3960 0 1 210
box -4 -6 68 206
use DFFPOSX1  _3421_
timestamp 1596991774
transform -1 0 4152 0 1 210
box -4 -6 196 206
use NOR2X1  _3418_
timestamp 1596991774
transform 1 0 4136 0 -1 210
box -4 -6 52 206
use NOR2X1  _3414_
timestamp 1596991774
transform -1 0 4232 0 -1 210
box -4 -6 52 206
use AOI21X1  _3407_
timestamp 1596991774
transform 1 0 4152 0 1 210
box -4 -6 68 206
use OAI21X1  _3408_
timestamp 1596991774
transform -1 0 4280 0 1 210
box -4 -6 68 206
use INVX1  _3404_
timestamp 1596991774
transform -1 0 4264 0 -1 210
box -4 -6 36 206
use INVX1  _3409_
timestamp 1596991774
transform -1 0 4296 0 -1 210
box -4 -6 36 206
use DFFPOSX1  _3419_
timestamp 1596991774
transform 1 0 4296 0 -1 210
box -4 -6 196 206
use OAI21X1  _3405_
timestamp 1596991774
transform 1 0 4280 0 1 210
box -4 -6 68 206
use INVX1  _3417_
timestamp 1596991774
transform -1 0 4376 0 1 210
box -4 -6 36 206
use OAI21X1  _3416_
timestamp 1596991774
transform 1 0 4376 0 1 210
box -4 -6 68 206
use FILL  SFILL44880x2100
timestamp 1596991774
transform 1 0 4488 0 1 210
box -4 -6 20 206
use FILL  SFILL44720x2100
timestamp 1596991774
transform 1 0 4472 0 1 210
box -4 -6 20 206
use FILL  SFILL44560x2100
timestamp 1596991774
transform 1 0 4456 0 1 210
box -4 -6 20 206
use FILL  SFILL44400x2100
timestamp 1596991774
transform 1 0 4440 0 1 210
box -4 -6 20 206
use FILL  SFILL45040x100
timestamp 1596991774
transform -1 0 4520 0 -1 210
box -4 -6 20 206
use FILL  SFILL44880x100
timestamp 1596991774
transform -1 0 4504 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_insert127
timestamp 1596991774
transform 1 0 4504 0 1 210
box -4 -6 52 206
use FILL  SFILL45360x100
timestamp 1596991774
transform -1 0 4552 0 -1 210
box -4 -6 20 206
use FILL  SFILL45200x100
timestamp 1596991774
transform -1 0 4536 0 -1 210
box -4 -6 20 206
use AOI21X1  _3613_
timestamp 1596991774
transform 1 0 4600 0 1 210
box -4 -6 68 206
use NAND2X1  _3611_
timestamp 1596991774
transform 1 0 4552 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3631_
timestamp 1596991774
transform 1 0 4552 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert191
timestamp 1596991774
transform 1 0 4744 0 -1 210
box -4 -6 52 206
use NAND2X1  _2123_
timestamp 1596991774
transform 1 0 4792 0 -1 210
box -4 -6 52 206
use NAND2X1  _3612_
timestamp 1596991774
transform -1 0 4712 0 1 210
box -4 -6 52 206
use NAND2X1  _3608_
timestamp 1596991774
transform 1 0 4712 0 1 210
box -4 -6 52 206
use AOI21X1  _3610_
timestamp 1596991774
transform -1 0 4824 0 1 210
box -4 -6 68 206
use BUFX2  _2095_
timestamp 1596991774
transform -1 0 4888 0 -1 210
box -4 -6 52 206
use OAI21X1  _2139_
timestamp 1596991774
transform -1 0 4952 0 -1 210
box -4 -6 68 206
use OAI21X1  _2124_
timestamp 1596991774
transform -1 0 5016 0 -1 210
box -4 -6 68 206
use BUFX2  _2090_
timestamp 1596991774
transform 1 0 5016 0 -1 210
box -4 -6 52 206
use NAND2X1  _3609_
timestamp 1596991774
transform -1 0 4872 0 1 210
box -4 -6 52 206
use NAND2X1  _2138_
timestamp 1596991774
transform 1 0 4872 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3630_
timestamp 1596991774
transform 1 0 4920 0 1 210
box -4 -6 196 206
use BUFX2  _2091_
timestamp 1596991774
transform -1 0 5112 0 -1 210
box -4 -6 52 206
use OAI21X1  _2127_
timestamp 1596991774
transform -1 0 5176 0 -1 210
box -4 -6 68 206
use INVX1  _2125_
timestamp 1596991774
transform -1 0 5208 0 -1 210
box -4 -6 36 206
use BUFX2  _2083_
timestamp 1596991774
transform 1 0 5208 0 -1 210
box -4 -6 52 206
use NAND2X1  _2126_
timestamp 1596991774
transform -1 0 5160 0 1 210
box -4 -6 52 206
use NAND2X1  _2120_
timestamp 1596991774
transform 1 0 5160 0 1 210
box -4 -6 52 206
use OAI21X1  _2121_
timestamp 1596991774
transform -1 0 5272 0 1 210
box -4 -6 68 206
use OAI21X1  _2136_
timestamp 1596991774
transform 1 0 5256 0 -1 210
box -4 -6 68 206
use BUFX2  _2094_
timestamp 1596991774
transform 1 0 5320 0 -1 210
box -4 -6 52 206
use BUFX2  _2097_
timestamp 1596991774
transform 1 0 5368 0 -1 210
box -4 -6 52 206
use OAI21X1  _2145_
timestamp 1596991774
transform -1 0 5480 0 -1 210
box -4 -6 68 206
use INVX1  _2122_
timestamp 1596991774
transform -1 0 5304 0 1 210
box -4 -6 36 206
use NAND2X1  _2135_
timestamp 1596991774
transform -1 0 5352 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert192
timestamp 1596991774
transform 1 0 5352 0 1 210
box -4 -6 52 206
use NAND2X1  _2144_
timestamp 1596991774
transform 1 0 5400 0 1 210
box -4 -6 52 206
use OAI21X1  _2133_
timestamp 1596991774
transform 1 0 5480 0 -1 210
box -4 -6 68 206
use BUFX2  _2082_
timestamp 1596991774
transform 1 0 5544 0 -1 210
box -4 -6 52 206
use BUFX2  _2093_
timestamp 1596991774
transform 1 0 5592 0 -1 210
box -4 -6 52 206
use NAND2X1  _2117_
timestamp 1596991774
transform 1 0 5448 0 1 210
box -4 -6 52 206
use NAND2X1  _2132_
timestamp 1596991774
transform 1 0 5496 0 1 210
box -4 -6 52 206
use OAI21X1  _2118_
timestamp 1596991774
transform -1 0 5608 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_insert194
timestamp 1596991774
transform -1 0 5656 0 1 210
box -4 -6 52 206
use INVX1  _2137_
timestamp 1596991774
transform -1 0 5672 0 -1 210
box -4 -6 36 206
use INVX1  _2131_
timestamp 1596991774
transform -1 0 5704 0 -1 210
box -4 -6 36 206
use BUFX2  _2096_
timestamp 1596991774
transform -1 0 5752 0 -1 210
box -4 -6 52 206
use BUFX2  _2092_
timestamp 1596991774
transform -1 0 5800 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _4572_
timestamp 1596991774
transform -1 0 5992 0 -1 210
box -4 -6 196 206
use INVX1  _2116_
timestamp 1596991774
transform -1 0 5688 0 1 210
box -4 -6 36 206
use AOI22X1  _4487_
timestamp 1596991774
transform 1 0 5688 0 1 210
box -4 -6 84 206
use OAI21X1  _2142_
timestamp 1596991774
transform -1 0 5832 0 1 210
box -4 -6 68 206
use AOI22X1  _4514_
timestamp 1596991774
transform 1 0 5832 0 1 210
box -4 -6 84 206
use AOI21X1  _4488_
timestamp 1596991774
transform 1 0 5976 0 1 210
box -4 -6 68 206
use FILL  SFILL59920x100
timestamp 1596991774
transform -1 0 6008 0 -1 210
box -4 -6 20 206
use FILL  SFILL60080x100
timestamp 1596991774
transform -1 0 6024 0 -1 210
box -4 -6 20 206
use FILL  SFILL59120x2100
timestamp 1596991774
transform 1 0 5912 0 1 210
box -4 -6 20 206
use FILL  SFILL59280x2100
timestamp 1596991774
transform 1 0 5928 0 1 210
box -4 -6 20 206
use FILL  SFILL59440x2100
timestamp 1596991774
transform 1 0 5944 0 1 210
box -4 -6 20 206
use FILL  SFILL59600x2100
timestamp 1596991774
transform 1 0 5960 0 1 210
box -4 -6 20 206
use FILL  SFILL60400x100
timestamp 1596991774
transform -1 0 6056 0 -1 210
box -4 -6 20 206
use FILL  SFILL60240x100
timestamp 1596991774
transform -1 0 6040 0 -1 210
box -4 -6 20 206
use NAND3X1  _4486_
timestamp 1596991774
transform 1 0 6120 0 1 210
box -4 -6 68 206
use AOI22X1  _4501_
timestamp 1596991774
transform 1 0 6040 0 1 210
box -4 -6 84 206
use BUFX2  _2086_
timestamp 1596991774
transform 1 0 6104 0 -1 210
box -4 -6 52 206
use BUFX2  _2087_
timestamp 1596991774
transform -1 0 6104 0 -1 210
box -4 -6 52 206
use INVX1  _4485_
timestamp 1596991774
transform -1 0 6248 0 1 210
box -4 -6 36 206
use INVX2  _4482_
timestamp 1596991774
transform -1 0 6216 0 1 210
box -4 -6 36 206
use AOI21X1  _4502_
timestamp 1596991774
transform -1 0 6216 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _4574_
timestamp 1596991774
transform 1 0 6216 0 -1 210
box -4 -6 196 206
use INVX1  _2134_
timestamp 1596991774
transform -1 0 6440 0 -1 210
box -4 -6 36 206
use NOR2X1  _4484_
timestamp 1596991774
transform -1 0 6296 0 1 210
box -4 -6 52 206
use OAI21X1  _4490_
timestamp 1596991774
transform 1 0 6296 0 1 210
box -4 -6 68 206
use NOR3X1  _4498_
timestamp 1596991774
transform 1 0 6360 0 1 210
box -4 -6 132 206
use NAND3X1  _4500_
timestamp 1596991774
transform -1 0 6504 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _4576_
timestamp 1596991774
transform -1 0 6696 0 -1 210
box -4 -6 196 206
use NAND3X1  _4493_
timestamp 1596991774
transform 1 0 6488 0 1 210
box -4 -6 68 206
use OAI21X1  _4497_
timestamp 1596991774
transform 1 0 6552 0 1 210
box -4 -6 68 206
use INVX1  _4496_
timestamp 1596991774
transform 1 0 6616 0 1 210
box -4 -6 36 206
use AOI21X1  _4515_
timestamp 1596991774
transform -1 0 6760 0 -1 210
box -4 -6 68 206
use INVX1  _2143_
timestamp 1596991774
transform -1 0 6792 0 -1 210
box -4 -6 36 206
use INVX1  _4503_
timestamp 1596991774
transform 1 0 6792 0 -1 210
box -4 -6 36 206
use OAI21X1  _4510_
timestamp 1596991774
transform 1 0 6824 0 -1 210
box -4 -6 68 206
use NAND2X1  _4499_
timestamp 1596991774
transform 1 0 6648 0 1 210
box -4 -6 52 206
use NAND3X1  _4505_
timestamp 1596991774
transform 1 0 6696 0 1 210
box -4 -6 68 206
use NAND3X1  _4506_
timestamp 1596991774
transform 1 0 6760 0 1 210
box -4 -6 68 206
use OAI21X1  _4504_
timestamp 1596991774
transform -1 0 6888 0 1 210
box -4 -6 68 206
use NAND3X1  _4513_
timestamp 1596991774
transform 1 0 6888 0 -1 210
box -4 -6 68 206
use INVX2  _4509_
timestamp 1596991774
transform -1 0 6984 0 -1 210
box -4 -6 36 206
use AND2X2  _4525_
timestamp 1596991774
transform -1 0 7048 0 -1 210
box -4 -6 68 206
use NOR3X1  _4518_
timestamp 1596991774
transform 1 0 6888 0 1 210
box -4 -6 132 206
use INVX1  _2140_
timestamp 1596991774
transform -1 0 7048 0 1 210
box -4 -6 36 206
use OAI21X1  _4524_
timestamp 1596991774
transform -1 0 7112 0 -1 210
box -4 -6 68 206
use INVX1  _4516_
timestamp 1596991774
transform 1 0 7112 0 -1 210
box -4 -6 36 206
use INVX1  _4512_
timestamp 1596991774
transform -1 0 7176 0 -1 210
box -4 -6 36 206
use DFFPOSX1  _4578_
timestamp 1596991774
transform 1 0 7176 0 -1 210
box -4 -6 196 206
use NAND3X1  _4519_
timestamp 1596991774
transform 1 0 7048 0 1 210
box -4 -6 68 206
use OAI21X1  _4526_
timestamp 1596991774
transform 1 0 7112 0 1 210
box -4 -6 68 206
use AOI21X1  _4528_
timestamp 1596991774
transform 1 0 7176 0 1 210
box -4 -6 68 206
use NOR3X1  _4529_
timestamp 1596991774
transform 1 0 7240 0 1 210
box -4 -6 132 206
use FILL  FILL71120x100
timestamp 1596991774
transform -1 0 7384 0 -1 210
box -4 -6 20 206
use FILL  FILL71280x100
timestamp 1596991774
transform -1 0 7400 0 -1 210
box -4 -6 20 206
use FILL  FILL71120x2100
timestamp 1596991774
transform 1 0 7368 0 1 210
box -4 -6 20 206
use FILL  FILL71280x2100
timestamp 1596991774
transform 1 0 7384 0 1 210
box -4 -6 20 206
use XNOR2X1  _2484_
timestamp 1596991774
transform -1 0 120 0 -1 610
box -4 -6 116 206
use AOI21X1  _2493_
timestamp 1596991774
transform -1 0 184 0 -1 610
box -4 -6 68 206
use XNOR2X1  _2485_
timestamp 1596991774
transform -1 0 296 0 -1 610
box -4 -6 116 206
use NOR2X1  _2483_
timestamp 1596991774
transform 1 0 296 0 -1 610
box -4 -6 52 206
use AOI21X1  _2495_
timestamp 1596991774
transform -1 0 408 0 -1 610
box -4 -6 68 206
use XNOR2X1  _2486_
timestamp 1596991774
transform -1 0 520 0 -1 610
box -4 -6 116 206
use BUFX2  BUFX2_insert35
timestamp 1596991774
transform -1 0 568 0 -1 610
box -4 -6 52 206
use INVX1  _3152_
timestamp 1596991774
transform 1 0 568 0 -1 610
box -4 -6 36 206
use INVX1  _2889_
timestamp 1596991774
transform 1 0 600 0 -1 610
box -4 -6 36 206
use AOI22X1  _2890_
timestamp 1596991774
transform -1 0 712 0 -1 610
box -4 -6 84 206
use INVX1  _2888_
timestamp 1596991774
transform -1 0 744 0 -1 610
box -4 -6 36 206
use INVX1  _3123_
timestamp 1596991774
transform 1 0 744 0 -1 610
box -4 -6 36 206
use OAI22X1  _3154_
timestamp 1596991774
transform 1 0 776 0 -1 610
box -4 -6 84 206
use INVX1  _3153_
timestamp 1596991774
transform -1 0 888 0 -1 610
box -4 -6 36 206
use OAI22X1  _3125_
timestamp 1596991774
transform 1 0 888 0 -1 610
box -4 -6 84 206
use INVX1  _3124_
timestamp 1596991774
transform -1 0 1000 0 -1 610
box -4 -6 36 206
use NOR2X1  _3129_
timestamp 1596991774
transform -1 0 1048 0 -1 610
box -4 -6 52 206
use NOR2X1  _3136_
timestamp 1596991774
transform 1 0 1048 0 -1 610
box -4 -6 52 206
use OR2X2  _2345_
timestamp 1596991774
transform -1 0 1160 0 -1 610
box -4 -6 68 206
use INVX1  _3133_
timestamp 1596991774
transform 1 0 1160 0 -1 610
box -4 -6 36 206
use OAI21X1  _3135_
timestamp 1596991774
transform 1 0 1192 0 -1 610
box -4 -6 68 206
use NAND2X1  _3134_
timestamp 1596991774
transform 1 0 1256 0 -1 610
box -4 -6 52 206
use INVX1  _2702_
timestamp 1596991774
transform 1 0 1304 0 -1 610
box -4 -6 36 206
use NAND2X1  _2703_
timestamp 1596991774
transform 1 0 1336 0 -1 610
box -4 -6 52 206
use FILL  SFILL13840x4100
timestamp 1596991774
transform -1 0 1400 0 -1 610
box -4 -6 20 206
use FILL  SFILL14000x4100
timestamp 1596991774
transform -1 0 1416 0 -1 610
box -4 -6 20 206
use OAI22X1  _2724_
timestamp 1596991774
transform -1 0 1528 0 -1 610
box -4 -6 84 206
use NAND2X1  _2701_
timestamp 1596991774
transform 1 0 1528 0 -1 610
box -4 -6 52 206
use INVX1  _2700_
timestamp 1596991774
transform -1 0 1608 0 -1 610
box -4 -6 36 206
use OR2X2  _2346_
timestamp 1596991774
transform 1 0 1608 0 -1 610
box -4 -6 68 206
use FILL  SFILL14160x4100
timestamp 1596991774
transform -1 0 1432 0 -1 610
box -4 -6 20 206
use FILL  SFILL14320x4100
timestamp 1596991774
transform -1 0 1448 0 -1 610
box -4 -6 20 206
use INVX1  _3097_
timestamp 1596991774
transform 1 0 1672 0 -1 610
box -4 -6 36 206
use NAND2X1  _3004_
timestamp 1596991774
transform -1 0 1752 0 -1 610
box -4 -6 52 206
use NAND2X1  _3290_
timestamp 1596991774
transform 1 0 1752 0 -1 610
box -4 -6 52 206
use INVX1  _3055_
timestamp 1596991774
transform 1 0 1800 0 -1 610
box -4 -6 36 206
use OAI21X1  _3057_
timestamp 1596991774
transform 1 0 1832 0 -1 610
box -4 -6 68 206
use INVX1  _3053_
timestamp 1596991774
transform 1 0 1896 0 -1 610
box -4 -6 36 206
use OAI22X1  _3054_
timestamp 1596991774
transform -1 0 2008 0 -1 610
box -4 -6 84 206
use INVX1  _3052_
timestamp 1596991774
transform 1 0 2008 0 -1 610
box -4 -6 36 206
use NOR2X1  _3058_
timestamp 1596991774
transform 1 0 2040 0 -1 610
box -4 -6 52 206
use NOR2X1  _3051_
timestamp 1596991774
transform 1 0 2088 0 -1 610
box -4 -6 52 206
use OAI22X1  _3047_
timestamp 1596991774
transform 1 0 2136 0 -1 610
box -4 -6 84 206
use INVX1  _3046_
timestamp 1596991774
transform -1 0 2248 0 -1 610
box -4 -6 36 206
use INVX1  _3049_
timestamp 1596991774
transform 1 0 2248 0 -1 610
box -4 -6 36 206
use OAI22X1  _3050_
timestamp 1596991774
transform -1 0 2360 0 -1 610
box -4 -6 84 206
use INVX1  _3045_
timestamp 1596991774
transform -1 0 2392 0 -1 610
box -4 -6 36 206
use OR2X2  _2344_
timestamp 1596991774
transform -1 0 2456 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert258
timestamp 1596991774
transform -1 0 2504 0 -1 610
box -4 -6 52 206
use INVX1  _2706_
timestamp 1596991774
transform 1 0 2504 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert257
timestamp 1596991774
transform 1 0 2536 0 -1 610
box -4 -6 52 206
use AOI22X1  _2708_
timestamp 1596991774
transform 1 0 2584 0 -1 610
box -4 -6 84 206
use INVX1  _2707_
timestamp 1596991774
transform -1 0 2696 0 -1 610
box -4 -6 36 206
use NOR2X1  _2721_
timestamp 1596991774
transform -1 0 2744 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert80
timestamp 1596991774
transform -1 0 2792 0 -1 610
box -4 -6 52 206
use AOI22X1  _2902_
timestamp 1596991774
transform -1 0 2872 0 -1 610
box -4 -6 84 206
use INVX1  _2901_
timestamp 1596991774
transform -1 0 2904 0 -1 610
box -4 -6 36 206
use NOR2X1  _2911_
timestamp 1596991774
transform -1 0 3016 0 -1 610
box -4 -6 52 206
use FILL  SFILL29040x4100
timestamp 1596991774
transform -1 0 2920 0 -1 610
box -4 -6 20 206
use FILL  SFILL29200x4100
timestamp 1596991774
transform -1 0 2936 0 -1 610
box -4 -6 20 206
use FILL  SFILL29360x4100
timestamp 1596991774
transform -1 0 2952 0 -1 610
box -4 -6 20 206
use FILL  SFILL29520x4100
timestamp 1596991774
transform -1 0 2968 0 -1 610
box -4 -6 20 206
use NAND2X1  _2903_
timestamp 1596991774
transform 1 0 3016 0 -1 610
box -4 -6 52 206
use AOI21X1  _2913_
timestamp 1596991774
transform 1 0 3064 0 -1 610
box -4 -6 68 206
use NAND2X1  _2912_
timestamp 1596991774
transform -1 0 3176 0 -1 610
box -4 -6 52 206
use NOR2X1  _2910_
timestamp 1596991774
transform -1 0 3224 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert84
timestamp 1596991774
transform -1 0 3272 0 -1 610
box -4 -6 52 206
use NOR2X1  _2628_
timestamp 1596991774
transform 1 0 3272 0 -1 610
box -4 -6 52 206
use NAND2X1  _2630_
timestamp 1596991774
transform 1 0 3320 0 -1 610
box -4 -6 52 206
use INVX1  _3394_
timestamp 1596991774
transform 1 0 3368 0 -1 610
box -4 -6 36 206
use INVX1  _2615_
timestamp 1596991774
transform 1 0 3400 0 -1 610
box -4 -6 36 206
use NAND2X1  _3397_
timestamp 1596991774
transform 1 0 3432 0 -1 610
box -4 -6 52 206
use NOR2X1  _3385_
timestamp 1596991774
transform 1 0 3480 0 -1 610
box -4 -6 52 206
use AOI22X1  _3398_
timestamp 1596991774
transform 1 0 3528 0 -1 610
box -4 -6 84 206
use NAND3X1  _3406_
timestamp 1596991774
transform 1 0 3608 0 -1 610
box -4 -6 68 206
use INVX1  _3386_
timestamp 1596991774
transform 1 0 3672 0 -1 610
box -4 -6 36 206
use NOR2X1  _3387_
timestamp 1596991774
transform 1 0 3704 0 -1 610
box -4 -6 52 206
use AOI21X1  _3598_
timestamp 1596991774
transform -1 0 3816 0 -1 610
box -4 -6 68 206
use NAND2X1  _3596_
timestamp 1596991774
transform -1 0 3864 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _3641_
timestamp 1596991774
transform -1 0 4056 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _3422_
timestamp 1596991774
transform 1 0 4056 0 -1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert128
timestamp 1596991774
transform -1 0 4296 0 -1 610
box -4 -6 52 206
use AND2X2  _3415_
timestamp 1596991774
transform 1 0 4296 0 -1 610
box -4 -6 68 206
use FILL  SFILL43600x4100
timestamp 1596991774
transform -1 0 4376 0 -1 610
box -4 -6 20 206
use FILL  SFILL43760x4100
timestamp 1596991774
transform -1 0 4392 0 -1 610
box -4 -6 20 206
use FILL  SFILL43920x4100
timestamp 1596991774
transform -1 0 4408 0 -1 610
box -4 -6 20 206
use FILL  SFILL44080x4100
timestamp 1596991774
transform -1 0 4424 0 -1 610
box -4 -6 20 206
use DFFPOSX1  _3634_
timestamp 1596991774
transform 1 0 4424 0 -1 610
box -4 -6 196 206
use NAND2X1  _3576_
timestamp 1596991774
transform -1 0 4664 0 -1 610
box -4 -6 52 206
use NAND2X1  _3573_
timestamp 1596991774
transform 1 0 4664 0 -1 610
box -4 -6 52 206
use NAND2X1  _3626_
timestamp 1596991774
transform 1 0 4712 0 -1 610
box -4 -6 52 206
use AOI21X1  _3628_
timestamp 1596991774
transform 1 0 4760 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _3629_
timestamp 1596991774
transform 1 0 4824 0 -1 610
box -4 -6 196 206
use INVX1  _3543_
timestamp 1596991774
transform 1 0 5016 0 -1 610
box -4 -6 36 206
use NOR2X1  _3544_
timestamp 1596991774
transform -1 0 5096 0 -1 610
box -4 -6 52 206
use NAND2X1  _4595_
timestamp 1596991774
transform 1 0 5096 0 -1 610
box -4 -6 52 206
use OAI21X1  _4596_
timestamp 1596991774
transform -1 0 5208 0 -1 610
box -4 -6 68 206
use INVX1  _4594_
timestamp 1596991774
transform -1 0 5240 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert170
timestamp 1596991774
transform -1 0 5288 0 -1 610
box -4 -6 52 206
use AND2X2  _3559_
timestamp 1596991774
transform 1 0 5288 0 -1 610
box -4 -6 68 206
use INVX1  _4609_
timestamp 1596991774
transform 1 0 5352 0 -1 610
box -4 -6 36 206
use INVX1  _2119_
timestamp 1596991774
transform -1 0 5416 0 -1 610
box -4 -6 36 206
use NAND2X1  _4586_
timestamp 1596991774
transform 1 0 5416 0 -1 610
box -4 -6 52 206
use INVX1  _4585_
timestamp 1596991774
transform 1 0 5464 0 -1 610
box -4 -6 36 206
use OAI21X1  _4587_
timestamp 1596991774
transform -1 0 5560 0 -1 610
box -4 -6 68 206
use OAI21X1  _4611_
timestamp 1596991774
transform 1 0 5560 0 -1 610
box -4 -6 68 206
use NAND3X1  _4478_
timestamp 1596991774
transform -1 0 5688 0 -1 610
box -4 -6 68 206
use AOI22X1  _4468_
timestamp 1596991774
transform 1 0 5688 0 -1 610
box -4 -6 84 206
use INVX1  _4470_
timestamp 1596991774
transform 1 0 5768 0 -1 610
box -4 -6 36 206
use INVX1  _4476_
timestamp 1596991774
transform 1 0 5800 0 -1 610
box -4 -6 36 206
use OAI21X1  _4477_
timestamp 1596991774
transform -1 0 5896 0 -1 610
box -4 -6 68 206
use INVX1  _4461_
timestamp 1596991774
transform 1 0 5896 0 -1 610
box -4 -6 36 206
use NAND3X1  _4479_
timestamp 1596991774
transform -1 0 6056 0 -1 610
box -4 -6 68 206
use FILL  SFILL59280x4100
timestamp 1596991774
transform -1 0 5944 0 -1 610
box -4 -6 20 206
use FILL  SFILL59440x4100
timestamp 1596991774
transform -1 0 5960 0 -1 610
box -4 -6 20 206
use FILL  SFILL59600x4100
timestamp 1596991774
transform -1 0 5976 0 -1 610
box -4 -6 20 206
use FILL  SFILL59760x4100
timestamp 1596991774
transform -1 0 5992 0 -1 610
box -4 -6 20 206
use NAND2X1  _4471_
timestamp 1596991774
transform -1 0 6104 0 -1 610
box -4 -6 52 206
use OAI21X1  _4483_
timestamp 1596991774
transform 1 0 6104 0 -1 610
box -4 -6 68 206
use NAND2X1  _4464_
timestamp 1596991774
transform -1 0 6216 0 -1 610
box -4 -6 52 206
use AOI21X1  _4469_
timestamp 1596991774
transform 1 0 6216 0 -1 610
box -4 -6 68 206
use INVX1  _4491_
timestamp 1596991774
transform 1 0 6280 0 -1 610
box -4 -6 36 206
use NAND3X1  _4492_
timestamp 1596991774
transform 1 0 6312 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4569_
timestamp 1596991774
transform -1 0 6568 0 -1 610
box -4 -6 196 206
use INVX1  _4489_
timestamp 1596991774
transform -1 0 6600 0 -1 610
box -4 -6 36 206
use AOI22X1  _4507_
timestamp 1596991774
transform 1 0 6600 0 -1 610
box -4 -6 84 206
use AOI21X1  _4508_
timestamp 1596991774
transform -1 0 6744 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4575_
timestamp 1596991774
transform -1 0 6936 0 -1 610
box -4 -6 196 206
use AOI22X1  _4521_
timestamp 1596991774
transform 1 0 6936 0 -1 610
box -4 -6 84 206
use INVX2  _4523_
timestamp 1596991774
transform 1 0 7016 0 -1 610
box -4 -6 36 206
use AOI21X1  _4522_
timestamp 1596991774
transform -1 0 7112 0 -1 610
box -4 -6 68 206
use NAND3X1  _4520_
timestamp 1596991774
transform 1 0 7112 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4577_
timestamp 1596991774
transform -1 0 7368 0 -1 610
box -4 -6 196 206
use FILL  FILL71120x4100
timestamp 1596991774
transform -1 0 7384 0 -1 610
box -4 -6 20 206
use FILL  FILL71280x4100
timestamp 1596991774
transform -1 0 7400 0 -1 610
box -4 -6 20 206
use XOR2X1  _2538_
timestamp 1596991774
transform -1 0 120 0 1 610
box -4 -6 116 206
use NOR2X1  _2492_
timestamp 1596991774
transform 1 0 120 0 1 610
box -4 -6 52 206
use INVX1  _2491_
timestamp 1596991774
transform -1 0 200 0 1 610
box -4 -6 36 206
use INVX1  _2479_
timestamp 1596991774
transform 1 0 200 0 1 610
box -4 -6 36 206
use NOR2X1  _2480_
timestamp 1596991774
transform -1 0 280 0 1 610
box -4 -6 52 206
use OAI21X1  _2916_
timestamp 1596991774
transform -1 0 344 0 1 610
box -4 -6 68 206
use INVX1  _2891_
timestamp 1596991774
transform -1 0 376 0 1 610
box -4 -6 36 206
use OAI22X1  _2915_
timestamp 1596991774
transform 1 0 376 0 1 610
box -4 -6 84 206
use NAND2X1  _2892_
timestamp 1596991774
transform -1 0 504 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert177
timestamp 1596991774
transform -1 0 552 0 1 610
box -4 -6 52 206
use INVX1  _2893_
timestamp 1596991774
transform 1 0 552 0 1 610
box -4 -6 36 206
use NAND2X1  _2894_
timestamp 1596991774
transform -1 0 632 0 1 610
box -4 -6 52 206
use NAND3X1  _2895_
timestamp 1596991774
transform 1 0 632 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert286
timestamp 1596991774
transform -1 0 744 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert181
timestamp 1596991774
transform 1 0 744 0 1 610
box -4 -6 52 206
use NOR2X1  _3155_
timestamp 1596991774
transform 1 0 792 0 1 610
box -4 -6 52 206
use INVX1  _3150_
timestamp 1596991774
transform 1 0 840 0 1 610
box -4 -6 36 206
use OAI22X1  _3151_
timestamp 1596991774
transform -1 0 952 0 1 610
box -4 -6 84 206
use INVX1  _3130_
timestamp 1596991774
transform 1 0 952 0 1 610
box -4 -6 36 206
use OAI22X1  _3132_
timestamp 1596991774
transform 1 0 984 0 1 610
box -4 -6 84 206
use INVX1  _3131_
timestamp 1596991774
transform -1 0 1096 0 1 610
box -4 -6 36 206
use NAND3X1  _3148_
timestamp 1596991774
transform 1 0 1096 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert289
timestamp 1596991774
transform 1 0 1160 0 1 610
box -4 -6 52 206
use INVX1  _2698_
timestamp 1596991774
transform 1 0 1208 0 1 610
box -4 -6 36 206
use AOI22X1  _2699_
timestamp 1596991774
transform -1 0 1320 0 1 610
box -4 -6 84 206
use INVX1  _2697_
timestamp 1596991774
transform -1 0 1352 0 1 610
box -4 -6 36 206
use OAI21X1  _2725_
timestamp 1596991774
transform 1 0 1352 0 1 610
box -4 -6 68 206
use NAND3X1  _2704_
timestamp 1596991774
transform -1 0 1544 0 1 610
box -4 -6 68 206
use INVX1  _3467_
timestamp 1596991774
transform 1 0 1544 0 1 610
box -4 -6 36 206
use INVX1  _3460_
timestamp 1596991774
transform 1 0 1576 0 1 610
box -4 -6 36 206
use INVX1  _3003_
timestamp 1596991774
transform 1 0 1608 0 1 610
box -4 -6 36 206
use FILL  SFILL14160x6100
timestamp 1596991774
transform 1 0 1416 0 1 610
box -4 -6 20 206
use FILL  SFILL14320x6100
timestamp 1596991774
transform 1 0 1432 0 1 610
box -4 -6 20 206
use FILL  SFILL14480x6100
timestamp 1596991774
transform 1 0 1448 0 1 610
box -4 -6 20 206
use FILL  SFILL14640x6100
timestamp 1596991774
transform 1 0 1464 0 1 610
box -4 -6 20 206
use OAI21X1  _3005_
timestamp 1596991774
transform 1 0 1640 0 1 610
box -4 -6 68 206
use INVX1  _3289_
timestamp 1596991774
transform 1 0 1704 0 1 610
box -4 -6 36 206
use OAI21X1  _3291_
timestamp 1596991774
transform 1 0 1736 0 1 610
box -4 -6 68 206
use INVX1  _3000_
timestamp 1596991774
transform 1 0 1800 0 1 610
box -4 -6 36 206
use OAI22X1  _3002_
timestamp 1596991774
transform 1 0 1832 0 1 610
box -4 -6 84 206
use INVX1  _3001_
timestamp 1596991774
transform -1 0 1944 0 1 610
box -4 -6 36 206
use INVX1  _3287_
timestamp 1596991774
transform -1 0 1976 0 1 610
box -4 -6 36 206
use NOR2X1  _3006_
timestamp 1596991774
transform -1 0 2024 0 1 610
box -4 -6 52 206
use NOR2X1  _2304_
timestamp 1596991774
transform 1 0 2024 0 1 610
box -4 -6 52 206
use NAND3X1  _3070_
timestamp 1596991774
transform -1 0 2136 0 1 610
box -4 -6 68 206
use AND2X2  _2303_
timestamp 1596991774
transform -1 0 2200 0 1 610
box -4 -6 68 206
use NOR2X1  _2302_
timestamp 1596991774
transform -1 0 2248 0 1 610
box -4 -6 52 206
use INVX1  _2801_
timestamp 1596991774
transform 1 0 2248 0 1 610
box -4 -6 36 206
use NOR2X1  _2807_
timestamp 1596991774
transform 1 0 2280 0 1 610
box -4 -6 52 206
use NAND2X1  _2805_
timestamp 1596991774
transform -1 0 2376 0 1 610
box -4 -6 52 206
use OAI22X1  _2803_
timestamp 1596991774
transform 1 0 2376 0 1 610
box -4 -6 84 206
use NOR2X1  _2804_
timestamp 1596991774
transform -1 0 2504 0 1 610
box -4 -6 52 206
use INVX1  _2798_
timestamp 1596991774
transform 1 0 2504 0 1 610
box -4 -6 36 206
use OAI22X1  _2800_
timestamp 1596991774
transform 1 0 2536 0 1 610
box -4 -6 84 206
use INVX1  _2709_
timestamp 1596991774
transform 1 0 2616 0 1 610
box -4 -6 36 206
use INVX1  _2802_
timestamp 1596991774
transform -1 0 2680 0 1 610
box -4 -6 36 206
use NAND3X1  _2758_
timestamp 1596991774
transform 1 0 2680 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert56
timestamp 1596991774
transform -1 0 2792 0 1 610
box -4 -6 52 206
use NAND2X1  _2712_
timestamp 1596991774
transform 1 0 2792 0 1 610
box -4 -6 52 206
use NOR2X1  _2719_
timestamp 1596991774
transform 1 0 2840 0 1 610
box -4 -6 52 206
use AOI21X1  _2722_
timestamp 1596991774
transform -1 0 2952 0 1 610
box -4 -6 68 206
use FILL  SFILL29520x6100
timestamp 1596991774
transform 1 0 2952 0 1 610
box -4 -6 20 206
use FILL  SFILL29680x6100
timestamp 1596991774
transform 1 0 2968 0 1 610
box -4 -6 20 206
use FILL  SFILL29840x6100
timestamp 1596991774
transform 1 0 2984 0 1 610
box -4 -6 20 206
use FILL  SFILL30000x6100
timestamp 1596991774
transform 1 0 3000 0 1 610
box -4 -6 20 206
use NAND2X1  _2720_
timestamp 1596991774
transform -1 0 3064 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert82
timestamp 1596991774
transform -1 0 3112 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert183
timestamp 1596991774
transform -1 0 3160 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert185
timestamp 1596991774
transform -1 0 3208 0 1 610
box -4 -6 52 206
use AOI22X1  _2711_
timestamp 1596991774
transform 1 0 3208 0 1 610
box -4 -6 84 206
use INVX1  _2710_
timestamp 1596991774
transform -1 0 3320 0 1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert83
timestamp 1596991774
transform -1 0 3368 0 1 610
box -4 -6 52 206
use OAI21X1  _2631_
timestamp 1596991774
transform -1 0 3432 0 1 610
box -4 -6 68 206
use NOR2X1  _2629_
timestamp 1596991774
transform -1 0 3480 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert53
timestamp 1596991774
transform -1 0 3528 0 1 610
box -4 -6 52 206
use INVX1  _3446_
timestamp 1596991774
transform 1 0 3528 0 1 610
box -4 -6 36 206
use INVX1  _3395_
timestamp 1596991774
transform 1 0 3560 0 1 610
box -4 -6 36 206
use NOR2X1  _3396_
timestamp 1596991774
transform -1 0 3640 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert182
timestamp 1596991774
transform 1 0 3640 0 1 610
box -4 -6 52 206
use DFFPOSX1  _3639_
timestamp 1596991774
transform -1 0 3880 0 1 610
box -4 -6 196 206
use NAND2X1  _3597_
timestamp 1596991774
transform 1 0 3880 0 1 610
box -4 -6 52 206
use AOI21X1  _3601_
timestamp 1596991774
transform -1 0 3992 0 1 610
box -4 -6 68 206
use NAND2X1  _3600_
timestamp 1596991774
transform -1 0 4040 0 1 610
box -4 -6 52 206
use NAND2X1  _3599_
timestamp 1596991774
transform -1 0 4088 0 1 610
box -4 -6 52 206
use NAND2X1  _3602_
timestamp 1596991774
transform -1 0 4136 0 1 610
box -4 -6 52 206
use NAND2X1  _3606_
timestamp 1596991774
transform 1 0 4136 0 1 610
box -4 -6 52 206
use AOI21X1  _3607_
timestamp 1596991774
transform -1 0 4248 0 1 610
box -4 -6 68 206
use NAND2X1  _3605_
timestamp 1596991774
transform -1 0 4296 0 1 610
box -4 -6 52 206
use DFFPOSX1  _3423_
timestamp 1596991774
transform 1 0 4296 0 1 610
box -4 -6 196 206
use AOI21X1  _3619_
timestamp 1596991774
transform -1 0 4616 0 1 610
box -4 -6 68 206
use INVX1  _3441_
timestamp 1596991774
transform 1 0 4616 0 1 610
box -4 -6 36 206
use FILL  SFILL44880x6100
timestamp 1596991774
transform 1 0 4488 0 1 610
box -4 -6 20 206
use FILL  SFILL45040x6100
timestamp 1596991774
transform 1 0 4504 0 1 610
box -4 -6 20 206
use FILL  SFILL45200x6100
timestamp 1596991774
transform 1 0 4520 0 1 610
box -4 -6 20 206
use FILL  SFILL45360x6100
timestamp 1596991774
transform 1 0 4536 0 1 610
box -4 -6 20 206
use INVX1  _3462_
timestamp 1596991774
transform 1 0 4648 0 1 610
box -4 -6 36 206
use NAND3X1  _3463_
timestamp 1596991774
transform 1 0 4680 0 1 610
box -4 -6 68 206
use INVX1  _3455_
timestamp 1596991774
transform 1 0 4744 0 1 610
box -4 -6 36 206
use NAND3X1  _3456_
timestamp 1596991774
transform 1 0 4776 0 1 610
box -4 -6 68 206
use NAND2X1  _3618_
timestamp 1596991774
transform -1 0 4888 0 1 610
box -4 -6 52 206
use NAND2X1  _3627_
timestamp 1596991774
transform -1 0 4936 0 1 610
box -4 -6 52 206
use AOI21X1  _3617_
timestamp 1596991774
transform -1 0 5000 0 1 610
box -4 -6 68 206
use NAND2X1  _3616_
timestamp 1596991774
transform -1 0 5048 0 1 610
box -4 -6 52 206
use DFFPOSX1  _3633_
timestamp 1596991774
transform 1 0 5048 0 1 610
box -4 -6 196 206
use INVX1  _3545_
timestamp 1596991774
transform -1 0 5272 0 1 610
box -4 -6 36 206
use AND2X2  _3560_
timestamp 1596991774
transform 1 0 5272 0 1 610
box -4 -6 68 206
use INVX1  _3549_
timestamp 1596991774
transform 1 0 5336 0 1 610
box -4 -6 36 206
use NOR2X1  _3550_
timestamp 1596991774
transform -1 0 5416 0 1 610
box -4 -6 52 206
use INVX1  _4612_
timestamp 1596991774
transform 1 0 5416 0 1 610
box -4 -6 36 206
use NAND2X1  _4613_
timestamp 1596991774
transform -1 0 5496 0 1 610
box -4 -6 52 206
use OAI21X1  _4614_
timestamp 1596991774
transform 1 0 5496 0 1 610
box -4 -6 68 206
use NAND2X1  _4604_
timestamp 1596991774
transform -1 0 5608 0 1 610
box -4 -6 52 206
use NAND2X1  _4610_
timestamp 1596991774
transform 1 0 5608 0 1 610
box -4 -6 52 206
use OAI21X1  _4605_
timestamp 1596991774
transform 1 0 5656 0 1 610
box -4 -6 68 206
use NAND2X1  _2141_
timestamp 1596991774
transform 1 0 5720 0 1 610
box -4 -6 52 206
use NAND2X1  _4592_
timestamp 1596991774
transform -1 0 5816 0 1 610
box -4 -6 52 206
use OAI21X1  _2130_
timestamp 1596991774
transform -1 0 5880 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert176
timestamp 1596991774
transform -1 0 5928 0 1 610
box -4 -6 52 206
use AOI21X1  _4481_
timestamp 1596991774
transform -1 0 6056 0 1 610
box -4 -6 68 206
use FILL  SFILL59280x6100
timestamp 1596991774
transform 1 0 5928 0 1 610
box -4 -6 20 206
use FILL  SFILL59440x6100
timestamp 1596991774
transform 1 0 5944 0 1 610
box -4 -6 20 206
use FILL  SFILL59600x6100
timestamp 1596991774
transform 1 0 5960 0 1 610
box -4 -6 20 206
use FILL  SFILL59760x6100
timestamp 1596991774
transform 1 0 5976 0 1 610
box -4 -6 20 206
use NAND3X1  _4473_
timestamp 1596991774
transform -1 0 6120 0 1 610
box -4 -6 68 206
use NAND2X1  _4472_
timestamp 1596991774
transform -1 0 6168 0 1 610
box -4 -6 52 206
use DFFPOSX1  _4571_
timestamp 1596991774
transform -1 0 6360 0 1 610
box -4 -6 196 206
use INVX1  _2128_
timestamp 1596991774
transform -1 0 6392 0 1 610
box -4 -6 36 206
use BUFX2  _2089_
timestamp 1596991774
transform 1 0 6392 0 1 610
box -4 -6 52 206
use AOI22X1  _4494_
timestamp 1596991774
transform 1 0 6440 0 1 610
box -4 -6 84 206
use AOI21X1  _4495_
timestamp 1596991774
transform 1 0 6520 0 1 610
box -4 -6 68 206
use DFFPOSX1  _4573_
timestamp 1596991774
transform -1 0 6776 0 1 610
box -4 -6 196 206
use NOR2X1  _4466_
timestamp 1596991774
transform 1 0 6776 0 1 610
box -4 -6 52 206
use INVX1  _4462_
timestamp 1596991774
transform 1 0 6824 0 1 610
box -4 -6 36 206
use INVX1  _4465_
timestamp 1596991774
transform -1 0 6888 0 1 610
box -4 -6 36 206
use NOR2X1  _4467_
timestamp 1596991774
transform -1 0 6936 0 1 610
box -4 -6 52 206
use NOR2X1  _4463_
timestamp 1596991774
transform -1 0 6984 0 1 610
box -4 -6 52 206
use AOI22X1  _4527_
timestamp 1596991774
transform 1 0 6984 0 1 610
box -4 -6 84 206
use NOR3X1  _4538_
timestamp 1596991774
transform 1 0 7064 0 1 610
box -4 -6 132 206
use NAND3X1  _4533_
timestamp 1596991774
transform 1 0 7192 0 1 610
box -4 -6 68 206
use OAI21X1  _4532_
timestamp 1596991774
transform 1 0 7256 0 1 610
box -4 -6 68 206
use INVX1  _4531_
timestamp 1596991774
transform -1 0 7352 0 1 610
box -4 -6 36 206
use INVX1  _4536_
timestamp 1596991774
transform -1 0 7384 0 1 610
box -4 -6 36 206
use FILL  FILL71280x6100
timestamp 1596991774
transform 1 0 7384 0 1 610
box -4 -6 20 206
use BUFX2  _2111_
timestamp 1596991774
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use INVX1  _2885_
timestamp 1596991774
transform 1 0 56 0 -1 1010
box -4 -6 36 206
use NOR2X1  _2918_
timestamp 1596991774
transform -1 0 136 0 -1 1010
box -4 -6 52 206
use AOI21X1  _2920_
timestamp 1596991774
transform 1 0 136 0 -1 1010
box -4 -6 68 206
use NOR2X1  _2917_
timestamp 1596991774
transform 1 0 200 0 -1 1010
box -4 -6 52 206
use AOI22X1  _2886_
timestamp 1596991774
transform 1 0 248 0 -1 1010
box -4 -6 84 206
use BUFX2  BUFX2_insert71
timestamp 1596991774
transform -1 0 376 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2887_
timestamp 1596991774
transform -1 0 424 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert68
timestamp 1596991774
transform 1 0 424 0 -1 1010
box -4 -6 52 206
use INVX1  _2813_
timestamp 1596991774
transform -1 0 504 0 -1 1010
box -4 -6 36 206
use INVX1  _2882_
timestamp 1596991774
transform 1 0 504 0 -1 1010
box -4 -6 36 206
use AOI22X1  _2883_
timestamp 1596991774
transform -1 0 616 0 -1 1010
box -4 -6 84 206
use INVX1  _2881_
timestamp 1596991774
transform -1 0 648 0 -1 1010
box -4 -6 36 206
use NOR2X1  _2896_
timestamp 1596991774
transform 1 0 648 0 -1 1010
box -4 -6 52 206
use OR2X2  _2347_
timestamp 1596991774
transform 1 0 696 0 -1 1010
box -4 -6 68 206
use INVX1  _2599_
timestamp 1596991774
transform 1 0 760 0 -1 1010
box -4 -6 36 206
use AOI22X1  _2601_
timestamp 1596991774
transform -1 0 872 0 -1 1010
box -4 -6 84 206
use INVX1  _2600_
timestamp 1596991774
transform 1 0 872 0 -1 1010
box -4 -6 36 206
use NOR2X1  _2821_
timestamp 1596991774
transform 1 0 904 0 -1 1010
box -4 -6 52 206
use INVX1  _2817_
timestamp 1596991774
transform -1 0 984 0 -1 1010
box -4 -6 36 206
use INVX1  _3149_
timestamp 1596991774
transform -1 0 1016 0 -1 1010
box -4 -6 36 206
use AOI21X1  _2822_
timestamp 1596991774
transform -1 0 1080 0 -1 1010
box -4 -6 68 206
use INVX1  _2820_
timestamp 1596991774
transform -1 0 1112 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert157
timestamp 1596991774
transform -1 0 1160 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert156
timestamp 1596991774
transform 1 0 1160 0 -1 1010
box -4 -6 52 206
use INVX1  _2597_
timestamp 1596991774
transform 1 0 1208 0 -1 1010
box -4 -6 36 206
use AOI22X1  _2598_
timestamp 1596991774
transform -1 0 1320 0 -1 1010
box -4 -6 84 206
use NOR2X1  _2633_
timestamp 1596991774
transform 1 0 1320 0 -1 1010
box -4 -6 52 206
use INVX1  _2596_
timestamp 1596991774
transform -1 0 1400 0 -1 1010
box -4 -6 36 206
use FILL  SFILL14000x8100
timestamp 1596991774
transform -1 0 1416 0 -1 1010
box -4 -6 20 206
use NAND2X1  _2602_
timestamp 1596991774
transform -1 0 1512 0 -1 1010
box -4 -6 52 206
use OAI22X1  _2636_
timestamp 1596991774
transform 1 0 1512 0 -1 1010
box -4 -6 84 206
use NOR2X1  _2610_
timestamp 1596991774
transform 1 0 1592 0 -1 1010
box -4 -6 52 206
use FILL  SFILL14160x8100
timestamp 1596991774
transform -1 0 1432 0 -1 1010
box -4 -6 20 206
use FILL  SFILL14320x8100
timestamp 1596991774
transform -1 0 1448 0 -1 1010
box -4 -6 20 206
use FILL  SFILL14480x8100
timestamp 1596991774
transform -1 0 1464 0 -1 1010
box -4 -6 20 206
use BUFX2  BUFX2_insert36
timestamp 1596991774
transform -1 0 1688 0 -1 1010
box -4 -6 52 206
use OAI21X1  _2730_
timestamp 1596991774
transform -1 0 1752 0 -1 1010
box -4 -6 68 206
use NOR2X1  _3292_
timestamp 1596991774
transform -1 0 1800 0 -1 1010
box -4 -6 52 206
use AOI21X1  _2731_
timestamp 1596991774
transform -1 0 1864 0 -1 1010
box -4 -6 68 206
use NOR2X1  _2705_
timestamp 1596991774
transform -1 0 1912 0 -1 1010
box -4 -6 52 206
use OAI22X1  _3288_
timestamp 1596991774
transform -1 0 1992 0 -1 1010
box -4 -6 84 206
use INVX1  _3286_
timestamp 1596991774
transform -1 0 2024 0 -1 1010
box -4 -6 36 206
use NOR3X1  _2759_
timestamp 1596991774
transform 1 0 2024 0 -1 1010
box -4 -6 132 206
use AOI21X1  _2637_
timestamp 1596991774
transform -1 0 2216 0 -1 1010
box -4 -6 68 206
use AND2X2  _2625_
timestamp 1596991774
transform -1 0 2280 0 -1 1010
box -4 -6 68 206
use NAND3X1  _3018_
timestamp 1596991774
transform -1 0 2344 0 -1 1010
box -4 -6 68 206
use INVX1  _2994_
timestamp 1596991774
transform -1 0 2376 0 -1 1010
box -4 -6 36 206
use OAI22X1  _2995_
timestamp 1596991774
transform -1 0 2456 0 -1 1010
box -4 -6 84 206
use NOR2X1  _2999_
timestamp 1596991774
transform -1 0 2504 0 -1 1010
box -4 -6 52 206
use INVX1  _2997_
timestamp 1596991774
transform -1 0 2536 0 -1 1010
box -4 -6 36 206
use OAI22X1  _2998_
timestamp 1596991774
transform -1 0 2616 0 -1 1010
box -4 -6 84 206
use OAI21X1  _2808_
timestamp 1596991774
transform -1 0 2680 0 -1 1010
box -4 -6 68 206
use NAND2X1  _2806_
timestamp 1596991774
transform -1 0 2728 0 -1 1010
box -4 -6 52 206
use INVX1  _2799_
timestamp 1596991774
transform -1 0 2760 0 -1 1010
box -4 -6 36 206
use NOR2X1  _2299_
timestamp 1596991774
transform 1 0 2760 0 -1 1010
box -4 -6 52 206
use AND2X2  _2300_
timestamp 1596991774
transform -1 0 2872 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert54
timestamp 1596991774
transform -1 0 2920 0 -1 1010
box -4 -6 52 206
use OAI21X1  _2723_
timestamp 1596991774
transform -1 0 3048 0 -1 1010
box -4 -6 68 206
use FILL  SFILL29200x8100
timestamp 1596991774
transform -1 0 2936 0 -1 1010
box -4 -6 20 206
use FILL  SFILL29360x8100
timestamp 1596991774
transform -1 0 2952 0 -1 1010
box -4 -6 20 206
use FILL  SFILL29520x8100
timestamp 1596991774
transform -1 0 2968 0 -1 1010
box -4 -6 20 206
use FILL  SFILL29680x8100
timestamp 1596991774
transform -1 0 2984 0 -1 1010
box -4 -6 20 206
use AOI21X1  _2718_
timestamp 1596991774
transform 1 0 3048 0 -1 1010
box -4 -6 68 206
use NOR2X1  _2714_
timestamp 1596991774
transform 1 0 3112 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2717_
timestamp 1596991774
transform -1 0 3208 0 -1 1010
box -4 -6 52 206
use INVX1  _2713_
timestamp 1596991774
transform -1 0 3240 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert298
timestamp 1596991774
transform 1 0 3240 0 -1 1010
box -4 -6 52 206
use OAI22X1  _2623_
timestamp 1596991774
transform 1 0 3288 0 -1 1010
box -4 -6 84 206
use INVX1  _2620_
timestamp 1596991774
transform 1 0 3368 0 -1 1010
box -4 -6 36 206
use NAND2X1  _2621_
timestamp 1596991774
transform -1 0 3448 0 -1 1010
box -4 -6 52 206
use OAI21X1  _2632_
timestamp 1596991774
transform -1 0 3512 0 -1 1010
box -4 -6 68 206
use NOR3X1  _2624_
timestamp 1596991774
transform 1 0 3512 0 -1 1010
box -4 -6 132 206
use INVX1  _3453_
timestamp 1596991774
transform 1 0 3640 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert300
timestamp 1596991774
transform -1 0 3720 0 -1 1010
box -4 -6 52 206
use OAI21X1  _3447_
timestamp 1596991774
transform -1 0 3784 0 -1 1010
box -4 -6 68 206
use OAI21X1  _3461_
timestamp 1596991774
transform -1 0 3848 0 -1 1010
box -4 -6 68 206
use OAI21X1  _3468_
timestamp 1596991774
transform -1 0 3912 0 -1 1010
box -4 -6 68 206
use NAND3X1  _3403_
timestamp 1596991774
transform 1 0 3912 0 -1 1010
box -4 -6 68 206
use OAI21X1  _3402_
timestamp 1596991774
transform -1 0 4040 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3401_
timestamp 1596991774
transform -1 0 4088 0 -1 1010
box -4 -6 52 206
use NOR2X1  _3412_
timestamp 1596991774
transform 1 0 4088 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3604_
timestamp 1596991774
transform -1 0 4200 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3603_
timestamp 1596991774
transform 1 0 4200 0 -1 1010
box -4 -6 52 206
use OAI21X1  _3454_
timestamp 1596991774
transform -1 0 4312 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _3650_
timestamp 1596991774
transform 1 0 4312 0 -1 1010
box -4 -6 196 206
use AOI21X1  _3577_
timestamp 1596991774
transform -1 0 4632 0 -1 1010
box -4 -6 68 206
use FILL  SFILL45040x8100
timestamp 1596991774
transform -1 0 4520 0 -1 1010
box -4 -6 20 206
use FILL  SFILL45200x8100
timestamp 1596991774
transform -1 0 4536 0 -1 1010
box -4 -6 20 206
use FILL  SFILL45360x8100
timestamp 1596991774
transform -1 0 4552 0 -1 1010
box -4 -6 20 206
use FILL  SFILL45520x8100
timestamp 1596991774
transform -1 0 4568 0 -1 1010
box -4 -6 20 206
use NAND2X1  _3575_
timestamp 1596991774
transform -1 0 4680 0 -1 1010
box -4 -6 52 206
use NAND3X1  _3464_
timestamp 1596991774
transform -1 0 4744 0 -1 1010
box -4 -6 68 206
use NAND3X1  _3457_
timestamp 1596991774
transform 1 0 4744 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3458_
timestamp 1596991774
transform -1 0 4856 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert113
timestamp 1596991774
transform -1 0 4904 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3465_
timestamp 1596991774
transform -1 0 4952 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert114
timestamp 1596991774
transform 1 0 4952 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3459_
timestamp 1596991774
transform -1 0 5048 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3452_
timestamp 1596991774
transform 1 0 5048 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3438_
timestamp 1596991774
transform 1 0 5096 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4608_
timestamp 1596991774
transform -1 0 5208 0 -1 1010
box -4 -6 68 206
use INVX1  _4606_
timestamp 1596991774
transform -1 0 5240 0 -1 1010
box -4 -6 36 206
use NOR2X1  _3546_
timestamp 1596991774
transform -1 0 5288 0 -1 1010
box -4 -6 52 206
use INVX1  _4588_
timestamp 1596991774
transform 1 0 5288 0 -1 1010
box -4 -6 36 206
use NAND2X1  _4589_
timestamp 1596991774
transform -1 0 5368 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4590_
timestamp 1596991774
transform -1 0 5432 0 -1 1010
box -4 -6 68 206
use AND2X2  _3562_
timestamp 1596991774
transform 1 0 5432 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert172
timestamp 1596991774
transform -1 0 5544 0 -1 1010
box -4 -6 52 206
use INVX1  _4597_
timestamp 1596991774
transform 1 0 5544 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4599_
timestamp 1596991774
transform 1 0 5576 0 -1 1010
box -4 -6 68 206
use INVX1  _4618_
timestamp 1596991774
transform 1 0 5640 0 -1 1010
box -4 -6 36 206
use INVX1  _4603_
timestamp 1596991774
transform -1 0 5704 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4620_
timestamp 1596991774
transform 1 0 5704 0 -1 1010
box -4 -6 68 206
use OAI21X1  _4593_
timestamp 1596991774
transform 1 0 5768 0 -1 1010
box -4 -6 68 206
use INVX1  _4591_
timestamp 1596991774
transform -1 0 5864 0 -1 1010
box -4 -6 36 206
use AOI22X1  _4480_
timestamp 1596991774
transform 1 0 5864 0 -1 1010
box -4 -6 84 206
use AOI22X1  _4474_
timestamp 1596991774
transform 1 0 6008 0 -1 1010
box -4 -6 84 206
use FILL  SFILL59440x8100
timestamp 1596991774
transform -1 0 5960 0 -1 1010
box -4 -6 20 206
use FILL  SFILL59600x8100
timestamp 1596991774
transform -1 0 5976 0 -1 1010
box -4 -6 20 206
use FILL  SFILL59760x8100
timestamp 1596991774
transform -1 0 5992 0 -1 1010
box -4 -6 20 206
use FILL  SFILL59920x8100
timestamp 1596991774
transform -1 0 6008 0 -1 1010
box -4 -6 20 206
use AOI21X1  _4475_
timestamp 1596991774
transform 1 0 6088 0 -1 1010
box -4 -6 68 206
use OAI21X1  _2154_
timestamp 1596991774
transform -1 0 6216 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert193
timestamp 1596991774
transform 1 0 6216 0 -1 1010
box -4 -6 52 206
use INVX1  _2152_
timestamp 1596991774
transform -1 0 6296 0 -1 1010
box -4 -6 36 206
use OAI21X1  _2157_
timestamp 1596991774
transform -1 0 6360 0 -1 1010
box -4 -6 68 206
use INVX1  _2155_
timestamp 1596991774
transform -1 0 6392 0 -1 1010
box -4 -6 36 206
use DFFPOSX1  _4584_
timestamp 1596991774
transform -1 0 6584 0 -1 1010
box -4 -6 196 206
use AOI21X1  _4568_
timestamp 1596991774
transform -1 0 6648 0 -1 1010
box -4 -6 68 206
use INVX1  _4563_
timestamp 1596991774
transform 1 0 6648 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4564_
timestamp 1596991774
transform -1 0 6744 0 -1 1010
box -4 -6 68 206
use NAND3X1  _4567_
timestamp 1596991774
transform 1 0 6744 0 -1 1010
box -4 -6 68 206
use NAND3X1  _4566_
timestamp 1596991774
transform 1 0 6808 0 -1 1010
box -4 -6 68 206
use AOI22X1  _4540_
timestamp 1596991774
transform 1 0 6872 0 -1 1010
box -4 -6 84 206
use INVX1  _4543_
timestamp 1596991774
transform 1 0 6952 0 -1 1010
box -4 -6 36 206
use AOI22X1  _4534_
timestamp 1596991774
transform 1 0 6984 0 -1 1010
box -4 -6 84 206
use OAI21X1  _4539_
timestamp 1596991774
transform 1 0 7064 0 -1 1010
box -4 -6 68 206
use AOI21X1  _4535_
timestamp 1596991774
transform -1 0 7192 0 -1 1010
box -4 -6 68 206
use OAI21X1  _4541_
timestamp 1596991774
transform -1 0 7256 0 -1 1010
box -4 -6 68 206
use AND2X2  _4542_
timestamp 1596991774
transform 1 0 7256 0 -1 1010
box -4 -6 68 206
use NOR2X1  _4537_
timestamp 1596991774
transform -1 0 7368 0 -1 1010
box -4 -6 52 206
use FILL  FILL71120x8100
timestamp 1596991774
transform -1 0 7384 0 -1 1010
box -4 -6 20 206
use FILL  FILL71280x8100
timestamp 1596991774
transform -1 0 7400 0 -1 1010
box -4 -6 20 206
use BUFX2  BUFX2_insert139
timestamp 1596991774
transform 1 0 8 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert243
timestamp 1596991774
transform -1 0 104 0 1 1010
box -4 -6 52 206
use INVX1  _2884_
timestamp 1596991774
transform 1 0 104 0 1 1010
box -4 -6 36 206
use NAND2X1  _2919_
timestamp 1596991774
transform -1 0 184 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert269
timestamp 1596991774
transform -1 0 232 0 1 1010
box -4 -6 52 206
use OAI21X1  _2921_
timestamp 1596991774
transform -1 0 296 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert138
timestamp 1596991774
transform 1 0 296 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert272
timestamp 1596991774
transform 1 0 344 0 1 1010
box -4 -6 52 206
use INVX1  _2814_
timestamp 1596991774
transform 1 0 392 0 1 1010
box -4 -6 36 206
use OAI22X1  _2815_
timestamp 1596991774
transform -1 0 504 0 1 1010
box -4 -6 84 206
use NAND2X1  _2824_
timestamp 1596991774
transform 1 0 504 0 1 1010
box -4 -6 52 206
use OAI22X1  _2812_
timestamp 1596991774
transform 1 0 552 0 1 1010
box -4 -6 84 206
use INVX1  _2811_
timestamp 1596991774
transform -1 0 664 0 1 1010
box -4 -6 36 206
use NOR2X1  _2816_
timestamp 1596991774
transform -1 0 712 0 1 1010
box -4 -6 52 206
use AOI22X1  _2826_
timestamp 1596991774
transform 1 0 712 0 1 1010
box -4 -6 84 206
use NOR2X1  _2825_
timestamp 1596991774
transform 1 0 792 0 1 1010
box -4 -6 52 206
use INVX1  _2818_
timestamp 1596991774
transform 1 0 840 0 1 1010
box -4 -6 36 206
use AOI22X1  _2819_
timestamp 1596991774
transform 1 0 872 0 1 1010
box -4 -6 84 206
use NAND3X1  _2823_
timestamp 1596991774
transform -1 0 1016 0 1 1010
box -4 -6 68 206
use OR2X2  _2348_
timestamp 1596991774
transform -1 0 1080 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert67
timestamp 1596991774
transform 1 0 1080 0 1 1010
box -4 -6 52 206
use INVX1  _2604_
timestamp 1596991774
transform 1 0 1128 0 1 1010
box -4 -6 36 206
use AOI22X1  _2605_
timestamp 1596991774
transform -1 0 1240 0 1 1010
box -4 -6 84 206
use INVX1  _2603_
timestamp 1596991774
transform -1 0 1272 0 1 1010
box -4 -6 36 206
use OAI21X1  _2635_
timestamp 1596991774
transform 1 0 1272 0 1 1010
box -4 -6 68 206
use NAND2X1  _2609_
timestamp 1596991774
transform 1 0 1336 0 1 1010
box -4 -6 52 206
use INVX1  _2690_
timestamp 1596991774
transform 1 0 1384 0 1 1010
box -4 -6 36 206
use NAND2X1  _2727_
timestamp 1596991774
transform 1 0 1480 0 1 1010
box -4 -6 52 206
use NOR2X1  _2726_
timestamp 1596991774
transform -1 0 1576 0 1 1010
box -4 -6 52 206
use AOI21X1  _2729_
timestamp 1596991774
transform -1 0 1640 0 1 1010
box -4 -6 68 206
use FILL  SFILL14160x10100
timestamp 1596991774
transform 1 0 1416 0 1 1010
box -4 -6 20 206
use FILL  SFILL14320x10100
timestamp 1596991774
transform 1 0 1432 0 1 1010
box -4 -6 20 206
use FILL  SFILL14480x10100
timestamp 1596991774
transform 1 0 1448 0 1 1010
box -4 -6 20 206
use FILL  SFILL14640x10100
timestamp 1596991774
transform 1 0 1464 0 1 1010
box -4 -6 20 206
use NOR2X1  _2728_
timestamp 1596991774
transform 1 0 1640 0 1 1010
box -4 -6 52 206
use INVX1  _2693_
timestamp 1596991774
transform -1 0 1720 0 1 1010
box -4 -6 36 206
use OAI21X1  _2827_
timestamp 1596991774
transform -1 0 1784 0 1 1010
box -4 -6 68 206
use AOI22X1  _2692_
timestamp 1596991774
transform 1 0 1784 0 1 1010
box -4 -6 84 206
use NAND2X1  _2696_
timestamp 1596991774
transform 1 0 1864 0 1 1010
box -4 -6 52 206
use INVX1  _2691_
timestamp 1596991774
transform -1 0 1944 0 1 1010
box -4 -6 36 206
use INVX1  _2694_
timestamp 1596991774
transform 1 0 1944 0 1 1010
box -4 -6 36 206
use AOI22X1  _2695_
timestamp 1596991774
transform -1 0 2056 0 1 1010
box -4 -6 84 206
use NOR2X1  _3043_
timestamp 1596991774
transform 1 0 2056 0 1 1010
box -4 -6 52 206
use NOR2X1  _3069_
timestamp 1596991774
transform 1 0 2104 0 1 1010
box -4 -6 52 206
use NOR3X1  _2845_
timestamp 1596991774
transform 1 0 2152 0 1 1010
box -4 -6 132 206
use INVX1  _2840_
timestamp 1596991774
transform -1 0 2312 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert271
timestamp 1596991774
transform 1 0 2312 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert180
timestamp 1596991774
transform -1 0 2408 0 1 1010
box -4 -6 52 206
use AOI21X1  _2809_
timestamp 1596991774
transform 1 0 2408 0 1 1010
box -4 -6 68 206
use OAI21X1  _2844_
timestamp 1596991774
transform -1 0 2536 0 1 1010
box -4 -6 68 206
use INVX1  _2841_
timestamp 1596991774
transform -1 0 2568 0 1 1010
box -4 -6 36 206
use OR2X2  _2755_
timestamp 1596991774
transform 1 0 2568 0 1 1010
box -4 -6 68 206
use NAND2X1  _2756_
timestamp 1596991774
transform 1 0 2632 0 1 1010
box -4 -6 52 206
use AOI22X1  _2757_
timestamp 1596991774
transform -1 0 2760 0 1 1010
box -4 -6 84 206
use NOR2X1  _2301_
timestamp 1596991774
transform -1 0 2808 0 1 1010
box -4 -6 52 206
use NAND2X1  _2754_
timestamp 1596991774
transform -1 0 2856 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert97
timestamp 1596991774
transform -1 0 2904 0 1 1010
box -4 -6 52 206
use NAND2X1  _2716_
timestamp 1596991774
transform 1 0 2968 0 1 1010
box -4 -6 52 206
use FILL  SFILL29040x10100
timestamp 1596991774
transform 1 0 2904 0 1 1010
box -4 -6 20 206
use FILL  SFILL29200x10100
timestamp 1596991774
transform 1 0 2920 0 1 1010
box -4 -6 20 206
use FILL  SFILL29360x10100
timestamp 1596991774
transform 1 0 2936 0 1 1010
box -4 -6 20 206
use FILL  SFILL29520x10100
timestamp 1596991774
transform 1 0 2952 0 1 1010
box -4 -6 20 206
use INVX1  _2715_
timestamp 1596991774
transform -1 0 3048 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert96
timestamp 1596991774
transform 1 0 3048 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert137
timestamp 1596991774
transform 1 0 3096 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert164
timestamp 1596991774
transform 1 0 3144 0 1 1010
box -4 -6 52 206
use INVX1  _2618_
timestamp 1596991774
transform 1 0 3192 0 1 1010
box -4 -6 36 206
use NOR2X1  _2626_
timestamp 1596991774
transform -1 0 3272 0 1 1010
box -4 -6 52 206
use NAND2X1  _2619_
timestamp 1596991774
transform 1 0 3272 0 1 1010
box -4 -6 52 206
use AOI21X1  _2627_
timestamp 1596991774
transform -1 0 3384 0 1 1010
box -4 -6 68 206
use NAND2X1  _2622_
timestamp 1596991774
transform 1 0 3384 0 1 1010
box -4 -6 52 206
use INVX1  _3439_
timestamp 1596991774
transform 1 0 3432 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert70
timestamp 1596991774
transform 1 0 3464 0 1 1010
box -4 -6 52 206
use INVX1  _3474_
timestamp 1596991774
transform 1 0 3512 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert179
timestamp 1596991774
transform -1 0 3592 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert246
timestamp 1596991774
transform -1 0 3640 0 1 1010
box -4 -6 52 206
use OR2X2  _3427_
timestamp 1596991774
transform 1 0 3640 0 1 1010
box -4 -6 68 206
use OAI21X1  _3440_
timestamp 1596991774
transform -1 0 3768 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _3640_
timestamp 1596991774
transform -1 0 3960 0 1 1010
box -4 -6 196 206
use INVX1  _3518_
timestamp 1596991774
transform 1 0 3960 0 1 1010
box -4 -6 36 206
use INVX1  _3413_
timestamp 1596991774
transform 1 0 3992 0 1 1010
box -4 -6 36 206
use NAND3X1  _3519_
timestamp 1596991774
transform 1 0 4024 0 1 1010
box -4 -6 68 206
use INVX1  _3532_
timestamp 1596991774
transform 1 0 4088 0 1 1010
box -4 -6 36 206
use NAND3X1  _3533_
timestamp 1596991774
transform 1 0 4120 0 1 1010
box -4 -6 68 206
use NAND3X1  _3540_
timestamp 1596991774
transform -1 0 4248 0 1 1010
box -4 -6 68 206
use INVX1  _3539_
timestamp 1596991774
transform -1 0 4280 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert201
timestamp 1596991774
transform -1 0 4328 0 1 1010
box -4 -6 52 206
use NAND3X1  _3470_
timestamp 1596991774
transform -1 0 4392 0 1 1010
box -4 -6 68 206
use NAND3X1  _3471_
timestamp 1596991774
transform -1 0 4456 0 1 1010
box -4 -6 68 206
use INVX1  _3469_
timestamp 1596991774
transform -1 0 4552 0 1 1010
box -4 -6 36 206
use NAND3X1  _3477_
timestamp 1596991774
transform -1 0 4616 0 1 1010
box -4 -6 68 206
use INVX1  _3476_
timestamp 1596991774
transform -1 0 4648 0 1 1010
box -4 -6 36 206
use FILL  SFILL44560x10100
timestamp 1596991774
transform 1 0 4456 0 1 1010
box -4 -6 20 206
use FILL  SFILL44720x10100
timestamp 1596991774
transform 1 0 4472 0 1 1010
box -4 -6 20 206
use FILL  SFILL44880x10100
timestamp 1596991774
transform 1 0 4488 0 1 1010
box -4 -6 20 206
use FILL  SFILL45040x10100
timestamp 1596991774
transform 1 0 4504 0 1 1010
box -4 -6 20 206
use NAND3X1  _3442_
timestamp 1596991774
transform 1 0 4648 0 1 1010
box -4 -6 68 206
use NAND3X1  _3443_
timestamp 1596991774
transform -1 0 4776 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert202
timestamp 1596991774
transform 1 0 4776 0 1 1010
box -4 -6 52 206
use INVX1  _3431_
timestamp 1596991774
transform 1 0 4824 0 1 1010
box -4 -6 36 206
use INVX4  _3667_
timestamp 1596991774
transform -1 0 4904 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert124
timestamp 1596991774
transform 1 0 4904 0 1 1010
box -4 -6 52 206
use INVX4  _3425_
timestamp 1596991774
transform 1 0 4952 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert175
timestamp 1596991774
transform 1 0 5000 0 1 1010
box -4 -6 52 206
use NAND2X1  _4607_
timestamp 1596991774
transform 1 0 5048 0 1 1010
box -4 -6 52 206
use NAND2X1  _3444_
timestamp 1596991774
transform -1 0 5144 0 1 1010
box -4 -6 52 206
use AND2X2  _3563_
timestamp 1596991774
transform 1 0 5144 0 1 1010
box -4 -6 68 206
use INVX1  _3551_
timestamp 1596991774
transform 1 0 5208 0 1 1010
box -4 -6 36 206
use NOR2X1  _3552_
timestamp 1596991774
transform -1 0 5288 0 1 1010
box -4 -6 52 206
use INVX4  _3658_
timestamp 1596991774
transform 1 0 5288 0 1 1010
box -4 -6 52 206
use INVX1  _4621_
timestamp 1596991774
transform 1 0 5336 0 1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert174
timestamp 1596991774
transform 1 0 5368 0 1 1010
box -4 -6 52 206
use OAI21X1  _4623_
timestamp 1596991774
transform 1 0 5416 0 1 1010
box -4 -6 68 206
use NAND2X1  _4622_
timestamp 1596991774
transform -1 0 5528 0 1 1010
box -4 -6 52 206
use NAND2X1  _4601_
timestamp 1596991774
transform -1 0 5576 0 1 1010
box -4 -6 52 206
use NAND2X1  _4598_
timestamp 1596991774
transform 1 0 5576 0 1 1010
box -4 -6 52 206
use OAI21X1  _4602_
timestamp 1596991774
transform -1 0 5688 0 1 1010
box -4 -6 68 206
use INVX1  _4600_
timestamp 1596991774
transform -1 0 5720 0 1 1010
box -4 -6 36 206
use NAND2X1  _2153_
timestamp 1596991774
transform -1 0 5768 0 1 1010
box -4 -6 52 206
use NAND2X1  _2129_
timestamp 1596991774
transform -1 0 5816 0 1 1010
box -4 -6 52 206
use NOR2X1  _3548_
timestamp 1596991774
transform 1 0 5816 0 1 1010
box -4 -6 52 206
use NAND2X1  _2156_
timestamp 1596991774
transform -1 0 5912 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _4570_
timestamp 1596991774
transform -1 0 6168 0 1 1010
box -4 -6 196 206
use FILL  SFILL59120x10100
timestamp 1596991774
transform 1 0 5912 0 1 1010
box -4 -6 20 206
use FILL  SFILL59280x10100
timestamp 1596991774
transform 1 0 5928 0 1 1010
box -4 -6 20 206
use FILL  SFILL59440x10100
timestamp 1596991774
transform 1 0 5944 0 1 1010
box -4 -6 20 206
use FILL  SFILL59600x10100
timestamp 1596991774
transform 1 0 5960 0 1 1010
box -4 -6 20 206
use BUFX2  BUFX2_insert190
timestamp 1596991774
transform 1 0 6168 0 1 1010
box -4 -6 52 206
use AOI22X1  _4546_
timestamp 1596991774
transform 1 0 6216 0 1 1010
box -4 -6 84 206
use OAI21X1  _2163_
timestamp 1596991774
transform -1 0 6360 0 1 1010
box -4 -6 68 206
use INVX1  _2161_
timestamp 1596991774
transform -1 0 6392 0 1 1010
box -4 -6 36 206
use NAND2X1  _4562_
timestamp 1596991774
transform 1 0 6392 0 1 1010
box -4 -6 52 206
use OAI21X1  _4552_
timestamp 1596991774
transform -1 0 6504 0 1 1010
box -4 -6 68 206
use NAND3X1  _4556_
timestamp 1596991774
transform -1 0 6568 0 1 1010
box -4 -6 68 206
use NAND3X1  _4559_
timestamp 1596991774
transform -1 0 6632 0 1 1010
box -4 -6 68 206
use OAI21X1  _4558_
timestamp 1596991774
transform -1 0 6696 0 1 1010
box -4 -6 68 206
use NOR3X1  _4565_
timestamp 1596991774
transform -1 0 6824 0 1 1010
box -4 -6 132 206
use OAI21X1  _4547_
timestamp 1596991774
transform -1 0 6888 0 1 1010
box -4 -6 68 206
use OAI21X1  _4545_
timestamp 1596991774
transform -1 0 6952 0 1 1010
box -4 -6 68 206
use NOR3X1  _4544_
timestamp 1596991774
transform 1 0 6952 0 1 1010
box -4 -6 132 206
use DFFPOSX1  _4579_
timestamp 1596991774
transform 1 0 7080 0 1 1010
box -4 -6 196 206
use INVX1  _2146_
timestamp 1596991774
transform 1 0 7272 0 1 1010
box -4 -6 36 206
use OAI21X1  _2148_
timestamp 1596991774
transform 1 0 7304 0 1 1010
box -4 -6 68 206
use FILL  FILL71120x10100
timestamp 1596991774
transform 1 0 7368 0 1 1010
box -4 -6 20 206
use FILL  FILL71280x10100
timestamp 1596991774
transform 1 0 7384 0 1 1010
box -4 -6 20 206
use BUFX2  _2108_
timestamp 1596991774
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use NAND2X1  _2191_
timestamp 1596991774
transform -1 0 104 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert245
timestamp 1596991774
transform 1 0 104 0 -1 1410
box -4 -6 52 206
use AND2X2  _2205_
timestamp 1596991774
transform -1 0 216 0 -1 1410
box -4 -6 68 206
use AND2X2  _2312_
timestamp 1596991774
transform 1 0 216 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert273
timestamp 1596991774
transform 1 0 280 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert69
timestamp 1596991774
transform -1 0 376 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert136
timestamp 1596991774
transform 1 0 376 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert244
timestamp 1596991774
transform 1 0 424 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert38
timestamp 1596991774
transform -1 0 520 0 -1 1410
box -4 -6 52 206
use INVX1  _2810_
timestamp 1596991774
transform 1 0 520 0 -1 1410
box -4 -6 36 206
use BUFX2  BUFX2_insert178
timestamp 1596991774
transform 1 0 552 0 -1 1410
box -4 -6 52 206
use AND2X2  _2309_
timestamp 1596991774
transform 1 0 600 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert39
timestamp 1596991774
transform 1 0 664 0 -1 1410
box -4 -6 52 206
use AND2X2  _2362_
timestamp 1596991774
transform 1 0 712 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3117_
timestamp 1596991774
transform 1 0 776 0 -1 1410
box -4 -6 52 206
use INVX1  _3159_
timestamp 1596991774
transform 1 0 824 0 -1 1410
box -4 -6 36 206
use OAI21X1  _3161_
timestamp 1596991774
transform 1 0 856 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3160_
timestamp 1596991774
transform -1 0 968 0 -1 1410
box -4 -6 52 206
use AOI21X1  _2922_
timestamp 1596991774
transform -1 0 1032 0 -1 1410
box -4 -6 68 206
use NOR2X1  _3162_
timestamp 1596991774
transform -1 0 1080 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3174_
timestamp 1596991774
transform 1 0 1080 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3143_
timestamp 1596991774
transform -1 0 1192 0 -1 1410
box -4 -6 52 206
use AND2X2  _2363_
timestamp 1596991774
transform -1 0 1256 0 -1 1410
box -4 -6 68 206
use AND2X2  _2938_
timestamp 1596991774
transform -1 0 1320 0 -1 1410
box -4 -6 68 206
use INVX1  _2607_
timestamp 1596991774
transform -1 0 1352 0 -1 1410
box -4 -6 36 206
use AOI22X1  _2608_
timestamp 1596991774
transform -1 0 1432 0 -1 1410
box -4 -6 84 206
use OAI22X1  _2634_
timestamp 1596991774
transform -1 0 1576 0 -1 1410
box -4 -6 84 206
use BUFX2  BUFX2_insert270
timestamp 1596991774
transform 1 0 1576 0 -1 1410
box -4 -6 52 206
use FILL  SFILL14320x12100
timestamp 1596991774
transform -1 0 1448 0 -1 1410
box -4 -6 20 206
use FILL  SFILL14480x12100
timestamp 1596991774
transform -1 0 1464 0 -1 1410
box -4 -6 20 206
use FILL  SFILL14640x12100
timestamp 1596991774
transform -1 0 1480 0 -1 1410
box -4 -6 20 206
use FILL  SFILL14800x12100
timestamp 1596991774
transform -1 0 1496 0 -1 1410
box -4 -6 20 206
use AND2X2  _2364_
timestamp 1596991774
transform -1 0 1688 0 -1 1410
box -4 -6 68 206
use INVX1  _2606_
timestamp 1596991774
transform -1 0 1720 0 -1 1410
box -4 -6 36 206
use NAND2X1  _3059_
timestamp 1596991774
transform 1 0 1720 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3064_
timestamp 1596991774
transform 1 0 1768 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3033_
timestamp 1596991774
transform 1 0 1832 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3038_
timestamp 1596991774
transform 1 0 1880 0 -1 1410
box -4 -6 68 206
use NAND3X1  _3060_
timestamp 1596991774
transform -1 0 2008 0 -1 1410
box -4 -6 68 206
use NAND3X1  _3034_
timestamp 1596991774
transform -1 0 2072 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3007_
timestamp 1596991774
transform -1 0 2120 0 -1 1410
box -4 -6 52 206
use XOR2X1  _2374_
timestamp 1596991774
transform 1 0 2120 0 -1 1410
box -4 -6 116 206
use NAND3X1  _3042_
timestamp 1596991774
transform 1 0 2232 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3039_
timestamp 1596991774
transform -1 0 2344 0 -1 1410
box -4 -6 52 206
use INVX1  _3481_
timestamp 1596991774
transform 1 0 2344 0 -1 1410
box -4 -6 36 206
use NAND2X1  _3013_
timestamp 1596991774
transform -1 0 2424 0 -1 1410
box -4 -6 52 206
use INVX1  _2993_
timestamp 1596991774
transform -1 0 2456 0 -1 1410
box -4 -6 36 206
use AND2X2  _2358_
timestamp 1596991774
transform -1 0 2520 0 -1 1410
box -4 -6 68 206
use OR2X2  _2342_
timestamp 1596991774
transform -1 0 2584 0 -1 1410
box -4 -6 68 206
use AND2X2  _2359_
timestamp 1596991774
transform -1 0 2648 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2843_
timestamp 1596991774
transform -1 0 2696 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2797_
timestamp 1596991774
transform 1 0 2696 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2796_
timestamp 1596991774
transform 1 0 2760 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2842_
timestamp 1596991774
transform 1 0 2808 0 -1 1410
box -4 -6 68 206
use OR2X2  _2753_
timestamp 1596991774
transform -1 0 2936 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert267
timestamp 1596991774
transform -1 0 3048 0 -1 1410
box -4 -6 52 206
use FILL  SFILL29360x12100
timestamp 1596991774
transform -1 0 2952 0 -1 1410
box -4 -6 20 206
use FILL  SFILL29520x12100
timestamp 1596991774
transform -1 0 2968 0 -1 1410
box -4 -6 20 206
use FILL  SFILL29680x12100
timestamp 1596991774
transform -1 0 2984 0 -1 1410
box -4 -6 20 206
use FILL  SFILL29840x12100
timestamp 1596991774
transform -1 0 3000 0 -1 1410
box -4 -6 20 206
use NOR2X1  _2937_
timestamp 1596991774
transform 1 0 3048 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2914_
timestamp 1596991774
transform -1 0 3160 0 -1 1410
box -4 -6 68 206
use XNOR2X1  _2935_
timestamp 1596991774
transform -1 0 3272 0 -1 1410
box -4 -6 116 206
use NAND2X1  _2936_
timestamp 1596991774
transform -1 0 3320 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert266
timestamp 1596991774
transform 1 0 3320 0 -1 1410
box -4 -6 52 206
use XNOR2X1  _2420_
timestamp 1596991774
transform -1 0 3480 0 -1 1410
box -4 -6 116 206
use DFFPOSX1  _4451_
timestamp 1596991774
transform -1 0 3672 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _4450_
timestamp 1596991774
transform -1 0 3864 0 -1 1410
box -4 -6 196 206
use OAI21X1  _3482_
timestamp 1596991774
transform -1 0 3928 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3429_
timestamp 1596991774
transform 1 0 3928 0 -1 1410
box -4 -6 52 206
use INVX1  _3428_
timestamp 1596991774
transform -1 0 4008 0 -1 1410
box -4 -6 36 206
use DFFPOSX1  _4434_
timestamp 1596991774
transform -1 0 4200 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _4435_
timestamp 1596991774
transform -1 0 4392 0 -1 1410
box -4 -6 196 206
use NAND3X1  _3520_
timestamp 1596991774
transform -1 0 4456 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3521_
timestamp 1596991774
transform -1 0 4568 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3475_
timestamp 1596991774
transform -1 0 4632 0 -1 1410
box -4 -6 68 206
use FILL  SFILL44560x12100
timestamp 1596991774
transform -1 0 4472 0 -1 1410
box -4 -6 20 206
use FILL  SFILL44720x12100
timestamp 1596991774
transform -1 0 4488 0 -1 1410
box -4 -6 20 206
use FILL  SFILL44880x12100
timestamp 1596991774
transform -1 0 4504 0 -1 1410
box -4 -6 20 206
use FILL  SFILL45040x12100
timestamp 1596991774
transform -1 0 4520 0 -1 1410
box -4 -6 20 206
use NAND3X1  _3485_
timestamp 1596991774
transform 1 0 4632 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3486_
timestamp 1596991774
transform -1 0 4744 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3478_
timestamp 1596991774
transform -1 0 4808 0 -1 1410
box -4 -6 68 206
use NAND3X1  _3484_
timestamp 1596991774
transform -1 0 4872 0 -1 1410
box -4 -6 68 206
use INVX1  _3483_
timestamp 1596991774
transform -1 0 4904 0 -1 1410
box -4 -6 36 206
use BUFX2  BUFX2_insert129
timestamp 1596991774
transform 1 0 4904 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3582_
timestamp 1596991774
transform -1 0 5000 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3585_
timestamp 1596991774
transform -1 0 5048 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3579_
timestamp 1596991774
transform -1 0 5096 0 -1 1410
box -4 -6 52 206
use INVX8  _3568_
timestamp 1596991774
transform 1 0 5096 0 -1 1410
box -4 -6 84 206
use NAND2X1  _3480_
timestamp 1596991774
transform -1 0 5224 0 -1 1410
box -4 -6 52 206
use INVX1  _3557_
timestamp 1596991774
transform 1 0 5224 0 -1 1410
box -4 -6 36 206
use NOR2X1  _3558_
timestamp 1596991774
transform -1 0 5304 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3515_
timestamp 1596991774
transform -1 0 5352 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3487_
timestamp 1596991774
transform -1 0 5400 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3494_
timestamp 1596991774
transform -1 0 5448 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3424_
timestamp 1596991774
transform 1 0 5448 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert123
timestamp 1596991774
transform -1 0 5544 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert126
timestamp 1596991774
transform 1 0 5544 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3508_
timestamp 1596991774
transform -1 0 5640 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _3635_
timestamp 1596991774
transform 1 0 5640 0 -1 1410
box -4 -6 196 206
use NAND2X1  _3473_
timestamp 1596991774
transform -1 0 5880 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3479_
timestamp 1596991774
transform 1 0 5880 0 -1 1410
box -4 -6 52 206
use INVX1  _3553_
timestamp 1596991774
transform 1 0 5992 0 -1 1410
box -4 -6 36 206
use FILL  SFILL59280x12100
timestamp 1596991774
transform -1 0 5944 0 -1 1410
box -4 -6 20 206
use FILL  SFILL59440x12100
timestamp 1596991774
transform -1 0 5960 0 -1 1410
box -4 -6 20 206
use FILL  SFILL59600x12100
timestamp 1596991774
transform -1 0 5976 0 -1 1410
box -4 -6 20 206
use FILL  SFILL59760x12100
timestamp 1596991774
transform -1 0 5992 0 -1 1410
box -4 -6 20 206
use NOR2X1  _3554_
timestamp 1596991774
transform -1 0 6072 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3466_
timestamp 1596991774
transform -1 0 6120 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3472_
timestamp 1596991774
transform 1 0 6120 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3445_
timestamp 1596991774
transform 1 0 6168 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert173
timestamp 1596991774
transform -1 0 6264 0 -1 1410
box -4 -6 52 206
use INVX1  _3547_
timestamp 1596991774
transform -1 0 6296 0 -1 1410
box -4 -6 36 206
use BUFX2  BUFX2_insert171
timestamp 1596991774
transform 1 0 6296 0 -1 1410
box -4 -6 52 206
use INVX1  _4615_
timestamp 1596991774
transform 1 0 6344 0 -1 1410
box -4 -6 36 206
use OAI21X1  _4617_
timestamp 1596991774
transform -1 0 6440 0 -1 1410
box -4 -6 68 206
use INVX1  _4627_
timestamp 1596991774
transform 1 0 6440 0 -1 1410
box -4 -6 36 206
use OAI21X1  _4629_
timestamp 1596991774
transform 1 0 6472 0 -1 1410
box -4 -6 68 206
use AOI22X1  _4553_
timestamp 1596991774
transform 1 0 6536 0 -1 1410
box -4 -6 84 206
use AOI21X1  _4561_
timestamp 1596991774
transform -1 0 6680 0 -1 1410
box -4 -6 68 206
use AOI22X1  _4560_
timestamp 1596991774
transform 1 0 6680 0 -1 1410
box -4 -6 84 206
use INVX1  _4557_
timestamp 1596991774
transform -1 0 6792 0 -1 1410
box -4 -6 36 206
use INVX1  _4549_
timestamp 1596991774
transform 1 0 6792 0 -1 1410
box -4 -6 36 206
use NOR2X1  _4551_
timestamp 1596991774
transform 1 0 6824 0 -1 1410
box -4 -6 52 206
use OAI21X1  _4554_
timestamp 1596991774
transform 1 0 6872 0 -1 1410
box -4 -6 68 206
use AND2X2  _4555_
timestamp 1596991774
transform 1 0 6936 0 -1 1410
box -4 -6 68 206
use NAND3X1  _4550_
timestamp 1596991774
transform 1 0 7000 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _4581_
timestamp 1596991774
transform -1 0 7256 0 -1 1410
box -4 -6 196 206
use NAND2X1  _3570_
timestamp 1596991774
transform -1 0 7304 0 -1 1410
box -4 -6 52 206
use OAI21X1  _4517_
timestamp 1596991774
transform -1 0 7368 0 -1 1410
box -4 -6 68 206
use FILL  FILL71120x12100
timestamp 1596991774
transform -1 0 7384 0 -1 1410
box -4 -6 20 206
use FILL  FILL71280x12100
timestamp 1596991774
transform -1 0 7400 0 -1 1410
box -4 -6 20 206
use NOR2X1  _2200_
timestamp 1596991774
transform 1 0 8 0 1 1410
box -4 -6 52 206
use NOR2X1  _2199_
timestamp 1596991774
transform -1 0 104 0 1 1410
box -4 -6 52 206
use AND2X2  _2196_
timestamp 1596991774
transform -1 0 168 0 1 1410
box -4 -6 68 206
use OR2X2  _2192_
timestamp 1596991774
transform -1 0 232 0 1 1410
box -4 -6 68 206
use NOR2X1  _2206_
timestamp 1596991774
transform 1 0 232 0 1 1410
box -4 -6 52 206
use NOR2X1  _2313_
timestamp 1596991774
transform -1 0 328 0 1 1410
box -4 -6 52 206
use NOR2X1  _2311_
timestamp 1596991774
transform -1 0 376 0 1 1410
box -4 -6 52 206
use XNOR2X1  _2203_
timestamp 1596991774
transform -1 0 488 0 1 1410
box -4 -6 116 206
use NOR2X1  _2308_
timestamp 1596991774
transform 1 0 488 0 1 1410
box -4 -6 52 206
use AND2X2  _2315_
timestamp 1596991774
transform 1 0 536 0 1 1410
box -4 -6 68 206
use NOR2X1  _2316_
timestamp 1596991774
transform -1 0 648 0 1 1410
box -4 -6 52 206
use NOR2X1  _2310_
timestamp 1596991774
transform 1 0 648 0 1 1410
box -4 -6 52 206
use NAND3X1  _3164_
timestamp 1596991774
transform 1 0 696 0 1 1410
box -4 -6 68 206
use NAND3X1  _3112_
timestamp 1596991774
transform 1 0 760 0 1 1410
box -4 -6 68 206
use NAND3X1  _3138_
timestamp 1596991774
transform 1 0 824 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert288
timestamp 1596991774
transform -1 0 936 0 1 1410
box -4 -6 52 206
use NAND3X1  _3120_
timestamp 1596991774
transform -1 0 1000 0 1 1410
box -4 -6 68 206
use NOR2X1  _3121_
timestamp 1596991774
transform 1 0 1000 0 1 1410
box -4 -6 52 206
use AOI22X1  _3119_
timestamp 1596991774
transform -1 0 1128 0 1 1410
box -4 -6 84 206
use NOR2X1  _3147_
timestamp 1596991774
transform 1 0 1128 0 1 1410
box -4 -6 52 206
use NAND3X1  _3146_
timestamp 1596991774
transform -1 0 1240 0 1 1410
box -4 -6 68 206
use NOR2X1  _3173_
timestamp 1596991774
transform 1 0 1240 0 1 1410
box -4 -6 52 206
use NAND3X1  _3144_
timestamp 1596991774
transform 1 0 1288 0 1 1410
box -4 -6 68 206
use NAND3X1  _3172_
timestamp 1596991774
transform 1 0 1352 0 1 1410
box -4 -6 68 206
use INVX1  _3157_
timestamp 1596991774
transform 1 0 1480 0 1 1410
box -4 -6 36 206
use OAI22X1  _3158_
timestamp 1596991774
transform -1 0 1592 0 1 1410
box -4 -6 84 206
use NAND2X1  _3169_
timestamp 1596991774
transform -1 0 1640 0 1 1410
box -4 -6 52 206
use FILL  SFILL14160x14100
timestamp 1596991774
transform 1 0 1416 0 1 1410
box -4 -6 20 206
use FILL  SFILL14320x14100
timestamp 1596991774
transform 1 0 1432 0 1 1410
box -4 -6 20 206
use FILL  SFILL14480x14100
timestamp 1596991774
transform 1 0 1448 0 1 1410
box -4 -6 20 206
use FILL  SFILL14640x14100
timestamp 1596991774
transform 1 0 1464 0 1 1410
box -4 -6 20 206
use INVX1  _3156_
timestamp 1596991774
transform -1 0 1672 0 1 1410
box -4 -6 36 206
use INVX1  _3365_
timestamp 1596991774
transform 1 0 1672 0 1 1410
box -4 -6 36 206
use OAI22X1  _3366_
timestamp 1596991774
transform -1 0 1784 0 1 1410
box -4 -6 84 206
use INVX1  _3364_
timestamp 1596991774
transform -1 0 1816 0 1 1410
box -4 -6 36 206
use AND2X2  _3063_
timestamp 1596991774
transform -1 0 1880 0 1 1410
box -4 -6 68 206
use AND2X2  _3037_
timestamp 1596991774
transform 1 0 1880 0 1 1410
box -4 -6 68 206
use XOR2X1  _2373_
timestamp 1596991774
transform 1 0 1944 0 1 1410
box -4 -6 116 206
use AND2X2  _3011_
timestamp 1596991774
transform 1 0 2056 0 1 1410
box -4 -6 68 206
use NOR2X1  _2375_
timestamp 1596991774
transform 1 0 2120 0 1 1410
box -4 -6 52 206
use NAND3X1  _3012_
timestamp 1596991774
transform 1 0 2168 0 1 1410
box -4 -6 68 206
use NAND3X1  _3008_
timestamp 1596991774
transform -1 0 2296 0 1 1410
box -4 -6 68 206
use NOR2X1  _3017_
timestamp 1596991774
transform 1 0 2296 0 1 1410
box -4 -6 52 206
use NAND3X1  _3014_
timestamp 1596991774
transform -1 0 2408 0 1 1410
box -4 -6 68 206
use NAND3X1  _3016_
timestamp 1596991774
transform 1 0 2408 0 1 1410
box -4 -6 68 206
use AOI22X1  _3041_
timestamp 1596991774
transform -1 0 2552 0 1 1410
box -4 -6 84 206
use AOI22X1  _3015_
timestamp 1596991774
transform 1 0 2552 0 1 1410
box -4 -6 84 206
use NOR2X1  _2167_
timestamp 1596991774
transform -1 0 2680 0 1 1410
box -4 -6 52 206
use AND2X2  _2297_
timestamp 1596991774
transform 1 0 2680 0 1 1410
box -4 -6 68 206
use NOR2X1  _2298_
timestamp 1596991774
transform -1 0 2792 0 1 1410
box -4 -6 52 206
use NOR2X1  _2296_
timestamp 1596991774
transform -1 0 2840 0 1 1410
box -4 -6 52 206
use NAND2X1  _2793_
timestamp 1596991774
transform 1 0 2840 0 1 1410
box -4 -6 52 206
use NOR2X1  _2794_
timestamp 1596991774
transform -1 0 2936 0 1 1410
box -4 -6 52 206
use OR2X2  _2413_
timestamp 1596991774
transform -1 0 3064 0 1 1410
box -4 -6 68 206
use FILL  SFILL29360x14100
timestamp 1596991774
transform 1 0 2936 0 1 1410
box -4 -6 20 206
use FILL  SFILL29520x14100
timestamp 1596991774
transform 1 0 2952 0 1 1410
box -4 -6 20 206
use FILL  SFILL29680x14100
timestamp 1596991774
transform 1 0 2968 0 1 1410
box -4 -6 20 206
use FILL  SFILL29840x14100
timestamp 1596991774
transform 1 0 2984 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_insert162
timestamp 1596991774
transform -1 0 3112 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert297
timestamp 1596991774
transform -1 0 3160 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert163
timestamp 1596991774
transform -1 0 3208 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert37
timestamp 1596991774
transform -1 0 3256 0 1 1410
box -4 -6 52 206
use XNOR2X1  _2419_
timestamp 1596991774
transform 1 0 3256 0 1 1410
box -4 -6 116 206
use NAND2X1  _2421_
timestamp 1596991774
transform 1 0 3368 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _4449_
timestamp 1596991774
transform -1 0 3608 0 1 1410
box -4 -6 196 206
use OAI21X1  _3999_
timestamp 1596991774
transform 1 0 3608 0 1 1410
box -4 -6 68 206
use AOI21X1  _4000_
timestamp 1596991774
transform -1 0 3736 0 1 1410
box -4 -6 68 206
use OAI21X1  _3988_
timestamp 1596991774
transform 1 0 3736 0 1 1410
box -4 -6 68 206
use AOI21X1  _3989_
timestamp 1596991774
transform -1 0 3864 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert184
timestamp 1596991774
transform -1 0 3912 0 1 1410
box -4 -6 52 206
use OAI21X1  _3517_
timestamp 1596991774
transform -1 0 3976 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _4430_
timestamp 1596991774
transform -1 0 4168 0 1 1410
box -4 -6 196 206
use DFFPOSX1  _4433_
timestamp 1596991774
transform -1 0 4360 0 1 1410
box -4 -6 196 206
use OAI21X1  _4177_
timestamp 1596991774
transform 1 0 4360 0 1 1410
box -4 -6 68 206
use AOI21X1  _4178_
timestamp 1596991774
transform -1 0 4552 0 1 1410
box -4 -6 68 206
use INVX1  _3525_
timestamp 1596991774
transform 1 0 4552 0 1 1410
box -4 -6 36 206
use NAND3X1  _3526_
timestamp 1596991774
transform 1 0 4584 0 1 1410
box -4 -6 68 206
use FILL  SFILL44240x14100
timestamp 1596991774
transform 1 0 4424 0 1 1410
box -4 -6 20 206
use FILL  SFILL44400x14100
timestamp 1596991774
transform 1 0 4440 0 1 1410
box -4 -6 20 206
use FILL  SFILL44560x14100
timestamp 1596991774
transform 1 0 4456 0 1 1410
box -4 -6 20 206
use FILL  SFILL44720x14100
timestamp 1596991774
transform 1 0 4472 0 1 1410
box -4 -6 20 206
use INVX4  _3676_
timestamp 1596991774
transform -1 0 4696 0 1 1410
box -4 -6 52 206
use OAI21X1  _4166_
timestamp 1596991774
transform 1 0 4696 0 1 1410
box -4 -6 68 206
use AOI21X1  _4167_
timestamp 1596991774
transform -1 0 4824 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _3637_
timestamp 1596991774
transform 1 0 4824 0 1 1410
box -4 -6 196 206
use AOI21X1  _3625_
timestamp 1596991774
transform -1 0 5080 0 1 1410
box -4 -6 68 206
use INVX1  _3490_
timestamp 1596991774
transform 1 0 5080 0 1 1410
box -4 -6 36 206
use NAND3X1  _3491_
timestamp 1596991774
transform 1 0 5112 0 1 1410
box -4 -6 68 206
use NAND2X1  _3624_
timestamp 1596991774
transform -1 0 5224 0 1 1410
box -4 -6 52 206
use AND2X2  _3566_
timestamp 1596991774
transform 1 0 5224 0 1 1410
box -4 -6 68 206
use NAND3X1  _3435_
timestamp 1596991774
transform 1 0 5288 0 1 1410
box -4 -6 68 206
use NAND3X1  _3450_
timestamp 1596991774
transform 1 0 5352 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert111
timestamp 1596991774
transform 1 0 5416 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert130
timestamp 1596991774
transform 1 0 5464 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert125
timestamp 1596991774
transform 1 0 5512 0 1 1410
box -4 -6 52 206
use AOI21X1  _3621_
timestamp 1596991774
transform -1 0 5624 0 1 1410
box -4 -6 68 206
use NAND2X1  _3620_
timestamp 1596991774
transform -1 0 5672 0 1 1410
box -4 -6 52 206
use AND2X2  _3564_
timestamp 1596991774
transform -1 0 5736 0 1 1410
box -4 -6 68 206
use NAND2X1  _4619_
timestamp 1596991774
transform -1 0 5784 0 1 1410
box -4 -6 52 206
use INVX1  _4624_
timestamp 1596991774
transform 1 0 5784 0 1 1410
box -4 -6 36 206
use NOR2X1  _3556_
timestamp 1596991774
transform 1 0 5816 0 1 1410
box -4 -6 52 206
use NAND2X1  _4625_
timestamp 1596991774
transform 1 0 5864 0 1 1410
box -4 -6 52 206
use INVX1  _3555_
timestamp 1596991774
transform -1 0 5944 0 1 1410
box -4 -6 36 206
use OAI21X1  _4626_
timestamp 1596991774
transform -1 0 6072 0 1 1410
box -4 -6 68 206
use FILL  SFILL59440x14100
timestamp 1596991774
transform 1 0 5944 0 1 1410
box -4 -6 20 206
use FILL  SFILL59600x14100
timestamp 1596991774
transform 1 0 5960 0 1 1410
box -4 -6 20 206
use FILL  SFILL59760x14100
timestamp 1596991774
transform 1 0 5976 0 1 1410
box -4 -6 20 206
use FILL  SFILL59920x14100
timestamp 1596991774
transform 1 0 5992 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_insert112
timestamp 1596991774
transform 1 0 6072 0 1 1410
box -4 -6 52 206
use INVX1  _4630_
timestamp 1596991774
transform 1 0 6120 0 1 1410
box -4 -6 36 206
use AND2X2  _3565_
timestamp 1596991774
transform 1 0 6152 0 1 1410
box -4 -6 68 206
use NAND2X1  _2162_
timestamp 1596991774
transform 1 0 6216 0 1 1410
box -4 -6 52 206
use AND2X2  _3561_
timestamp 1596991774
transform -1 0 6328 0 1 1410
box -4 -6 68 206
use NAND2X1  _4616_
timestamp 1596991774
transform 1 0 6328 0 1 1410
box -4 -6 52 206
use OAI21X1  _4632_
timestamp 1596991774
transform 1 0 6376 0 1 1410
box -4 -6 68 206
use NAND2X1  _4631_
timestamp 1596991774
transform -1 0 6488 0 1 1410
box -4 -6 52 206
use NAND2X1  _4628_
timestamp 1596991774
transform 1 0 6488 0 1 1410
box -4 -6 52 206
use NAND2X1  _2159_
timestamp 1596991774
transform 1 0 6536 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _4583_
timestamp 1596991774
transform 1 0 6584 0 1 1410
box -4 -6 196 206
use DFFPOSX1  _4582_
timestamp 1596991774
transform -1 0 6968 0 1 1410
box -4 -6 196 206
use INVX1  _2158_
timestamp 1596991774
transform 1 0 6968 0 1 1410
box -4 -6 36 206
use OAI21X1  _2160_
timestamp 1596991774
transform -1 0 7064 0 1 1410
box -4 -6 68 206
use AND2X2  _4548_
timestamp 1596991774
transform 1 0 7064 0 1 1410
box -4 -6 68 206
use INVX4  _4460_
timestamp 1596991774
transform -1 0 7176 0 1 1410
box -4 -6 52 206
use NAND2X1  _2150_
timestamp 1596991774
transform -1 0 7224 0 1 1410
box -4 -6 52 206
use OAI21X1  _2151_
timestamp 1596991774
transform 1 0 7224 0 1 1410
box -4 -6 68 206
use INVX1  _2149_
timestamp 1596991774
transform -1 0 7320 0 1 1410
box -4 -6 36 206
use NAND2X1  _2147_
timestamp 1596991774
transform -1 0 7368 0 1 1410
box -4 -6 52 206
use FILL  FILL71120x14100
timestamp 1596991774
transform 1 0 7368 0 1 1410
box -4 -6 20 206
use FILL  FILL71280x14100
timestamp 1596991774
transform 1 0 7384 0 1 1410
box -4 -6 20 206
use NAND2X1  _2201_
timestamp 1596991774
transform -1 0 56 0 -1 1810
box -4 -6 52 206
use NOR2X1  _2198_
timestamp 1596991774
transform 1 0 56 0 -1 1810
box -4 -6 52 206
use AOI21X1  _2197_
timestamp 1596991774
transform -1 0 168 0 -1 1810
box -4 -6 68 206
use NAND2X1  _2193_
timestamp 1596991774
transform 1 0 168 0 -1 1810
box -4 -6 52 206
use NOR2X1  _2207_
timestamp 1596991774
transform 1 0 216 0 -1 1810
box -4 -6 52 206
use AOI21X1  _2215_
timestamp 1596991774
transform 1 0 264 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2211_
timestamp 1596991774
transform -1 0 376 0 -1 1810
box -4 -6 52 206
use NOR2X1  _2210_
timestamp 1596991774
transform 1 0 376 0 -1 1810
box -4 -6 52 206
use AND2X2  _2209_
timestamp 1596991774
transform -1 0 488 0 -1 1810
box -4 -6 68 206
use XNOR2X1  _2277_
timestamp 1596991774
transform -1 0 600 0 -1 1810
box -4 -6 116 206
use NOR2X1  _2314_
timestamp 1596991774
transform 1 0 600 0 -1 1810
box -4 -6 52 206
use AND2X2  _2195_
timestamp 1596991774
transform 1 0 648 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3163_
timestamp 1596991774
transform 1 0 712 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3168_
timestamp 1596991774
transform 1 0 760 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3142_
timestamp 1596991774
transform -1 0 888 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3137_
timestamp 1596991774
transform -1 0 936 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3116_
timestamp 1596991774
transform -1 0 1000 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3111_
timestamp 1596991774
transform -1 0 1048 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3118_
timestamp 1596991774
transform 1 0 1048 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert154
timestamp 1596991774
transform -1 0 1160 0 -1 1810
box -4 -6 52 206
use AOI22X1  _3145_
timestamp 1596991774
transform 1 0 1160 0 -1 1810
box -4 -6 84 206
use AND2X2  _2361_
timestamp 1596991774
transform -1 0 1304 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3170_
timestamp 1596991774
transform -1 0 1368 0 -1 1810
box -4 -6 68 206
use AOI22X1  _3171_
timestamp 1596991774
transform -1 0 1448 0 -1 1810
box -4 -6 84 206
use BUFX2  BUFX2_insert240
timestamp 1596991774
transform 1 0 1512 0 -1 1810
box -4 -6 52 206
use AND2X2  _2975_
timestamp 1596991774
transform -1 0 1624 0 -1 1810
box -4 -6 68 206
use FILL  SFILL14480x16100
timestamp 1596991774
transform -1 0 1464 0 -1 1810
box -4 -6 20 206
use FILL  SFILL14640x16100
timestamp 1596991774
transform -1 0 1480 0 -1 1810
box -4 -6 20 206
use FILL  SFILL14800x16100
timestamp 1596991774
transform -1 0 1496 0 -1 1810
box -4 -6 20 206
use FILL  SFILL14960x16100
timestamp 1596991774
transform -1 0 1512 0 -1 1810
box -4 -6 20 206
use NOR2X1  _2977_
timestamp 1596991774
transform -1 0 1672 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3010_
timestamp 1596991774
transform -1 0 1736 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3062_
timestamp 1596991774
transform -1 0 1800 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3036_
timestamp 1596991774
transform -1 0 1864 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert231
timestamp 1596991774
transform 1 0 1864 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3035_
timestamp 1596991774
transform -1 0 1976 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3061_
timestamp 1596991774
transform -1 0 2040 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3009_
timestamp 1596991774
transform -1 0 2104 0 -1 1810
box -4 -6 68 206
use XNOR2X1  _2179_
timestamp 1596991774
transform -1 0 2216 0 -1 1810
box -4 -6 116 206
use NAND3X1  _3040_
timestamp 1596991774
transform 1 0 2216 0 -1 1810
box -4 -6 68 206
use INVX1  _3516_
timestamp 1596991774
transform 1 0 2280 0 -1 1810
box -4 -6 36 206
use NAND3X1  _3068_
timestamp 1596991774
transform 1 0 2312 0 -1 1810
box -4 -6 68 206
use AOI22X1  _3067_
timestamp 1596991774
transform -1 0 2456 0 -1 1810
box -4 -6 84 206
use NOR2X1  _2178_
timestamp 1596991774
transform -1 0 2504 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3065_
timestamp 1596991774
transform -1 0 2552 0 -1 1810
box -4 -6 52 206
use XNOR2X1  _2169_
timestamp 1596991774
transform 1 0 2552 0 -1 1810
box -4 -6 116 206
use OAI21X1  _2170_
timestamp 1596991774
transform 1 0 2664 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2168_
timestamp 1596991774
transform 1 0 2728 0 -1 1810
box -4 -6 52 206
use INVX1  _2795_
timestamp 1596991774
transform 1 0 2776 0 -1 1810
box -4 -6 36 206
use INVX1  _2166_
timestamp 1596991774
transform -1 0 2840 0 -1 1810
box -4 -6 36 206
use NAND2X1  _2165_
timestamp 1596991774
transform -1 0 2888 0 -1 1810
box -4 -6 52 206
use INVX1  _2792_
timestamp 1596991774
transform -1 0 2920 0 -1 1810
box -4 -6 36 206
use OR2X2  _2415_
timestamp 1596991774
transform 1 0 2984 0 -1 1810
box -4 -6 68 206
use FILL  SFILL29200x16100
timestamp 1596991774
transform -1 0 2936 0 -1 1810
box -4 -6 20 206
use FILL  SFILL29360x16100
timestamp 1596991774
transform -1 0 2952 0 -1 1810
box -4 -6 20 206
use FILL  SFILL29520x16100
timestamp 1596991774
transform -1 0 2968 0 -1 1810
box -4 -6 20 206
use FILL  SFILL29680x16100
timestamp 1596991774
transform -1 0 2984 0 -1 1810
box -4 -6 20 206
use AOI22X1  _2416_
timestamp 1596991774
transform 1 0 3048 0 -1 1810
box -4 -6 84 206
use NAND2X1  _2414_
timestamp 1596991774
transform -1 0 3176 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert299
timestamp 1596991774
transform 1 0 3176 0 -1 1810
box -4 -6 52 206
use NAND2X1  _2412_
timestamp 1596991774
transform 1 0 3224 0 -1 1810
box -4 -6 52 206
use XNOR2X1  _2934_
timestamp 1596991774
transform 1 0 3272 0 -1 1810
box -4 -6 116 206
use AND2X2  _2396_
timestamp 1596991774
transform -1 0 3448 0 -1 1810
box -4 -6 68 206
use AOI21X1  _2909_
timestamp 1596991774
transform 1 0 3448 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2905_
timestamp 1596991774
transform 1 0 3512 0 -1 1810
box -4 -6 52 206
use INVX1  _2904_
timestamp 1596991774
transform 1 0 3560 0 -1 1810
box -4 -6 36 206
use NAND2X1  _2908_
timestamp 1596991774
transform -1 0 3640 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert287
timestamp 1596991774
transform 1 0 3640 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert296
timestamp 1596991774
transform 1 0 3688 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert301
timestamp 1596991774
transform 1 0 3736 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _4429_
timestamp 1596991774
transform -1 0 3976 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_insert165
timestamp 1596991774
transform 1 0 3976 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert216
timestamp 1596991774
transform -1 0 4072 0 -1 1810
box -4 -6 52 206
use INVX1  _3426_
timestamp 1596991774
transform -1 0 4104 0 -1 1810
box -4 -6 36 206
use OAI21X1  _4122_
timestamp 1596991774
transform 1 0 4104 0 -1 1810
box -4 -6 68 206
use AOI21X1  _4123_
timestamp 1596991774
transform -1 0 4232 0 -1 1810
box -4 -6 68 206
use NOR2X1  _3434_
timestamp 1596991774
transform 1 0 4232 0 -1 1810
box -4 -6 52 206
use INVX1  _3433_
timestamp 1596991774
transform -1 0 4312 0 -1 1810
box -4 -6 36 206
use BUFX2  BUFX2_insert217
timestamp 1596991774
transform 1 0 4312 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert293
timestamp 1596991774
transform -1 0 4408 0 -1 1810
box -4 -6 52 206
use FILL  SFILL44080x16100
timestamp 1596991774
transform -1 0 4424 0 -1 1810
box -4 -6 20 206
use BUFX2  BUFX2_insert295
timestamp 1596991774
transform 1 0 4472 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3534_
timestamp 1596991774
transform -1 0 4584 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3535_
timestamp 1596991774
transform -1 0 4632 0 -1 1810
box -4 -6 52 206
use FILL  SFILL44240x16100
timestamp 1596991774
transform -1 0 4440 0 -1 1810
box -4 -6 20 206
use FILL  SFILL44400x16100
timestamp 1596991774
transform -1 0 4456 0 -1 1810
box -4 -6 20 206
use FILL  SFILL44560x16100
timestamp 1596991774
transform -1 0 4472 0 -1 1810
box -4 -6 20 206
use OAI21X1  _3430_
timestamp 1596991774
transform -1 0 4696 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3541_
timestamp 1596991774
transform -1 0 4760 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3542_
timestamp 1596991774
transform -1 0 4808 0 -1 1810
box -4 -6 52 206
use INVX8  _3567_
timestamp 1596991774
transform 1 0 4808 0 -1 1810
box -4 -6 84 206
use NAND3X1  _3492_
timestamp 1596991774
transform 1 0 4888 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3493_
timestamp 1596991774
transform -1 0 5000 0 -1 1810
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert15
timestamp 1596991774
transform -1 0 5144 0 -1 1810
box -4 -6 148 206
use NAND2X1  _3584_
timestamp 1596991774
transform 1 0 5144 0 -1 1810
box -4 -6 52 206
use AOI21X1  _3586_
timestamp 1596991774
transform 1 0 5192 0 -1 1810
box -4 -6 68 206
use AOI21X1  _3574_
timestamp 1596991774
transform -1 0 5320 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3436_
timestamp 1596991774
transform -1 0 5384 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3449_
timestamp 1596991774
transform -1 0 5448 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert203
timestamp 1596991774
transform -1 0 5496 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3437_
timestamp 1596991774
transform 1 0 5496 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3536_
timestamp 1596991774
transform -1 0 5592 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3522_
timestamp 1596991774
transform 1 0 5592 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3529_
timestamp 1596991774
transform 1 0 5640 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3501_
timestamp 1596991774
transform 1 0 5688 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert200
timestamp 1596991774
transform 1 0 5736 0 -1 1810
box -4 -6 52 206
use AOI21X1  _3580_
timestamp 1596991774
transform -1 0 5848 0 -1 1810
box -4 -6 68 206
use AOI21X1  _3623_
timestamp 1596991774
transform -1 0 5912 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3622_
timestamp 1596991774
transform -1 0 6024 0 -1 1810
box -4 -6 52 206
use FILL  SFILL59120x16100
timestamp 1596991774
transform -1 0 5928 0 -1 1810
box -4 -6 20 206
use FILL  SFILL59280x16100
timestamp 1596991774
transform -1 0 5944 0 -1 1810
box -4 -6 20 206
use FILL  SFILL59440x16100
timestamp 1596991774
transform -1 0 5960 0 -1 1810
box -4 -6 20 206
use FILL  SFILL59600x16100
timestamp 1596991774
transform -1 0 5976 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  _3636_
timestamp 1596991774
transform 1 0 6024 0 -1 1810
box -4 -6 196 206
use NAND2X1  _3451_
timestamp 1596991774
transform -1 0 6264 0 -1 1810
box -4 -6 52 206
use INVX1  _3448_
timestamp 1596991774
transform -1 0 6296 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  _3646_
timestamp 1596991774
transform -1 0 6488 0 -1 1810
box -4 -6 196 206
use AOI21X1  _3583_
timestamp 1596991774
transform -1 0 6552 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3581_
timestamp 1596991774
transform -1 0 6600 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _4381_
timestamp 1596991774
transform 1 0 6600 0 -1 1810
box -4 -6 196 206
use DFFPOSX1  _4382_
timestamp 1596991774
transform -1 0 6984 0 -1 1810
box -4 -6 196 206
use DFFPOSX1  _3632_
timestamp 1596991774
transform 1 0 6984 0 -1 1810
box -4 -6 196 206
use NAND2X1  _3614_
timestamp 1596991774
transform -1 0 7224 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3787_
timestamp 1596991774
transform -1 0 7272 0 -1 1810
box -4 -6 52 206
use AOI21X1  _3615_
timestamp 1596991774
transform 1 0 7272 0 -1 1810
box -4 -6 68 206
use NOR2X1  _4511_
timestamp 1596991774
transform 1 0 7336 0 -1 1810
box -4 -6 52 206
use FILL  FILL71280x16100
timestamp 1596991774
transform -1 0 7400 0 -1 1810
box -4 -6 20 206
use NOR2X1  _2214_
timestamp 1596991774
transform 1 0 8 0 1 1810
box -4 -6 52 206
use OAI21X1  _2202_
timestamp 1596991774
transform 1 0 56 0 1 1810
box -4 -6 68 206
use OAI21X1  _2216_
timestamp 1596991774
transform 1 0 120 0 1 1810
box -4 -6 68 206
use NAND2X1  _2213_
timestamp 1596991774
transform -1 0 232 0 1 1810
box -4 -6 52 206
use AOI21X1  _2208_
timestamp 1596991774
transform 1 0 232 0 1 1810
box -4 -6 68 206
use XNOR2X1  _2212_
timestamp 1596991774
transform 1 0 296 0 1 1810
box -4 -6 116 206
use NOR2X1  _2278_
timestamp 1596991774
transform 1 0 408 0 1 1810
box -4 -6 52 206
use XNOR2X1  _2204_
timestamp 1596991774
transform -1 0 568 0 1 1810
box -4 -6 116 206
use NAND3X1  _3165_
timestamp 1596991774
transform 1 0 568 0 1 1810
box -4 -6 68 206
use NAND3X1  _3139_
timestamp 1596991774
transform 1 0 632 0 1 1810
box -4 -6 68 206
use AND2X2  _3167_
timestamp 1596991774
transform 1 0 696 0 1 1810
box -4 -6 68 206
use AND2X2  _3141_
timestamp 1596991774
transform -1 0 824 0 1 1810
box -4 -6 68 206
use AND2X2  _3115_
timestamp 1596991774
transform -1 0 888 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert215
timestamp 1596991774
transform 1 0 888 0 1 1810
box -4 -6 52 206
use NAND2X1  _2951_
timestamp 1596991774
transform -1 0 984 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert229
timestamp 1596991774
transform 1 0 984 0 1 1810
box -4 -6 52 206
use NOR2X1  _3095_
timestamp 1596991774
transform 1 0 1032 0 1 1810
box -4 -6 52 206
use NAND3X1  _3092_
timestamp 1596991774
transform -1 0 1144 0 1 1810
box -4 -6 68 206
use NAND3X1  _3094_
timestamp 1596991774
transform 1 0 1144 0 1 1810
box -4 -6 68 206
use NAND2X1  _3091_
timestamp 1596991774
transform -1 0 1256 0 1 1810
box -4 -6 52 206
use AOI22X1  _3093_
timestamp 1596991774
transform -1 0 1336 0 1 1810
box -4 -6 84 206
use NAND2X1  _2957_
timestamp 1596991774
transform -1 0 1384 0 1 1810
box -4 -6 52 206
use NAND2X1  _3368_
timestamp 1596991774
transform 1 0 1384 0 1 1810
box -4 -6 52 206
use INVX1  _3367_
timestamp 1596991774
transform 1 0 1496 0 1 1810
box -4 -6 36 206
use OAI21X1  _3369_
timestamp 1596991774
transform 1 0 1528 0 1 1810
box -4 -6 68 206
use AND2X2  _2974_
timestamp 1596991774
transform -1 0 1656 0 1 1810
box -4 -6 68 206
use FILL  SFILL14320x18100
timestamp 1596991774
transform 1 0 1432 0 1 1810
box -4 -6 20 206
use FILL  SFILL14480x18100
timestamp 1596991774
transform 1 0 1448 0 1 1810
box -4 -6 20 206
use FILL  SFILL14640x18100
timestamp 1596991774
transform 1 0 1464 0 1 1810
box -4 -6 20 206
use FILL  SFILL14800x18100
timestamp 1596991774
transform 1 0 1480 0 1 1810
box -4 -6 20 206
use NAND2X1  _2964_
timestamp 1596991774
transform 1 0 1656 0 1 1810
box -4 -6 52 206
use NOR2X1  _3370_
timestamp 1596991774
transform -1 0 1752 0 1 1810
box -4 -6 52 206
use NAND2X1  _2971_
timestamp 1596991774
transform 1 0 1752 0 1 1810
box -4 -6 52 206
use NOR2X1  _2950_
timestamp 1596991774
transform -1 0 1848 0 1 1810
box -4 -6 52 206
use INVX1  _2946_
timestamp 1596991774
transform -1 0 1880 0 1 1810
box -4 -6 36 206
use NAND2X1  _2947_
timestamp 1596991774
transform -1 0 1928 0 1 1810
box -4 -6 52 206
use INVX1  _2948_
timestamp 1596991774
transform 1 0 1928 0 1 1810
box -4 -6 36 206
use NAND2X1  _2949_
timestamp 1596991774
transform -1 0 2008 0 1 1810
box -4 -6 52 206
use NAND2X1  _2956_
timestamp 1596991774
transform -1 0 2056 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert214
timestamp 1596991774
transform -1 0 2104 0 1 1810
box -4 -6 52 206
use NAND3X1  _2180_
timestamp 1596991774
transform -1 0 2168 0 1 1810
box -4 -6 68 206
use XOR2X1  _2174_
timestamp 1596991774
transform -1 0 2280 0 1 1810
box -4 -6 116 206
use AOI21X1  _2175_
timestamp 1596991774
transform 1 0 2280 0 1 1810
box -4 -6 68 206
use NOR2X1  _2173_
timestamp 1596991774
transform -1 0 2392 0 1 1810
box -4 -6 52 206
use AOI21X1  _2182_
timestamp 1596991774
transform 1 0 2392 0 1 1810
box -4 -6 68 206
use INVX1  _2181_
timestamp 1596991774
transform -1 0 2488 0 1 1810
box -4 -6 36 206
use AND2X2  _2176_
timestamp 1596991774
transform -1 0 2552 0 1 1810
box -4 -6 68 206
use NOR2X1  _2177_
timestamp 1596991774
transform -1 0 2600 0 1 1810
box -4 -6 52 206
use AND2X2  _2360_
timestamp 1596991774
transform -1 0 2664 0 1 1810
box -4 -6 68 206
use NAND2X1  _2164_
timestamp 1596991774
transform -1 0 2712 0 1 1810
box -4 -6 52 206
use NOR2X1  _2172_
timestamp 1596991774
transform 1 0 2712 0 1 1810
box -4 -6 52 206
use AND2X2  _2171_
timestamp 1596991774
transform -1 0 2824 0 1 1810
box -4 -6 68 206
use INVX1  _2941_
timestamp 1596991774
transform -1 0 2856 0 1 1810
box -4 -6 36 206
use OR2X2  _2341_
timestamp 1596991774
transform -1 0 2920 0 1 1810
box -4 -6 68 206
use XOR2X1  _2380_
timestamp 1596991774
transform 1 0 2984 0 1 1810
box -4 -6 116 206
use FILL  SFILL29200x18100
timestamp 1596991774
transform 1 0 2920 0 1 1810
box -4 -6 20 206
use FILL  SFILL29360x18100
timestamp 1596991774
transform 1 0 2936 0 1 1810
box -4 -6 20 206
use FILL  SFILL29520x18100
timestamp 1596991774
transform 1 0 2952 0 1 1810
box -4 -6 20 206
use FILL  SFILL29680x18100
timestamp 1596991774
transform 1 0 2968 0 1 1810
box -4 -6 20 206
use INVX1  _2906_
timestamp 1596991774
transform 1 0 3096 0 1 1810
box -4 -6 36 206
use NAND2X1  _2907_
timestamp 1596991774
transform 1 0 3128 0 1 1810
box -4 -6 52 206
use XNOR2X1  _2408_
timestamp 1596991774
transform -1 0 3288 0 1 1810
box -4 -6 116 206
use NOR2X1  _2397_
timestamp 1596991774
transform -1 0 3336 0 1 1810
box -4 -6 52 206
use OAI22X1  _2398_
timestamp 1596991774
transform -1 0 3416 0 1 1810
box -4 -6 84 206
use NOR2X1  _2395_
timestamp 1596991774
transform 1 0 3416 0 1 1810
box -4 -6 52 206
use AND2X2  _2394_
timestamp 1596991774
transform -1 0 3528 0 1 1810
box -4 -6 68 206
use OAI21X1  _3977_
timestamp 1596991774
transform 1 0 3528 0 1 1810
box -4 -6 68 206
use AOI21X1  _3978_
timestamp 1596991774
transform -1 0 3656 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert55
timestamp 1596991774
transform 1 0 3656 0 1 1810
box -4 -6 52 206
use OAI21X1  _3944_
timestamp 1596991774
transform 1 0 3704 0 1 1810
box -4 -6 68 206
use OAI21X1  _4111_
timestamp 1596991774
transform 1 0 3768 0 1 1810
box -4 -6 68 206
use AOI21X1  _4112_
timestamp 1596991774
transform -1 0 3896 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _4446_
timestamp 1596991774
transform -1 0 4088 0 1 1810
box -4 -6 196 206
use AOI21X1  _3945_
timestamp 1596991774
transform -1 0 4152 0 1 1810
box -4 -6 68 206
use INVX1  _3920_
timestamp 1596991774
transform 1 0 4152 0 1 1810
box -4 -6 36 206
use NOR2X1  _3921_
timestamp 1596991774
transform -1 0 4232 0 1 1810
box -4 -6 52 206
use NAND3X1  _3653_
timestamp 1596991774
transform -1 0 4296 0 1 1810
box -4 -6 68 206
use OAI21X1  _3933_
timestamp 1596991774
transform 1 0 4296 0 1 1810
box -4 -6 68 206
use AOI21X1  _3934_
timestamp 1596991774
transform -1 0 4424 0 1 1810
box -4 -6 68 206
use OAI21X1  _3531_
timestamp 1596991774
transform -1 0 4552 0 1 1810
box -4 -6 68 206
use OAI21X1  _3489_
timestamp 1596991774
transform -1 0 4616 0 1 1810
box -4 -6 68 206
use OAI21X1  _3538_
timestamp 1596991774
transform -1 0 4680 0 1 1810
box -4 -6 68 206
use FILL  SFILL44240x18100
timestamp 1596991774
transform 1 0 4424 0 1 1810
box -4 -6 20 206
use FILL  SFILL44400x18100
timestamp 1596991774
transform 1 0 4440 0 1 1810
box -4 -6 20 206
use FILL  SFILL44560x18100
timestamp 1596991774
transform 1 0 4456 0 1 1810
box -4 -6 20 206
use FILL  SFILL44720x18100
timestamp 1596991774
transform 1 0 4472 0 1 1810
box -4 -6 20 206
use NAND3X1  _3527_
timestamp 1596991774
transform -1 0 4744 0 1 1810
box -4 -6 68 206
use OAI21X1  _4155_
timestamp 1596991774
transform 1 0 4744 0 1 1810
box -4 -6 68 206
use AOI21X1  _4156_
timestamp 1596991774
transform -1 0 4872 0 1 1810
box -4 -6 68 206
use INVX8  _3909_
timestamp 1596991774
transform 1 0 4872 0 1 1810
box -4 -6 84 206
use INVX4  _3679_
timestamp 1596991774
transform 1 0 4952 0 1 1810
box -4 -6 52 206
use INVX8  _4089_
timestamp 1596991774
transform -1 0 5080 0 1 1810
box -4 -6 84 206
use DFFPOSX1  _3647_
timestamp 1596991774
transform -1 0 5272 0 1 1810
box -4 -6 196 206
use NAND2X1  _3572_
timestamp 1596991774
transform 1 0 5272 0 1 1810
box -4 -6 52 206
use NAND3X1  _3505_
timestamp 1596991774
transform -1 0 5384 0 1 1810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert11
timestamp 1596991774
transform -1 0 5528 0 1 1810
box -4 -6 148 206
use DFFPOSX1  _3645_
timestamp 1596991774
transform -1 0 5720 0 1 1810
box -4 -6 196 206
use DFFPOSX1  _4317_
timestamp 1596991774
transform 1 0 5720 0 1 1810
box -4 -6 196 206
use NAND2X1  _3578_
timestamp 1596991774
transform -1 0 6024 0 1 1810
box -4 -6 52 206
use FILL  SFILL59120x18100
timestamp 1596991774
transform 1 0 5912 0 1 1810
box -4 -6 20 206
use FILL  SFILL59280x18100
timestamp 1596991774
transform 1 0 5928 0 1 1810
box -4 -6 20 206
use FILL  SFILL59440x18100
timestamp 1596991774
transform 1 0 5944 0 1 1810
box -4 -6 20 206
use FILL  SFILL59600x18100
timestamp 1596991774
transform 1 0 5960 0 1 1810
box -4 -6 20 206
use BUFX2  BUFX2_insert211
timestamp 1596991774
transform 1 0 6024 0 1 1810
box -4 -6 52 206
use OAI21X1  _3746_
timestamp 1596991774
transform 1 0 6072 0 1 1810
box -4 -6 68 206
use NAND2X1  _3745_
timestamp 1596991774
transform -1 0 6184 0 1 1810
box -4 -6 52 206
use INVX4  _3670_
timestamp 1596991774
transform 1 0 6184 0 1 1810
box -4 -6 52 206
use INVX4  _3661_
timestamp 1596991774
transform 1 0 6232 0 1 1810
box -4 -6 52 206
use MUX2X1  _4113_
timestamp 1596991774
transform -1 0 6376 0 1 1810
box -4 -6 100 206
use MUX2X1  _3935_
timestamp 1596991774
transform -1 0 6472 0 1 1810
box -4 -6 100 206
use NOR2X1  _3812_
timestamp 1596991774
transform -1 0 6520 0 1 1810
box -4 -6 52 206
use AOI21X1  _3813_
timestamp 1596991774
transform -1 0 6584 0 1 1810
box -4 -6 68 206
use NOR2X1  _3814_
timestamp 1596991774
transform 1 0 6584 0 1 1810
box -4 -6 52 206
use AOI21X1  _3815_
timestamp 1596991774
transform -1 0 6696 0 1 1810
box -4 -6 68 206
use OAI21X1  _3782_
timestamp 1596991774
transform 1 0 6696 0 1 1810
box -4 -6 68 206
use NAND2X1  _3781_
timestamp 1596991774
transform -1 0 6808 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _4350_
timestamp 1596991774
transform -1 0 7000 0 1 1810
box -4 -6 196 206
use INVX1  _3504_
timestamp 1596991774
transform -1 0 7032 0 1 1810
box -4 -6 36 206
use NAND2X1  _3590_
timestamp 1596991774
transform 1 0 7032 0 1 1810
box -4 -6 52 206
use NAND2X1  _3591_
timestamp 1596991774
transform 1 0 7080 0 1 1810
box -4 -6 52 206
use AOI21X1  _3592_
timestamp 1596991774
transform 1 0 7128 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _3643_
timestamp 1596991774
transform -1 0 7384 0 1 1810
box -4 -6 196 206
use FILL  FILL71280x18100
timestamp 1596991774
transform 1 0 7384 0 1 1810
box -4 -6 20 206
use AOI21X1  _2217_
timestamp 1596991774
transform 1 0 8 0 -1 2210
box -4 -6 68 206
use OAI21X1  _2190_
timestamp 1596991774
transform 1 0 72 0 -1 2210
box -4 -6 68 206
use INVX1  _2188_
timestamp 1596991774
transform -1 0 168 0 -1 2210
box -4 -6 36 206
use XNOR2X1  _2194_
timestamp 1596991774
transform 1 0 168 0 -1 2210
box -4 -6 116 206
use NOR2X1  _2276_
timestamp 1596991774
transform -1 0 328 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2279_
timestamp 1596991774
transform 1 0 328 0 -1 2210
box -4 -6 52 206
use AOI21X1  _2280_
timestamp 1596991774
transform 1 0 376 0 -1 2210
box -4 -6 68 206
use NAND2X1  _2183_
timestamp 1596991774
transform -1 0 488 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3085_
timestamp 1596991774
transform 1 0 488 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3090_
timestamp 1596991774
transform 1 0 536 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3113_
timestamp 1596991774
transform 1 0 600 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3166_
timestamp 1596991774
transform -1 0 728 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3140_
timestamp 1596991774
transform 1 0 728 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3114_
timestamp 1596991774
transform -1 0 856 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert49
timestamp 1596991774
transform -1 0 904 0 -1 2210
box -4 -6 52 206
use INVX1  _3260_
timestamp 1596991774
transform 1 0 904 0 -1 2210
box -4 -6 36 206
use OAI22X1  _3262_
timestamp 1596991774
transform 1 0 936 0 -1 2210
box -4 -6 84 206
use INVX1  _3261_
timestamp 1596991774
transform -1 0 1048 0 -1 2210
box -4 -6 36 206
use NAND2X1  _3238_
timestamp 1596991774
transform -1 0 1096 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3212_
timestamp 1596991774
transform -1 0 1144 0 -1 2210
box -4 -6 52 206
use INVX1  _3509_
timestamp 1596991774
transform 1 0 1144 0 -1 2210
box -4 -6 36 206
use INVX1  _3183_
timestamp 1596991774
transform 1 0 1176 0 -1 2210
box -4 -6 36 206
use OAI22X1  _3184_
timestamp 1596991774
transform -1 0 1288 0 -1 2210
box -4 -6 84 206
use INVX1  _3182_
timestamp 1596991774
transform -1 0 1320 0 -1 2210
box -4 -6 36 206
use NAND2X1  _3316_
timestamp 1596991774
transform 1 0 1320 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3186_
timestamp 1596991774
transform -1 0 1416 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert108
timestamp 1596991774
transform -1 0 1528 0 -1 2210
box -4 -6 52 206
use INVX1  _3488_
timestamp 1596991774
transform 1 0 1528 0 -1 2210
box -4 -6 36 206
use BUFX2  BUFX2_insert274
timestamp 1596991774
transform 1 0 1560 0 -1 2210
box -4 -6 52 206
use NOR3X1  _2988_
timestamp 1596991774
transform -1 0 1736 0 -1 2210
box -4 -6 132 206
use FILL  SFILL14160x20100
timestamp 1596991774
transform -1 0 1432 0 -1 2210
box -4 -6 20 206
use FILL  SFILL14320x20100
timestamp 1596991774
transform -1 0 1448 0 -1 2210
box -4 -6 20 206
use FILL  SFILL14480x20100
timestamp 1596991774
transform -1 0 1464 0 -1 2210
box -4 -6 20 206
use FILL  SFILL14640x20100
timestamp 1596991774
transform -1 0 1480 0 -1 2210
box -4 -6 20 206
use NAND2X1  _2828_
timestamp 1596991774
transform -1 0 1784 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert51
timestamp 1596991774
transform 1 0 1784 0 -1 2210
box -4 -6 52 206
use NOR2X1  _2968_
timestamp 1596991774
transform 1 0 1832 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2967_
timestamp 1596991774
transform -1 0 1928 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2963_
timestamp 1596991774
transform 1 0 1928 0 -1 2210
box -4 -6 52 206
use AND2X2  _2970_
timestamp 1596991774
transform -1 0 2040 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert110
timestamp 1596991774
transform 1 0 2040 0 -1 2210
box -4 -6 52 206
use INVX8  _2945_
timestamp 1596991774
transform -1 0 2168 0 -1 2210
box -4 -6 84 206
use NOR2X1  _2984_
timestamp 1596991774
transform 1 0 2168 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2983_
timestamp 1596991774
transform -1 0 2264 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3066_
timestamp 1596991774
transform -1 0 2328 0 -1 2210
box -4 -6 68 206
use AOI22X1  _3301_
timestamp 1596991774
transform -1 0 2408 0 -1 2210
box -4 -6 84 206
use NAND3X1  _2992_
timestamp 1596991774
transform -1 0 2472 0 -1 2210
box -4 -6 68 206
use INVX1  _2942_
timestamp 1596991774
transform 1 0 2472 0 -1 2210
box -4 -6 36 206
use NOR2X1  _2959_
timestamp 1596991774
transform 1 0 2504 0 -1 2210
box -4 -6 52 206
use OAI22X1  _2952_
timestamp 1596991774
transform -1 0 2632 0 -1 2210
box -4 -6 84 206
use NOR2X1  _2293_
timestamp 1596991774
transform 1 0 2632 0 -1 2210
box -4 -6 52 206
use XOR2X1  _2435_
timestamp 1596991774
transform 1 0 2680 0 -1 2210
box -4 -6 116 206
use XOR2X1  _2379_
timestamp 1596991774
transform -1 0 2904 0 -1 2210
box -4 -6 116 206
use BUFX2  BUFX2_insert94
timestamp 1596991774
transform -1 0 3016 0 -1 2210
box -4 -6 52 206
use FILL  SFILL29040x20100
timestamp 1596991774
transform -1 0 2920 0 -1 2210
box -4 -6 20 206
use FILL  SFILL29200x20100
timestamp 1596991774
transform -1 0 2936 0 -1 2210
box -4 -6 20 206
use FILL  SFILL29360x20100
timestamp 1596991774
transform -1 0 2952 0 -1 2210
box -4 -6 20 206
use FILL  SFILL29520x20100
timestamp 1596991774
transform -1 0 2968 0 -1 2210
box -4 -6 20 206
use INVX1  _3523_
timestamp 1596991774
transform 1 0 3016 0 -1 2210
box -4 -6 36 206
use BUFX2  BUFX2_insert268
timestamp 1596991774
transform -1 0 3096 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert259
timestamp 1596991774
transform -1 0 3144 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2409_
timestamp 1596991774
transform -1 0 3192 0 -1 2210
box -4 -6 52 206
use XNOR2X1  _2407_
timestamp 1596991774
transform 1 0 3192 0 -1 2210
box -4 -6 116 206
use DFFPOSX1  _4447_
timestamp 1596991774
transform -1 0 3496 0 -1 2210
box -4 -6 196 206
use OAI21X1  _3955_
timestamp 1596991774
transform 1 0 3496 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert81
timestamp 1596991774
transform -1 0 3608 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4431_
timestamp 1596991774
transform -1 0 3800 0 -1 2210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert12
timestamp 1596991774
transform 1 0 3800 0 -1 2210
box -4 -6 148 206
use OAI21X1  _3510_
timestamp 1596991774
transform -1 0 4008 0 -1 2210
box -4 -6 68 206
use NOR2X1  _3432_
timestamp 1596991774
transform 1 0 4008 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4445_
timestamp 1596991774
transform -1 0 4248 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  _4341_
timestamp 1596991774
transform 1 0 4248 0 -1 2210
box -4 -6 196 206
use OAI21X1  _3496_
timestamp 1596991774
transform -1 0 4568 0 -1 2210
box -4 -6 68 206
use INVX1  _3537_
timestamp 1596991774
transform 1 0 4568 0 -1 2210
box -4 -6 36 206
use OAI21X1  _3524_
timestamp 1596991774
transform -1 0 4664 0 -1 2210
box -4 -6 68 206
use FILL  SFILL44400x20100
timestamp 1596991774
transform -1 0 4456 0 -1 2210
box -4 -6 20 206
use FILL  SFILL44560x20100
timestamp 1596991774
transform -1 0 4472 0 -1 2210
box -4 -6 20 206
use FILL  SFILL44720x20100
timestamp 1596991774
transform -1 0 4488 0 -1 2210
box -4 -6 20 206
use FILL  SFILL44880x20100
timestamp 1596991774
transform -1 0 4504 0 -1 2210
box -4 -6 20 206
use OAI21X1  _3503_
timestamp 1596991774
transform 1 0 4664 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert284
timestamp 1596991774
transform -1 0 4776 0 -1 2210
box -4 -6 52 206
use INVX4  _3664_
timestamp 1596991774
transform -1 0 4824 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3528_
timestamp 1596991774
transform -1 0 4872 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _3649_
timestamp 1596991774
transform -1 0 5064 0 -1 2210
box -4 -6 196 206
use NAND3X1  _3513_
timestamp 1596991774
transform 1 0 5064 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3512_
timestamp 1596991774
transform 1 0 5128 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3506_
timestamp 1596991774
transform -1 0 5256 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3507_
timestamp 1596991774
transform -1 0 5304 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3499_
timestamp 1596991774
transform 1 0 5304 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3500_
timestamp 1596991774
transform -1 0 5416 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3498_
timestamp 1596991774
transform -1 0 5480 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3514_
timestamp 1596991774
transform -1 0 5528 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert279
timestamp 1596991774
transform 1 0 5528 0 -1 2210
box -4 -6 52 206
use MUX2X1  _3943_
timestamp 1596991774
transform 1 0 5576 0 -1 2210
box -4 -6 100 206
use DFFPOSX1  _4389_
timestamp 1596991774
transform -1 0 5864 0 -1 2210
box -4 -6 196 206
use OAI22X1  _4116_
timestamp 1596991774
transform 1 0 5864 0 -1 2210
box -4 -6 84 206
use MUX2X1  _4121_
timestamp 1596991774
transform 1 0 6008 0 -1 2210
box -4 -6 100 206
use FILL  SFILL59440x20100
timestamp 1596991774
transform -1 0 5960 0 -1 2210
box -4 -6 20 206
use FILL  SFILL59600x20100
timestamp 1596991774
transform -1 0 5976 0 -1 2210
box -4 -6 20 206
use FILL  SFILL59760x20100
timestamp 1596991774
transform -1 0 5992 0 -1 2210
box -4 -6 20 206
use FILL  SFILL59920x20100
timestamp 1596991774
transform -1 0 6008 0 -1 2210
box -4 -6 20 206
use MUX2X1  _3932_
timestamp 1596991774
transform 1 0 6104 0 -1 2210
box -4 -6 100 206
use OAI21X1  _3926_
timestamp 1596991774
transform 1 0 6200 0 -1 2210
box -4 -6 68 206
use OAI22X1  _3927_
timestamp 1596991774
transform 1 0 6264 0 -1 2210
box -4 -6 84 206
use MUX2X1  _4110_
timestamp 1596991774
transform 1 0 6344 0 -1 2210
box -4 -6 100 206
use OAI21X1  _4104_
timestamp 1596991774
transform 1 0 6440 0 -1 2210
box -4 -6 68 206
use OAI22X1  _4105_
timestamp 1596991774
transform 1 0 6504 0 -1 2210
box -4 -6 84 206
use BUFX2  BUFX2_insert119
timestamp 1596991774
transform -1 0 6632 0 -1 2210
box -4 -6 52 206
use MUX2X1  _4102_
timestamp 1596991774
transform -1 0 6728 0 -1 2210
box -4 -6 100 206
use MUX2X1  _3924_
timestamp 1596991774
transform 1 0 6728 0 -1 2210
box -4 -6 100 206
use INVX1  _3497_
timestamp 1596991774
transform -1 0 6856 0 -1 2210
box -4 -6 36 206
use OAI21X1  _3780_
timestamp 1596991774
transform 1 0 6856 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3779_
timestamp 1596991774
transform -1 0 6968 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4349_
timestamp 1596991774
transform -1 0 7160 0 -1 2210
box -4 -6 196 206
use NAND2X1  _3569_
timestamp 1596991774
transform 1 0 7160 0 -1 2210
box -4 -6 52 206
use AOI21X1  _3571_
timestamp 1596991774
transform 1 0 7208 0 -1 2210
box -4 -6 68 206
use AOI21X1  _3595_
timestamp 1596991774
transform -1 0 7336 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3593_
timestamp 1596991774
transform -1 0 7384 0 -1 2210
box -4 -6 52 206
use FILL  FILL71280x20100
timestamp 1596991774
transform -1 0 7400 0 -1 2210
box -4 -6 20 206
use NOR2X1  _2189_
timestamp 1596991774
transform 1 0 8 0 1 2210
box -4 -6 52 206
use NAND2X1  _2184_
timestamp 1596991774
transform -1 0 104 0 1 2210
box -4 -6 52 206
use NAND2X1  _2186_
timestamp 1596991774
transform 1 0 104 0 1 2210
box -4 -6 52 206
use OR2X2  _2185_
timestamp 1596991774
transform -1 0 216 0 1 2210
box -4 -6 68 206
use XNOR2X1  _2187_
timestamp 1596991774
transform 1 0 216 0 1 2210
box -4 -6 116 206
use NAND3X1  _3087_
timestamp 1596991774
transform 1 0 328 0 1 2210
box -4 -6 68 206
use AND2X2  _3089_
timestamp 1596991774
transform 1 0 392 0 1 2210
box -4 -6 68 206
use NAND3X1  _3088_
timestamp 1596991774
transform 1 0 456 0 1 2210
box -4 -6 68 206
use OAI21X1  _2543_
timestamp 1596991774
transform -1 0 584 0 1 2210
box -4 -6 68 206
use NAND3X1  _3192_
timestamp 1596991774
transform 1 0 584 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert241
timestamp 1596991774
transform 1 0 648 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert276
timestamp 1596991774
transform -1 0 744 0 1 2210
box -4 -6 52 206
use NOR2X1  _3266_
timestamp 1596991774
transform 1 0 744 0 1 2210
box -4 -6 52 206
use INVX1  _3263_
timestamp 1596991774
transform 1 0 792 0 1 2210
box -4 -6 36 206
use OAI21X1  _3265_
timestamp 1596991774
transform 1 0 824 0 1 2210
box -4 -6 68 206
use NAND2X1  _3264_
timestamp 1596991774
transform -1 0 936 0 1 2210
box -4 -6 52 206
use NAND3X1  _3200_
timestamp 1596991774
transform -1 0 1000 0 1 2210
box -4 -6 68 206
use INVX1  _3211_
timestamp 1596991774
transform 1 0 1000 0 1 2210
box -4 -6 36 206
use OAI21X1  _3213_
timestamp 1596991774
transform 1 0 1032 0 1 2210
box -4 -6 68 206
use NOR2X1  _3188_
timestamp 1596991774
transform -1 0 1144 0 1 2210
box -4 -6 52 206
use OAI21X1  _3187_
timestamp 1596991774
transform -1 0 1208 0 1 2210
box -4 -6 68 206
use INVX1  _3185_
timestamp 1596991774
transform -1 0 1240 0 1 2210
box -4 -6 36 206
use INVX1  _3315_
timestamp 1596991774
transform 1 0 1240 0 1 2210
box -4 -6 36 206
use OAI21X1  _3317_
timestamp 1596991774
transform 1 0 1272 0 1 2210
box -4 -6 68 206
use INVX1  _2961_
timestamp 1596991774
transform 1 0 1336 0 1 2210
box -4 -6 36 206
use OAI22X1  _2965_
timestamp 1596991774
transform -1 0 1448 0 1 2210
box -4 -6 84 206
use INVX1  _2960_
timestamp 1596991774
transform -1 0 1544 0 1 2210
box -4 -6 36 206
use NOR2X1  _2973_
timestamp 1596991774
transform 1 0 1544 0 1 2210
box -4 -6 52 206
use OAI21X1  _2972_
timestamp 1596991774
transform -1 0 1656 0 1 2210
box -4 -6 68 206
use FILL  SFILL14480x22100
timestamp 1596991774
transform 1 0 1448 0 1 2210
box -4 -6 20 206
use FILL  SFILL14640x22100
timestamp 1596991774
transform 1 0 1464 0 1 2210
box -4 -6 20 206
use FILL  SFILL14800x22100
timestamp 1596991774
transform 1 0 1480 0 1 2210
box -4 -6 20 206
use FILL  SFILL14960x22100
timestamp 1596991774
transform 1 0 1496 0 1 2210
box -4 -6 20 206
use INVX1  _2966_
timestamp 1596991774
transform -1 0 1688 0 1 2210
box -4 -6 36 206
use AOI22X1  _2846_
timestamp 1596991774
transform -1 0 1768 0 1 2210
box -4 -6 84 206
use BUFX2  BUFX2_insert228
timestamp 1596991774
transform -1 0 1816 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert277
timestamp 1596991774
transform 1 0 1816 0 1 2210
box -4 -6 52 206
use NOR2X1  _2962_
timestamp 1596991774
transform -1 0 1912 0 1 2210
box -4 -6 52 206
use NOR2X1  _2955_
timestamp 1596991774
transform 1 0 1912 0 1 2210
box -4 -6 52 206
use INVX1  _2943_
timestamp 1596991774
transform 1 0 1960 0 1 2210
box -4 -6 36 206
use NOR3X1  _2987_
timestamp 1596991774
transform -1 0 2120 0 1 2210
box -4 -6 132 206
use NAND2X1  _2944_
timestamp 1596991774
transform 1 0 2120 0 1 2210
box -4 -6 52 206
use NOR2X1  _2991_
timestamp 1596991774
transform 1 0 2168 0 1 2210
box -4 -6 52 206
use NAND3X1  _3302_
timestamp 1596991774
transform 1 0 2216 0 1 2210
box -4 -6 68 206
use NAND3X1  _2387_
timestamp 1596991774
transform 1 0 2280 0 1 2210
box -4 -6 68 206
use NAND2X1  _3299_
timestamp 1596991774
transform -1 0 2392 0 1 2210
box -4 -6 52 206
use OAI22X1  _2958_
timestamp 1596991774
transform -1 0 2472 0 1 2210
box -4 -6 84 206
use INVX1  _2953_
timestamp 1596991774
transform -1 0 2504 0 1 2210
box -4 -6 36 206
use NOR2X1  _2295_
timestamp 1596991774
transform -1 0 2552 0 1 2210
box -4 -6 52 206
use AND2X2  _2294_
timestamp 1596991774
transform -1 0 2616 0 1 2210
box -4 -6 68 206
use AND2X2  _2369_
timestamp 1596991774
transform -1 0 2680 0 1 2210
box -4 -6 68 206
use XNOR2X1  _2422_
timestamp 1596991774
transform 1 0 2680 0 1 2210
box -4 -6 116 206
use NOR3X1  _2386_
timestamp 1596991774
transform 1 0 2792 0 1 2210
box -4 -6 132 206
use BUFX2  BUFX2_insert95
timestamp 1596991774
transform -1 0 3032 0 1 2210
box -4 -6 52 206
use FILL  SFILL29200x22100
timestamp 1596991774
transform 1 0 2920 0 1 2210
box -4 -6 20 206
use FILL  SFILL29360x22100
timestamp 1596991774
transform 1 0 2936 0 1 2210
box -4 -6 20 206
use FILL  SFILL29520x22100
timestamp 1596991774
transform 1 0 2952 0 1 2210
box -4 -6 20 206
use FILL  SFILL29680x22100
timestamp 1596991774
transform 1 0 2968 0 1 2210
box -4 -6 20 206
use BUFX2  BUFX2_insert155
timestamp 1596991774
transform 1 0 3032 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert265
timestamp 1596991774
transform 1 0 3080 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _4428_
timestamp 1596991774
transform -1 0 3320 0 1 2210
box -4 -6 196 206
use OAI21X1  _4100_
timestamp 1596991774
transform 1 0 3320 0 1 2210
box -4 -6 68 206
use AOI21X1  _4101_
timestamp 1596991774
transform -1 0 3448 0 1 2210
box -4 -6 68 206
use AOI21X1  _3956_
timestamp 1596991774
transform 1 0 3448 0 1 2210
box -4 -6 68 206
use OAI21X1  _4133_
timestamp 1596991774
transform 1 0 3512 0 1 2210
box -4 -6 68 206
use AOI21X1  _4134_
timestamp 1596991774
transform -1 0 3640 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert221
timestamp 1596991774
transform -1 0 3688 0 1 2210
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert14
timestamp 1596991774
transform -1 0 3832 0 1 2210
box -4 -6 148 206
use BUFX2  BUFX2_insert220
timestamp 1596991774
transform -1 0 3880 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _4355_
timestamp 1596991774
transform 1 0 3880 0 1 2210
box -4 -6 196 206
use OAI21X1  _3792_
timestamp 1596991774
transform 1 0 4072 0 1 2210
box -4 -6 68 206
use NAND2X1  _3791_
timestamp 1596991774
transform -1 0 4184 0 1 2210
box -4 -6 52 206
use INVX4  _3700_
timestamp 1596991774
transform -1 0 4232 0 1 2210
box -4 -6 52 206
use AOI21X1  _3896_
timestamp 1596991774
transform 1 0 4232 0 1 2210
box -4 -6 68 206
use NOR2X1  _3895_
timestamp 1596991774
transform -1 0 4344 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _4323_
timestamp 1596991774
transform 1 0 4408 0 1 2210
box -4 -6 196 206
use FILL  SFILL43440x22100
timestamp 1596991774
transform 1 0 4344 0 1 2210
box -4 -6 20 206
use FILL  SFILL43600x22100
timestamp 1596991774
transform 1 0 4360 0 1 2210
box -4 -6 20 206
use FILL  SFILL43760x22100
timestamp 1596991774
transform 1 0 4376 0 1 2210
box -4 -6 20 206
use FILL  SFILL43920x22100
timestamp 1596991774
transform 1 0 4392 0 1 2210
box -4 -6 20 206
use NAND2X1  _3757_
timestamp 1596991774
transform 1 0 4600 0 1 2210
box -4 -6 52 206
use OAI21X1  _3758_
timestamp 1596991774
transform -1 0 4712 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4339_
timestamp 1596991774
transform -1 0 4904 0 1 2210
box -4 -6 196 206
use OAI21X1  _4174_
timestamp 1596991774
transform 1 0 4904 0 1 2210
box -4 -6 68 206
use NOR2X1  _3891_
timestamp 1596991774
transform 1 0 4968 0 1 2210
box -4 -6 52 206
use AOI21X1  _3892_
timestamp 1596991774
transform -1 0 5080 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert204
timestamp 1596991774
transform -1 0 5128 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert122
timestamp 1596991774
transform 1 0 5128 0 1 2210
box -4 -6 52 206
use INVX4  _3685_
timestamp 1596991774
transform -1 0 5224 0 1 2210
box -4 -6 52 206
use OAI21X1  _4115_
timestamp 1596991774
transform -1 0 5288 0 1 2210
box -4 -6 68 206
use INVX4  _3682_
timestamp 1596991774
transform -1 0 5336 0 1 2210
box -4 -6 52 206
use NOR2X1  _3828_
timestamp 1596991774
transform 1 0 5336 0 1 2210
box -4 -6 52 206
use AOI21X1  _3829_
timestamp 1596991774
transform 1 0 5384 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert73
timestamp 1596991774
transform 1 0 5448 0 1 2210
box -4 -6 52 206
use OAI21X1  _3937_
timestamp 1596991774
transform 1 0 5496 0 1 2210
box -4 -6 68 206
use OAI22X1  _3938_
timestamp 1596991774
transform 1 0 5560 0 1 2210
box -4 -6 84 206
use NOR2X1  _3936_
timestamp 1596991774
transform -1 0 5688 0 1 2210
box -4 -6 52 206
use OAI21X1  _3941_
timestamp 1596991774
transform -1 0 5752 0 1 2210
box -4 -6 68 206
use OAI22X1  _3942_
timestamp 1596991774
transform 1 0 5752 0 1 2210
box -4 -6 84 206
use NOR2X1  _4114_
timestamp 1596991774
transform 1 0 5832 0 1 2210
box -4 -6 52 206
use OAI21X1  _4119_
timestamp 1596991774
transform 1 0 5880 0 1 2210
box -4 -6 68 206
use OAI22X1  _4120_
timestamp 1596991774
transform 1 0 6008 0 1 2210
box -4 -6 84 206
use FILL  SFILL59440x22100
timestamp 1596991774
transform 1 0 5944 0 1 2210
box -4 -6 20 206
use FILL  SFILL59600x22100
timestamp 1596991774
transform 1 0 5960 0 1 2210
box -4 -6 20 206
use FILL  SFILL59760x22100
timestamp 1596991774
transform 1 0 5976 0 1 2210
box -4 -6 20 206
use FILL  SFILL59920x22100
timestamp 1596991774
transform 1 0 5992 0 1 2210
box -4 -6 20 206
use DFFPOSX1  _4366_
timestamp 1596991774
transform -1 0 6280 0 1 2210
box -4 -6 196 206
use NOR2X1  _3925_
timestamp 1596991774
transform -1 0 6328 0 1 2210
box -4 -6 52 206
use MUX2X1  _4117_
timestamp 1596991774
transform -1 0 6424 0 1 2210
box -4 -6 100 206
use MUX2X1  _3939_
timestamp 1596991774
transform -1 0 6520 0 1 2210
box -4 -6 100 206
use NOR2X1  _4103_
timestamp 1596991774
transform -1 0 6568 0 1 2210
box -4 -6 52 206
use NOR2X1  _4272_
timestamp 1596991774
transform 1 0 6568 0 1 2210
box -4 -6 52 206
use AOI21X1  _4273_
timestamp 1596991774
transform -1 0 6680 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4414_
timestamp 1596991774
transform -1 0 6872 0 1 2210
box -4 -6 196 206
use DFFPOSX1  _3648_
timestamp 1596991774
transform -1 0 7064 0 1 2210
box -4 -6 196 206
use DFFPOSX1  _3644_
timestamp 1596991774
transform -1 0 7256 0 1 2210
box -4 -6 196 206
use NAND2X1  _3594_
timestamp 1596991774
transform 1 0 7256 0 1 2210
box -4 -6 52 206
use AOI21X1  _3589_
timestamp 1596991774
transform -1 0 7368 0 1 2210
box -4 -6 68 206
use FILL  FILL71120x22100
timestamp 1596991774
transform 1 0 7368 0 1 2210
box -4 -6 20 206
use FILL  FILL71280x22100
timestamp 1596991774
transform 1 0 7384 0 1 2210
box -4 -6 20 206
use AND2X2  _2306_
timestamp 1596991774
transform -1 0 72 0 -1 2610
box -4 -6 68 206
use NOR2X1  _2307_
timestamp 1596991774
transform -1 0 120 0 -1 2610
box -4 -6 52 206
use NOR2X1  _2305_
timestamp 1596991774
transform -1 0 168 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert290
timestamp 1596991774
transform -1 0 216 0 -1 2610
box -4 -6 52 206
use NAND3X1  _3191_
timestamp 1596991774
transform 1 0 216 0 -1 2610
box -4 -6 68 206
use NAND3X1  _3086_
timestamp 1596991774
transform 1 0 280 0 -1 2610
box -4 -6 68 206
use AND2X2  _3193_
timestamp 1596991774
transform 1 0 344 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert233
timestamp 1596991774
transform -1 0 456 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert212
timestamp 1596991774
transform 1 0 456 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert242
timestamp 1596991774
transform -1 0 552 0 -1 2610
box -4 -6 52 206
use INVX1  _3235_
timestamp 1596991774
transform 1 0 552 0 -1 2610
box -4 -6 36 206
use INVX1  _3234_
timestamp 1596991774
transform 1 0 584 0 -1 2610
box -4 -6 36 206
use OAI22X1  _3236_
timestamp 1596991774
transform -1 0 696 0 -1 2610
box -4 -6 84 206
use NAND3X1  _3278_
timestamp 1596991774
transform -1 0 760 0 -1 2610
box -4 -6 68 206
use NOR2X1  _3240_
timestamp 1596991774
transform 1 0 760 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3239_
timestamp 1596991774
transform 1 0 808 0 -1 2610
box -4 -6 68 206
use INVX1  _3208_
timestamp 1596991774
transform 1 0 872 0 -1 2610
box -4 -6 36 206
use OAI22X1  _3210_
timestamp 1596991774
transform 1 0 904 0 -1 2610
box -4 -6 84 206
use INVX1  _3209_
timestamp 1596991774
transform -1 0 1016 0 -1 2610
box -4 -6 36 206
use NOR2X1  _3214_
timestamp 1596991774
transform 1 0 1016 0 -1 2610
box -4 -6 52 206
use INVX1  _3313_
timestamp 1596991774
transform 1 0 1064 0 -1 2610
box -4 -6 36 206
use OAI22X1  _3314_
timestamp 1596991774
transform -1 0 1176 0 -1 2610
box -4 -6 84 206
use INVX1  _3312_
timestamp 1596991774
transform -1 0 1208 0 -1 2610
box -4 -6 36 206
use NOR2X1  _3318_
timestamp 1596991774
transform -1 0 1256 0 -1 2610
box -4 -6 52 206
use INVX1  _3341_
timestamp 1596991774
transform 1 0 1256 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3343_
timestamp 1596991774
transform 1 0 1288 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3342_
timestamp 1596991774
transform -1 0 1400 0 -1 2610
box -4 -6 52 206
use FILL  SFILL14000x24100
timestamp 1596991774
transform -1 0 1416 0 -1 2610
box -4 -6 20 206
use NOR2X1  _3344_
timestamp 1596991774
transform -1 0 1512 0 -1 2610
box -4 -6 52 206
use NAND2X1  _2969_
timestamp 1596991774
transform 1 0 1512 0 -1 2610
box -4 -6 52 206
use INVX1  _3339_
timestamp 1596991774
transform 1 0 1560 0 -1 2610
box -4 -6 36 206
use OAI22X1  _3340_
timestamp 1596991774
transform -1 0 1672 0 -1 2610
box -4 -6 84 206
use FILL  SFILL14160x24100
timestamp 1596991774
transform -1 0 1432 0 -1 2610
box -4 -6 20 206
use FILL  SFILL14320x24100
timestamp 1596991774
transform -1 0 1448 0 -1 2610
box -4 -6 20 206
use FILL  SFILL14480x24100
timestamp 1596991774
transform -1 0 1464 0 -1 2610
box -4 -6 20 206
use INVX1  _3338_
timestamp 1596991774
transform -1 0 1704 0 -1 2610
box -4 -6 36 206
use BUFX2  BUFX2_insert213
timestamp 1596991774
transform 1 0 1704 0 -1 2610
box -4 -6 52 206
use NAND3X1  _3304_
timestamp 1596991774
transform 1 0 1752 0 -1 2610
box -4 -6 68 206
use NOR2X1  _3303_
timestamp 1596991774
transform 1 0 1816 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3371_
timestamp 1596991774
transform -1 0 1912 0 -1 2610
box -4 -6 52 206
use NAND2X1  _2976_
timestamp 1596991774
transform -1 0 1960 0 -1 2610
box -4 -6 52 206
use NAND3X1  _2982_
timestamp 1596991774
transform 1 0 1960 0 -1 2610
box -4 -6 68 206
use NAND3X1  _2978_
timestamp 1596991774
transform -1 0 2088 0 -1 2610
box -4 -6 68 206
use NAND3X1  _3300_
timestamp 1596991774
transform -1 0 2152 0 -1 2610
box -4 -6 68 206
use NAND3X1  _2990_
timestamp 1596991774
transform -1 0 2216 0 -1 2610
box -4 -6 68 206
use NAND2X1  _2985_
timestamp 1596991774
transform -1 0 2264 0 -1 2610
box -4 -6 52 206
use NAND3X1  _3382_
timestamp 1596991774
transform -1 0 2328 0 -1 2610
box -4 -6 68 206
use AND2X2  _2357_
timestamp 1596991774
transform -1 0 2392 0 -1 2610
box -4 -6 68 206
use INVX1  _2954_
timestamp 1596991774
transform -1 0 2424 0 -1 2610
box -4 -6 36 206
use XOR2X1  _2391_
timestamp 1596991774
transform -1 0 2536 0 -1 2610
box -4 -6 116 206
use XOR2X1  _2399_
timestamp 1596991774
transform 1 0 2536 0 -1 2610
box -4 -6 116 206
use NOR3X1  _2401_
timestamp 1596991774
transform 1 0 2648 0 -1 2610
box -4 -6 132 206
use XNOR2X1  _2423_
timestamp 1596991774
transform 1 0 2776 0 -1 2610
box -4 -6 116 206
use NAND2X1  _2424_
timestamp 1596991774
transform 1 0 2888 0 -1 2610
box -4 -6 52 206
use INVX1  _3495_
timestamp 1596991774
transform 1 0 3000 0 -1 2610
box -4 -6 36 206
use FILL  SFILL29360x24100
timestamp 1596991774
transform -1 0 2952 0 -1 2610
box -4 -6 20 206
use FILL  SFILL29520x24100
timestamp 1596991774
transform -1 0 2968 0 -1 2610
box -4 -6 20 206
use FILL  SFILL29680x24100
timestamp 1596991774
transform -1 0 2984 0 -1 2610
box -4 -6 20 206
use FILL  SFILL29840x24100
timestamp 1596991774
transform -1 0 3000 0 -1 2610
box -4 -6 20 206
use XNOR2X1  _2431_
timestamp 1596991774
transform 1 0 3032 0 -1 2610
box -4 -6 116 206
use DFFPOSX1  _4444_
timestamp 1596991774
transform -1 0 3336 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  _4432_
timestamp 1596991774
transform -1 0 3528 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_insert291
timestamp 1596991774
transform -1 0 3576 0 -1 2610
box -4 -6 52 206
use INVX1  _3530_
timestamp 1596991774
transform 1 0 3576 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  _4405_
timestamp 1596991774
transform 1 0 3608 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  _4387_
timestamp 1596991774
transform 1 0 3800 0 -1 2610
box -4 -6 196 206
use NOR2X1  _3824_
timestamp 1596991774
transform 1 0 3992 0 -1 2610
box -4 -6 52 206
use AOI21X1  _3825_
timestamp 1596991774
transform -1 0 4104 0 -1 2610
box -4 -6 68 206
use INVX1  _3502_
timestamp 1596991774
transform 1 0 4104 0 -1 2610
box -4 -6 36 206
use MUX2X1  _4168_
timestamp 1596991774
transform -1 0 4232 0 -1 2610
box -4 -6 100 206
use MUX2X1  _3990_
timestamp 1596991774
transform -1 0 4328 0 -1 2610
box -4 -6 100 206
use OAI21X1  _4196_
timestamp 1596991774
transform -1 0 4392 0 -1 2610
box -4 -6 68 206
use OAI21X1  _4018_
timestamp 1596991774
transform 1 0 4392 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3992_
timestamp 1596991774
transform -1 0 4584 0 -1 2610
box -4 -6 68 206
use OAI22X1  _3993_
timestamp 1596991774
transform -1 0 4664 0 -1 2610
box -4 -6 84 206
use FILL  SFILL44560x24100
timestamp 1596991774
transform -1 0 4472 0 -1 2610
box -4 -6 20 206
use FILL  SFILL44720x24100
timestamp 1596991774
transform -1 0 4488 0 -1 2610
box -4 -6 20 206
use FILL  SFILL44880x24100
timestamp 1596991774
transform -1 0 4504 0 -1 2610
box -4 -6 20 206
use FILL  SFILL45040x24100
timestamp 1596991774
transform -1 0 4520 0 -1 2610
box -4 -6 20 206
use MUX2X1  _3998_
timestamp 1596991774
transform 1 0 4664 0 -1 2610
box -4 -6 100 206
use OAI21X1  _4170_
timestamp 1596991774
transform 1 0 4760 0 -1 2610
box -4 -6 68 206
use OAI22X1  _4171_
timestamp 1596991774
transform -1 0 4904 0 -1 2610
box -4 -6 84 206
use OAI21X1  _3996_
timestamp 1596991774
transform -1 0 4968 0 -1 2610
box -4 -6 68 206
use MUX2X1  _4176_
timestamp 1596991774
transform 1 0 4968 0 -1 2610
box -4 -6 100 206
use OAI22X1  _4175_
timestamp 1596991774
transform 1 0 5064 0 -1 2610
box -4 -6 84 206
use MUX2X1  _4172_
timestamp 1596991774
transform -1 0 5240 0 -1 2610
box -4 -6 100 206
use DFFPOSX1  _4419_
timestamp 1596991774
transform -1 0 5432 0 -1 2610
box -4 -6 196 206
use OAI21X1  _4014_
timestamp 1596991774
transform 1 0 5432 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert76
timestamp 1596991774
transform -1 0 5544 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _4325_
timestamp 1596991774
transform -1 0 5736 0 -1 2610
box -4 -6 196 206
use NAND2X1  _3761_
timestamp 1596991774
transform 1 0 5736 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3762_
timestamp 1596991774
transform -1 0 5848 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4318_
timestamp 1596991774
transform 1 0 5912 0 -1 2610
box -4 -6 196 206
use FILL  SFILL58480x24100
timestamp 1596991774
transform -1 0 5864 0 -1 2610
box -4 -6 20 206
use FILL  SFILL58640x24100
timestamp 1596991774
transform -1 0 5880 0 -1 2610
box -4 -6 20 206
use FILL  SFILL58800x24100
timestamp 1596991774
transform -1 0 5896 0 -1 2610
box -4 -6 20 206
use FILL  SFILL58960x24100
timestamp 1596991774
transform -1 0 5912 0 -1 2610
box -4 -6 20 206
use NAND2X1  _3747_
timestamp 1596991774
transform 1 0 6104 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3748_
timestamp 1596991774
transform -1 0 6216 0 -1 2610
box -4 -6 68 206
use AOI21X1  _3880_
timestamp 1596991774
transform 1 0 6216 0 -1 2610
box -4 -6 68 206
use NOR2X1  _3879_
timestamp 1596991774
transform -1 0 6328 0 -1 2610
box -4 -6 52 206
use OAI21X1  _4108_
timestamp 1596991774
transform 1 0 6328 0 -1 2610
box -4 -6 68 206
use OAI22X1  _4109_
timestamp 1596991774
transform 1 0 6392 0 -1 2610
box -4 -6 84 206
use NOR2X1  _3940_
timestamp 1596991774
transform -1 0 6520 0 -1 2610
box -4 -6 52 206
use NOR2X1  _4118_
timestamp 1596991774
transform -1 0 6568 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3714_
timestamp 1596991774
transform -1 0 6632 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3715_
timestamp 1596991774
transform -1 0 6696 0 -1 2610
box -4 -6 68 206
use MUX2X1  _4106_
timestamp 1596991774
transform 1 0 6696 0 -1 2610
box -4 -6 100 206
use DFFPOSX1  _4398_
timestamp 1596991774
transform -1 0 6984 0 -1 2610
box -4 -6 196 206
use NOR2X1  _4270_
timestamp 1596991774
transform 1 0 6984 0 -1 2610
box -4 -6 52 206
use NOR2X1  _3659_
timestamp 1596991774
transform -1 0 7080 0 -1 2610
box -4 -6 52 206
use AOI21X1  _4271_
timestamp 1596991774
transform -1 0 7144 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3713_
timestamp 1596991774
transform 1 0 7144 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3712_
timestamp 1596991774
transform 1 0 7208 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3588_
timestamp 1596991774
transform 1 0 7272 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3587_
timestamp 1596991774
transform 1 0 7320 0 -1 2610
box -4 -6 52 206
use FILL  FILL71120x24100
timestamp 1596991774
transform -1 0 7384 0 -1 2610
box -4 -6 20 206
use FILL  FILL71280x24100
timestamp 1596991774
transform -1 0 7400 0 -1 2610
box -4 -6 20 206
use XNOR2X1  _2222_
timestamp 1596991774
transform 1 0 8 0 1 2610
box -4 -6 116 206
use OAI21X1  _2282_
timestamp 1596991774
transform -1 0 184 0 1 2610
box -4 -6 68 206
use NAND2X1  _3215_
timestamp 1596991774
transform 1 0 184 0 1 2610
box -4 -6 52 206
use NAND3X1  _3220_
timestamp 1596991774
transform 1 0 232 0 1 2610
box -4 -6 68 206
use AND2X2  _3219_
timestamp 1596991774
transform -1 0 360 0 1 2610
box -4 -6 68 206
use NAND3X1  _3218_
timestamp 1596991774
transform 1 0 360 0 1 2610
box -4 -6 68 206
use NAND3X1  _3270_
timestamp 1596991774
transform -1 0 488 0 1 2610
box -4 -6 68 206
use NAND3X1  _3244_
timestamp 1596991774
transform -1 0 552 0 1 2610
box -4 -6 68 206
use NAND3X1  _3194_
timestamp 1596991774
transform -1 0 616 0 1 2610
box -4 -6 68 206
use NAND2X1  _3189_
timestamp 1596991774
transform -1 0 664 0 1 2610
box -4 -6 52 206
use NOR2X1  _3277_
timestamp 1596991774
transform 1 0 664 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert275
timestamp 1596991774
transform -1 0 760 0 1 2610
box -4 -6 52 206
use NOR2X1  _3199_
timestamp 1596991774
transform 1 0 760 0 1 2610
box -4 -6 52 206
use INVX1  _3237_
timestamp 1596991774
transform -1 0 840 0 1 2610
box -4 -6 36 206
use BUFX2  BUFX2_insert52
timestamp 1596991774
transform -1 0 888 0 1 2610
box -4 -6 52 206
use AOI22X1  _3197_
timestamp 1596991774
transform -1 0 968 0 1 2610
box -4 -6 84 206
use NOR2X1  _3225_
timestamp 1596991774
transform 1 0 968 0 1 2610
box -4 -6 52 206
use NAND3X1  _3226_
timestamp 1596991774
transform -1 0 1080 0 1 2610
box -4 -6 68 206
use NAND3X1  _2980_
timestamp 1596991774
transform -1 0 1144 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert239
timestamp 1596991774
transform -1 0 1192 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert107
timestamp 1596991774
transform -1 0 1240 0 1 2610
box -4 -6 52 206
use NAND3X1  _3330_
timestamp 1596991774
transform 1 0 1240 0 1 2610
box -4 -6 68 206
use NOR2X1  _3329_
timestamp 1596991774
transform -1 0 1352 0 1 2610
box -4 -6 52 206
use NAND3X1  _3296_
timestamp 1596991774
transform 1 0 1352 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert50
timestamp 1596991774
transform -1 0 1528 0 1 2610
box -4 -6 52 206
use NAND3X1  _3322_
timestamp 1596991774
transform -1 0 1592 0 1 2610
box -4 -6 68 206
use NAND3X1  _3374_
timestamp 1596991774
transform -1 0 1656 0 1 2610
box -4 -6 68 206
use FILL  SFILL14160x26100
timestamp 1596991774
transform 1 0 1416 0 1 2610
box -4 -6 20 206
use FILL  SFILL14320x26100
timestamp 1596991774
transform 1 0 1432 0 1 2610
box -4 -6 20 206
use FILL  SFILL14480x26100
timestamp 1596991774
transform 1 0 1448 0 1 2610
box -4 -6 20 206
use FILL  SFILL14640x26100
timestamp 1596991774
transform 1 0 1464 0 1 2610
box -4 -6 20 206
use NAND3X1  _3348_
timestamp 1596991774
transform -1 0 1720 0 1 2610
box -4 -6 68 206
use AND2X2  _2981_
timestamp 1596991774
transform 1 0 1720 0 1 2610
box -4 -6 68 206
use NAND3X1  _2979_
timestamp 1596991774
transform -1 0 1848 0 1 2610
box -4 -6 68 206
use AND2X2  _3375_
timestamp 1596991774
transform 1 0 1848 0 1 2610
box -4 -6 68 206
use NAND3X1  _3376_
timestamp 1596991774
transform -1 0 1976 0 1 2610
box -4 -6 68 206
use NAND3X1  _3372_
timestamp 1596991774
transform -1 0 2040 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert109
timestamp 1596991774
transform 1 0 2040 0 1 2610
box -4 -6 52 206
use NAND3X1  _3352_
timestamp 1596991774
transform -1 0 2152 0 1 2610
box -4 -6 68 206
use NAND3X1  _2986_
timestamp 1596991774
transform -1 0 2216 0 1 2610
box -4 -6 68 206
use NAND3X1  _3378_
timestamp 1596991774
transform -1 0 2280 0 1 2610
box -4 -6 68 206
use NOR2X1  _3381_
timestamp 1596991774
transform 1 0 2280 0 1 2610
box -4 -6 52 206
use NOR2X1  _2403_
timestamp 1596991774
transform 1 0 2328 0 1 2610
box -4 -6 52 206
use XOR2X1  _2292_
timestamp 1596991774
transform -1 0 2488 0 1 2610
box -4 -6 116 206
use NAND3X1  _2402_
timestamp 1596991774
transform -1 0 2552 0 1 2610
box -4 -6 68 206
use NOR2X1  _2393_
timestamp 1596991774
transform 1 0 2552 0 1 2610
box -4 -6 52 206
use XOR2X1  _2392_
timestamp 1596991774
transform -1 0 2712 0 1 2610
box -4 -6 116 206
use XOR2X1  _2400_
timestamp 1596991774
transform 1 0 2712 0 1 2610
box -4 -6 116 206
use NAND2X1  _2434_
timestamp 1596991774
transform 1 0 2824 0 1 2610
box -4 -6 52 206
use NOR3X1  _2433_
timestamp 1596991774
transform -1 0 3064 0 1 2610
box -4 -6 132 206
use FILL  SFILL28720x26100
timestamp 1596991774
transform 1 0 2872 0 1 2610
box -4 -6 20 206
use FILL  SFILL28880x26100
timestamp 1596991774
transform 1 0 2888 0 1 2610
box -4 -6 20 206
use FILL  SFILL29040x26100
timestamp 1596991774
transform 1 0 2904 0 1 2610
box -4 -6 20 206
use FILL  SFILL29200x26100
timestamp 1596991774
transform 1 0 2920 0 1 2610
box -4 -6 20 206
use NAND3X1  _2432_
timestamp 1596991774
transform -1 0 3128 0 1 2610
box -4 -6 68 206
use XNOR2X1  _2430_
timestamp 1596991774
transform -1 0 3240 0 1 2610
box -4 -6 116 206
use OAI21X1  _3922_
timestamp 1596991774
transform 1 0 3240 0 1 2610
box -4 -6 68 206
use AOI21X1  _3923_
timestamp 1596991774
transform -1 0 3368 0 1 2610
box -4 -6 68 206
use OAI21X1  _4144_
timestamp 1596991774
transform 1 0 3368 0 1 2610
box -4 -6 68 206
use AOI21X1  _4145_
timestamp 1596991774
transform -1 0 3496 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4335_
timestamp 1596991774
transform -1 0 3688 0 1 2610
box -4 -6 196 206
use NOR2X1  _3683_
timestamp 1596991774
transform 1 0 3688 0 1 2610
box -4 -6 52 206
use AOI21X1  _3684_
timestamp 1596991774
transform -1 0 3800 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4309_
timestamp 1596991774
transform 1 0 3800 0 1 2610
box -4 -6 196 206
use NAND2X1  _3862_
timestamp 1596991774
transform 1 0 3992 0 1 2610
box -4 -6 52 206
use OAI21X1  _3863_
timestamp 1596991774
transform -1 0 4104 0 1 2610
box -4 -6 68 206
use MUX2X1  _4194_
timestamp 1596991774
transform -1 0 4200 0 1 2610
box -4 -6 100 206
use MUX2X1  _4016_
timestamp 1596991774
transform -1 0 4296 0 1 2610
box -4 -6 100 206
use OAI22X1  _4197_
timestamp 1596991774
transform -1 0 4376 0 1 2610
box -4 -6 84 206
use NOR2X1  _4195_
timestamp 1596991774
transform -1 0 4424 0 1 2610
box -4 -6 52 206
use NOR2X1  _4017_
timestamp 1596991774
transform 1 0 4488 0 1 2610
box -4 -6 52 206
use OAI22X1  _4019_
timestamp 1596991774
transform 1 0 4536 0 1 2610
box -4 -6 84 206
use NOR2X1  _3991_
timestamp 1596991774
transform 1 0 4616 0 1 2610
box -4 -6 52 206
use FILL  SFILL44240x26100
timestamp 1596991774
transform 1 0 4424 0 1 2610
box -4 -6 20 206
use FILL  SFILL44400x26100
timestamp 1596991774
transform 1 0 4440 0 1 2610
box -4 -6 20 206
use FILL  SFILL44560x26100
timestamp 1596991774
transform 1 0 4456 0 1 2610
box -4 -6 20 206
use FILL  SFILL44720x26100
timestamp 1596991774
transform 1 0 4472 0 1 2610
box -4 -6 20 206
use MUX2X1  _4020_
timestamp 1596991774
transform -1 0 4760 0 1 2610
box -4 -6 100 206
use NOR2X1  _4169_
timestamp 1596991774
transform 1 0 4760 0 1 2610
box -4 -6 52 206
use OAI22X1  _3997_
timestamp 1596991774
transform -1 0 4888 0 1 2610
box -4 -6 84 206
use NOR2X1  _3995_
timestamp 1596991774
transform -1 0 4936 0 1 2610
box -4 -6 52 206
use NOR2X1  _4173_
timestamp 1596991774
transform -1 0 4984 0 1 2610
box -4 -6 52 206
use MUX2X1  _3994_
timestamp 1596991774
transform -1 0 5080 0 1 2610
box -4 -6 100 206
use NOR2X1  _4013_
timestamp 1596991774
transform -1 0 5128 0 1 2610
box -4 -6 52 206
use OAI22X1  _4015_
timestamp 1596991774
transform 1 0 5128 0 1 2610
box -4 -6 84 206
use OAI21X1  _4192_
timestamp 1596991774
transform -1 0 5272 0 1 2610
box -4 -6 68 206
use NOR2X1  _4282_
timestamp 1596991774
transform 1 0 5272 0 1 2610
box -4 -6 52 206
use AOI21X1  _4283_
timestamp 1596991774
transform -1 0 5384 0 1 2610
box -4 -6 68 206
use MUX2X1  _4190_
timestamp 1596991774
transform 1 0 5384 0 1 2610
box -4 -6 100 206
use MUX2X1  _4012_
timestamp 1596991774
transform 1 0 5480 0 1 2610
box -4 -6 100 206
use DFFPOSX1  _4373_
timestamp 1596991774
transform -1 0 5768 0 1 2610
box -4 -6 196 206
use OAI21X1  _3729_
timestamp 1596991774
transform 1 0 5768 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4333_
timestamp 1596991774
transform 1 0 5832 0 1 2610
box -4 -6 196 206
use OAI21X1  _3930_
timestamp 1596991774
transform 1 0 6088 0 1 2610
box -4 -6 68 206
use OAI22X1  _3931_
timestamp 1596991774
transform 1 0 6152 0 1 2610
box -4 -6 84 206
use FILL  SFILL60240x26100
timestamp 1596991774
transform 1 0 6024 0 1 2610
box -4 -6 20 206
use FILL  SFILL60400x26100
timestamp 1596991774
transform 1 0 6040 0 1 2610
box -4 -6 20 206
use FILL  SFILL60560x26100
timestamp 1596991774
transform 1 0 6056 0 1 2610
box -4 -6 20 206
use FILL  SFILL60720x26100
timestamp 1596991774
transform 1 0 6072 0 1 2610
box -4 -6 20 206
use NOR2X1  _3881_
timestamp 1596991774
transform -1 0 6280 0 1 2610
box -4 -6 52 206
use AOI21X1  _3882_
timestamp 1596991774
transform 1 0 6280 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4334_
timestamp 1596991774
transform -1 0 6536 0 1 2610
box -4 -6 196 206
use BUFX2  BUFX2_insert143
timestamp 1596991774
transform -1 0 6584 0 1 2610
box -4 -6 52 206
use MUX2X1  _3928_
timestamp 1596991774
transform -1 0 6680 0 1 2610
box -4 -6 100 206
use AOI21X1  _3663_
timestamp 1596991774
transform 1 0 6680 0 1 2610
box -4 -6 68 206
use NOR2X1  _3662_
timestamp 1596991774
transform 1 0 6744 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _4413_
timestamp 1596991774
transform -1 0 6984 0 1 2610
box -4 -6 196 206
use DFFPOSX1  _4397_
timestamp 1596991774
transform -1 0 7176 0 1 2610
box -4 -6 196 206
use DFFPOSX1  _3642_
timestamp 1596991774
transform -1 0 7368 0 1 2610
box -4 -6 196 206
use FILL  FILL71120x26100
timestamp 1596991774
transform 1 0 7368 0 1 2610
box -4 -6 20 206
use FILL  FILL71280x26100
timestamp 1596991774
transform 1 0 7384 0 1 2610
box -4 -6 20 206
use NOR2X1  _2226_
timestamp 1596991774
transform 1 0 8 0 -1 3010
box -4 -6 52 206
use INVX1  _2225_
timestamp 1596991774
transform -1 0 88 0 -1 3010
box -4 -6 36 206
use NOR2X1  _2228_
timestamp 1596991774
transform -1 0 136 0 -1 3010
box -4 -6 52 206
use NOR2X1  _2227_
timestamp 1596991774
transform -1 0 184 0 -1 3010
box -4 -6 52 206
use NOR2X1  _2320_
timestamp 1596991774
transform -1 0 232 0 -1 3010
box -4 -6 52 206
use NOR2X1  _2322_
timestamp 1596991774
transform 1 0 232 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3216_
timestamp 1596991774
transform 1 0 280 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3217_
timestamp 1596991774
transform 1 0 344 0 -1 3010
box -4 -6 68 206
use AND2X2  _3271_
timestamp 1596991774
transform 1 0 408 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3272_
timestamp 1596991774
transform -1 0 536 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3267_
timestamp 1596991774
transform -1 0 584 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3190_
timestamp 1596991774
transform 1 0 584 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3274_
timestamp 1596991774
transform -1 0 712 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3276_
timestamp 1596991774
transform 1 0 712 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3196_
timestamp 1596991774
transform -1 0 840 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3198_
timestamp 1596991774
transform 1 0 840 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3252_
timestamp 1596991774
transform 1 0 904 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3275_
timestamp 1596991774
transform -1 0 1048 0 -1 3010
box -4 -6 84 206
use NAND3X1  _3224_
timestamp 1596991774
transform -1 0 1112 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3222_
timestamp 1596991774
transform 1 0 1112 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert232
timestamp 1596991774
transform -1 0 1224 0 -1 3010
box -4 -6 52 206
use AOI22X1  _3223_
timestamp 1596991774
transform -1 0 1304 0 -1 3010
box -4 -6 84 206
use NAND3X1  _3326_
timestamp 1596991774
transform -1 0 1368 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3328_
timestamp 1596991774
transform 1 0 1368 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3327_
timestamp 1596991774
transform -1 0 1576 0 -1 3010
box -4 -6 84 206
use AND2X2  _3323_
timestamp 1596991774
transform 1 0 1576 0 -1 3010
box -4 -6 68 206
use FILL  SFILL14320x28100
timestamp 1596991774
transform -1 0 1448 0 -1 3010
box -4 -6 20 206
use FILL  SFILL14480x28100
timestamp 1596991774
transform -1 0 1464 0 -1 3010
box -4 -6 20 206
use FILL  SFILL14640x28100
timestamp 1596991774
transform -1 0 1480 0 -1 3010
box -4 -6 20 206
use FILL  SFILL14800x28100
timestamp 1596991774
transform -1 0 1496 0 -1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert230
timestamp 1596991774
transform 1 0 1640 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3319_
timestamp 1596991774
transform 1 0 1688 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3324_
timestamp 1596991774
transform 1 0 1736 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3298_
timestamp 1596991774
transform -1 0 1864 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3373_
timestamp 1596991774
transform 1 0 1864 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3347_
timestamp 1596991774
transform 1 0 1928 0 -1 3010
box -4 -6 68 206
use AND2X2  _3349_
timestamp 1596991774
transform 1 0 1992 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3353_
timestamp 1596991774
transform 1 0 2056 0 -1 3010
box -4 -6 84 206
use NAND3X1  _3354_
timestamp 1596991774
transform 1 0 2136 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3355_
timestamp 1596991774
transform 1 0 2200 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3356_
timestamp 1596991774
transform -1 0 2312 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3380_
timestamp 1596991774
transform 1 0 2312 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3379_
timestamp 1596991774
transform -1 0 2456 0 -1 3010
box -4 -6 84 206
use OAI22X1  _3362_
timestamp 1596991774
transform 1 0 2456 0 -1 3010
box -4 -6 84 206
use INVX1  _3361_
timestamp 1596991774
transform -1 0 2568 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3377_
timestamp 1596991774
transform -1 0 2616 0 -1 3010
box -4 -6 52 206
use AND2X2  _2372_
timestamp 1596991774
transform -1 0 2680 0 -1 3010
box -4 -6 68 206
use XNOR2X1  _2410_
timestamp 1596991774
transform 1 0 2680 0 -1 3010
box -4 -6 116 206
use NAND3X1  _2417_
timestamp 1596991774
transform 1 0 2792 0 -1 3010
box -4 -6 68 206
use NOR3X1  _2418_
timestamp 1596991774
transform 1 0 2856 0 -1 3010
box -4 -6 132 206
use FILL  SFILL29840x28100
timestamp 1596991774
transform -1 0 3000 0 -1 3010
box -4 -6 20 206
use FILL  SFILL30000x28100
timestamp 1596991774
transform -1 0 3016 0 -1 3010
box -4 -6 20 206
use DFFPOSX1  _4448_
timestamp 1596991774
transform -1 0 3240 0 -1 3010
box -4 -6 196 206
use FILL  SFILL30160x28100
timestamp 1596991774
transform -1 0 3032 0 -1 3010
box -4 -6 20 206
use FILL  SFILL30320x28100
timestamp 1596991774
transform -1 0 3048 0 -1 3010
box -4 -6 20 206
use NAND2X1  _2427_
timestamp 1596991774
transform -1 0 3288 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3966_
timestamp 1596991774
transform 1 0 3288 0 -1 3010
box -4 -6 68 206
use AOI21X1  _3967_
timestamp 1596991774
transform -1 0 3416 0 -1 3010
box -4 -6 68 206
use OAI21X1  _4021_
timestamp 1596991774
transform 1 0 3416 0 -1 3010
box -4 -6 68 206
use AOI21X1  _4022_
timestamp 1596991774
transform -1 0 3544 0 -1 3010
box -4 -6 68 206
use OAI21X1  _4199_
timestamp 1596991774
transform -1 0 3608 0 -1 3010
box -4 -6 68 206
use AOI21X1  _4200_
timestamp 1596991774
transform -1 0 3672 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3883_
timestamp 1596991774
transform 1 0 3672 0 -1 3010
box -4 -6 52 206
use AOI21X1  _3884_
timestamp 1596991774
transform -1 0 3784 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _4388_
timestamp 1596991774
transform -1 0 3976 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  _4421_
timestamp 1596991774
transform 1 0 3976 0 -1 3010
box -4 -6 196 206
use NOR2X1  _4286_
timestamp 1596991774
transform 1 0 4168 0 -1 3010
box -4 -6 52 206
use AOI21X1  _4287_
timestamp 1596991774
transform -1 0 4280 0 -1 3010
box -4 -6 68 206
use MUX2X1  _4198_
timestamp 1596991774
transform -1 0 4376 0 -1 3010
box -4 -6 100 206
use FILL  SFILL43760x28100
timestamp 1596991774
transform -1 0 4392 0 -1 3010
box -4 -6 20 206
use FILL  SFILL43920x28100
timestamp 1596991774
transform -1 0 4408 0 -1 3010
box -4 -6 20 206
use FILL  SFILL44080x28100
timestamp 1596991774
transform -1 0 4424 0 -1 3010
box -4 -6 20 206
use DFFPOSX1  _4371_
timestamp 1596991774
transform 1 0 4440 0 -1 3010
box -4 -6 196 206
use FILL  SFILL44240x28100
timestamp 1596991774
transform -1 0 4440 0 -1 3010
box -4 -6 20 206
use OAI21X1  _3725_
timestamp 1596991774
transform 1 0 4632 0 -1 3010
box -4 -6 68 206
use OAI21X1  _3724_
timestamp 1596991774
transform 1 0 4696 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _4307_
timestamp 1596991774
transform 1 0 4760 0 -1 3010
box -4 -6 196 206
use NAND2X1  _3858_
timestamp 1596991774
transform 1 0 4952 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3859_
timestamp 1596991774
transform -1 0 5064 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert149
timestamp 1596991774
transform -1 0 5112 0 -1 3010
box -4 -6 52 206
use NOR2X1  _4191_
timestamp 1596991774
transform -1 0 5160 0 -1 3010
box -4 -6 52 206
use OAI22X1  _4193_
timestamp 1596991774
transform 1 0 5160 0 -1 3010
box -4 -6 84 206
use DFFPOSX1  _4403_
timestamp 1596991774
transform -1 0 5432 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  _4357_
timestamp 1596991774
transform -1 0 5624 0 -1 3010
box -4 -6 196 206
use NAND2X1  _3795_
timestamp 1596991774
transform 1 0 5624 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3796_
timestamp 1596991774
transform -1 0 5736 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert133
timestamp 1596991774
transform 1 0 5736 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3728_
timestamp 1596991774
transform -1 0 5848 0 -1 3010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert20
timestamp 1596991774
transform -1 0 5992 0 -1 3010
box -4 -6 148 206
use FILL  SFILL59920x28100
timestamp 1596991774
transform -1 0 6008 0 -1 3010
box -4 -6 20 206
use FILL  SFILL60080x28100
timestamp 1596991774
transform -1 0 6024 0 -1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert224
timestamp 1596991774
transform -1 0 6104 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3929_
timestamp 1596991774
transform -1 0 6152 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4301_
timestamp 1596991774
transform -1 0 6344 0 -1 3010
box -4 -6 196 206
use FILL  SFILL60240x28100
timestamp 1596991774
transform -1 0 6040 0 -1 3010
box -4 -6 20 206
use FILL  SFILL60400x28100
timestamp 1596991774
transform -1 0 6056 0 -1 3010
box -4 -6 20 206
use NOR2X1  _4107_
timestamp 1596991774
transform 1 0 6344 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3846_
timestamp 1596991774
transform 1 0 6392 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3847_
timestamp 1596991774
transform -1 0 6504 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert254
timestamp 1596991774
transform 1 0 6504 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3848_
timestamp 1596991774
transform -1 0 6600 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3849_
timestamp 1596991774
transform -1 0 6664 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _4302_
timestamp 1596991774
transform -1 0 6856 0 -1 3010
box -4 -6 196 206
use NAND2X1  _3742_
timestamp 1596991774
transform -1 0 6904 0 -1 3010
box -4 -6 52 206
use AND2X2  _4267_
timestamp 1596991774
transform -1 0 6968 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3707_
timestamp 1596991774
transform -1 0 7016 0 -1 3010
box -4 -6 52 206
use INVX1  _3706_
timestamp 1596991774
transform -1 0 7048 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3709_
timestamp 1596991774
transform -1 0 7096 0 -1 3010
box -4 -6 52 206
use INVX1  _3703_
timestamp 1596991774
transform -1 0 7128 0 -1 3010
box -4 -6 36 206
use BUFX2  BUFX2_insert152
timestamp 1596991774
transform 1 0 7128 0 -1 3010
box -4 -6 52 206
use AND2X2  _3655_
timestamp 1596991774
transform -1 0 7240 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3652_
timestamp 1596991774
transform -1 0 7288 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3654_
timestamp 1596991774
transform 1 0 7288 0 -1 3010
box -4 -6 52 206
use BUFX2  _2084_
timestamp 1596991774
transform 1 0 7336 0 -1 3010
box -4 -6 52 206
use FILL  FILL71280x28100
timestamp 1596991774
transform -1 0 7400 0 -1 3010
box -4 -6 20 206
use OAI21X1  _2231_
timestamp 1596991774
transform 1 0 8 0 1 3010
box -4 -6 68 206
use OAI21X1  _2230_
timestamp 1596991774
transform -1 0 136 0 1 3010
box -4 -6 68 206
use INVX1  _2224_
timestamp 1596991774
transform -1 0 168 0 1 3010
box -4 -6 36 206
use XOR2X1  _2229_
timestamp 1596991774
transform -1 0 280 0 1 3010
box -4 -6 116 206
use AND2X2  _2321_
timestamp 1596991774
transform -1 0 344 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert238
timestamp 1596991774
transform 1 0 344 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert58
timestamp 1596991774
transform -1 0 440 0 1 3010
box -4 -6 52 206
use NAND3X1  _3269_
timestamp 1596991774
transform 1 0 440 0 1 3010
box -4 -6 68 206
use NAND3X1  _3268_
timestamp 1596991774
transform 1 0 504 0 1 3010
box -4 -6 68 206
use AND2X2  _3245_
timestamp 1596991774
transform 1 0 568 0 1 3010
box -4 -6 68 206
use NAND3X1  _3242_
timestamp 1596991774
transform 1 0 632 0 1 3010
box -4 -6 68 206
use NAND2X1  _3273_
timestamp 1596991774
transform 1 0 696 0 1 3010
box -4 -6 52 206
use NAND3X1  _3246_
timestamp 1596991774
transform -1 0 808 0 1 3010
box -4 -6 68 206
use NAND2X1  _3241_
timestamp 1596991774
transform -1 0 856 0 1 3010
box -4 -6 52 206
use NAND2X1  _3195_
timestamp 1596991774
transform 1 0 856 0 1 3010
box -4 -6 52 206
use NOR2X1  _3251_
timestamp 1596991774
transform 1 0 904 0 1 3010
box -4 -6 52 206
use AND2X2  _2366_
timestamp 1596991774
transform 1 0 952 0 1 3010
box -4 -6 68 206
use NAND2X1  _3221_
timestamp 1596991774
transform 1 0 1016 0 1 3010
box -4 -6 52 206
use NAND3X1  _3248_
timestamp 1596991774
transform -1 0 1128 0 1 3010
box -4 -6 68 206
use NAND3X1  _3250_
timestamp 1596991774
transform 1 0 1128 0 1 3010
box -4 -6 68 206
use AOI22X1  _3249_
timestamp 1596991774
transform -1 0 1272 0 1 3010
box -4 -6 84 206
use NAND2X1  _3247_
timestamp 1596991774
transform -1 0 1320 0 1 3010
box -4 -6 52 206
use NAND2X1  _3325_
timestamp 1596991774
transform -1 0 1368 0 1 3010
box -4 -6 52 206
use AND2X2  _3297_
timestamp 1596991774
transform 1 0 1368 0 1 3010
box -4 -6 68 206
use OAI22X1  _3284_
timestamp 1596991774
transform 1 0 1496 0 1 3010
box -4 -6 84 206
use INVX1  _3283_
timestamp 1596991774
transform -1 0 1608 0 1 3010
box -4 -6 36 206
use XNOR2X1  _2275_
timestamp 1596991774
transform 1 0 1608 0 1 3010
box -4 -6 116 206
use FILL  SFILL14320x30100
timestamp 1596991774
transform 1 0 1432 0 1 3010
box -4 -6 20 206
use FILL  SFILL14480x30100
timestamp 1596991774
transform 1 0 1448 0 1 3010
box -4 -6 20 206
use FILL  SFILL14640x30100
timestamp 1596991774
transform 1 0 1464 0 1 3010
box -4 -6 20 206
use FILL  SFILL14800x30100
timestamp 1596991774
transform 1 0 1480 0 1 3010
box -4 -6 20 206
use NOR2X1  _3285_
timestamp 1596991774
transform 1 0 1720 0 1 3010
box -4 -6 52 206
use INVX1  _3279_
timestamp 1596991774
transform 1 0 1768 0 1 3010
box -4 -6 36 206
use OAI22X1  _3281_
timestamp 1596991774
transform 1 0 1800 0 1 3010
box -4 -6 84 206
use INVX1  _3280_
timestamp 1596991774
transform -1 0 1912 0 1 3010
box -4 -6 36 206
use NAND3X1  _3320_
timestamp 1596991774
transform 1 0 1912 0 1 3010
box -4 -6 68 206
use NAND2X1  _3293_
timestamp 1596991774
transform -1 0 2024 0 1 3010
box -4 -6 52 206
use NAND3X1  _3350_
timestamp 1596991774
transform -1 0 2088 0 1 3010
box -4 -6 68 206
use NAND2X1  _3345_
timestamp 1596991774
transform -1 0 2136 0 1 3010
box -4 -6 52 206
use AOI22X1  _2989_
timestamp 1596991774
transform 1 0 2136 0 1 3010
box -4 -6 84 206
use NAND2X1  _3351_
timestamp 1596991774
transform -1 0 2264 0 1 3010
box -4 -6 52 206
use AND2X2  _2371_
timestamp 1596991774
transform -1 0 2328 0 1 3010
box -4 -6 68 206
use OAI22X1  _3359_
timestamp 1596991774
transform 1 0 2328 0 1 3010
box -4 -6 84 206
use INVX1  _3358_
timestamp 1596991774
transform -1 0 2440 0 1 3010
box -4 -6 36 206
use NOR2X1  _3363_
timestamp 1596991774
transform -1 0 2488 0 1 3010
box -4 -6 52 206
use XNOR2X1  _2411_
timestamp 1596991774
transform 1 0 2488 0 1 3010
box -4 -6 116 206
use NOR2X1  _2384_
timestamp 1596991774
transform -1 0 2648 0 1 3010
box -4 -6 52 206
use AND2X2  _2383_
timestamp 1596991774
transform 1 0 2648 0 1 3010
box -4 -6 68 206
use OAI22X1  _2385_
timestamp 1596991774
transform -1 0 2792 0 1 3010
box -4 -6 84 206
use NOR2X1  _2382_
timestamp 1596991774
transform 1 0 2792 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert234
timestamp 1596991774
transform -1 0 2888 0 1 3010
box -4 -6 52 206
use NAND2X1  _2425_
timestamp 1596991774
transform 1 0 2888 0 1 3010
box -4 -6 52 206
use OR2X2  _2426_
timestamp 1596991774
transform 1 0 3000 0 1 3010
box -4 -6 68 206
use FILL  SFILL29360x30100
timestamp 1596991774
transform 1 0 2936 0 1 3010
box -4 -6 20 206
use FILL  SFILL29520x30100
timestamp 1596991774
transform 1 0 2952 0 1 3010
box -4 -6 20 206
use FILL  SFILL29680x30100
timestamp 1596991774
transform 1 0 2968 0 1 3010
box -4 -6 20 206
use FILL  SFILL29840x30100
timestamp 1596991774
transform 1 0 2984 0 1 3010
box -4 -6 20 206
use AOI22X1  _2429_
timestamp 1596991774
transform 1 0 3064 0 1 3010
box -4 -6 84 206
use OR2X2  _2428_
timestamp 1596991774
transform -1 0 3208 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert60
timestamp 1596991774
transform 1 0 3208 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4437_
timestamp 1596991774
transform -1 0 3448 0 1 3010
box -4 -6 196 206
use OAI22X1  _4131_
timestamp 1596991774
transform -1 0 3528 0 1 3010
box -4 -6 84 206
use OAI21X1  _4130_
timestamp 1596991774
transform -1 0 3592 0 1 3010
box -4 -6 68 206
use MUX2X1  _4132_
timestamp 1596991774
transform -1 0 3688 0 1 3010
box -4 -6 100 206
use NAND2X1  _3785_
timestamp 1596991774
transform 1 0 3688 0 1 3010
box -4 -6 52 206
use OAI21X1  _3786_
timestamp 1596991774
transform -1 0 3800 0 1 3010
box -4 -6 68 206
use NOR2X1  _4129_
timestamp 1596991774
transform 1 0 3800 0 1 3010
box -4 -6 52 206
use NOR2X1  _3826_
timestamp 1596991774
transform -1 0 3896 0 1 3010
box -4 -6 52 206
use AOI21X1  _3827_
timestamp 1596991774
transform -1 0 3960 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert25
timestamp 1596991774
transform -1 0 4008 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert142
timestamp 1596991774
transform 1 0 4008 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert91
timestamp 1596991774
transform -1 0 4104 0 1 3010
box -4 -6 52 206
use INVX4  _3697_
timestamp 1596991774
transform -1 0 4152 0 1 3010
box -4 -6 52 206
use OAI21X1  _3794_
timestamp 1596991774
transform 1 0 4152 0 1 3010
box -4 -6 68 206
use NAND2X1  _3793_
timestamp 1596991774
transform -1 0 4264 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4356_
timestamp 1596991774
transform 1 0 4264 0 1 3010
box -4 -6 196 206
use MUX2X1  _4179_
timestamp 1596991774
transform -1 0 4616 0 1 3010
box -4 -6 100 206
use MUX2X1  _4001_
timestamp 1596991774
transform -1 0 4712 0 1 3010
box -4 -6 100 206
use FILL  SFILL44560x30100
timestamp 1596991774
transform 1 0 4456 0 1 3010
box -4 -6 20 206
use FILL  SFILL44720x30100
timestamp 1596991774
transform 1 0 4472 0 1 3010
box -4 -6 20 206
use FILL  SFILL44880x30100
timestamp 1596991774
transform 1 0 4488 0 1 3010
box -4 -6 20 206
use FILL  SFILL45040x30100
timestamp 1596991774
transform 1 0 4504 0 1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert207
timestamp 1596991774
transform -1 0 4760 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert117
timestamp 1596991774
transform -1 0 4808 0 1 3010
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert18
timestamp 1596991774
transform -1 0 4952 0 1 3010
box -4 -6 148 206
use OAI21X1  _3853_
timestamp 1596991774
transform 1 0 4952 0 1 3010
box -4 -6 68 206
use NAND2X1  _3852_
timestamp 1596991774
transform -1 0 5064 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert101
timestamp 1596991774
transform -1 0 5112 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert63
timestamp 1596991774
transform -1 0 5160 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4304_
timestamp 1596991774
transform -1 0 5352 0 1 3010
box -4 -6 196 206
use AOI21X1  _3678_
timestamp 1596991774
transform 1 0 5352 0 1 3010
box -4 -6 68 206
use NOR2X1  _3677_
timestamp 1596991774
transform 1 0 5416 0 1 3010
box -4 -6 52 206
use AOI21X1  _3886_
timestamp 1596991774
transform 1 0 5464 0 1 3010
box -4 -6 68 206
use INVX4  _3651_
timestamp 1596991774
transform -1 0 5576 0 1 3010
box -4 -6 52 206
use NOR2X1  _3885_
timestamp 1596991774
transform 1 0 5576 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4336_
timestamp 1596991774
transform -1 0 5816 0 1 3010
box -4 -6 196 206
use BUFX2  BUFX2_insert150
timestamp 1596991774
transform -1 0 5864 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert65
timestamp 1596991774
transform 1 0 5864 0 1 3010
box -4 -6 52 206
use NOR2X1  _4184_
timestamp 1596991774
transform -1 0 6024 0 1 3010
box -4 -6 52 206
use FILL  SFILL59120x30100
timestamp 1596991774
transform 1 0 5912 0 1 3010
box -4 -6 20 206
use FILL  SFILL59280x30100
timestamp 1596991774
transform 1 0 5928 0 1 3010
box -4 -6 20 206
use FILL  SFILL59440x30100
timestamp 1596991774
transform 1 0 5944 0 1 3010
box -4 -6 20 206
use FILL  SFILL59600x30100
timestamp 1596991774
transform 1 0 5960 0 1 3010
box -4 -6 20 206
use NOR2X1  _4006_
timestamp 1596991774
transform -1 0 6072 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert22
timestamp 1596991774
transform -1 0 6120 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert90
timestamp 1596991774
transform -1 0 6168 0 1 3010
box -4 -6 52 206
use INVX4  _3673_
timestamp 1596991774
transform 1 0 6168 0 1 3010
box -4 -6 52 206
use NAND2X1  _3860_
timestamp 1596991774
transform 1 0 6216 0 1 3010
box -4 -6 52 206
use OAI21X1  _3861_
timestamp 1596991774
transform -1 0 6328 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4308_
timestamp 1596991774
transform -1 0 6520 0 1 3010
box -4 -6 196 206
use BUFX2  BUFX2_insert99
timestamp 1596991774
transform 1 0 6520 0 1 3010
box -4 -6 52 206
use NAND2X1  _3776_
timestamp 1596991774
transform -1 0 6616 0 1 3010
box -4 -6 52 206
use NAND2X1  _3843_
timestamp 1596991774
transform -1 0 6664 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert24
timestamp 1596991774
transform 1 0 6664 0 1 3010
box -4 -6 52 206
use AND2X2  _3809_
timestamp 1596991774
transform -1 0 6776 0 1 3010
box -4 -6 68 206
use AND2X2  _3876_
timestamp 1596991774
transform -1 0 6840 0 1 3010
box -4 -6 68 206
use NAND2X1  _3708_
timestamp 1596991774
transform -1 0 6888 0 1 3010
box -4 -6 52 206
use NOR2X1  _3775_
timestamp 1596991774
transform 1 0 6888 0 1 3010
box -4 -6 52 206
use NOR2X1  _3705_
timestamp 1596991774
transform 1 0 6936 0 1 3010
box -4 -6 52 206
use INVX1  _3704_
timestamp 1596991774
transform 1 0 6984 0 1 3010
box -4 -6 36 206
use NOR2X1  _3842_
timestamp 1596991774
transform -1 0 7064 0 1 3010
box -4 -6 52 206
use NOR2X1  _3887_
timestamp 1596991774
transform 1 0 7064 0 1 3010
box -4 -6 52 206
use AOI21X1  _3888_
timestamp 1596991774
transform 1 0 7112 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4337_
timestamp 1596991774
transform -1 0 7368 0 1 3010
box -4 -6 196 206
use FILL  FILL71120x30100
timestamp 1596991774
transform 1 0 7368 0 1 3010
box -4 -6 20 206
use FILL  FILL71280x30100
timestamp 1596991774
transform 1 0 7384 0 1 3010
box -4 -6 20 206
use INVX1  _2219_
timestamp 1596991774
transform 1 0 8 0 -1 3410
box -4 -6 36 206
use NOR2X1  _2221_
timestamp 1596991774
transform -1 0 88 0 -1 3410
box -4 -6 52 206
use NAND2X1  _2233_
timestamp 1596991774
transform 1 0 88 0 -1 3410
box -4 -6 52 206
use OAI21X1  _2223_
timestamp 1596991774
transform 1 0 136 0 -1 3410
box -4 -6 68 206
use NAND2X1  _2218_
timestamp 1596991774
transform -1 0 248 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2220_
timestamp 1596991774
transform 1 0 248 0 -1 3410
box -4 -6 52 206
use AND2X2  _2318_
timestamp 1596991774
transform 1 0 296 0 -1 3410
box -4 -6 68 206
use NOR2X1  _2319_
timestamp 1596991774
transform -1 0 408 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2317_
timestamp 1596991774
transform -1 0 456 0 -1 3410
box -4 -6 52 206
use AND2X2  _2365_
timestamp 1596991774
transform 1 0 456 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3243_
timestamp 1596991774
transform 1 0 520 0 -1 3410
box -4 -6 68 206
use INVX1  _3179_
timestamp 1596991774
transform 1 0 584 0 -1 3410
box -4 -6 36 206
use OAI22X1  _3180_
timestamp 1596991774
transform -1 0 696 0 -1 3410
box -4 -6 84 206
use NOR2X1  _3259_
timestamp 1596991774
transform 1 0 696 0 -1 3410
box -4 -6 52 206
use OAI22X1  _3255_
timestamp 1596991774
transform 1 0 744 0 -1 3410
box -4 -6 84 206
use INVX1  _3254_
timestamp 1596991774
transform -1 0 856 0 -1 3410
box -4 -6 36 206
use OAI22X1  _3206_
timestamp 1596991774
transform 1 0 856 0 -1 3410
box -4 -6 84 206
use INVX1  _3205_
timestamp 1596991774
transform 1 0 936 0 -1 3410
box -4 -6 36 206
use NOR2X1  _3181_
timestamp 1596991774
transform 1 0 968 0 -1 3410
box -4 -6 52 206
use NOR2X1  _3207_
timestamp 1596991774
transform 1 0 1016 0 -1 3410
box -4 -6 52 206
use OAI22X1  _3203_
timestamp 1596991774
transform 1 0 1064 0 -1 3410
box -4 -6 84 206
use INVX1  _3202_
timestamp 1596991774
transform -1 0 1176 0 -1 3410
box -4 -6 36 206
use INVX1  _3282_
timestamp 1596991774
transform 1 0 1176 0 -1 3410
box -4 -6 36 206
use INVX1  _3309_
timestamp 1596991774
transform -1 0 1240 0 -1 3410
box -4 -6 36 206
use NAND3X1  _3321_
timestamp 1596991774
transform -1 0 1304 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3295_
timestamp 1596991774
transform -1 0 1368 0 -1 3410
box -4 -6 68 206
use AND2X2  _2370_
timestamp 1596991774
transform -1 0 1432 0 -1 3410
box -4 -6 68 206
use OR2X2  _2354_
timestamp 1596991774
transform -1 0 1560 0 -1 3410
box -4 -6 68 206
use INVX1  _2288_
timestamp 1596991774
transform -1 0 1592 0 -1 3410
box -4 -6 36 206
use OAI21X1  _2289_
timestamp 1596991774
transform 1 0 1592 0 -1 3410
box -4 -6 68 206
use FILL  SFILL14320x32100
timestamp 1596991774
transform -1 0 1448 0 -1 3410
box -4 -6 20 206
use FILL  SFILL14480x32100
timestamp 1596991774
transform -1 0 1464 0 -1 3410
box -4 -6 20 206
use FILL  SFILL14640x32100
timestamp 1596991774
transform -1 0 1480 0 -1 3410
box -4 -6 20 206
use FILL  SFILL14800x32100
timestamp 1596991774
transform -1 0 1496 0 -1 3410
box -4 -6 20 206
use NAND2X1  _2290_
timestamp 1596991774
transform -1 0 1704 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3294_
timestamp 1596991774
transform 1 0 1704 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3346_
timestamp 1596991774
transform -1 0 1832 0 -1 3410
box -4 -6 68 206
use NOR2X1  _2332_
timestamp 1596991774
transform -1 0 1880 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2334_
timestamp 1596991774
transform 1 0 1880 0 -1 3410
box -4 -6 52 206
use AND2X2  _2333_
timestamp 1596991774
transform -1 0 1992 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert250
timestamp 1596991774
transform -1 0 2040 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2337_
timestamp 1596991774
transform -1 0 2088 0 -1 3410
box -4 -6 52 206
use AND2X2  _2336_
timestamp 1596991774
transform -1 0 2152 0 -1 3410
box -4 -6 68 206
use INVX1  _3357_
timestamp 1596991774
transform -1 0 2184 0 -1 3410
box -4 -6 36 206
use OR2X2  _2356_
timestamp 1596991774
transform -1 0 2248 0 -1 3410
box -4 -6 68 206
use NOR2X1  _2338_
timestamp 1596991774
transform 1 0 2248 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2340_
timestamp 1596991774
transform 1 0 2296 0 -1 3410
box -4 -6 52 206
use AND2X2  _2339_
timestamp 1596991774
transform -1 0 2408 0 -1 3410
box -4 -6 68 206
use XOR2X1  _2389_
timestamp 1596991774
transform -1 0 2520 0 -1 3410
box -4 -6 116 206
use NOR2X1  _2390_
timestamp 1596991774
transform -1 0 2568 0 -1 3410
box -4 -6 52 206
use AND2X2  _2381_
timestamp 1596991774
transform 1 0 2568 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert42
timestamp 1596991774
transform 1 0 2632 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert146
timestamp 1596991774
transform 1 0 2680 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert219
timestamp 1596991774
transform -1 0 2776 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert251
timestamp 1596991774
transform 1 0 2776 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4399_
timestamp 1596991774
transform 1 0 2824 0 -1 3410
box -4 -6 196 206
use NOR2X1  _3665_
timestamp 1596991774
transform 1 0 3080 0 -1 3410
box -4 -6 52 206
use AOI21X1  _3666_
timestamp 1596991774
transform -1 0 3192 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4352_
timestamp 1596991774
transform 1 0 3192 0 -1 3410
box -4 -6 196 206
use FILL  SFILL30160x32100
timestamp 1596991774
transform -1 0 3032 0 -1 3410
box -4 -6 20 206
use FILL  SFILL30320x32100
timestamp 1596991774
transform -1 0 3048 0 -1 3410
box -4 -6 20 206
use FILL  SFILL30480x32100
timestamp 1596991774
transform -1 0 3064 0 -1 3410
box -4 -6 20 206
use FILL  SFILL30640x32100
timestamp 1596991774
transform -1 0 3080 0 -1 3410
box -4 -6 20 206
use MUX2X1  _4128_
timestamp 1596991774
transform -1 0 3480 0 -1 3410
box -4 -6 100 206
use MUX2X1  _3954_
timestamp 1596991774
transform -1 0 3576 0 -1 3410
box -4 -6 100 206
use AOI21X1  _3819_
timestamp 1596991774
transform 1 0 3576 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3818_
timestamp 1596991774
transform -1 0 3688 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4384_
timestamp 1596991774
transform -1 0 3880 0 -1 3410
box -4 -6 196 206
use MUX2X1  _4143_
timestamp 1596991774
transform -1 0 3976 0 -1 3410
box -4 -6 100 206
use MUX2X1  _3965_
timestamp 1596991774
transform -1 0 4072 0 -1 3410
box -4 -6 100 206
use DFFPOSX1  _4372_
timestamp 1596991774
transform 1 0 4072 0 -1 3410
box -4 -6 196 206
use OAI21X1  _3727_
timestamp 1596991774
transform 1 0 4264 0 -1 3410
box -4 -6 68 206
use OAI21X1  _3726_
timestamp 1596991774
transform -1 0 4392 0 -1 3410
box -4 -6 68 206
use NOR2X1  _4180_
timestamp 1596991774
transform -1 0 4440 0 -1 3410
box -4 -6 52 206
use OAI22X1  _4182_
timestamp 1596991774
transform 1 0 4504 0 -1 3410
box -4 -6 84 206
use OAI21X1  _4181_
timestamp 1596991774
transform -1 0 4648 0 -1 3410
box -4 -6 68 206
use FILL  SFILL44400x32100
timestamp 1596991774
transform -1 0 4456 0 -1 3410
box -4 -6 20 206
use FILL  SFILL44560x32100
timestamp 1596991774
transform -1 0 4472 0 -1 3410
box -4 -6 20 206
use FILL  SFILL44720x32100
timestamp 1596991774
transform -1 0 4488 0 -1 3410
box -4 -6 20 206
use FILL  SFILL44880x32100
timestamp 1596991774
transform -1 0 4504 0 -1 3410
box -4 -6 20 206
use BUFX2  BUFX2_insert135
timestamp 1596991774
transform -1 0 4696 0 -1 3410
box -4 -6 52 206
use NAND2X1  _3759_
timestamp 1596991774
transform 1 0 4696 0 -1 3410
box -4 -6 52 206
use OAI22X1  _3964_
timestamp 1596991774
transform -1 0 4824 0 -1 3410
box -4 -6 84 206
use NOR2X1  _3962_
timestamp 1596991774
transform -1 0 4872 0 -1 3410
box -4 -6 52 206
use NOR2X1  _4140_
timestamp 1596991774
transform 1 0 4872 0 -1 3410
box -4 -6 52 206
use OAI22X1  _4142_
timestamp 1596991774
transform 1 0 4920 0 -1 3410
box -4 -6 84 206
use MUX2X1  _4139_
timestamp 1596991774
transform 1 0 5000 0 -1 3410
box -4 -6 100 206
use MUX2X1  _3961_
timestamp 1596991774
transform -1 0 5192 0 -1 3410
box -4 -6 100 206
use DFFPOSX1  _4416_
timestamp 1596991774
transform -1 0 5384 0 -1 3410
box -4 -6 196 206
use OAI21X1  _4141_
timestamp 1596991774
transform -1 0 5448 0 -1 3410
box -4 -6 68 206
use INVX8  _4091_
timestamp 1596991774
transform -1 0 5528 0 -1 3410
box -4 -6 84 206
use BUFX2  BUFX2_insert48
timestamp 1596991774
transform 1 0 5528 0 -1 3410
box -4 -6 52 206
use OAI21X1  _3963_
timestamp 1596991774
transform -1 0 5640 0 -1 3410
box -4 -6 68 206
use OAI22X1  _4186_
timestamp 1596991774
transform -1 0 5720 0 -1 3410
box -4 -6 84 206
use MUX2X1  _4183_
timestamp 1596991774
transform 1 0 5720 0 -1 3410
box -4 -6 100 206
use MUX2X1  _4005_
timestamp 1596991774
transform 1 0 5816 0 -1 3410
box -4 -6 100 206
use OAI22X1  _4008_
timestamp 1596991774
transform 1 0 5976 0 -1 3410
box -4 -6 84 206
use FILL  SFILL59120x32100
timestamp 1596991774
transform -1 0 5928 0 -1 3410
box -4 -6 20 206
use FILL  SFILL59280x32100
timestamp 1596991774
transform -1 0 5944 0 -1 3410
box -4 -6 20 206
use FILL  SFILL59440x32100
timestamp 1596991774
transform -1 0 5960 0 -1 3410
box -4 -6 20 206
use FILL  SFILL59600x32100
timestamp 1596991774
transform -1 0 5976 0 -1 3410
box -4 -6 20 206
use MUX2X1  _3976_
timestamp 1596991774
transform 1 0 6056 0 -1 3410
box -4 -6 100 206
use OAI22X1  _3975_
timestamp 1596991774
transform -1 0 6232 0 -1 3410
box -4 -6 84 206
use OAI21X1  _3974_
timestamp 1596991774
transform -1 0 6296 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3973_
timestamp 1596991774
transform 1 0 6296 0 -1 3410
box -4 -6 52 206
use NOR2X1  _4151_
timestamp 1596991774
transform -1 0 6392 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4420_
timestamp 1596991774
transform -1 0 6584 0 -1 3410
box -4 -6 196 206
use MUX2X1  _3972_
timestamp 1596991774
transform 1 0 6584 0 -1 3410
box -4 -6 100 206
use NAND2X1  _3854_
timestamp 1596991774
transform -1 0 6728 0 -1 3410
box -4 -6 52 206
use OAI21X1  _3855_
timestamp 1596991774
transform -1 0 6792 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4305_
timestamp 1596991774
transform -1 0 6984 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  _4306_
timestamp 1596991774
transform -1 0 7176 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  _4401_
timestamp 1596991774
transform -1 0 7368 0 -1 3410
box -4 -6 196 206
use FILL  FILL71120x32100
timestamp 1596991774
transform -1 0 7384 0 -1 3410
box -4 -6 20 206
use FILL  FILL71280x32100
timestamp 1596991774
transform -1 0 7400 0 -1 3410
box -4 -6 20 206
use INVX1  _2232_
timestamp 1596991774
transform 1 0 8 0 1 3410
box -4 -6 36 206
use OAI21X1  _2234_
timestamp 1596991774
transform -1 0 104 0 1 3410
box -4 -6 68 206
use NOR2X1  _2281_
timestamp 1596991774
transform -1 0 152 0 1 3410
box -4 -6 52 206
use OR2X2  _2252_
timestamp 1596991774
transform 1 0 152 0 1 3410
box -4 -6 68 206
use AOI21X1  _2256_
timestamp 1596991774
transform 1 0 8 0 -1 3810
box -4 -6 68 206
use INVX1  _3178_
timestamp 1596991774
transform 1 0 72 0 -1 3810
box -4 -6 36 206
use INVX1  _2253_
timestamp 1596991774
transform -1 0 136 0 -1 3810
box -4 -6 36 206
use NAND2X1  _2251_
timestamp 1596991774
transform -1 0 184 0 -1 3810
box -4 -6 52 206
use INVX1  _2246_
timestamp 1596991774
transform 1 0 184 0 -1 3810
box -4 -6 36 206
use OAI21X1  _2257_
timestamp 1596991774
transform 1 0 216 0 1 3410
box -4 -6 68 206
use AND2X2  _2238_
timestamp 1596991774
transform -1 0 344 0 1 3410
box -4 -6 68 206
use NAND2X1  _2250_
timestamp 1596991774
transform 1 0 344 0 1 3410
box -4 -6 52 206
use NOR2X1  _2239_
timestamp 1596991774
transform -1 0 440 0 1 3410
box -4 -6 52 206
use NAND2X1  _2249_
timestamp 1596991774
transform 1 0 216 0 -1 3810
box -4 -6 52 206
use NOR2X1  _2248_
timestamp 1596991774
transform -1 0 312 0 -1 3810
box -4 -6 52 206
use OAI21X1  _2247_
timestamp 1596991774
transform -1 0 376 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert28
timestamp 1596991774
transform 1 0 376 0 -1 3810
box -4 -6 52 206
use NOR2X1  _2240_
timestamp 1596991774
transform -1 0 488 0 1 3410
box -4 -6 52 206
use AOI21X1  _2283_
timestamp 1596991774
transform 1 0 488 0 1 3410
box -4 -6 68 206
use INVX1  _3257_
timestamp 1596991774
transform 1 0 552 0 1 3410
box -4 -6 36 206
use OAI22X1  _3258_
timestamp 1596991774
transform -1 0 664 0 1 3410
box -4 -6 84 206
use INVX1  _3230_
timestamp 1596991774
transform -1 0 456 0 -1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert167
timestamp 1596991774
transform -1 0 504 0 -1 3810
box -4 -6 52 206
use OR2X2  _2352_
timestamp 1596991774
transform 1 0 504 0 -1 3810
box -4 -6 68 206
use INVX1  _3253_
timestamp 1596991774
transform 1 0 568 0 -1 3810
box -4 -6 36 206
use AND2X2  _2544_
timestamp 1596991774
transform 1 0 600 0 -1 3810
box -4 -6 68 206
use OAI22X1  _3232_
timestamp 1596991774
transform 1 0 664 0 1 3410
box -4 -6 84 206
use INVX1  _3231_
timestamp 1596991774
transform -1 0 776 0 1 3410
box -4 -6 36 206
use NOR2X1  _3233_
timestamp 1596991774
transform 1 0 776 0 1 3410
box -4 -6 52 206
use AOI21X1  _2560_
timestamp 1596991774
transform 1 0 664 0 -1 3810
box -4 -6 68 206
use INVX1  _3227_
timestamp 1596991774
transform 1 0 728 0 -1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert236
timestamp 1596991774
transform 1 0 760 0 -1 3810
box -4 -6 52 206
use OAI21X1  _2545_
timestamp 1596991774
transform 1 0 808 0 -1 3810
box -4 -6 68 206
use OAI22X1  _3229_
timestamp 1596991774
transform 1 0 824 0 1 3410
box -4 -6 84 206
use INVX1  _3228_
timestamp 1596991774
transform -1 0 936 0 1 3410
box -4 -6 36 206
use INVX1  _3176_
timestamp 1596991774
transform 1 0 936 0 1 3410
box -4 -6 36 206
use OAI22X1  _3177_
timestamp 1596991774
transform -1 0 1048 0 1 3410
box -4 -6 84 206
use INVX1  _3175_
timestamp 1596991774
transform 1 0 872 0 -1 3810
box -4 -6 36 206
use XNOR2X1  _2551_
timestamp 1596991774
transform 1 0 904 0 -1 3810
box -4 -6 116 206
use OR2X2  _2350_
timestamp 1596991774
transform 1 0 1048 0 1 3410
box -4 -6 68 206
use INVX1  _3201_
timestamp 1596991774
transform -1 0 1144 0 1 3410
box -4 -6 36 206
use OAI22X1  _3310_
timestamp 1596991774
transform 1 0 1144 0 1 3410
box -4 -6 84 206
use NOR2X1  _2552_
timestamp 1596991774
transform -1 0 1064 0 -1 3810
box -4 -6 52 206
use INVX1  _3308_
timestamp 1596991774
transform 1 0 1064 0 -1 3810
box -4 -6 36 206
use XNOR2X1  _2536_
timestamp 1596991774
transform 1 0 1096 0 -1 3810
box -4 -6 116 206
use NAND2X1  _2535_
timestamp 1596991774
transform -1 0 1256 0 -1 3810
box -4 -6 52 206
use NOR2X1  _3311_
timestamp 1596991774
transform 1 0 1224 0 1 3410
box -4 -6 52 206
use OAI22X1  _3307_
timestamp 1596991774
transform 1 0 1272 0 1 3410
box -4 -6 84 206
use INVX1  _3306_
timestamp 1596991774
transform -1 0 1384 0 1 3410
box -4 -6 36 206
use INVX1  _3305_
timestamp 1596991774
transform -1 0 1416 0 1 3410
box -4 -6 36 206
use XNOR2X1  _2264_
timestamp 1596991774
transform -1 0 1368 0 -1 3810
box -4 -6 116 206
use AOI21X1  _2262_
timestamp 1596991774
transform 1 0 1368 0 -1 3810
box -4 -6 68 206
use FILL  SFILL14160x34100
timestamp 1596991774
transform 1 0 1416 0 1 3410
box -4 -6 20 206
use FILL  SFILL14320x34100
timestamp 1596991774
transform 1 0 1432 0 1 3410
box -4 -6 20 206
use FILL  SFILL14480x34100
timestamp 1596991774
transform 1 0 1448 0 1 3410
box -4 -6 20 206
use FILL  SFILL14320x36100
timestamp 1596991774
transform -1 0 1448 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14480x36100
timestamp 1596991774
transform -1 0 1464 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14640x34100
timestamp 1596991774
transform 1 0 1464 0 1 3410
box -4 -6 20 206
use FILL  SFILL14640x36100
timestamp 1596991774
transform -1 0 1480 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14800x36100
timestamp 1596991774
transform -1 0 1496 0 -1 3810
box -4 -6 20 206
use NAND2X1  _2265_
timestamp 1596991774
transform -1 0 1528 0 1 3410
box -4 -6 52 206
use NOR2X1  _2260_
timestamp 1596991774
transform -1 0 1544 0 -1 3810
box -4 -6 52 206
use OAI21X1  _2270_
timestamp 1596991774
transform -1 0 1672 0 -1 3810
box -4 -6 68 206
use OAI21X1  _2269_
timestamp 1596991774
transform -1 0 1608 0 -1 3810
box -4 -6 68 206
use XOR2X1  _2261_
timestamp 1596991774
transform -1 0 1640 0 1 3410
box -4 -6 116 206
use INVX1  _2266_
timestamp 1596991774
transform 1 0 1640 0 1 3410
box -4 -6 36 206
use AOI21X1  _2271_
timestamp 1596991774
transform 1 0 1672 0 1 3410
box -4 -6 68 206
use OAI21X1  _2284_
timestamp 1596991774
transform 1 0 1736 0 1 3410
box -4 -6 68 206
use NAND2X1  _2291_
timestamp 1596991774
transform -1 0 1848 0 1 3410
box -4 -6 52 206
use INVX1  _2267_
timestamp 1596991774
transform 1 0 1672 0 -1 3810
box -4 -6 36 206
use NOR2X1  _2331_
timestamp 1596991774
transform -1 0 1752 0 -1 3810
box -4 -6 52 206
use AND2X2  _2330_
timestamp 1596991774
transform -1 0 1816 0 -1 3810
box -4 -6 68 206
use NAND3X1  _2287_
timestamp 1596991774
transform -1 0 1912 0 1 3410
box -4 -6 68 206
use INVX1  _2286_
timestamp 1596991774
transform -1 0 1944 0 1 3410
box -4 -6 36 206
use AND2X2  _2274_
timestamp 1596991774
transform 1 0 1944 0 1 3410
box -4 -6 68 206
use NAND2X1  _2272_
timestamp 1596991774
transform -1 0 2056 0 1 3410
box -4 -6 52 206
use NOR2X1  _2329_
timestamp 1596991774
transform -1 0 1864 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert1
timestamp 1596991774
transform 1 0 1864 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert189
timestamp 1596991774
transform 1 0 1912 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert187
timestamp 1596991774
transform 1 0 1960 0 -1 3810
box -4 -6 52 206
use OR2X2  _2273_
timestamp 1596991774
transform -1 0 2072 0 -1 3810
box -4 -6 68 206
use NOR2X1  _2335_
timestamp 1596991774
transform -1 0 2104 0 1 3410
box -4 -6 52 206
use INVX1  _3335_
timestamp 1596991774
transform 1 0 2104 0 1 3410
box -4 -6 36 206
use OAI22X1  _3336_
timestamp 1596991774
transform -1 0 2216 0 1 3410
box -4 -6 84 206
use XNOR2X1  _2555_
timestamp 1596991774
transform -1 0 2184 0 -1 3810
box -4 -6 116 206
use INVX1  _3334_
timestamp 1596991774
transform -1 0 2216 0 -1 3810
box -4 -6 36 206
use NOR2X1  _3337_
timestamp 1596991774
transform 1 0 2216 0 1 3410
box -4 -6 52 206
use OR2X2  _2355_
timestamp 1596991774
transform 1 0 2264 0 1 3410
box -4 -6 68 206
use INVX1  _3331_
timestamp 1596991774
transform 1 0 2328 0 1 3410
box -4 -6 36 206
use OAI22X1  _3333_
timestamp 1596991774
transform 1 0 2360 0 1 3410
box -4 -6 84 206
use INVX1  _3360_
timestamp 1596991774
transform 1 0 2216 0 -1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert61
timestamp 1596991774
transform -1 0 2296 0 -1 3810
box -4 -6 52 206
use XNOR2X1  _2285_
timestamp 1596991774
transform -1 0 2408 0 -1 3810
box -4 -6 116 206
use BUFX2  BUFX2_insert86
timestamp 1596991774
transform -1 0 2456 0 -1 3810
box -4 -6 52 206
use INVX1  _3332_
timestamp 1596991774
transform -1 0 2472 0 1 3410
box -4 -6 36 206
use BUFX2  BUFX2_insert148
timestamp 1596991774
transform -1 0 2520 0 1 3410
box -4 -6 52 206
use XOR2X1  _2388_
timestamp 1596991774
transform -1 0 2632 0 1 3410
box -4 -6 116 206
use DFFPOSX1  _4452_
timestamp 1596991774
transform -1 0 2648 0 -1 3810
box -4 -6 196 206
use AND2X2  _2367_
timestamp 1596991774
transform -1 0 2696 0 1 3410
box -4 -6 68 206
use XNOR2X1  _2405_
timestamp 1596991774
transform 1 0 2696 0 1 3410
box -4 -6 116 206
use NAND2X1  _2406_
timestamp 1596991774
transform -1 0 2856 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4436_
timestamp 1596991774
transform -1 0 2840 0 -1 3810
box -4 -6 196 206
use FILL  SFILL29040x36100
timestamp 1596991774
transform -1 0 2920 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29040x34100
timestamp 1596991774
transform 1 0 2904 0 1 3410
box -4 -6 20 206
use FILL  SFILL28880x34100
timestamp 1596991774
transform 1 0 2888 0 1 3410
box -4 -6 20 206
use FILL  SFILL28720x34100
timestamp 1596991774
transform 1 0 2872 0 1 3410
box -4 -6 20 206
use FILL  SFILL28560x34100
timestamp 1596991774
transform 1 0 2856 0 1 3410
box -4 -6 20 206
use AOI21X1  _4189_
timestamp 1596991774
transform -1 0 2904 0 -1 3810
box -4 -6 68 206
use FILL  SFILL29520x36100
timestamp 1596991774
transform -1 0 2968 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29360x36100
timestamp 1596991774
transform -1 0 2952 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29200x36100
timestamp 1596991774
transform -1 0 2936 0 -1 3810
box -4 -6 20 206
use DFFPOSX1  _4351_
timestamp 1596991774
transform 1 0 2968 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  _4453_
timestamp 1596991774
transform -1 0 3112 0 1 3410
box -4 -6 196 206
use DFFPOSX1  _4415_
timestamp 1596991774
transform 1 0 3112 0 1 3410
box -4 -6 196 206
use OAI21X1  _3784_
timestamp 1596991774
transform 1 0 3160 0 -1 3810
box -4 -6 68 206
use AOI21X1  _4275_
timestamp 1596991774
transform 1 0 3304 0 1 3410
box -4 -6 68 206
use NOR2X1  _4274_
timestamp 1596991774
transform -1 0 3416 0 1 3410
box -4 -6 52 206
use MUX2X1  _3950_
timestamp 1596991774
transform -1 0 3512 0 1 3410
box -4 -6 100 206
use NAND2X1  _3783_
timestamp 1596991774
transform -1 0 3272 0 -1 3810
box -4 -6 52 206
use AOI21X1  _4297_
timestamp 1596991774
transform 1 0 3272 0 -1 3810
box -4 -6 68 206
use NOR2X1  _4296_
timestamp 1596991774
transform -1 0 3384 0 -1 3810
box -4 -6 52 206
use MUX2X1  _4124_
timestamp 1596991774
transform -1 0 3480 0 -1 3810
box -4 -6 100 206
use OAI22X1  _4127_
timestamp 1596991774
transform -1 0 3592 0 1 3410
box -4 -6 84 206
use OAI22X1  _3953_
timestamp 1596991774
transform -1 0 3672 0 1 3410
box -4 -6 84 206
use MUX2X1  _3946_
timestamp 1596991774
transform -1 0 3576 0 -1 3810
box -4 -6 100 206
use OAI21X1  _4126_
timestamp 1596991774
transform 1 0 3576 0 -1 3810
box -4 -6 68 206
use OAI21X1  _3952_
timestamp 1596991774
transform 1 0 3672 0 1 3410
box -4 -6 68 206
use NOR2X1  _3951_
timestamp 1596991774
transform 1 0 3736 0 1 3410
box -4 -6 52 206
use NOR2X1  _3698_
timestamp 1596991774
transform -1 0 3832 0 1 3410
box -4 -6 52 206
use OAI22X1  _3949_
timestamp 1596991774
transform -1 0 3720 0 -1 3810
box -4 -6 84 206
use NAND2X1  _3850_
timestamp 1596991774
transform 1 0 3720 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3851_
timestamp 1596991774
transform -1 0 3832 0 -1 3810
box -4 -6 68 206
use AOI21X1  _3699_
timestamp 1596991774
transform -1 0 3896 0 1 3410
box -4 -6 68 206
use MUX2X1  _4135_
timestamp 1596991774
transform 1 0 3896 0 1 3410
box -4 -6 100 206
use MUX2X1  _3957_
timestamp 1596991774
transform 1 0 3992 0 1 3410
box -4 -6 100 206
use DFFPOSX1  _4303_
timestamp 1596991774
transform -1 0 4024 0 -1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert74
timestamp 1596991774
transform -1 0 4136 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4410_
timestamp 1596991774
transform -1 0 4328 0 1 3410
box -4 -6 196 206
use OAI22X1  _4138_
timestamp 1596991774
transform -1 0 4104 0 -1 3810
box -4 -6 84 206
use OAI22X1  _3960_
timestamp 1596991774
transform -1 0 4184 0 -1 3810
box -4 -6 84 206
use NOR2X1  _3958_
timestamp 1596991774
transform -1 0 4232 0 -1 3810
box -4 -6 52 206
use MUX2X1  _4009_
timestamp 1596991774
transform -1 0 4424 0 1 3410
box -4 -6 100 206
use NOR2X1  _4136_
timestamp 1596991774
transform 1 0 4232 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3959_
timestamp 1596991774
transform -1 0 4344 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4368_
timestamp 1596991774
transform -1 0 4600 0 -1 3810
box -4 -6 196 206
use FILL  SFILL43440x36100
timestamp 1596991774
transform -1 0 4360 0 -1 3810
box -4 -6 20 206
use FILL  SFILL43600x36100
timestamp 1596991774
transform -1 0 4376 0 -1 3810
box -4 -6 20 206
use FILL  SFILL43760x36100
timestamp 1596991774
transform -1 0 4392 0 -1 3810
box -4 -6 20 206
use FILL  SFILL43920x36100
timestamp 1596991774
transform -1 0 4408 0 -1 3810
box -4 -6 20 206
use NOR2X1  _4002_
timestamp 1596991774
transform 1 0 4488 0 1 3410
box -4 -6 52 206
use OAI22X1  _4004_
timestamp 1596991774
transform -1 0 4616 0 1 3410
box -4 -6 84 206
use OAI21X1  _4003_
timestamp 1596991774
transform -1 0 4680 0 1 3410
box -4 -6 68 206
use OAI21X1  _3718_
timestamp 1596991774
transform -1 0 4664 0 -1 3810
box -4 -6 68 206
use FILL  SFILL44240x34100
timestamp 1596991774
transform 1 0 4424 0 1 3410
box -4 -6 20 206
use FILL  SFILL44400x34100
timestamp 1596991774
transform 1 0 4440 0 1 3410
box -4 -6 20 206
use FILL  SFILL44560x34100
timestamp 1596991774
transform 1 0 4456 0 1 3410
box -4 -6 20 206
use FILL  SFILL44720x34100
timestamp 1596991774
transform 1 0 4472 0 1 3410
box -4 -6 20 206
use BUFX2  BUFX2_insert227
timestamp 1596991774
transform -1 0 4728 0 1 3410
box -4 -6 52 206
use MUX2X1  _4187_
timestamp 1596991774
transform 1 0 4728 0 1 3410
box -4 -6 100 206
use OAI21X1  _3719_
timestamp 1596991774
transform -1 0 4728 0 -1 3810
box -4 -6 68 206
use NAND2X1  _3751_
timestamp 1596991774
transform 1 0 4728 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3752_
timestamp 1596991774
transform -1 0 4840 0 -1 3810
box -4 -6 68 206
use OAI21X1  _3760_
timestamp 1596991774
transform -1 0 4888 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert45
timestamp 1596991774
transform -1 0 4936 0 1 3410
box -4 -6 52 206
use AOI21X1  _3669_
timestamp 1596991774
transform 1 0 4936 0 1 3410
box -4 -6 68 206
use NOR2X1  _3668_
timestamp 1596991774
transform -1 0 5048 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4324_
timestamp 1596991774
transform -1 0 5032 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  _4400_
timestamp 1596991774
transform 1 0 5048 0 1 3410
box -4 -6 196 206
use NOR2X1  _4261_
timestamp 1596991774
transform 1 0 5032 0 -1 3810
box -4 -6 52 206
use OAI22X1  _4263_
timestamp 1596991774
transform -1 0 5160 0 -1 3810
box -4 -6 84 206
use OAI21X1  _4262_
timestamp 1596991774
transform -1 0 5224 0 -1 3810
box -4 -6 68 206
use NOR2X1  _4276_
timestamp 1596991774
transform 1 0 5240 0 1 3410
box -4 -6 52 206
use AOI21X1  _4277_
timestamp 1596991774
transform -1 0 5352 0 1 3410
box -4 -6 68 206
use NOR2X1  _3701_
timestamp 1596991774
transform 1 0 5352 0 1 3410
box -4 -6 52 206
use AOI21X1  _3702_
timestamp 1596991774
transform -1 0 5464 0 1 3410
box -4 -6 68 206
use MUX2X1  _4082_
timestamp 1596991774
transform 1 0 5224 0 -1 3810
box -4 -6 100 206
use MUX2X1  _4260_
timestamp 1596991774
transform -1 0 5416 0 -1 3810
box -4 -6 100 206
use BUFX2  BUFX2_insert210
timestamp 1596991774
transform -1 0 5464 0 -1 3810
box -4 -6 52 206
use DFFPOSX1  _4411_
timestamp 1596991774
transform -1 0 5656 0 1 3410
box -4 -6 196 206
use AOI21X1  _4299_
timestamp 1596991774
transform 1 0 5464 0 -1 3810
box -4 -6 68 206
use NOR2X1  _4298_
timestamp 1596991774
transform 1 0 5528 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert280
timestamp 1596991774
transform 1 0 5576 0 -1 3810
box -4 -6 52 206
use OAI21X1  _4185_
timestamp 1596991774
transform -1 0 5720 0 1 3410
box -4 -6 68 206
use NOR2X1  _3893_
timestamp 1596991774
transform -1 0 5768 0 1 3410
box -4 -6 52 206
use AOI21X1  _3894_
timestamp 1596991774
transform -1 0 5832 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert93
timestamp 1596991774
transform -1 0 5672 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert205
timestamp 1596991774
transform 1 0 5672 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert64
timestamp 1596991774
transform 1 0 5720 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert253
timestamp 1596991774
transform -1 0 5816 0 -1 3810
box -4 -6 52 206
use MUX2X1  _3987_
timestamp 1596991774
transform 1 0 5816 0 -1 3810
box -4 -6 100 206
use DFFPOSX1  _4340_
timestamp 1596991774
transform 1 0 5832 0 1 3410
box -4 -6 196 206
use MUX2X1  _4165_
timestamp 1596991774
transform -1 0 6072 0 -1 3810
box -4 -6 100 206
use FILL  SFILL59120x36100
timestamp 1596991774
transform -1 0 5928 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59280x36100
timestamp 1596991774
transform -1 0 5944 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59440x36100
timestamp 1596991774
transform -1 0 5960 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59600x36100
timestamp 1596991774
transform -1 0 5976 0 -1 3810
box -4 -6 20 206
use OAI21X1  _4007_
timestamp 1596991774
transform 1 0 6088 0 1 3410
box -4 -6 68 206
use MUX2X1  _4154_
timestamp 1596991774
transform 1 0 6152 0 1 3410
box -4 -6 100 206
use NOR2X1  _3984_
timestamp 1596991774
transform -1 0 6120 0 -1 3810
box -4 -6 52 206
use OAI22X1  _3986_
timestamp 1596991774
transform 1 0 6120 0 -1 3810
box -4 -6 84 206
use OAI21X1  _3985_
timestamp 1596991774
transform -1 0 6264 0 -1 3810
box -4 -6 68 206
use FILL  SFILL60240x34100
timestamp 1596991774
transform 1 0 6024 0 1 3410
box -4 -6 20 206
use FILL  SFILL60400x34100
timestamp 1596991774
transform 1 0 6040 0 1 3410
box -4 -6 20 206
use FILL  SFILL60560x34100
timestamp 1596991774
transform 1 0 6056 0 1 3410
box -4 -6 20 206
use FILL  SFILL60720x34100
timestamp 1596991774
transform 1 0 6072 0 1 3410
box -4 -6 20 206
use BUFX2  BUFX2_insert75
timestamp 1596991774
transform 1 0 6248 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert255
timestamp 1596991774
transform 1 0 6296 0 1 3410
box -4 -6 52 206
use OAI22X1  _4153_
timestamp 1596991774
transform 1 0 6344 0 1 3410
box -4 -6 84 206
use NOR2X1  _4162_
timestamp 1596991774
transform -1 0 6312 0 -1 3810
box -4 -6 52 206
use OAI22X1  _4164_
timestamp 1596991774
transform 1 0 6312 0 -1 3810
box -4 -6 84 206
use OAI21X1  _4163_
timestamp 1596991774
transform -1 0 6456 0 -1 3810
box -4 -6 68 206
use OAI21X1  _4152_
timestamp 1596991774
transform -1 0 6488 0 1 3410
box -4 -6 68 206
use NOR2X1  _4284_
timestamp 1596991774
transform 1 0 6488 0 1 3410
box -4 -6 52 206
use AOI21X1  _4285_
timestamp 1596991774
transform -1 0 6600 0 1 3410
box -4 -6 68 206
use MUX2X1  _4150_
timestamp 1596991774
transform 1 0 6600 0 1 3410
box -4 -6 100 206
use MUX2X1  _4161_
timestamp 1596991774
transform -1 0 6552 0 -1 3810
box -4 -6 100 206
use MUX2X1  _3983_
timestamp 1596991774
transform 1 0 6552 0 -1 3810
box -4 -6 100 206
use AOI21X1  _3681_
timestamp 1596991774
transform 1 0 6696 0 1 3410
box -4 -6 68 206
use NOR2X1  _3680_
timestamp 1596991774
transform -1 0 6808 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4404_
timestamp 1596991774
transform -1 0 7000 0 1 3410
box -4 -6 196 206
use DFFPOSX1  _4422_
timestamp 1596991774
transform -1 0 6840 0 -1 3810
box -4 -6 196 206
use AOI21X1  _3833_
timestamp 1596991774
transform -1 0 7064 0 1 3410
box -4 -6 68 206
use NOR2X1  _3674_
timestamp 1596991774
transform -1 0 6888 0 -1 3810
box -4 -6 52 206
use AOI21X1  _3675_
timestamp 1596991774
transform -1 0 6952 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4402_
timestamp 1596991774
transform -1 0 7144 0 -1 3810
box -4 -6 196 206
use OAI21X1  _3857_
timestamp 1596991774
transform 1 0 7064 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert23
timestamp 1596991774
transform 1 0 7128 0 1 3410
box -4 -6 52 206
use NOR2X1  _3671_
timestamp 1596991774
transform -1 0 7224 0 1 3410
box -4 -6 52 206
use AOI21X1  _3672_
timestamp 1596991774
transform -1 0 7288 0 1 3410
box -4 -6 68 206
use AOI21X1  _4281_
timestamp 1596991774
transform 1 0 7144 0 -1 3810
box -4 -6 68 206
use NOR2X1  _4280_
timestamp 1596991774
transform 1 0 7208 0 -1 3810
box -4 -6 52 206
use AOI21X1  _4279_
timestamp 1596991774
transform 1 0 7288 0 1 3410
box -4 -6 68 206
use NOR2X1  _4278_
timestamp 1596991774
transform -1 0 7400 0 1 3410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert17
timestamp 1596991774
transform -1 0 7400 0 -1 3810
box -4 -6 148 206
use XNOR2X1  _2500_
timestamp 1596991774
transform 1 0 8 0 1 3810
box -4 -6 116 206
use OAI21X1  _2255_
timestamp 1596991774
transform -1 0 184 0 1 3810
box -4 -6 68 206
use NOR2X1  _2243_
timestamp 1596991774
transform 1 0 184 0 1 3810
box -4 -6 52 206
use NOR2X1  _2245_
timestamp 1596991774
transform -1 0 280 0 1 3810
box -4 -6 52 206
use INVX1  _2241_
timestamp 1596991774
transform -1 0 312 0 1 3810
box -4 -6 36 206
use INVX1  _2242_
timestamp 1596991774
transform -1 0 344 0 1 3810
box -4 -6 36 206
use NOR2X1  _2244_
timestamp 1596991774
transform 1 0 344 0 1 3810
box -4 -6 52 206
use OAI21X1  _2254_
timestamp 1596991774
transform -1 0 456 0 1 3810
box -4 -6 68 206
use NOR2X1  _2237_
timestamp 1596991774
transform -1 0 504 0 1 3810
box -4 -6 52 206
use AND2X2  _2235_
timestamp 1596991774
transform -1 0 568 0 1 3810
box -4 -6 68 206
use NOR2X1  _2236_
timestamp 1596991774
transform 1 0 568 0 1 3810
box -4 -6 52 206
use AND2X2  _2368_
timestamp 1596991774
transform 1 0 616 0 1 3810
box -4 -6 68 206
use OR2X2  _2351_
timestamp 1596991774
transform 1 0 680 0 1 3810
box -4 -6 68 206
use INVX1  _2559_
timestamp 1596991774
transform -1 0 776 0 1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert168
timestamp 1596991774
transform 1 0 776 0 1 3810
box -4 -6 52 206
use INVX1  _2876_
timestamp 1596991774
transform 1 0 824 0 1 3810
box -4 -6 36 206
use OR2X2  _2349_
timestamp 1596991774
transform -1 0 920 0 1 3810
box -4 -6 68 206
use OAI21X1  _2932_
timestamp 1596991774
transform 1 0 920 0 1 3810
box -4 -6 68 206
use NAND2X1  _2940_
timestamp 1596991774
transform -1 0 1032 0 1 3810
box -4 -6 52 206
use NAND2X1  _2550_
timestamp 1596991774
transform -1 0 1080 0 1 3810
box -4 -6 52 206
use INVX1  _2548_
timestamp 1596991774
transform -1 0 1112 0 1 3810
box -4 -6 36 206
use OAI21X1  _2553_
timestamp 1596991774
transform 1 0 1112 0 1 3810
box -4 -6 68 206
use AOI21X1  _2554_
timestamp 1596991774
transform 1 0 1176 0 1 3810
box -4 -6 68 206
use OR2X2  _2534_
timestamp 1596991774
transform -1 0 1304 0 1 3810
box -4 -6 68 206
use NAND2X1  _2533_
timestamp 1596991774
transform -1 0 1352 0 1 3810
box -4 -6 52 206
use INVX1  _2532_
timestamp 1596991774
transform -1 0 1384 0 1 3810
box -4 -6 36 206
use AND2X2  _2258_
timestamp 1596991774
transform 1 0 1384 0 1 3810
box -4 -6 68 206
use NOR2X1  _2259_
timestamp 1596991774
transform -1 0 1560 0 1 3810
box -4 -6 52 206
use OAI21X1  _2561_
timestamp 1596991774
transform 1 0 1560 0 1 3810
box -4 -6 68 206
use FILL  SFILL14480x38100
timestamp 1596991774
transform 1 0 1448 0 1 3810
box -4 -6 20 206
use FILL  SFILL14640x38100
timestamp 1596991774
transform 1 0 1464 0 1 3810
box -4 -6 20 206
use FILL  SFILL14800x38100
timestamp 1596991774
transform 1 0 1480 0 1 3810
box -4 -6 20 206
use FILL  SFILL14960x38100
timestamp 1596991774
transform 1 0 1496 0 1 3810
box -4 -6 20 206
use INVX1  _2268_
timestamp 1596991774
transform 1 0 1624 0 1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert248
timestamp 1596991774
transform -1 0 1704 0 1 3810
box -4 -6 52 206
use OR2X2  _2353_
timestamp 1596991774
transform 1 0 1704 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert104
timestamp 1596991774
transform -1 0 1816 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert41
timestamp 1596991774
transform -1 0 1864 0 1 3810
box -4 -6 52 206
use XNOR2X1  _2556_
timestamp 1596991774
transform 1 0 1864 0 1 3810
box -4 -6 116 206
use INVX1  _2565_
timestamp 1596991774
transform 1 0 1976 0 1 3810
box -4 -6 36 206
use OAI21X1  _2566_
timestamp 1596991774
transform 1 0 2008 0 1 3810
box -4 -6 68 206
use NAND3X1  _2564_
timestamp 1596991774
transform 1 0 2072 0 1 3810
box -4 -6 68 206
use NAND2X1  _2568_
timestamp 1596991774
transform 1 0 2136 0 1 3810
box -4 -6 52 206
use NAND2X1  _2567_
timestamp 1596991774
transform -1 0 2232 0 1 3810
box -4 -6 52 206
use INVX1  _2563_
timestamp 1596991774
transform -1 0 2264 0 1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert106
timestamp 1596991774
transform 1 0 2264 0 1 3810
box -4 -6 52 206
use XOR2X1  _2562_
timestamp 1596991774
transform -1 0 2424 0 1 3810
box -4 -6 116 206
use BUFX2  BUFX2_insert88
timestamp 1596991774
transform -1 0 2472 0 1 3810
box -4 -6 52 206
use XNOR2X1  _2404_
timestamp 1596991774
transform 1 0 2472 0 1 3810
box -4 -6 116 206
use BUFX2  BUFX2_insert166
timestamp 1596991774
transform 1 0 2584 0 1 3810
box -4 -6 52 206
use OAI21X1  _4010_
timestamp 1596991774
transform -1 0 2696 0 1 3810
box -4 -6 68 206
use AOI21X1  _4011_
timestamp 1596991774
transform -1 0 2760 0 1 3810
box -4 -6 68 206
use OAI21X1  _4188_
timestamp 1596991774
transform 1 0 2760 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4319_
timestamp 1596991774
transform 1 0 2824 0 1 3810
box -4 -6 196 206
use NAND2X1  _3749_
timestamp 1596991774
transform 1 0 3080 0 1 3810
box -4 -6 52 206
use OAI21X1  _3750_
timestamp 1596991774
transform -1 0 3192 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4426_
timestamp 1596991774
transform 1 0 3192 0 1 3810
box -4 -6 196 206
use FILL  SFILL30160x38100
timestamp 1596991774
transform 1 0 3016 0 1 3810
box -4 -6 20 206
use FILL  SFILL30320x38100
timestamp 1596991774
transform 1 0 3032 0 1 3810
box -4 -6 20 206
use FILL  SFILL30480x38100
timestamp 1596991774
transform 1 0 3048 0 1 3810
box -4 -6 20 206
use FILL  SFILL30640x38100
timestamp 1596991774
transform 1 0 3064 0 1 3810
box -4 -6 20 206
use MUX2X1  _4249_
timestamp 1596991774
transform -1 0 3480 0 1 3810
box -4 -6 100 206
use MUX2X1  _4071_
timestamp 1596991774
transform -1 0 3576 0 1 3810
box -4 -6 100 206
use OAI21X1  _3948_
timestamp 1596991774
transform 1 0 3576 0 1 3810
box -4 -6 68 206
use NOR2X1  _4125_
timestamp 1596991774
transform -1 0 3688 0 1 3810
box -4 -6 52 206
use NOR2X1  _3947_
timestamp 1596991774
transform 1 0 3688 0 1 3810
box -4 -6 52 206
use MUX2X1  _4086_
timestamp 1596991774
transform 1 0 3736 0 1 3810
box -4 -6 100 206
use DFFPOSX1  _4367_
timestamp 1596991774
transform -1 0 4024 0 1 3810
box -4 -6 196 206
use OAI21X1  _3717_
timestamp 1596991774
transform 1 0 4024 0 1 3810
box -4 -6 68 206
use OAI21X1  _3716_
timestamp 1596991774
transform -1 0 4152 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert281
timestamp 1596991774
transform 1 0 4152 0 1 3810
box -4 -6 52 206
use INVX4  _3691_
timestamp 1596991774
transform -1 0 4248 0 1 3810
box -4 -6 52 206
use OAI21X1  _4137_
timestamp 1596991774
transform -1 0 4312 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert100
timestamp 1596991774
transform -1 0 4360 0 1 3810
box -4 -6 52 206
use FILL  SFILL43600x38100
timestamp 1596991774
transform 1 0 4360 0 1 3810
box -4 -6 20 206
use FILL  SFILL43760x38100
timestamp 1596991774
transform 1 0 4376 0 1 3810
box -4 -6 20 206
use FILL  SFILL43920x38100
timestamp 1596991774
transform 1 0 4392 0 1 3810
box -4 -6 20 206
use FILL  SFILL44080x38100
timestamp 1596991774
transform 1 0 4408 0 1 3810
box -4 -6 20 206
use DFFPOSX1  _4320_
timestamp 1596991774
transform -1 0 4616 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert131
timestamp 1596991774
transform -1 0 4664 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert285
timestamp 1596991774
transform 1 0 4664 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert72
timestamp 1596991774
transform 1 0 4712 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert62
timestamp 1596991774
transform -1 0 4808 0 1 3810
box -4 -6 52 206
use INVX4  _3694_
timestamp 1596991774
transform -1 0 4856 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert115
timestamp 1596991774
transform 1 0 4856 0 1 3810
box -4 -6 52 206
use NOR2X1  _4083_
timestamp 1596991774
transform -1 0 4952 0 1 3810
box -4 -6 52 206
use OAI22X1  _4085_
timestamp 1596991774
transform -1 0 5032 0 1 3810
box -4 -6 84 206
use OAI21X1  _4084_
timestamp 1596991774
transform -1 0 5096 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4347_
timestamp 1596991774
transform -1 0 5288 0 1 3810
box -4 -6 196 206
use NOR2X1  _3907_
timestamp 1596991774
transform 1 0 5288 0 1 3810
box -4 -6 52 206
use AOI21X1  _3908_
timestamp 1596991774
transform -1 0 5400 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4427_
timestamp 1596991774
transform -1 0 5592 0 1 3810
box -4 -6 196 206
use NOR2X1  _3897_
timestamp 1596991774
transform 1 0 5592 0 1 3810
box -4 -6 52 206
use AOI21X1  _3898_
timestamp 1596991774
transform -1 0 5704 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4342_
timestamp 1596991774
transform -1 0 5896 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert66
timestamp 1596991774
transform 1 0 5896 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert98
timestamp 1596991774
transform -1 0 6056 0 1 3810
box -4 -6 52 206
use FILL  SFILL59440x38100
timestamp 1596991774
transform 1 0 5944 0 1 3810
box -4 -6 20 206
use FILL  SFILL59600x38100
timestamp 1596991774
transform 1 0 5960 0 1 3810
box -4 -6 20 206
use FILL  SFILL59760x38100
timestamp 1596991774
transform 1 0 5976 0 1 3810
box -4 -6 20 206
use FILL  SFILL59920x38100
timestamp 1596991774
transform 1 0 5992 0 1 3810
box -4 -6 20 206
use MUX2X1  _4027_
timestamp 1596991774
transform -1 0 6152 0 1 3810
box -4 -6 100 206
use MUX2X1  _4205_
timestamp 1596991774
transform -1 0 6248 0 1 3810
box -4 -6 100 206
use BUFX2  BUFX2_insert116
timestamp 1596991774
transform -1 0 6296 0 1 3810
box -4 -6 52 206
use NOR2X1  _4268_
timestamp 1596991774
transform -1 0 6344 0 1 3810
box -4 -6 52 206
use AOI21X1  _4269_
timestamp 1596991774
transform -1 0 6408 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4412_
timestamp 1596991774
transform -1 0 6600 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert252
timestamp 1596991774
transform -1 0 6648 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert102
timestamp 1596991774
transform 1 0 6648 0 1 3810
box -4 -6 52 206
use NOR2X1  _4288_
timestamp 1596991774
transform 1 0 6696 0 1 3810
box -4 -6 52 206
use AOI21X1  _4289_
timestamp 1596991774
transform -1 0 6808 0 1 3810
box -4 -6 68 206
use AOI21X1  _3687_
timestamp 1596991774
transform 1 0 6808 0 1 3810
box -4 -6 68 206
use NOR2X1  _3686_
timestamp 1596991774
transform 1 0 6872 0 1 3810
box -4 -6 52 206
use DFFPOSX1  _4406_
timestamp 1596991774
transform -1 0 7112 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert151
timestamp 1596991774
transform 1 0 7112 0 1 3810
box -4 -6 52 206
use AOI21X1  _3890_
timestamp 1596991774
transform 1 0 7160 0 1 3810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert9
timestamp 1596991774
transform -1 0 7368 0 1 3810
box -4 -6 148 206
use FILL  FILL71120x38100
timestamp 1596991774
transform 1 0 7368 0 1 3810
box -4 -6 20 206
use FILL  FILL71280x38100
timestamp 1596991774
transform 1 0 7384 0 1 3810
box -4 -6 20 206
use INVX1  _2510_
timestamp 1596991774
transform 1 0 8 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2512_
timestamp 1596991774
transform -1 0 104 0 -1 4210
box -4 -6 68 206
use OR2X2  _2526_
timestamp 1596991774
transform 1 0 104 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2542_
timestamp 1596991774
transform -1 0 216 0 -1 4210
box -4 -6 52 206
use OAI21X1  _2531_
timestamp 1596991774
transform 1 0 216 0 -1 4210
box -4 -6 68 206
use NAND2X1  _2514_
timestamp 1596991774
transform -1 0 328 0 -1 4210
box -4 -6 52 206
use OR2X2  _2515_
timestamp 1596991774
transform 1 0 328 0 -1 4210
box -4 -6 68 206
use AND2X2  _2516_
timestamp 1596991774
transform 1 0 392 0 -1 4210
box -4 -6 68 206
use INVX1  _3204_
timestamp 1596991774
transform 1 0 456 0 -1 4210
box -4 -6 36 206
use BUFX2  BUFX2_insert199
timestamp 1596991774
transform -1 0 536 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2323_
timestamp 1596991774
transform -1 0 584 0 -1 4210
box -4 -6 52 206
use INVX1  _3256_
timestamp 1596991774
transform 1 0 584 0 -1 4210
box -4 -6 36 206
use NOR2X1  _2325_
timestamp 1596991774
transform 1 0 616 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert264
timestamp 1596991774
transform -1 0 712 0 -1 4210
box -4 -6 52 206
use INVX1  _2872_
timestamp 1596991774
transform 1 0 712 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2924_
timestamp 1596991774
transform -1 0 808 0 -1 4210
box -4 -6 68 206
use OAI21X1  _2878_
timestamp 1596991774
transform 1 0 808 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2879_
timestamp 1596991774
transform -1 0 920 0 -1 4210
box -4 -6 52 206
use NAND3X1  _2880_
timestamp 1596991774
transform 1 0 920 0 -1 4210
box -4 -6 68 206
use AND2X2  _2933_
timestamp 1596991774
transform 1 0 984 0 -1 4210
box -4 -6 68 206
use NAND3X1  _2939_
timestamp 1596991774
transform 1 0 1048 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2547_
timestamp 1596991774
transform 1 0 1112 0 -1 4210
box -4 -6 52 206
use NAND2X1  _2549_
timestamp 1596991774
transform -1 0 1208 0 -1 4210
box -4 -6 52 206
use INVX1  _2546_
timestamp 1596991774
transform -1 0 1240 0 -1 4210
box -4 -6 36 206
use XOR2X1  _2263_
timestamp 1596991774
transform 1 0 1240 0 -1 4210
box -4 -6 116 206
use BUFX2  BUFX2_insert2
timestamp 1596991774
transform -1 0 1400 0 -1 4210
box -4 -6 52 206
use FILL  SFILL14000x40100
timestamp 1596991774
transform -1 0 1416 0 -1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert198
timestamp 1596991774
transform 1 0 1464 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2378_
timestamp 1596991774
transform -1 0 1560 0 -1 4210
box -4 -6 52 206
use XOR2X1  _2376_
timestamp 1596991774
transform 1 0 1560 0 -1 4210
box -4 -6 116 206
use FILL  SFILL14160x40100
timestamp 1596991774
transform -1 0 1432 0 -1 4210
box -4 -6 20 206
use FILL  SFILL14320x40100
timestamp 1596991774
transform -1 0 1448 0 -1 4210
box -4 -6 20 206
use FILL  SFILL14480x40100
timestamp 1596991774
transform -1 0 1464 0 -1 4210
box -4 -6 20 206
use INVX1  _2855_
timestamp 1596991774
transform 1 0 1672 0 -1 4210
box -4 -6 36 206
use INVX1  _2595_
timestamp 1596991774
transform 1 0 1704 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2655_
timestamp 1596991774
transform 1 0 1736 0 -1 4210
box -4 -6 68 206
use NAND2X1  _2656_
timestamp 1596991774
transform -1 0 1848 0 -1 4210
box -4 -6 52 206
use AOI22X1  _2657_
timestamp 1596991774
transform 1 0 1848 0 -1 4210
box -4 -6 84 206
use NAND2X1  _2570_
timestamp 1596991774
transform 1 0 1928 0 -1 4210
box -4 -6 52 206
use INVX1  _2557_
timestamp 1596991774
transform 1 0 1976 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2558_
timestamp 1596991774
transform -1 0 2056 0 -1 4210
box -4 -6 52 206
use OAI21X1  _2652_
timestamp 1596991774
transform -1 0 2120 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2650_
timestamp 1596991774
transform -1 0 2168 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2651_
timestamp 1596991774
transform 1 0 2168 0 -1 4210
box -4 -6 52 206
use NAND2X1  _2574_
timestamp 1596991774
transform -1 0 2264 0 -1 4210
box -4 -6 52 206
use INVX1  _2569_
timestamp 1596991774
transform -1 0 2296 0 -1 4210
box -4 -6 36 206
use BUFX2  BUFX2_insert27
timestamp 1596991774
transform 1 0 2296 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert34
timestamp 1596991774
transform -1 0 2392 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert33
timestamp 1596991774
transform -1 0 2440 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert147
timestamp 1596991774
transform -1 0 2488 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert32
timestamp 1596991774
transform 1 0 2488 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4087_
timestamp 1596991774
transform 1 0 2536 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert263
timestamp 1596991774
transform 1 0 2600 0 -1 4210
box -4 -6 52 206
use AOI21X1  _4088_
timestamp 1596991774
transform -1 0 2712 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert223
timestamp 1596991774
transform -1 0 2760 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4210_
timestamp 1596991774
transform 1 0 2760 0 -1 4210
box -4 -6 68 206
use AOI21X1  _4211_
timestamp 1596991774
transform -1 0 2888 0 -1 4210
box -4 -6 68 206
use OAI21X1  _4265_
timestamp 1596991774
transform 1 0 2888 0 -1 4210
box -4 -6 68 206
use FILL  SFILL29520x40100
timestamp 1596991774
transform -1 0 2968 0 -1 4210
box -4 -6 20 206
use FILL  SFILL29680x40100
timestamp 1596991774
transform -1 0 2984 0 -1 4210
box -4 -6 20 206
use FILL  SFILL29840x40100
timestamp 1596991774
transform -1 0 3000 0 -1 4210
box -4 -6 20 206
use FILL  SFILL30000x40100
timestamp 1596991774
transform -1 0 3016 0 -1 4210
box -4 -6 20 206
use AOI21X1  _4266_
timestamp 1596991774
transform -1 0 3080 0 -1 4210
box -4 -6 68 206
use AOI21X1  _3817_
timestamp 1596991774
transform -1 0 3144 0 -1 4210
box -4 -6 68 206
use NOR2X1  _3816_
timestamp 1596991774
transform -1 0 3192 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4363_
timestamp 1596991774
transform -1 0 3384 0 -1 4210
box -4 -6 196 206
use NAND2X1  _3807_
timestamp 1596991774
transform 1 0 3384 0 -1 4210
box -4 -6 52 206
use OAI21X1  _3808_
timestamp 1596991774
transform -1 0 3496 0 -1 4210
box -4 -6 68 206
use MUX2X1  _4078_
timestamp 1596991774
transform 1 0 3496 0 -1 4210
box -4 -6 100 206
use MUX2X1  _4264_
timestamp 1596991774
transform -1 0 3688 0 -1 4210
box -4 -6 100 206
use BUFX2  BUFX2_insert89
timestamp 1596991774
transform -1 0 3736 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4081_
timestamp 1596991774
transform -1 0 3816 0 -1 4210
box -4 -6 84 206
use NOR2X1  _4079_
timestamp 1596991774
transform 1 0 3816 0 -1 4210
box -4 -6 52 206
use NAND2X1  _3773_
timestamp 1596991774
transform -1 0 3912 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4080_
timestamp 1596991774
transform 1 0 3912 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4379_
timestamp 1596991774
transform -1 0 4168 0 -1 4210
box -4 -6 196 206
use OAI21X1  _3741_
timestamp 1596991774
transform -1 0 4232 0 -1 4210
box -4 -6 68 206
use MUX2X1  _4209_
timestamp 1596991774
transform -1 0 4328 0 -1 4210
box -4 -6 100 206
use NOR2X1  _4202_
timestamp 1596991774
transform 1 0 4328 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4204_
timestamp 1596991774
transform -1 0 4456 0 -1 4210
box -4 -6 84 206
use OAI21X1  _4203_
timestamp 1596991774
transform -1 0 4584 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4326_
timestamp 1596991774
transform -1 0 4776 0 -1 4210
box -4 -6 196 206
use FILL  SFILL44560x40100
timestamp 1596991774
transform -1 0 4472 0 -1 4210
box -4 -6 20 206
use FILL  SFILL44720x40100
timestamp 1596991774
transform -1 0 4488 0 -1 4210
box -4 -6 20 206
use FILL  SFILL44880x40100
timestamp 1596991774
transform -1 0 4504 0 -1 4210
box -4 -6 20 206
use FILL  SFILL45040x40100
timestamp 1596991774
transform -1 0 4520 0 -1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert44
timestamp 1596991774
transform -1 0 4824 0 -1 4210
box -4 -6 52 206
use INVX8  _3911_
timestamp 1596991774
transform -1 0 4904 0 -1 4210
box -4 -6 84 206
use OAI22X1  _4030_
timestamp 1596991774
transform -1 0 4984 0 -1 4210
box -4 -6 84 206
use NOR2X1  _4028_
timestamp 1596991774
transform -1 0 5032 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4029_
timestamp 1596991774
transform -1 0 5096 0 -1 4210
box -4 -6 68 206
use OAI21X1  _4207_
timestamp 1596991774
transform 1 0 5096 0 -1 4210
box -4 -6 68 206
use OAI22X1  _4208_
timestamp 1596991774
transform 1 0 5160 0 -1 4210
box -4 -6 84 206
use NOR2X1  _4206_
timestamp 1596991774
transform -1 0 5288 0 -1 4210
box -4 -6 52 206
use MUX2X1  _4099_
timestamp 1596991774
transform -1 0 5384 0 -1 4210
box -4 -6 100 206
use NAND2X1  _3753_
timestamp 1596991774
transform 1 0 5384 0 -1 4210
box -4 -6 52 206
use OAI21X1  _3754_
timestamp 1596991774
transform -1 0 5496 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4321_
timestamp 1596991774
transform 1 0 5496 0 -1 4210
box -4 -6 196 206
use OAI21X1  _4148_
timestamp 1596991774
transform 1 0 5688 0 -1 4210
box -4 -6 68 206
use NOR2X1  _4147_
timestamp 1596991774
transform -1 0 5800 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4149_
timestamp 1596991774
transform 1 0 5800 0 -1 4210
box -4 -6 84 206
use NOR2X1  _3980_
timestamp 1596991774
transform -1 0 5928 0 -1 4210
box -4 -6 52 206
use NOR2X1  _4158_
timestamp 1596991774
transform -1 0 6040 0 -1 4210
box -4 -6 52 206
use FILL  SFILL59280x40100
timestamp 1596991774
transform -1 0 5944 0 -1 4210
box -4 -6 20 206
use FILL  SFILL59440x40100
timestamp 1596991774
transform -1 0 5960 0 -1 4210
box -4 -6 20 206
use FILL  SFILL59600x40100
timestamp 1596991774
transform -1 0 5976 0 -1 4210
box -4 -6 20 206
use FILL  SFILL59760x40100
timestamp 1596991774
transform -1 0 5992 0 -1 4210
box -4 -6 20 206
use OAI22X1  _4160_
timestamp 1596991774
transform 1 0 6040 0 -1 4210
box -4 -6 84 206
use OAI21X1  _4159_
timestamp 1596991774
transform -1 0 6184 0 -1 4210
box -4 -6 68 206
use MUX2X1  _4095_
timestamp 1596991774
transform -1 0 6280 0 -1 4210
box -4 -6 100 206
use OAI22X1  _4098_
timestamp 1596991774
transform -1 0 6360 0 -1 4210
box -4 -6 84 206
use OAI21X1  _4097_
timestamp 1596991774
transform -1 0 6424 0 -1 4210
box -4 -6 68 206
use NAND2X1  _3864_
timestamp 1596991774
transform -1 0 6472 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4310_
timestamp 1596991774
transform -1 0 6664 0 -1 4210
box -4 -6 196 206
use OAI21X1  _3865_
timestamp 1596991774
transform -1 0 6728 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4396_
timestamp 1596991774
transform -1 0 6920 0 -1 4210
box -4 -6 196 206
use NOR2X1  _3656_
timestamp 1596991774
transform 1 0 6920 0 -1 4210
box -4 -6 52 206
use AOI21X1  _3657_
timestamp 1596991774
transform -1 0 7032 0 -1 4210
box -4 -6 68 206
use AOI21X1  _3878_
timestamp 1596991774
transform 1 0 7032 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4332_
timestamp 1596991774
transform -1 0 7288 0 -1 4210
box -4 -6 196 206
use NAND3X1  _4530_
timestamp 1596991774
transform 1 0 7288 0 -1 4210
box -4 -6 68 206
use FILL  FILL70960x40100
timestamp 1596991774
transform -1 0 7368 0 -1 4210
box -4 -6 20 206
use FILL  FILL71120x40100
timestamp 1596991774
transform -1 0 7384 0 -1 4210
box -4 -6 20 206
use FILL  FILL71280x40100
timestamp 1596991774
transform -1 0 7400 0 -1 4210
box -4 -6 20 206
use AND2X2  _2499_
timestamp 1596991774
transform 1 0 8 0 1 4210
box -4 -6 68 206
use OAI21X1  _2502_
timestamp 1596991774
transform -1 0 136 0 1 4210
box -4 -6 68 206
use INVX1  _2501_
timestamp 1596991774
transform -1 0 168 0 1 4210
box -4 -6 36 206
use NAND2X1  _2511_
timestamp 1596991774
transform 1 0 168 0 1 4210
box -4 -6 52 206
use XOR2X1  _2508_
timestamp 1596991774
transform -1 0 328 0 1 4210
box -4 -6 116 206
use AOI21X1  _2530_
timestamp 1596991774
transform 1 0 328 0 1 4210
box -4 -6 68 206
use INVX1  _2527_
timestamp 1596991774
transform 1 0 392 0 1 4210
box -4 -6 36 206
use NAND2X1  _2525_
timestamp 1596991774
transform -1 0 472 0 1 4210
box -4 -6 52 206
use NAND2X1  _2519_
timestamp 1596991774
transform -1 0 520 0 1 4210
box -4 -6 52 206
use XOR2X1  _2524_
timestamp 1596991774
transform -1 0 632 0 1 4210
box -4 -6 116 206
use XNOR2X1  _2513_
timestamp 1596991774
transform -1 0 744 0 1 4210
box -4 -6 116 206
use AND2X2  _2324_
timestamp 1596991774
transform -1 0 808 0 1 4210
box -4 -6 68 206
use OAI22X1  _2925_
timestamp 1596991774
transform -1 0 888 0 1 4210
box -4 -6 84 206
use BUFX2  BUFX2_insert6
timestamp 1596991774
transform -1 0 936 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert262
timestamp 1596991774
transform -1 0 984 0 1 4210
box -4 -6 52 206
use INVX1  _2588_
timestamp 1596991774
transform -1 0 1016 0 1 4210
box -4 -6 36 206
use INVX1  _2873_
timestamp 1596991774
transform 1 0 1016 0 1 4210
box -4 -6 36 206
use OAI22X1  _2875_
timestamp 1596991774
transform 1 0 1048 0 1 4210
box -4 -6 84 206
use NAND2X1  _2877_
timestamp 1596991774
transform 1 0 1128 0 1 4210
box -4 -6 52 206
use INVX1  _2874_
timestamp 1596991774
transform -1 0 1208 0 1 4210
box -4 -6 36 206
use AOI21X1  _2931_
timestamp 1596991774
transform 1 0 1208 0 1 4210
box -4 -6 68 206
use NOR2X1  _2593_
timestamp 1596991774
transform -1 0 1320 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert261
timestamp 1596991774
transform 1 0 1320 0 1 4210
box -4 -6 52 206
use INVX1  _2580_
timestamp 1596991774
transform -1 0 1400 0 1 4210
box -4 -6 36 206
use FILL  SFILL14000x42100
timestamp 1596991774
transform 1 0 1400 0 1 4210
box -4 -6 20 206
use XOR2X1  _2377_
timestamp 1596991774
transform -1 0 1576 0 1 4210
box -4 -6 116 206
use BUFX2  BUFX2_insert7
timestamp 1596991774
transform 1 0 1576 0 1 4210
box -4 -6 52 206
use FILL  SFILL14160x42100
timestamp 1596991774
transform 1 0 1416 0 1 4210
box -4 -6 20 206
use FILL  SFILL14320x42100
timestamp 1596991774
transform 1 0 1432 0 1 4210
box -4 -6 20 206
use FILL  SFILL14480x42100
timestamp 1596991774
transform 1 0 1448 0 1 4210
box -4 -6 20 206
use NOR2X1  _2863_
timestamp 1596991774
transform 1 0 1624 0 1 4210
box -4 -6 52 206
use OAI21X1  _2930_
timestamp 1596991774
transform 1 0 1672 0 1 4210
box -4 -6 68 206
use NAND2X1  _2594_
timestamp 1596991774
transform -1 0 1784 0 1 4210
box -4 -6 52 206
use AOI21X1  _2929_
timestamp 1596991774
transform 1 0 1784 0 1 4210
box -4 -6 68 206
use NAND2X1  _2850_
timestamp 1596991774
transform 1 0 1848 0 1 4210
box -4 -6 52 206
use INVX1  _2849_
timestamp 1596991774
transform -1 0 1928 0 1 4210
box -4 -6 36 206
use NAND3X1  _2854_
timestamp 1596991774
transform -1 0 1992 0 1 4210
box -4 -6 68 206
use AOI21X1  _2928_
timestamp 1596991774
transform -1 0 2056 0 1 4210
box -4 -6 68 206
use INVX1  _2851_
timestamp 1596991774
transform -1 0 2088 0 1 4210
box -4 -6 36 206
use INVX1  _2852_
timestamp 1596991774
transform 1 0 2088 0 1 4210
box -4 -6 36 206
use AOI22X1  _2853_
timestamp 1596991774
transform 1 0 2120 0 1 4210
box -4 -6 84 206
use NAND3X1  _2575_
timestamp 1596991774
transform -1 0 2264 0 1 4210
box -4 -6 68 206
use OR2X2  _2573_
timestamp 1596991774
transform -1 0 2328 0 1 4210
box -4 -6 68 206
use INVX1  _2572_
timestamp 1596991774
transform -1 0 2360 0 1 4210
box -4 -6 36 206
use NAND2X1  _2848_
timestamp 1596991774
transform 1 0 2360 0 1 4210
box -4 -6 52 206
use INVX1  _2847_
timestamp 1596991774
transform -1 0 2440 0 1 4210
box -4 -6 36 206
use XNOR2X1  _2571_
timestamp 1596991774
transform -1 0 2552 0 1 4210
box -4 -6 116 206
use DFFPOSX1  _4459_
timestamp 1596991774
transform -1 0 2744 0 1 4210
box -4 -6 196 206
use DFFPOSX1  _4438_
timestamp 1596991774
transform -1 0 2936 0 1 4210
box -4 -6 196 206
use BUFX2  BUFX2_insert294
timestamp 1596991774
transform -1 0 3048 0 1 4210
box -4 -6 52 206
use FILL  SFILL29360x42100
timestamp 1596991774
transform 1 0 2936 0 1 4210
box -4 -6 20 206
use FILL  SFILL29520x42100
timestamp 1596991774
transform 1 0 2952 0 1 4210
box -4 -6 20 206
use FILL  SFILL29680x42100
timestamp 1596991774
transform 1 0 2968 0 1 4210
box -4 -6 20 206
use FILL  SFILL29840x42100
timestamp 1596991774
transform 1 0 2984 0 1 4210
box -4 -6 20 206
use DFFPOSX1  _4383_
timestamp 1596991774
transform 1 0 3048 0 1 4210
box -4 -6 196 206
use DFFPOSX1  _4395_
timestamp 1596991774
transform -1 0 3432 0 1 4210
box -4 -6 196 206
use AOI21X1  _3841_
timestamp 1596991774
transform 1 0 3432 0 1 4210
box -4 -6 68 206
use NOR2X1  _3840_
timestamp 1596991774
transform 1 0 3496 0 1 4210
box -4 -6 52 206
use MUX2X1  _4256_
timestamp 1596991774
transform -1 0 3640 0 1 4210
box -4 -6 100 206
use OAI22X1  _4259_
timestamp 1596991774
transform -1 0 3720 0 1 4210
box -4 -6 84 206
use OAI21X1  _4258_
timestamp 1596991774
transform -1 0 3784 0 1 4210
box -4 -6 68 206
use NOR2X1  _4257_
timestamp 1596991774
transform -1 0 3832 0 1 4210
box -4 -6 52 206
use OAI21X1  _3774_
timestamp 1596991774
transform 1 0 3832 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4331_
timestamp 1596991774
transform -1 0 4088 0 1 4210
box -4 -6 196 206
use BUFX2  BUFX2_insert278
timestamp 1596991774
transform -1 0 4136 0 1 4210
box -4 -6 52 206
use OAI21X1  _3740_
timestamp 1596991774
transform -1 0 4200 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert225
timestamp 1596991774
transform -1 0 4248 0 1 4210
box -4 -6 52 206
use NOR2X1  _4024_
timestamp 1596991774
transform -1 0 4296 0 1 4210
box -4 -6 52 206
use OAI22X1  _4026_
timestamp 1596991774
transform 1 0 4296 0 1 4210
box -4 -6 84 206
use MUX2X1  _4031_
timestamp 1596991774
transform 1 0 4376 0 1 4210
box -4 -6 100 206
use OAI21X1  _4025_
timestamp 1596991774
transform -1 0 4600 0 1 4210
box -4 -6 68 206
use NAND2X1  _3763_
timestamp 1596991774
transform 1 0 4600 0 1 4210
box -4 -6 52 206
use FILL  SFILL44720x42100
timestamp 1596991774
transform 1 0 4472 0 1 4210
box -4 -6 20 206
use FILL  SFILL44880x42100
timestamp 1596991774
transform 1 0 4488 0 1 4210
box -4 -6 20 206
use FILL  SFILL45040x42100
timestamp 1596991774
transform 1 0 4504 0 1 4210
box -4 -6 20 206
use FILL  SFILL45200x42100
timestamp 1596991774
transform 1 0 4520 0 1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert134
timestamp 1596991774
transform 1 0 4648 0 1 4210
box -4 -6 52 206
use OAI21X1  _3764_
timestamp 1596991774
transform -1 0 4760 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert46
timestamp 1596991774
transform -1 0 4808 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4315_
timestamp 1596991774
transform 1 0 4808 0 1 4210
box -4 -6 196 206
use NAND2X1  _3874_
timestamp 1596991774
transform 1 0 5000 0 1 4210
box -4 -6 52 206
use OAI21X1  _3875_
timestamp 1596991774
transform -1 0 5112 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert153
timestamp 1596991774
transform 1 0 5112 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert78
timestamp 1596991774
transform 1 0 5160 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert283
timestamp 1596991774
transform 1 0 5208 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert120
timestamp 1596991774
transform -1 0 5304 0 1 4210
box -4 -6 52 206
use MUX2X1  _3919_
timestamp 1596991774
transform -1 0 5400 0 1 4210
box -4 -6 100 206
use INVX4  _3688_
timestamp 1596991774
transform 1 0 5400 0 1 4210
box -4 -6 52 206
use OAI21X1  _3970_
timestamp 1596991774
transform 1 0 5448 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert47
timestamp 1596991774
transform 1 0 5512 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert282
timestamp 1596991774
transform 1 0 5560 0 1 4210
box -4 -6 52 206
use OAI22X1  _3971_
timestamp 1596991774
transform 1 0 5608 0 1 4210
box -4 -6 84 206
use NOR2X1  _3969_
timestamp 1596991774
transform -1 0 5736 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert92
timestamp 1596991774
transform 1 0 5736 0 1 4210
box -4 -6 52 206
use OAI21X1  _3981_
timestamp 1596991774
transform -1 0 5848 0 1 4210
box -4 -6 68 206
use OAI22X1  _3982_
timestamp 1596991774
transform 1 0 5848 0 1 4210
box -4 -6 84 206
use OAI21X1  _3917_
timestamp 1596991774
transform -1 0 6056 0 1 4210
box -4 -6 68 206
use FILL  SFILL59280x42100
timestamp 1596991774
transform 1 0 5928 0 1 4210
box -4 -6 20 206
use FILL  SFILL59440x42100
timestamp 1596991774
transform 1 0 5944 0 1 4210
box -4 -6 20 206
use FILL  SFILL59600x42100
timestamp 1596991774
transform 1 0 5960 0 1 4210
box -4 -6 20 206
use FILL  SFILL59760x42100
timestamp 1596991774
transform 1 0 5976 0 1 4210
box -4 -6 20 206
use OAI22X1  _3918_
timestamp 1596991774
transform 1 0 6056 0 1 4210
box -4 -6 84 206
use NOR2X1  _3916_
timestamp 1596991774
transform -1 0 6184 0 1 4210
box -4 -6 52 206
use MUX2X1  _3915_
timestamp 1596991774
transform -1 0 6280 0 1 4210
box -4 -6 100 206
use NOR2X1  _4096_
timestamp 1596991774
transform -1 0 6328 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4322_
timestamp 1596991774
transform -1 0 6520 0 1 4210
box -4 -6 196 206
use NAND2X1  _3755_
timestamp 1596991774
transform 1 0 6520 0 1 4210
box -4 -6 52 206
use OAI21X1  _3756_
timestamp 1596991774
transform -1 0 6632 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert132
timestamp 1596991774
transform -1 0 6680 0 1 4210
box -4 -6 52 206
use MUX2X1  _3979_
timestamp 1596991774
transform 1 0 6680 0 1 4210
box -4 -6 100 206
use OAI21X1  _3845_
timestamp 1596991774
transform 1 0 6776 0 1 4210
box -4 -6 68 206
use NAND2X1  _3844_
timestamp 1596991774
transform -1 0 6888 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4300_
timestamp 1596991774
transform -1 0 7080 0 1 4210
box -4 -6 196 206
use NAND2X1  _3789_
timestamp 1596991774
transform 1 0 7080 0 1 4210
box -4 -6 52 206
use OAI21X1  _3790_
timestamp 1596991774
transform -1 0 7192 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4354_
timestamp 1596991774
transform -1 0 7384 0 1 4210
box -4 -6 196 206
use FILL  FILL71280x42100
timestamp 1596991774
transform 1 0 7384 0 1 4210
box -4 -6 20 206
use OR2X2  _2498_
timestamp 1596991774
transform -1 0 72 0 -1 4610
box -4 -6 68 206
use OAI21X1  _2509_
timestamp 1596991774
transform 1 0 72 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2507_
timestamp 1596991774
transform 1 0 136 0 -1 4610
box -4 -6 52 206
use INVX1  _2506_
timestamp 1596991774
transform 1 0 184 0 -1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert29
timestamp 1596991774
transform -1 0 264 0 -1 4610
box -4 -6 52 206
use INVX1  _2528_
timestamp 1596991774
transform -1 0 296 0 -1 4610
box -4 -6 36 206
use NOR2X1  _2523_
timestamp 1596991774
transform -1 0 344 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2529_
timestamp 1596991774
transform -1 0 408 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2326_
timestamp 1596991774
transform -1 0 456 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2328_
timestamp 1596991774
transform 1 0 456 0 -1 4610
box -4 -6 52 206
use NAND2X1  _2518_
timestamp 1596991774
transform 1 0 504 0 -1 4610
box -4 -6 52 206
use INVX1  _2517_
timestamp 1596991774
transform -1 0 584 0 -1 4610
box -4 -6 36 206
use INVX1  _2869_
timestamp 1596991774
transform 1 0 584 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2870_
timestamp 1596991774
transform -1 0 664 0 -1 4610
box -4 -6 52 206
use NAND3X1  _2871_
timestamp 1596991774
transform 1 0 664 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert169
timestamp 1596991774
transform -1 0 776 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert30
timestamp 1596991774
transform 1 0 776 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert5
timestamp 1596991774
transform -1 0 872 0 -1 4610
box -4 -6 52 206
use INVX1  _2590_
timestamp 1596991774
transform -1 0 904 0 -1 4610
box -4 -6 36 206
use AOI22X1  _2591_
timestamp 1596991774
transform 1 0 904 0 -1 4610
box -4 -6 84 206
use OR2X2  _2589_
timestamp 1596991774
transform 1 0 984 0 -1 4610
box -4 -6 68 206
use NAND3X1  _2592_
timestamp 1596991774
transform -1 0 1112 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert59
timestamp 1596991774
transform -1 0 1160 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert4
timestamp 1596991774
transform -1 0 1208 0 -1 4610
box -4 -6 52 206
use NAND2X1  _2581_
timestamp 1596991774
transform 1 0 1208 0 -1 4610
box -4 -6 52 206
use NAND3X1  _2585_
timestamp 1596991774
transform 1 0 1256 0 -1 4610
box -4 -6 68 206
use NAND3X1  _2643_
timestamp 1596991774
transform -1 0 1384 0 -1 4610
box -4 -6 68 206
use FILL  SFILL13840x44100
timestamp 1596991774
transform -1 0 1400 0 -1 4610
box -4 -6 20 206
use FILL  SFILL14000x44100
timestamp 1596991774
transform -1 0 1416 0 -1 4610
box -4 -6 20 206
use OAI22X1  _2644_
timestamp 1596991774
transform -1 0 1528 0 -1 4610
box -4 -6 84 206
use AOI22X1  _2639_
timestamp 1596991774
transform -1 0 1608 0 -1 4610
box -4 -6 84 206
use NOR2X1  _2640_
timestamp 1596991774
transform -1 0 1656 0 -1 4610
box -4 -6 52 206
use FILL  SFILL14160x44100
timestamp 1596991774
transform -1 0 1432 0 -1 4610
box -4 -6 20 206
use FILL  SFILL14320x44100
timestamp 1596991774
transform -1 0 1448 0 -1 4610
box -4 -6 20 206
use INVX1  _2638_
timestamp 1596991774
transform -1 0 1688 0 -1 4610
box -4 -6 36 206
use OAI21X1  _2927_
timestamp 1596991774
transform -1 0 1752 0 -1 4610
box -4 -6 68 206
use NAND3X1  _2862_
timestamp 1596991774
transform -1 0 1816 0 -1 4610
box -4 -6 68 206
use AOI21X1  _2654_
timestamp 1596991774
transform 1 0 1816 0 -1 4610
box -4 -6 68 206
use AOI22X1  _2857_
timestamp 1596991774
transform 1 0 1880 0 -1 4610
box -4 -6 84 206
use INVX1  _2856_
timestamp 1596991774
transform -1 0 1992 0 -1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert103
timestamp 1596991774
transform -1 0 2040 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2653_
timestamp 1596991774
transform -1 0 2104 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2579_
timestamp 1596991774
transform -1 0 2152 0 -1 4610
box -4 -6 52 206
use XNOR2X1  _2576_
timestamp 1596991774
transform -1 0 2264 0 -1 4610
box -4 -6 116 206
use BUFX2  BUFX2_insert87
timestamp 1596991774
transform -1 0 2312 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert85
timestamp 1596991774
transform -1 0 2360 0 -1 4610
box -4 -6 52 206
use DFFPOSX1  _4454_
timestamp 1596991774
transform -1 0 2552 0 -1 4610
box -4 -6 196 206
use OAI21X1  _4065_
timestamp 1596991774
transform 1 0 2552 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert145
timestamp 1596991774
transform 1 0 2616 0 -1 4610
box -4 -6 52 206
use OAI21X1  _4032_
timestamp 1596991774
transform -1 0 2728 0 -1 4610
box -4 -6 68 206
use AOI21X1  _4033_
timestamp 1596991774
transform -1 0 2792 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4442_
timestamp 1596991774
transform -1 0 2984 0 -1 4610
box -4 -6 196 206
use FILL  SFILL29840x44100
timestamp 1596991774
transform -1 0 3000 0 -1 4610
box -4 -6 20 206
use FILL  SFILL30000x44100
timestamp 1596991774
transform -1 0 3016 0 -1 4610
box -4 -6 20 206
use DFFPOSX1  _4443_
timestamp 1596991774
transform -1 0 3240 0 -1 4610
box -4 -6 196 206
use FILL  SFILL30160x44100
timestamp 1596991774
transform -1 0 3032 0 -1 4610
box -4 -6 20 206
use FILL  SFILL30320x44100
timestamp 1596991774
transform -1 0 3048 0 -1 4610
box -4 -6 20 206
use BUFX2  BUFX2_insert222
timestamp 1596991774
transform -1 0 3288 0 -1 4610
box -4 -6 52 206
use NAND2X1  _3797_
timestamp 1596991774
transform -1 0 3336 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3798_
timestamp 1596991774
transform -1 0 3400 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4358_
timestamp 1596991774
transform 1 0 3400 0 -1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert140
timestamp 1596991774
transform -1 0 3640 0 -1 4610
box -4 -6 52 206
use OAI22X1  _4252_
timestamp 1596991774
transform -1 0 3720 0 -1 4610
box -4 -6 84 206
use NOR2X1  _4250_
timestamp 1596991774
transform 1 0 3720 0 -1 4610
box -4 -6 52 206
use OAI21X1  _4251_
timestamp 1596991774
transform -1 0 3832 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4346_
timestamp 1596991774
transform -1 0 4024 0 -1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert141
timestamp 1596991774
transform 1 0 4024 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert79
timestamp 1596991774
transform -1 0 4120 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert206
timestamp 1596991774
transform -1 0 4168 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3831_
timestamp 1596991774
transform 1 0 4168 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3830_
timestamp 1596991774
transform -1 0 4280 0 -1 4610
box -4 -6 52 206
use MUX2X1  _4023_
timestamp 1596991774
transform 1 0 4280 0 -1 4610
box -4 -6 100 206
use MUX2X1  _4201_
timestamp 1596991774
transform -1 0 4472 0 -1 4610
box -4 -6 100 206
use OAI21X1  _3730_
timestamp 1596991774
transform 1 0 4536 0 -1 4610
box -4 -6 68 206
use OAI21X1  _3731_
timestamp 1596991774
transform -1 0 4664 0 -1 4610
box -4 -6 68 206
use FILL  SFILL44720x44100
timestamp 1596991774
transform -1 0 4488 0 -1 4610
box -4 -6 20 206
use FILL  SFILL44880x44100
timestamp 1596991774
transform -1 0 4504 0 -1 4610
box -4 -6 20 206
use FILL  SFILL45040x44100
timestamp 1596991774
transform -1 0 4520 0 -1 4610
box -4 -6 20 206
use FILL  SFILL45200x44100
timestamp 1596991774
transform -1 0 4536 0 -1 4610
box -4 -6 20 206
use DFFPOSX1  _4374_
timestamp 1596991774
transform -1 0 4856 0 -1 4610
box -4 -6 196 206
use DFFPOSX1  _4393_
timestamp 1596991774
transform 1 0 4856 0 -1 4610
box -4 -6 196 206
use AOI21X1  _3837_
timestamp 1596991774
transform 1 0 5048 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3836_
timestamp 1596991774
transform 1 0 5112 0 -1 4610
box -4 -6 52 206
use NOR2X1  _3810_
timestamp 1596991774
transform -1 0 5208 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3811_
timestamp 1596991774
transform -1 0 5272 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4380_
timestamp 1596991774
transform 1 0 5272 0 -1 4610
box -4 -6 196 206
use OAI21X1  _4093_
timestamp 1596991774
transform -1 0 5528 0 -1 4610
box -4 -6 68 206
use OAI22X1  _4094_
timestamp 1596991774
transform -1 0 5608 0 -1 4610
box -4 -6 84 206
use MUX2X1  _4090_
timestamp 1596991774
transform 1 0 5608 0 -1 4610
box -4 -6 100 206
use MUX2X1  _3910_
timestamp 1596991774
transform 1 0 5704 0 -1 4610
box -4 -6 100 206
use OAI21X1  _3913_
timestamp 1596991774
transform 1 0 5800 0 -1 4610
box -4 -6 68 206
use OAI22X1  _3914_
timestamp 1596991774
transform -1 0 5944 0 -1 4610
box -4 -6 84 206
use NOR2X1  _3912_
timestamp 1596991774
transform -1 0 6056 0 -1 4610
box -4 -6 52 206
use FILL  SFILL59440x44100
timestamp 1596991774
transform -1 0 5960 0 -1 4610
box -4 -6 20 206
use FILL  SFILL59600x44100
timestamp 1596991774
transform -1 0 5976 0 -1 4610
box -4 -6 20 206
use FILL  SFILL59760x44100
timestamp 1596991774
transform -1 0 5992 0 -1 4610
box -4 -6 20 206
use FILL  SFILL59920x44100
timestamp 1596991774
transform -1 0 6008 0 -1 4610
box -4 -6 20 206
use NOR2X1  _4092_
timestamp 1596991774
transform 1 0 6056 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3721_
timestamp 1596991774
transform 1 0 6104 0 -1 4610
box -4 -6 68 206
use OAI21X1  _3720_
timestamp 1596991774
transform -1 0 6232 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert226
timestamp 1596991774
transform 1 0 6232 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3722_
timestamp 1596991774
transform 1 0 6280 0 -1 4610
box -4 -6 68 206
use OAI21X1  _3723_
timestamp 1596991774
transform -1 0 6408 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4370_
timestamp 1596991774
transform -1 0 6600 0 -1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert77
timestamp 1596991774
transform -1 0 6648 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert256
timestamp 1596991774
transform 1 0 6648 0 -1 4610
box -4 -6 52 206
use MUX2X1  _4157_
timestamp 1596991774
transform 1 0 6696 0 -1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert144
timestamp 1596991774
transform 1 0 6792 0 -1 4610
box -4 -6 52 206
use MUX2X1  _3968_
timestamp 1596991774
transform 1 0 6840 0 -1 4610
box -4 -6 100 206
use MUX2X1  _4146_
timestamp 1596991774
transform 1 0 6936 0 -1 4610
box -4 -6 100 206
use AOI21X1  _3821_
timestamp 1596991774
transform 1 0 7032 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3820_
timestamp 1596991774
transform 1 0 7096 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3823_
timestamp 1596991774
transform 1 0 7144 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3822_
timestamp 1596991774
transform 1 0 7208 0 -1 4610
box -4 -6 52 206
use BUFX2  _2085_
timestamp 1596991774
transform 1 0 7256 0 -1 4610
box -4 -6 52 206
use BUFX2  _2088_
timestamp 1596991774
transform 1 0 7304 0 -1 4610
box -4 -6 52 206
use FILL  FILL70960x44100
timestamp 1596991774
transform -1 0 7368 0 -1 4610
box -4 -6 20 206
use FILL  FILL71120x44100
timestamp 1596991774
transform -1 0 7384 0 -1 4610
box -4 -6 20 206
use FILL  FILL71280x44100
timestamp 1596991774
transform -1 0 7400 0 -1 4610
box -4 -6 20 206
use NAND2X1  _2497_
timestamp 1596991774
transform 1 0 8 0 1 4610
box -4 -6 52 206
use INVX1  _2496_
timestamp 1596991774
transform -1 0 88 0 1 4610
box -4 -6 36 206
use NOR2X1  _2504_
timestamp 1596991774
transform 1 0 88 0 1 4610
box -4 -6 52 206
use INVX1  _2503_
timestamp 1596991774
transform -1 0 168 0 1 4610
box -4 -6 36 206
use NAND2X1  _2505_
timestamp 1596991774
transform -1 0 216 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert235
timestamp 1596991774
transform -1 0 264 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert57
timestamp 1596991774
transform -1 0 312 0 1 4610
box -4 -6 52 206
use AND2X2  _2522_
timestamp 1596991774
transform -1 0 376 0 1 4610
box -4 -6 68 206
use NOR2X1  _2521_
timestamp 1596991774
transform 1 0 376 0 1 4610
box -4 -6 52 206
use INVX1  _2520_
timestamp 1596991774
transform -1 0 456 0 1 4610
box -4 -6 36 206
use INVX1  _2777_
timestamp 1596991774
transform -1 0 488 0 1 4610
box -4 -6 36 206
use AND2X2  _2327_
timestamp 1596991774
transform -1 0 552 0 1 4610
box -4 -6 68 206
use INVX1  _2864_
timestamp 1596991774
transform 1 0 552 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert197
timestamp 1596991774
transform 1 0 584 0 1 4610
box -4 -6 52 206
use NAND2X1  _2868_
timestamp 1596991774
transform -1 0 680 0 1 4610
box -4 -6 52 206
use INVX1  _2865_
timestamp 1596991774
transform 1 0 680 0 1 4610
box -4 -6 36 206
use AOI22X1  _2866_
timestamp 1596991774
transform -1 0 792 0 1 4610
box -4 -6 84 206
use NOR2X1  _2923_
timestamp 1596991774
transform -1 0 840 0 1 4610
box -4 -6 52 206
use INVX1  _2682_
timestamp 1596991774
transform 1 0 840 0 1 4610
box -4 -6 36 206
use OAI22X1  _2683_
timestamp 1596991774
transform -1 0 952 0 1 4610
box -4 -6 84 206
use INVX1  _2681_
timestamp 1596991774
transform -1 0 984 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert237
timestamp 1596991774
transform 1 0 984 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert195
timestamp 1596991774
transform -1 0 1080 0 1 4610
box -4 -6 52 206
use INVX1  _2586_
timestamp 1596991774
transform 1 0 1080 0 1 4610
box -4 -6 36 206
use NAND2X1  _2587_
timestamp 1596991774
transform -1 0 1160 0 1 4610
box -4 -6 52 206
use AOI22X1  _2642_
timestamp 1596991774
transform -1 0 1240 0 1 4610
box -4 -6 84 206
use INVX1  _2641_
timestamp 1596991774
transform -1 0 1272 0 1 4610
box -4 -6 36 206
use XNOR2X1  _2584_
timestamp 1596991774
transform -1 0 1384 0 1 4610
box -4 -6 116 206
use INVX1  _2582_
timestamp 1596991774
transform 1 0 1384 0 1 4610
box -4 -6 36 206
use NAND2X1  _2583_
timestamp 1596991774
transform -1 0 1528 0 1 4610
box -4 -6 52 206
use NAND2X1  _2761_
timestamp 1596991774
transform -1 0 1576 0 1 4610
box -4 -6 52 206
use AOI22X1  _2760_
timestamp 1596991774
transform -1 0 1656 0 1 4610
box -4 -6 84 206
use FILL  SFILL14160x46100
timestamp 1596991774
transform 1 0 1416 0 1 4610
box -4 -6 20 206
use FILL  SFILL14320x46100
timestamp 1596991774
transform 1 0 1432 0 1 4610
box -4 -6 20 206
use FILL  SFILL14480x46100
timestamp 1596991774
transform 1 0 1448 0 1 4610
box -4 -6 20 206
use FILL  SFILL14640x46100
timestamp 1596991774
transform 1 0 1464 0 1 4610
box -4 -6 20 206
use OAI22X1  _2926_
timestamp 1596991774
transform 1 0 1656 0 1 4610
box -4 -6 84 206
use INVX1  _2860_
timestamp 1596991774
transform 1 0 1736 0 1 4610
box -4 -6 36 206
use NAND2X1  _2861_
timestamp 1596991774
transform 1 0 1768 0 1 4610
box -4 -6 52 206
use NAND2X1  _2859_
timestamp 1596991774
transform -1 0 1864 0 1 4610
box -4 -6 52 206
use INVX1  _2858_
timestamp 1596991774
transform -1 0 1896 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert0
timestamp 1596991774
transform -1 0 1944 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert247
timestamp 1596991774
transform -1 0 1992 0 1 4610
box -4 -6 52 206
use INVX1  _2762_
timestamp 1596991774
transform 1 0 1992 0 1 4610
box -4 -6 36 206
use XNOR2X1  _2577_
timestamp 1596991774
transform -1 0 2136 0 1 4610
box -4 -6 116 206
use NAND2X1  _2578_
timestamp 1596991774
transform -1 0 2184 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert3
timestamp 1596991774
transform 1 0 2184 0 1 4610
box -4 -6 52 206
use OAI21X1  _2649_
timestamp 1596991774
transform 1 0 2232 0 1 4610
box -4 -6 68 206
use INVX1  _2645_
timestamp 1596991774
transform -1 0 2328 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert31
timestamp 1596991774
transform -1 0 2376 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4457_
timestamp 1596991774
transform -1 0 2568 0 1 4610
box -4 -6 196 206
use AOI21X1  _4066_
timestamp 1596991774
transform -1 0 2632 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert249
timestamp 1596991774
transform -1 0 2680 0 1 4610
box -4 -6 52 206
use OAI21X1  _4254_
timestamp 1596991774
transform 1 0 2680 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert218
timestamp 1596991774
transform -1 0 2792 0 1 4610
box -4 -6 52 206
use OAI21X1  _4243_
timestamp 1596991774
transform 1 0 2792 0 1 4610
box -4 -6 68 206
use AOI21X1  _4255_
timestamp 1596991774
transform -1 0 2920 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert292
timestamp 1596991774
transform -1 0 3032 0 1 4610
box -4 -6 52 206
use FILL  SFILL29200x46100
timestamp 1596991774
transform 1 0 2920 0 1 4610
box -4 -6 20 206
use FILL  SFILL29360x46100
timestamp 1596991774
transform 1 0 2936 0 1 4610
box -4 -6 20 206
use FILL  SFILL29520x46100
timestamp 1596991774
transform 1 0 2952 0 1 4610
box -4 -6 20 206
use FILL  SFILL29680x46100
timestamp 1596991774
transform 1 0 2968 0 1 4610
box -4 -6 20 206
use DFFPOSX1  _4441_
timestamp 1596991774
transform -1 0 3224 0 1 4610
box -4 -6 196 206
use AOI21X1  _4244_
timestamp 1596991774
transform -1 0 3288 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4314_
timestamp 1596991774
transform 1 0 3288 0 1 4610
box -4 -6 196 206
use MUX2X1  _4253_
timestamp 1596991774
transform -1 0 3576 0 1 4610
box -4 -6 100 206
use NAND2X1  _3872_
timestamp 1596991774
transform 1 0 3576 0 1 4610
box -4 -6 52 206
use OAI21X1  _3873_
timestamp 1596991774
transform -1 0 3688 0 1 4610
box -4 -6 68 206
use OAI22X1  _4074_
timestamp 1596991774
transform -1 0 3768 0 1 4610
box -4 -6 84 206
use NOR2X1  _4072_
timestamp 1596991774
transform 1 0 3768 0 1 4610
box -4 -6 52 206
use OAI21X1  _4073_
timestamp 1596991774
transform -1 0 3880 0 1 4610
box -4 -6 68 206
use NOR2X1  _3905_
timestamp 1596991774
transform 1 0 3880 0 1 4610
box -4 -6 52 206
use AOI21X1  _3906_
timestamp 1596991774
transform -1 0 3992 0 1 4610
box -4 -6 68 206
use OAI21X1  _3869_
timestamp 1596991774
transform 1 0 3992 0 1 4610
box -4 -6 68 206
use NAND2X1  _3868_
timestamp 1596991774
transform -1 0 4104 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4312_
timestamp 1596991774
transform -1 0 4296 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4390_
timestamp 1596991774
transform 1 0 4296 0 1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert208
timestamp 1596991774
transform -1 0 4600 0 1 4610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert16
timestamp 1596991774
transform -1 0 4744 0 1 4610
box -4 -6 148 206
use FILL  SFILL44880x46100
timestamp 1596991774
transform 1 0 4488 0 1 4610
box -4 -6 20 206
use FILL  SFILL45040x46100
timestamp 1596991774
transform 1 0 4504 0 1 4610
box -4 -6 20 206
use FILL  SFILL45200x46100
timestamp 1596991774
transform 1 0 4520 0 1 4610
box -4 -6 20 206
use FILL  SFILL45360x46100
timestamp 1596991774
transform 1 0 4536 0 1 4610
box -4 -6 20 206
use BUFX2  BUFX2_insert121
timestamp 1596991774
transform -1 0 4792 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4329_
timestamp 1596991774
transform -1 0 4984 0 1 4610
box -4 -6 196 206
use NAND2X1  _3769_
timestamp 1596991774
transform 1 0 4984 0 1 4610
box -4 -6 52 206
use OAI21X1  _3770_
timestamp 1596991774
transform -1 0 5096 0 1 4610
box -4 -6 68 206
use MUX2X1  _4234_
timestamp 1596991774
transform 1 0 5096 0 1 4610
box -4 -6 100 206
use MUX2X1  _4056_
timestamp 1596991774
transform 1 0 5192 0 1 4610
box -4 -6 100 206
use OAI21X1  _3744_
timestamp 1596991774
transform 1 0 5288 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4316_
timestamp 1596991774
transform 1 0 5352 0 1 4610
box -4 -6 196 206
use NAND2X1  _3743_
timestamp 1596991774
transform -1 0 5592 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4348_
timestamp 1596991774
transform -1 0 5784 0 1 4610
box -4 -6 196 206
use NAND2X1  _3777_
timestamp 1596991774
transform 1 0 5784 0 1 4610
box -4 -6 52 206
use OAI21X1  _3778_
timestamp 1596991774
transform -1 0 5896 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert209
timestamp 1596991774
transform 1 0 5896 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4369_
timestamp 1596991774
transform -1 0 6200 0 1 4610
box -4 -6 196 206
use FILL  SFILL59440x46100
timestamp 1596991774
transform 1 0 5944 0 1 4610
box -4 -6 20 206
use FILL  SFILL59600x46100
timestamp 1596991774
transform 1 0 5960 0 1 4610
box -4 -6 20 206
use FILL  SFILL59760x46100
timestamp 1596991774
transform 1 0 5976 0 1 4610
box -4 -6 20 206
use FILL  SFILL59920x46100
timestamp 1596991774
transform 1 0 5992 0 1 4610
box -4 -6 20 206
use BUFX2  BUFX2_insert118
timestamp 1596991774
transform 1 0 6200 0 1 4610
box -4 -6 52 206
use OAI21X1  _3710_
timestamp 1596991774
transform 1 0 6248 0 1 4610
box -4 -6 68 206
use OAI21X1  _3711_
timestamp 1596991774
transform -1 0 6376 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4364_
timestamp 1596991774
transform -1 0 6568 0 1 4610
box -4 -6 196 206
use NAND2X1  _3765_
timestamp 1596991774
transform -1 0 6616 0 1 4610
box -4 -6 52 206
use OAI21X1  _3766_
timestamp 1596991774
transform -1 0 6680 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert26
timestamp 1596991774
transform -1 0 6728 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4327_
timestamp 1596991774
transform 1 0 6728 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4385_
timestamp 1596991774
transform -1 0 7112 0 1 4610
box -4 -6 196 206
use OAI21X1  _3788_
timestamp 1596991774
transform 1 0 7112 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4353_
timestamp 1596991774
transform -1 0 7368 0 1 4610
box -4 -6 196 206
use FILL  FILL71120x46100
timestamp 1596991774
transform 1 0 7368 0 1 4610
box -4 -6 20 206
use FILL  FILL71280x46100
timestamp 1596991774
transform 1 0 7384 0 1 4610
box -4 -6 20 206
use BUFX2  _2112_
timestamp 1596991774
transform -1 0 56 0 -1 5010
box -4 -6 52 206
use NAND2X1  _2785_
timestamp 1596991774
transform 1 0 56 0 -1 5010
box -4 -6 52 206
use INVX1  _2784_
timestamp 1596991774
transform -1 0 136 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2788_
timestamp 1596991774
transform -1 0 216 0 -1 5010
box -4 -6 84 206
use INVX1  _2787_
timestamp 1596991774
transform -1 0 248 0 -1 5010
box -4 -6 36 206
use INVX1  _2684_
timestamp 1596991774
transform 1 0 248 0 -1 5010
box -4 -6 36 206
use OR2X2  _2830_
timestamp 1596991774
transform -1 0 344 0 -1 5010
box -4 -6 68 206
use INVX1  _2776_
timestamp 1596991774
transform 1 0 344 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2778_
timestamp 1596991774
transform 1 0 376 0 -1 5010
box -4 -6 84 206
use NAND2X1  _2780_
timestamp 1596991774
transform -1 0 504 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert158
timestamp 1596991774
transform -1 0 552 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert159
timestamp 1596991774
transform -1 0 600 0 -1 5010
box -4 -6 52 206
use INVX1  _2867_
timestamp 1596991774
transform 1 0 600 0 -1 5010
box -4 -6 36 206
use OAI21X1  _2737_
timestamp 1596991774
transform 1 0 632 0 -1 5010
box -4 -6 68 206
use INVX1  _2685_
timestamp 1596991774
transform 1 0 696 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2686_
timestamp 1596991774
transform 1 0 728 0 -1 5010
box -4 -6 84 206
use INVX1  _2677_
timestamp 1596991774
transform -1 0 840 0 -1 5010
box -4 -6 36 206
use AOI22X1  _2732_
timestamp 1596991774
transform 1 0 840 0 -1 5010
box -4 -6 84 206
use INVX1  _2678_
timestamp 1596991774
transform -1 0 952 0 -1 5010
box -4 -6 36 206
use NOR2X1  _2687_
timestamp 1596991774
transform -1 0 1000 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert160
timestamp 1596991774
transform -1 0 1048 0 -1 5010
box -4 -6 52 206
use NAND2X1  _2751_
timestamp 1596991774
transform 1 0 1048 0 -1 5010
box -4 -6 52 206
use AND2X2  _2688_
timestamp 1596991774
transform 1 0 1096 0 -1 5010
box -4 -6 68 206
use OAI21X1  _2746_
timestamp 1596991774
transform -1 0 1224 0 -1 5010
box -4 -6 68 206
use NOR2X1  _2791_
timestamp 1596991774
transform -1 0 1272 0 -1 5010
box -4 -6 52 206
use INVX1  _2829_
timestamp 1596991774
transform 1 0 1272 0 -1 5010
box -4 -6 36 206
use AOI21X1  _2839_
timestamp 1596991774
transform 1 0 1304 0 -1 5010
box -4 -6 68 206
use INVX1  _2665_
timestamp 1596991774
transform 1 0 1368 0 -1 5010
box -4 -6 36 206
use FILL  SFILL14000x48100
timestamp 1596991774
transform -1 0 1416 0 -1 5010
box -4 -6 20 206
use NAND2X1  _2668_
timestamp 1596991774
transform -1 0 1512 0 -1 5010
box -4 -6 52 206
use AOI21X1  _2749_
timestamp 1596991774
transform 1 0 1512 0 -1 5010
box -4 -6 68 206
use OAI22X1  _2667_
timestamp 1596991774
transform 1 0 1576 0 -1 5010
box -4 -6 84 206
use FILL  SFILL14160x48100
timestamp 1596991774
transform -1 0 1432 0 -1 5010
box -4 -6 20 206
use FILL  SFILL14320x48100
timestamp 1596991774
transform -1 0 1448 0 -1 5010
box -4 -6 20 206
use FILL  SFILL14480x48100
timestamp 1596991774
transform -1 0 1464 0 -1 5010
box -4 -6 20 206
use NAND2X1  _2671_
timestamp 1596991774
transform -1 0 1704 0 -1 5010
box -4 -6 52 206
use OAI22X1  _2748_
timestamp 1596991774
transform 1 0 1704 0 -1 5010
box -4 -6 84 206
use INVX1  _2666_
timestamp 1596991774
transform -1 0 1816 0 -1 5010
box -4 -6 36 206
use INVX1  _2747_
timestamp 1596991774
transform -1 0 1848 0 -1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert43
timestamp 1596991774
transform -1 0 1896 0 -1 5010
box -4 -6 52 206
use OAI21X1  _2838_
timestamp 1596991774
transform -1 0 1960 0 -1 5010
box -4 -6 68 206
use INVX1  _2769_
timestamp 1596991774
transform -1 0 1992 0 -1 5010
box -4 -6 36 206
use NAND3X1  _2775_
timestamp 1596991774
transform 1 0 1992 0 -1 5010
box -4 -6 68 206
use OAI21X1  _2834_
timestamp 1596991774
transform -1 0 2120 0 -1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert105
timestamp 1596991774
transform 1 0 2120 0 -1 5010
box -4 -6 52 206
use INVX1  _2773_
timestamp 1596991774
transform 1 0 2168 0 -1 5010
box -4 -6 36 206
use AOI22X1  _2774_
timestamp 1596991774
transform -1 0 2280 0 -1 5010
box -4 -6 84 206
use INVX1  _2772_
timestamp 1596991774
transform -1 0 2312 0 -1 5010
box -4 -6 36 206
use INVX1  _2647_
timestamp 1596991774
transform 1 0 2312 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2648_
timestamp 1596991774
transform -1 0 2424 0 -1 5010
box -4 -6 84 206
use INVX1  _2646_
timestamp 1596991774
transform 1 0 2424 0 -1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert161
timestamp 1596991774
transform 1 0 2456 0 -1 5010
box -4 -6 52 206
use OAI21X1  _4043_
timestamp 1596991774
transform 1 0 2504 0 -1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert40
timestamp 1596991774
transform -1 0 2616 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4455_
timestamp 1596991774
transform -1 0 2808 0 -1 5010
box -4 -6 196 206
use AOI21X1  _4044_
timestamp 1596991774
transform -1 0 2872 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4232_
timestamp 1596991774
transform 1 0 2872 0 -1 5010
box -4 -6 68 206
use AOI21X1  _4233_
timestamp 1596991774
transform -1 0 3064 0 -1 5010
box -4 -6 68 206
use FILL  SFILL29360x48100
timestamp 1596991774
transform -1 0 2952 0 -1 5010
box -4 -6 20 206
use FILL  SFILL29520x48100
timestamp 1596991774
transform -1 0 2968 0 -1 5010
box -4 -6 20 206
use FILL  SFILL29680x48100
timestamp 1596991774
transform -1 0 2984 0 -1 5010
box -4 -6 20 206
use FILL  SFILL29840x48100
timestamp 1596991774
transform -1 0 3000 0 -1 5010
box -4 -6 20 206
use OAI21X1  _4221_
timestamp 1596991774
transform -1 0 3128 0 -1 5010
box -4 -6 68 206
use AOI21X1  _4222_
timestamp 1596991774
transform -1 0 3192 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4330_
timestamp 1596991774
transform 1 0 3192 0 -1 5010
box -4 -6 196 206
use OAI21X1  _3772_
timestamp 1596991774
transform -1 0 3448 0 -1 5010
box -4 -6 68 206
use NAND2X1  _3771_
timestamp 1596991774
transform -1 0 3496 0 -1 5010
box -4 -6 52 206
use OAI22X1  _4248_
timestamp 1596991774
transform -1 0 3576 0 -1 5010
box -4 -6 84 206
use OAI21X1  _4247_
timestamp 1596991774
transform -1 0 3640 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4069_
timestamp 1596991774
transform 1 0 3640 0 -1 5010
box -4 -6 68 206
use NOR2X1  _4246_
timestamp 1596991774
transform -1 0 3752 0 -1 5010
box -4 -6 52 206
use MUX2X1  _4231_
timestamp 1596991774
transform -1 0 3848 0 -1 5010
box -4 -6 100 206
use OAI22X1  _4226_
timestamp 1596991774
transform -1 0 3928 0 -1 5010
box -4 -6 84 206
use NOR2X1  _4224_
timestamp 1596991774
transform 1 0 3928 0 -1 5010
box -4 -6 52 206
use OAI21X1  _4225_
timestamp 1596991774
transform -1 0 4040 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4229_
timestamp 1596991774
transform 1 0 4040 0 -1 5010
box -4 -6 68 206
use NOR2X1  _4228_
timestamp 1596991774
transform 1 0 4104 0 -1 5010
box -4 -6 52 206
use OAI22X1  _4230_
timestamp 1596991774
transform -1 0 4232 0 -1 5010
box -4 -6 84 206
use DFFPOSX1  _4328_
timestamp 1596991774
transform -1 0 4424 0 -1 5010
box -4 -6 196 206
use OAI21X1  _3768_
timestamp 1596991774
transform 1 0 4488 0 -1 5010
box -4 -6 68 206
use NAND2X1  _3767_
timestamp 1596991774
transform 1 0 4552 0 -1 5010
box -4 -6 52 206
use MUX2X1  _4242_
timestamp 1596991774
transform -1 0 4696 0 -1 5010
box -4 -6 100 206
use FILL  SFILL44240x48100
timestamp 1596991774
transform -1 0 4440 0 -1 5010
box -4 -6 20 206
use FILL  SFILL44400x48100
timestamp 1596991774
transform -1 0 4456 0 -1 5010
box -4 -6 20 206
use FILL  SFILL44560x48100
timestamp 1596991774
transform -1 0 4472 0 -1 5010
box -4 -6 20 206
use FILL  SFILL44720x48100
timestamp 1596991774
transform -1 0 4488 0 -1 5010
box -4 -6 20 206
use NOR2X1  _4235_
timestamp 1596991774
transform 1 0 4696 0 -1 5010
box -4 -6 52 206
use OAI22X1  _4237_
timestamp 1596991774
transform 1 0 4744 0 -1 5010
box -4 -6 84 206
use OAI21X1  _4236_
timestamp 1596991774
transform -1 0 4888 0 -1 5010
box -4 -6 68 206
use NOR2X1  _4057_
timestamp 1596991774
transform -1 0 4936 0 -1 5010
box -4 -6 52 206
use MUX2X1  _4064_
timestamp 1596991774
transform -1 0 5032 0 -1 5010
box -4 -6 100 206
use OAI22X1  _4059_
timestamp 1596991774
transform 1 0 5032 0 -1 5010
box -4 -6 84 206
use OAI21X1  _4058_
timestamp 1596991774
transform -1 0 5176 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4408_
timestamp 1596991774
transform -1 0 5368 0 -1 5010
box -4 -6 196 206
use NOR2X1  _3692_
timestamp 1596991774
transform 1 0 5368 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3693_
timestamp 1596991774
transform -1 0 5480 0 -1 5010
box -4 -6 68 206
use AOI21X1  _3904_
timestamp 1596991774
transform 1 0 5480 0 -1 5010
box -4 -6 68 206
use NOR2X1  _3903_
timestamp 1596991774
transform -1 0 5592 0 -1 5010
box -4 -6 52 206
use OAI21X1  _4062_
timestamp 1596991774
transform 1 0 5592 0 -1 5010
box -4 -6 68 206
use OAI22X1  _4063_
timestamp 1596991774
transform 1 0 5656 0 -1 5010
box -4 -6 84 206
use NOR2X1  _4061_
timestamp 1596991774
transform -1 0 5784 0 -1 5010
box -4 -6 52 206
use NAND2X1  _3870_
timestamp 1596991774
transform 1 0 5784 0 -1 5010
box -4 -6 52 206
use MUX2X1  _4042_
timestamp 1596991774
transform -1 0 5928 0 -1 5010
box -4 -6 100 206
use NOR2X1  _4035_
timestamp 1596991774
transform -1 0 6040 0 -1 5010
box -4 -6 52 206
use FILL  SFILL59280x48100
timestamp 1596991774
transform -1 0 5944 0 -1 5010
box -4 -6 20 206
use FILL  SFILL59440x48100
timestamp 1596991774
transform -1 0 5960 0 -1 5010
box -4 -6 20 206
use FILL  SFILL59600x48100
timestamp 1596991774
transform -1 0 5976 0 -1 5010
box -4 -6 20 206
use FILL  SFILL59760x48100
timestamp 1596991774
transform -1 0 5992 0 -1 5010
box -4 -6 20 206
use OAI22X1  _4037_
timestamp 1596991774
transform 1 0 6040 0 -1 5010
box -4 -6 84 206
use MUX2X1  _4220_
timestamp 1596991774
transform 1 0 6120 0 -1 5010
box -4 -6 100 206
use OAI21X1  _4214_
timestamp 1596991774
transform -1 0 6280 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4036_
timestamp 1596991774
transform -1 0 6344 0 -1 5010
box -4 -6 68 206
use NOR2X1  _4039_
timestamp 1596991774
transform -1 0 6392 0 -1 5010
box -4 -6 52 206
use NOR2X1  _4217_
timestamp 1596991774
transform 1 0 6392 0 -1 5010
box -4 -6 52 206
use OAI22X1  _4041_
timestamp 1596991774
transform 1 0 6440 0 -1 5010
box -4 -6 84 206
use OAI21X1  _4040_
timestamp 1596991774
transform -1 0 6584 0 -1 5010
box -4 -6 68 206
use OAI22X1  _4219_
timestamp 1596991774
transform 1 0 6584 0 -1 5010
box -4 -6 84 206
use OAI21X1  _4218_
timestamp 1596991774
transform -1 0 6728 0 -1 5010
box -4 -6 68 206
use MUX2X1  _4038_
timestamp 1596991774
transform 1 0 6728 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4216_
timestamp 1596991774
transform 1 0 6824 0 -1 5010
box -4 -6 100 206
use NOR2X1  _4290_
timestamp 1596991774
transform -1 0 6968 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4423_
timestamp 1596991774
transform -1 0 7160 0 -1 5010
box -4 -6 196 206
use NOR2X1  _3877_
timestamp 1596991774
transform 1 0 7160 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3900_
timestamp 1596991774
transform 1 0 7208 0 -1 5010
box -4 -6 68 206
use NOR2X1  _3889_
timestamp 1596991774
transform -1 0 7320 0 -1 5010
box -4 -6 52 206
use NOR2X1  _3899_
timestamp 1596991774
transform -1 0 7368 0 -1 5010
box -4 -6 52 206
use FILL  FILL71120x48100
timestamp 1596991774
transform -1 0 7384 0 -1 5010
box -4 -6 20 206
use FILL  FILL71280x48100
timestamp 1596991774
transform -1 0 7400 0 -1 5010
box -4 -6 20 206
use INVX1  _2783_
timestamp 1596991774
transform -1 0 40 0 1 5010
box -4 -6 36 206
use OAI21X1  _2786_
timestamp 1596991774
transform 1 0 40 0 1 5010
box -4 -6 68 206
use NOR2X1  _2789_
timestamp 1596991774
transform -1 0 152 0 1 5010
box -4 -6 52 206
use OAI21X1  _2832_
timestamp 1596991774
transform -1 0 216 0 1 5010
box -4 -6 68 206
use NAND2X1  _2790_
timestamp 1596991774
transform -1 0 264 0 1 5010
box -4 -6 52 206
use OAI21X1  _2833_
timestamp 1596991774
transform 1 0 264 0 1 5010
box -4 -6 68 206
use NOR2X1  _2782_
timestamp 1596991774
transform -1 0 376 0 1 5010
box -4 -6 52 206
use OAI21X1  _2831_
timestamp 1596991774
transform -1 0 440 0 1 5010
box -4 -6 68 206
use OAI21X1  _2781_
timestamp 1596991774
transform 1 0 440 0 1 5010
box -4 -6 68 206
use INVX1  _2779_
timestamp 1596991774
transform 1 0 504 0 1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert196
timestamp 1596991774
transform 1 0 536 0 1 5010
box -4 -6 52 206
use INVX1  _2674_
timestamp 1596991774
transform -1 0 616 0 1 5010
box -4 -6 36 206
use OAI21X1  _2738_
timestamp 1596991774
transform 1 0 616 0 1 5010
box -4 -6 68 206
use OAI21X1  _2736_
timestamp 1596991774
transform -1 0 744 0 1 5010
box -4 -6 68 206
use NOR2X1  _2680_
timestamp 1596991774
transform 1 0 744 0 1 5010
box -4 -6 52 206
use OAI22X1  _2679_
timestamp 1596991774
transform 1 0 792 0 1 5010
box -4 -6 84 206
use AOI21X1  _2745_
timestamp 1596991774
transform 1 0 872 0 1 5010
box -4 -6 68 206
use NAND2X1  _2689_
timestamp 1596991774
transform 1 0 936 0 1 5010
box -4 -6 52 206
use INVX1  _2742_
timestamp 1596991774
transform 1 0 984 0 1 5010
box -4 -6 36 206
use OAI21X1  _2744_
timestamp 1596991774
transform 1 0 1016 0 1 5010
box -4 -6 68 206
use NOR2X1  _2752_
timestamp 1596991774
transform 1 0 1080 0 1 5010
box -4 -6 52 206
use NAND3X1  _2750_
timestamp 1596991774
transform 1 0 1128 0 1 5010
box -4 -6 68 206
use AOI22X1  _2741_
timestamp 1596991774
transform 1 0 1192 0 1 5010
box -4 -6 84 206
use NAND2X1  _2740_
timestamp 1596991774
transform -1 0 1320 0 1 5010
box -4 -6 52 206
use OAI21X1  _2743_
timestamp 1596991774
transform 1 0 1320 0 1 5010
box -4 -6 68 206
use NAND3X1  _2672_
timestamp 1596991774
transform 1 0 1384 0 1 5010
box -4 -6 68 206
use INVX1  _2669_
timestamp 1596991774
transform 1 0 1512 0 1 5010
box -4 -6 36 206
use NAND2X1  _2670_
timestamp 1596991774
transform -1 0 1592 0 1 5010
box -4 -6 52 206
use INVX1  _2766_
timestamp 1596991774
transform 1 0 1592 0 1 5010
box -4 -6 36 206
use FILL  SFILL14480x50100
timestamp 1596991774
transform 1 0 1448 0 1 5010
box -4 -6 20 206
use FILL  SFILL14640x50100
timestamp 1596991774
transform 1 0 1464 0 1 5010
box -4 -6 20 206
use FILL  SFILL14800x50100
timestamp 1596991774
transform 1 0 1480 0 1 5010
box -4 -6 20 206
use FILL  SFILL14960x50100
timestamp 1596991774
transform 1 0 1496 0 1 5010
box -4 -6 20 206
use NAND2X1  _2835_
timestamp 1596991774
transform -1 0 1672 0 1 5010
box -4 -6 52 206
use INVX2  _2662_
timestamp 1596991774
transform -1 0 1704 0 1 5010
box -4 -6 36 206
use AOI22X1  _2771_
timestamp 1596991774
transform -1 0 1784 0 1 5010
box -4 -6 84 206
use INVX1  _2770_
timestamp 1596991774
transform -1 0 1816 0 1 5010
box -4 -6 36 206
use AOI21X1  _2837_
timestamp 1596991774
transform 1 0 1816 0 1 5010
box -4 -6 68 206
use AOI21X1  _2836_
timestamp 1596991774
transform -1 0 1944 0 1 5010
box -4 -6 68 206
use OAI22X1  _2764_
timestamp 1596991774
transform 1 0 1944 0 1 5010
box -4 -6 84 206
use NOR2X1  _2768_
timestamp 1596991774
transform 1 0 2024 0 1 5010
box -4 -6 52 206
use INVX1  _2763_
timestamp 1596991774
transform -1 0 2104 0 1 5010
box -4 -6 36 206
use DFFPOSX1  _4456_
timestamp 1596991774
transform -1 0 2296 0 1 5010
box -4 -6 196 206
use OAI21X1  _4054_
timestamp 1596991774
transform 1 0 2296 0 1 5010
box -4 -6 68 206
use AOI21X1  _4055_
timestamp 1596991774
transform -1 0 2424 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4439_
timestamp 1596991774
transform -1 0 2616 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4440_
timestamp 1596991774
transform -1 0 2808 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4362_
timestamp 1596991774
transform 1 0 2808 0 1 5010
box -4 -6 196 206
use FILL  SFILL30000x50100
timestamp 1596991774
transform 1 0 3000 0 1 5010
box -4 -6 20 206
use NAND2X1  _3805_
timestamp 1596991774
transform 1 0 3064 0 1 5010
box -4 -6 52 206
use OAI21X1  _3806_
timestamp 1596991774
transform -1 0 3176 0 1 5010
box -4 -6 68 206
use MUX2X1  _4067_
timestamp 1596991774
transform 1 0 3176 0 1 5010
box -4 -6 100 206
use FILL  SFILL30160x50100
timestamp 1596991774
transform 1 0 3016 0 1 5010
box -4 -6 20 206
use FILL  SFILL30320x50100
timestamp 1596991774
transform 1 0 3032 0 1 5010
box -4 -6 20 206
use FILL  SFILL30480x50100
timestamp 1596991774
transform 1 0 3048 0 1 5010
box -4 -6 20 206
use MUX2X1  _4245_
timestamp 1596991774
transform -1 0 3368 0 1 5010
box -4 -6 100 206
use MUX2X1  _4075_
timestamp 1596991774
transform -1 0 3464 0 1 5010
box -4 -6 100 206
use OAI22X1  _4070_
timestamp 1596991774
transform -1 0 3544 0 1 5010
box -4 -6 84 206
use NOR2X1  _4068_
timestamp 1596991774
transform 1 0 3544 0 1 5010
box -4 -6 52 206
use NOR2X1  _4046_
timestamp 1596991774
transform -1 0 3640 0 1 5010
box -4 -6 52 206
use OAI22X1  _4048_
timestamp 1596991774
transform -1 0 3720 0 1 5010
box -4 -6 84 206
use MUX2X1  _4053_
timestamp 1596991774
transform 1 0 3720 0 1 5010
box -4 -6 100 206
use OAI21X1  _4047_
timestamp 1596991774
transform -1 0 3880 0 1 5010
box -4 -6 68 206
use OAI21X1  _4051_
timestamp 1596991774
transform 1 0 3880 0 1 5010
box -4 -6 68 206
use OAI22X1  _4052_
timestamp 1596991774
transform 1 0 3944 0 1 5010
box -4 -6 84 206
use NOR2X1  _4050_
timestamp 1596991774
transform -1 0 4072 0 1 5010
box -4 -6 52 206
use OAI21X1  _3739_
timestamp 1596991774
transform 1 0 4072 0 1 5010
box -4 -6 68 206
use OAI21X1  _3738_
timestamp 1596991774
transform -1 0 4200 0 1 5010
box -4 -6 68 206
use OAI21X1  _3734_
timestamp 1596991774
transform -1 0 4264 0 1 5010
box -4 -6 68 206
use OAI21X1  _3735_
timestamp 1596991774
transform -1 0 4328 0 1 5010
box -4 -6 68 206
use MUX2X1  _4049_
timestamp 1596991774
transform 1 0 4328 0 1 5010
box -4 -6 100 206
use MUX2X1  _4227_
timestamp 1596991774
transform -1 0 4584 0 1 5010
box -4 -6 100 206
use OAI21X1  _3736_
timestamp 1596991774
transform 1 0 4584 0 1 5010
box -4 -6 68 206
use FILL  SFILL44240x50100
timestamp 1596991774
transform 1 0 4424 0 1 5010
box -4 -6 20 206
use FILL  SFILL44400x50100
timestamp 1596991774
transform 1 0 4440 0 1 5010
box -4 -6 20 206
use FILL  SFILL44560x50100
timestamp 1596991774
transform 1 0 4456 0 1 5010
box -4 -6 20 206
use FILL  SFILL44720x50100
timestamp 1596991774
transform 1 0 4472 0 1 5010
box -4 -6 20 206
use OAI21X1  _3737_
timestamp 1596991774
transform -1 0 4712 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4377_
timestamp 1596991774
transform 1 0 4712 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4424_
timestamp 1596991774
transform -1 0 5096 0 1 5010
box -4 -6 196 206
use NOR2X1  _4292_
timestamp 1596991774
transform 1 0 5096 0 1 5010
box -4 -6 52 206
use AOI21X1  _4293_
timestamp 1596991774
transform -1 0 5208 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4345_
timestamp 1596991774
transform 1 0 5208 0 1 5010
box -4 -6 196 206
use OAI21X1  _4240_
timestamp 1596991774
transform 1 0 5400 0 1 5010
box -4 -6 68 206
use OAI22X1  _4241_
timestamp 1596991774
transform 1 0 5464 0 1 5010
box -4 -6 84 206
use NOR2X1  _4239_
timestamp 1596991774
transform -1 0 5592 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4313_
timestamp 1596991774
transform -1 0 5784 0 1 5010
box -4 -6 196 206
use OAI21X1  _3871_
timestamp 1596991774
transform 1 0 5784 0 1 5010
box -4 -6 68 206
use OAI21X1  _3733_
timestamp 1596991774
transform 1 0 5848 0 1 5010
box -4 -6 68 206
use OAI21X1  _3732_
timestamp 1596991774
transform 1 0 5976 0 1 5010
box -4 -6 68 206
use FILL  SFILL59120x50100
timestamp 1596991774
transform 1 0 5912 0 1 5010
box -4 -6 20 206
use FILL  SFILL59280x50100
timestamp 1596991774
transform 1 0 5928 0 1 5010
box -4 -6 20 206
use FILL  SFILL59440x50100
timestamp 1596991774
transform 1 0 5944 0 1 5010
box -4 -6 20 206
use FILL  SFILL59600x50100
timestamp 1596991774
transform 1 0 5960 0 1 5010
box -4 -6 20 206
use NOR2X1  _4213_
timestamp 1596991774
transform 1 0 6040 0 1 5010
box -4 -6 52 206
use OAI22X1  _4215_
timestamp 1596991774
transform 1 0 6088 0 1 5010
box -4 -6 84 206
use MUX2X1  _4212_
timestamp 1596991774
transform -1 0 6264 0 1 5010
box -4 -6 100 206
use MUX2X1  _4034_
timestamp 1596991774
transform -1 0 6360 0 1 5010
box -4 -6 100 206
use MUX2X1  _4060_
timestamp 1596991774
transform 1 0 6360 0 1 5010
box -4 -6 100 206
use MUX2X1  _4238_
timestamp 1596991774
transform -1 0 6552 0 1 5010
box -4 -6 100 206
use NOR2X1  _3689_
timestamp 1596991774
transform -1 0 6600 0 1 5010
box -4 -6 52 206
use AOI21X1  _3690_
timestamp 1596991774
transform -1 0 6664 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4407_
timestamp 1596991774
transform 1 0 6664 0 1 5010
box -4 -6 196 206
use NOR2X1  _3832_
timestamp 1596991774
transform -1 0 6904 0 1 5010
box -4 -6 52 206
use AOI21X1  _4291_
timestamp 1596991774
transform 1 0 6904 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4391_
timestamp 1596991774
transform -1 0 7160 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4386_
timestamp 1596991774
transform -1 0 7352 0 1 5010
box -4 -6 196 206
use FILL  FILL70960x50100
timestamp 1596991774
transform 1 0 7352 0 1 5010
box -4 -6 20 206
use FILL  FILL71120x50100
timestamp 1596991774
transform 1 0 7368 0 1 5010
box -4 -6 20 206
use FILL  FILL71280x50100
timestamp 1596991774
transform 1 0 7384 0 1 5010
box -4 -6 20 206
use BUFX2  _2113_
timestamp 1596991774
transform -1 0 56 0 -1 5410
box -4 -6 52 206
use BUFX2  _2101_
timestamp 1596991774
transform -1 0 104 0 -1 5410
box -4 -6 52 206
use NAND3X1  _2735_
timestamp 1596991774
transform -1 0 168 0 -1 5410
box -4 -6 68 206
use NAND2X1  _2734_
timestamp 1596991774
transform -1 0 216 0 -1 5410
box -4 -6 52 206
use NAND2X1  _2733_
timestamp 1596991774
transform -1 0 264 0 -1 5410
box -4 -6 52 206
use OAI22X1  _2676_
timestamp 1596991774
transform -1 0 344 0 -1 5410
box -4 -6 84 206
use INVX1  _2675_
timestamp 1596991774
transform -1 0 376 0 -1 5410
box -4 -6 36 206
use BUFX2  _2100_
timestamp 1596991774
transform 1 0 376 0 -1 5410
box -4 -6 52 206
use NOR3X1  _2673_
timestamp 1596991774
transform -1 0 552 0 -1 5410
box -4 -6 132 206
use BUFX2  _2103_
timestamp 1596991774
transform -1 0 600 0 -1 5410
box -4 -6 52 206
use NAND3X1  _2664_
timestamp 1596991774
transform 1 0 600 0 -1 5410
box -4 -6 68 206
use NAND2X1  _2659_
timestamp 1596991774
transform -1 0 712 0 -1 5410
box -4 -6 52 206
use NAND2X1  _2663_
timestamp 1596991774
transform -1 0 760 0 -1 5410
box -4 -6 52 206
use INVX1  _2660_
timestamp 1596991774
transform 1 0 760 0 -1 5410
box -4 -6 36 206
use NAND2X1  _2661_
timestamp 1596991774
transform -1 0 840 0 -1 5410
box -4 -6 52 206
use INVX1  _2658_
timestamp 1596991774
transform 1 0 840 0 -1 5410
box -4 -6 36 206
use NAND2X1  _2739_
timestamp 1596991774
transform 1 0 872 0 -1 5410
box -4 -6 52 206
use BUFX2  _2105_
timestamp 1596991774
transform -1 0 968 0 -1 5410
box -4 -6 52 206
use BUFX2  _2104_
timestamp 1596991774
transform -1 0 1016 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert186
timestamp 1596991774
transform -1 0 1064 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert188
timestamp 1596991774
transform 1 0 1064 0 -1 5410
box -4 -6 52 206
use INVX1  _2765_
timestamp 1596991774
transform 1 0 1112 0 -1 5410
box -4 -6 36 206
use OAI22X1  _2767_
timestamp 1596991774
transform 1 0 1144 0 -1 5410
box -4 -6 84 206
use BUFX2  _2102_
timestamp 1596991774
transform -1 0 1272 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4458_
timestamp 1596991774
transform -1 0 1464 0 -1 5410
box -4 -6 196 206
use AOI21X1  _4077_
timestamp 1596991774
transform -1 0 1592 0 -1 5410
box -4 -6 68 206
use OAI21X1  _4076_
timestamp 1596991774
transform 1 0 1592 0 -1 5410
box -4 -6 68 206
use FILL  SFILL14640x52100
timestamp 1596991774
transform -1 0 1480 0 -1 5410
box -4 -6 20 206
use FILL  SFILL14800x52100
timestamp 1596991774
transform -1 0 1496 0 -1 5410
box -4 -6 20 206
use FILL  SFILL14960x52100
timestamp 1596991774
transform -1 0 1512 0 -1 5410
box -4 -6 20 206
use FILL  SFILL15120x52100
timestamp 1596991774
transform -1 0 1528 0 -1 5410
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert13
timestamp 1596991774
transform -1 0 1800 0 -1 5410
box -4 -6 148 206
use CLKBUF1  CLKBUF1_insert10
timestamp 1596991774
transform 1 0 1800 0 -1 5410
box -4 -6 148 206
use DFFPOSX1  _4394_
timestamp 1596991774
transform 1 0 1944 0 -1 5410
box -4 -6 196 206
use NOR2X1  _3838_
timestamp 1596991774
transform 1 0 2136 0 -1 5410
box -4 -6 52 206
use AOI21X1  _3839_
timestamp 1596991774
transform -1 0 2248 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4392_
timestamp 1596991774
transform 1 0 2248 0 -1 5410
box -4 -6 196 206
use NOR2X1  _3834_
timestamp 1596991774
transform 1 0 2440 0 -1 5410
box -4 -6 52 206
use AOI21X1  _3835_
timestamp 1596991774
transform -1 0 2552 0 -1 5410
box -4 -6 68 206
use MUX2X1  _4223_
timestamp 1596991774
transform 1 0 2552 0 -1 5410
box -4 -6 100 206
use MUX2X1  _4045_
timestamp 1596991774
transform -1 0 2744 0 -1 5410
box -4 -6 100 206
use NAND2X1  _3801_
timestamp 1596991774
transform 1 0 2744 0 -1 5410
box -4 -6 52 206
use OAI21X1  _3802_
timestamp 1596991774
transform -1 0 2856 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4360_
timestamp 1596991774
transform -1 0 3112 0 -1 5410
box -4 -6 196 206
use FILL  SFILL28560x52100
timestamp 1596991774
transform -1 0 2872 0 -1 5410
box -4 -6 20 206
use FILL  SFILL28720x52100
timestamp 1596991774
transform -1 0 2888 0 -1 5410
box -4 -6 20 206
use FILL  SFILL28880x52100
timestamp 1596991774
transform -1 0 2904 0 -1 5410
box -4 -6 20 206
use FILL  SFILL29040x52100
timestamp 1596991774
transform -1 0 2920 0 -1 5410
box -4 -6 20 206
use DFFPOSX1  _4376_
timestamp 1596991774
transform 1 0 3112 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4378_
timestamp 1596991774
transform 1 0 3304 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4344_
timestamp 1596991774
transform 1 0 3496 0 -1 5410
box -4 -6 196 206
use AOI21X1  _3902_
timestamp 1596991774
transform 1 0 3688 0 -1 5410
box -4 -6 68 206
use NOR2X1  _3901_
timestamp 1596991774
transform 1 0 3752 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4361_
timestamp 1596991774
transform -1 0 3992 0 -1 5410
box -4 -6 196 206
use NAND2X1  _3803_
timestamp 1596991774
transform 1 0 3992 0 -1 5410
box -4 -6 52 206
use OAI21X1  _3804_
timestamp 1596991774
transform -1 0 4104 0 -1 5410
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert21
timestamp 1596991774
transform -1 0 4248 0 -1 5410
box -4 -6 148 206
use NAND2X1  _3799_
timestamp 1596991774
transform -1 0 4296 0 -1 5410
box -4 -6 52 206
use OAI21X1  _3800_
timestamp 1596991774
transform -1 0 4360 0 -1 5410
box -4 -6 68 206
use FILL  SFILL43600x52100
timestamp 1596991774
transform -1 0 4376 0 -1 5410
box -4 -6 20 206
use FILL  SFILL43760x52100
timestamp 1596991774
transform -1 0 4392 0 -1 5410
box -4 -6 20 206
use FILL  SFILL43920x52100
timestamp 1596991774
transform -1 0 4408 0 -1 5410
box -4 -6 20 206
use FILL  SFILL44080x52100
timestamp 1596991774
transform -1 0 4424 0 -1 5410
box -4 -6 20 206
use DFFPOSX1  _4359_
timestamp 1596991774
transform 1 0 4424 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4375_
timestamp 1596991774
transform 1 0 4616 0 -1 5410
box -4 -6 196 206
use OAI21X1  _3867_
timestamp 1596991774
transform 1 0 4808 0 -1 5410
box -4 -6 68 206
use NAND2X1  _3866_
timestamp 1596991774
transform -1 0 4920 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4311_
timestamp 1596991774
transform 1 0 4920 0 -1 5410
box -4 -6 196 206
use AOI21X1  _3696_
timestamp 1596991774
transform 1 0 5112 0 -1 5410
box -4 -6 68 206
use NOR2X1  _3695_
timestamp 1596991774
transform -1 0 5224 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4409_
timestamp 1596991774
transform 1 0 5224 0 -1 5410
box -4 -6 196 206
use NOR2X1  _4294_
timestamp 1596991774
transform -1 0 5464 0 -1 5410
box -4 -6 52 206
use AOI21X1  _4295_
timestamp 1596991774
transform -1 0 5528 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4425_
timestamp 1596991774
transform 1 0 5528 0 -1 5410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert19
timestamp 1596991774
transform -1 0 5864 0 -1 5410
box -4 -6 148 206
use AOI21X1  _3660_
timestamp 1596991774
transform -1 0 5928 0 -1 5410
box -4 -6 68 206
use INVX1  _3511_
timestamp 1596991774
transform -1 0 6024 0 -1 5410
box -4 -6 36 206
use FILL  SFILL59280x52100
timestamp 1596991774
transform -1 0 5944 0 -1 5410
box -4 -6 20 206
use FILL  SFILL59440x52100
timestamp 1596991774
transform -1 0 5960 0 -1 5410
box -4 -6 20 206
use FILL  SFILL59600x52100
timestamp 1596991774
transform -1 0 5976 0 -1 5410
box -4 -6 20 206
use FILL  SFILL59760x52100
timestamp 1596991774
transform -1 0 5992 0 -1 5410
box -4 -6 20 206
use NAND2X1  _3856_
timestamp 1596991774
transform -1 0 6072 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4580_
timestamp 1596991774
transform 1 0 6072 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4418_
timestamp 1596991774
transform -1 0 6456 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4417_
timestamp 1596991774
transform -1 0 6648 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4365_
timestamp 1596991774
transform -1 0 6840 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4338_
timestamp 1596991774
transform -1 0 7032 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4343_
timestamp 1596991774
transform -1 0 7224 0 -1 5410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert8
timestamp 1596991774
transform -1 0 7368 0 -1 5410
box -4 -6 148 206
use FILL  FILL71120x52100
timestamp 1596991774
transform -1 0 7384 0 -1 5410
box -4 -6 20 206
use FILL  FILL71280x52100
timestamp 1596991774
transform -1 0 7400 0 -1 5410
box -4 -6 20 206
<< labels >>
flabel metal4 s 2912 -10 2976 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 1408 -10 1472 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 6413 -23 6419 -17 7 FreeSans 24 270 0 0 adrs_bus[15]
port 2 nsew
flabel metal3 s 7437 4537 7443 4543 3 FreeSans 24 0 0 0 adrs_bus[14]
port 3 nsew
flabel metal2 s 6077 -23 6083 -17 7 FreeSans 24 270 0 0 adrs_bus[13]
port 4 nsew
flabel metal2 s 6125 -23 6131 -17 7 FreeSans 24 270 0 0 adrs_bus[12]
port 5 nsew
flabel metal3 s 7437 4497 7443 4503 3 FreeSans 24 0 0 0 adrs_bus[11]
port 6 nsew
flabel metal3 s 7437 2897 7443 2903 3 FreeSans 24 0 0 0 adrs_bus[10]
port 7 nsew
flabel metal2 s 5389 -23 5395 -17 7 FreeSans 24 270 0 0 adrs_bus[9]
port 8 nsew
flabel metal2 s 5725 -23 5731 -17 7 FreeSans 24 270 0 0 adrs_bus[8]
port 9 nsew
flabel metal2 s 4861 -23 4867 -17 7 FreeSans 24 270 0 0 adrs_bus[7]
port 10 nsew
flabel metal2 s 5341 -23 5347 -17 7 FreeSans 24 270 0 0 adrs_bus[6]
port 11 nsew
flabel metal2 s 5613 -23 5619 -17 7 FreeSans 24 270 0 0 adrs_bus[5]
port 12 nsew
flabel metal2 s 5773 -23 5779 -17 7 FreeSans 24 270 0 0 adrs_bus[4]
port 13 nsew
flabel metal2 s 5085 -23 5091 -17 7 FreeSans 24 270 0 0 adrs_bus[3]
port 14 nsew
flabel metal2 s 5037 -23 5043 -17 7 FreeSans 24 270 0 0 adrs_bus[2]
port 15 nsew
flabel metal2 s 5229 -23 5235 -17 7 FreeSans 24 270 0 0 adrs_bus[1]
port 16 nsew
flabel metal2 s 5565 -23 5571 -17 7 FreeSans 24 270 0 0 adrs_bus[0]
port 17 nsew
flabel metal3 s 7437 3737 7443 3743 3 FreeSans 24 0 0 0 clock
port 18 nsew
flabel metal2 s 4253 -23 4259 -17 7 FreeSans 24 270 0 0 data_in[15]
port 19 nsew
flabel metal2 s 4093 -23 4099 -17 7 FreeSans 24 270 0 0 data_in[14]
port 20 nsew
flabel metal2 s 4061 -23 4067 -17 7 FreeSans 24 270 0 0 data_in[13]
port 21 nsew
flabel metal2 s 3837 -23 3843 -17 7 FreeSans 24 270 0 0 data_in[12]
port 22 nsew
flabel metal3 s 7437 2957 7443 2963 3 FreeSans 24 0 0 0 data_in[11]
port 23 nsew
flabel metal3 s 7437 1897 7443 1903 3 FreeSans 24 0 0 0 data_in[10]
port 24 nsew
flabel metal3 s 7437 2497 7443 2503 3 FreeSans 24 0 0 0 data_in[9]
port 25 nsew
flabel metal2 s 4749 -23 4755 -17 7 FreeSans 24 270 0 0 data_in[8]
port 26 nsew
flabel metal2 s 4989 -23 4995 -17 7 FreeSans 24 270 0 0 data_in[7]
port 27 nsew
flabel metal2 s 4669 -23 4675 -17 7 FreeSans 24 270 0 0 data_in[6]
port 28 nsew
flabel metal2 s 4541 -23 4547 -17 7 FreeSans 24 270 0 0 data_in[5]
port 29 nsew
flabel metal2 s 4637 -23 4643 -17 7 FreeSans 24 270 0 0 data_in[4]
port 30 nsew
flabel metal2 s 4717 -23 4723 -17 7 FreeSans 24 270 0 0 data_in[3]
port 31 nsew
flabel metal3 s 7437 1697 7443 1703 3 FreeSans 24 0 0 0 data_in[2]
port 32 nsew
flabel metal2 s 4589 -23 4595 -17 7 FreeSans 24 270 0 0 data_in[1]
port 33 nsew
flabel metal2 s 4797 -23 4803 -17 7 FreeSans 24 270 0 0 data_in[0]
port 34 nsew
flabel metal2 s 941 5457 947 5463 3 FreeSans 24 90 0 0 data_out[15]
port 35 nsew
flabel metal2 s 989 5457 995 5463 3 FreeSans 24 90 0 0 data_out[14]
port 36 nsew
flabel metal2 s 573 5457 579 5463 3 FreeSans 24 90 0 0 data_out[13]
port 37 nsew
flabel metal2 s 1245 5457 1251 5463 3 FreeSans 24 90 0 0 data_out[12]
port 38 nsew
flabel metal3 s -35 5297 -29 5303 7 FreeSans 24 0 0 0 data_out[11]
port 39 nsew
flabel metal2 s 397 5457 403 5463 3 FreeSans 24 90 0 0 data_out[10]
port 40 nsew
flabel metal3 s -35 5337 -29 5343 7 FreeSans 24 0 0 0 data_out[9]
port 41 nsew
flabel metal3 s -35 4897 -29 4903 7 FreeSans 24 0 0 0 data_out[8]
port 42 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 data_out[7]
port 43 nsew
flabel metal3 s -35 97 -29 103 7 FreeSans 24 0 0 0 data_out[6]
port 44 nsew
flabel metal2 s 461 -23 467 -17 7 FreeSans 24 270 0 0 data_out[5]
port 45 nsew
flabel metal3 s -35 1297 -29 1303 7 FreeSans 24 0 0 0 data_out[4]
port 46 nsew
flabel metal2 s 3405 -23 3411 -17 7 FreeSans 24 270 0 0 data_out[3]
port 47 nsew
flabel metal2 s 3453 -23 3459 -17 7 FreeSans 24 270 0 0 data_out[2]
port 48 nsew
flabel metal2 s 3501 -23 3507 -17 7 FreeSans 24 270 0 0 data_out[1]
port 49 nsew
flabel metal2 s 2861 -23 2867 -17 7 FreeSans 24 270 0 0 data_out[0]
port 50 nsew
flabel metal2 s 3805 -23 3811 -17 7 FreeSans 24 270 0 0 mem_rd
port 51 nsew
flabel metal2 s 3741 -23 3747 -17 7 FreeSans 24 270 0 0 mem_wr
port 52 nsew
flabel metal2 s 3037 5457 3043 5463 3 FreeSans 24 90 0 0 reset
port 53 nsew
<< end >>
