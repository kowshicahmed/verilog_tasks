magic
tech scmos
magscale 1 2
timestamp 1589549099
<< metal1 >>
rect 762 2014 774 2016
rect 747 2006 749 2014
rect 757 2006 759 2014
rect 767 2006 769 2014
rect 777 2006 779 2014
rect 787 2006 789 2014
rect 762 2004 774 2006
rect 733 1977 796 1983
rect 2410 1936 2412 1944
rect 29 1917 44 1923
rect 829 1917 844 1923
rect 1140 1917 1155 1923
rect 1213 1917 1235 1923
rect 1597 1917 1612 1923
rect 1805 1917 1827 1923
rect 77 1903 83 1916
rect 77 1897 99 1903
rect 269 1897 300 1903
rect 493 1897 508 1903
rect 605 1897 627 1903
rect 605 1884 611 1897
rect 1284 1897 1315 1903
rect 1469 1897 1491 1903
rect 1533 1897 1555 1903
rect 1821 1897 1852 1903
rect 2237 1903 2243 1923
rect 2756 1916 2764 1924
rect 2836 1917 2851 1923
rect 2173 1897 2211 1903
rect 2237 1897 2332 1903
rect 61 1877 92 1883
rect 109 1877 147 1883
rect 141 1857 147 1877
rect 372 1877 387 1883
rect 877 1877 892 1883
rect 932 1877 947 1883
rect 1268 1877 1283 1883
rect 301 1857 348 1863
rect 1277 1857 1283 1877
rect 1757 1877 1772 1883
rect 2116 1877 2131 1883
rect 2205 1877 2211 1897
rect 2349 1897 2380 1903
rect 2797 1903 2803 1916
rect 2765 1897 2803 1903
rect 2276 1877 2323 1883
rect 2429 1877 2444 1883
rect 2573 1883 2579 1896
rect 2652 1892 2660 1896
rect 2972 1892 2980 1896
rect 2461 1877 2483 1883
rect 2557 1877 2579 1883
rect 2637 1877 2659 1883
rect 2157 1857 2179 1863
rect 2580 1857 2595 1863
rect 2637 1857 2643 1877
rect 3021 1877 3036 1883
rect 2884 1857 2899 1863
rect 586 1836 588 1844
rect 986 1836 988 1844
rect 1124 1836 1126 1844
rect 1162 1836 1164 1844
rect 1242 1836 1244 1844
rect 2228 1836 2230 1844
rect 2500 1836 2502 1844
rect 2266 1814 2278 1816
rect 2251 1806 2253 1814
rect 2261 1806 2263 1814
rect 2271 1806 2273 1814
rect 2281 1806 2283 1814
rect 2291 1806 2293 1814
rect 2266 1804 2278 1806
rect 2938 1776 2940 1784
rect 109 1744 115 1763
rect 708 1757 723 1763
rect 77 1737 108 1743
rect 237 1737 307 1743
rect 141 1717 172 1723
rect 276 1717 291 1723
rect 397 1723 403 1743
rect 733 1743 739 1763
rect 1085 1757 1100 1763
rect 733 1737 835 1743
rect 1117 1737 1132 1743
rect 372 1717 403 1723
rect 861 1717 892 1723
rect 1069 1717 1100 1723
rect 1149 1723 1155 1743
rect 1188 1737 1203 1743
rect 1485 1737 1500 1743
rect 1549 1737 1587 1743
rect 1885 1737 1923 1743
rect 2276 1737 2339 1743
rect 2356 1737 2371 1743
rect 1140 1717 1155 1723
rect 1165 1717 1196 1723
rect 1229 1717 1267 1723
rect 548 1696 556 1704
rect 1053 1697 1075 1703
rect 1229 1697 1235 1717
rect 1773 1717 1811 1723
rect 1773 1697 1779 1717
rect 2028 1717 2067 1723
rect 2028 1712 2036 1717
rect 2221 1697 2259 1703
rect 2685 1697 2700 1703
rect 2964 1697 2979 1703
rect 1228 1684 1236 1688
rect 829 1677 844 1683
rect 1021 1677 1036 1683
rect 2196 1676 2198 1684
rect 2253 1677 2284 1683
rect 2541 1677 2556 1683
rect 1748 1656 1750 1664
rect 2541 1657 2547 1677
rect 362 1636 364 1644
rect 420 1636 422 1644
rect 964 1636 966 1644
rect 1514 1636 1516 1644
rect 2068 1636 2070 1644
rect 2756 1636 2758 1644
rect 2836 1636 2838 1644
rect 2884 1636 2886 1644
rect 762 1614 774 1616
rect 747 1606 749 1614
rect 757 1606 759 1614
rect 767 1606 769 1614
rect 777 1606 779 1614
rect 787 1606 789 1614
rect 762 1604 774 1606
rect 948 1576 950 1584
rect 685 1537 723 1543
rect 532 1516 540 1524
rect 189 1497 236 1503
rect 324 1497 355 1503
rect 564 1497 579 1503
rect 717 1497 723 1537
rect 2676 1537 2707 1543
rect 3021 1537 3036 1543
rect 820 1517 835 1523
rect 2413 1517 2435 1523
rect 2477 1517 2492 1523
rect 2669 1517 2684 1523
rect 772 1497 851 1503
rect 1357 1497 1372 1503
rect 1412 1497 1427 1503
rect 1460 1497 1475 1503
rect 1508 1497 1539 1503
rect 1556 1497 1587 1503
rect 1773 1484 1779 1503
rect 2125 1497 2140 1503
rect 2349 1497 2364 1503
rect 2076 1492 2084 1496
rect 301 1477 371 1483
rect 477 1477 515 1483
rect 964 1477 979 1483
rect 1364 1477 1395 1483
rect 1741 1477 1772 1483
rect 1901 1477 1923 1483
rect 2036 1477 2051 1483
rect 2061 1477 2083 1483
rect 205 1457 220 1463
rect 317 1457 332 1463
rect 1284 1457 1299 1463
rect 1508 1457 1516 1463
rect 2061 1457 2067 1477
rect 2788 1477 2803 1483
rect 2612 1457 2627 1463
rect 1626 1436 1628 1444
rect 2154 1436 2156 1444
rect 2712 1436 2716 1444
rect 2266 1414 2278 1416
rect 2251 1406 2253 1414
rect 2261 1406 2263 1414
rect 2271 1406 2273 1414
rect 2281 1406 2283 1414
rect 2291 1406 2293 1414
rect 2266 1404 2278 1406
rect 1588 1376 1598 1384
rect 2948 1376 2950 1384
rect 84 1357 99 1363
rect 733 1357 748 1363
rect 109 1337 131 1343
rect 212 1337 243 1343
rect 269 1337 284 1343
rect 420 1337 435 1343
rect 980 1337 995 1343
rect 1101 1343 1107 1363
rect 1716 1357 1731 1363
rect 1965 1357 1980 1363
rect 2429 1357 2444 1363
rect 1092 1337 1107 1343
rect 1229 1337 1244 1343
rect 1629 1337 1699 1343
rect 1972 1337 2003 1343
rect 2045 1337 2067 1343
rect 2164 1337 2195 1343
rect 2317 1337 2364 1343
rect 2733 1337 2755 1343
rect 29 1317 44 1323
rect 141 1317 172 1323
rect 285 1317 316 1323
rect 436 1317 451 1323
rect 868 1317 899 1323
rect 916 1317 947 1323
rect 1005 1317 1043 1323
rect 1037 1297 1043 1317
rect 1197 1317 1212 1323
rect 1293 1317 1324 1323
rect 2292 1317 2307 1323
rect 2429 1317 2451 1323
rect 2893 1317 2908 1323
rect 2093 1297 2115 1303
rect 2221 1297 2284 1303
rect 2669 1297 2691 1303
rect 2957 1297 2972 1303
rect 109 1277 124 1283
rect 1172 1277 1187 1283
rect 2045 1277 2060 1283
rect 58 1236 60 1244
rect 538 1236 540 1244
rect 586 1236 588 1244
rect 1524 1236 1526 1244
rect 2714 1236 2716 1244
rect 762 1214 774 1216
rect 747 1206 749 1214
rect 757 1206 759 1214
rect 767 1206 769 1214
rect 777 1206 779 1214
rect 787 1206 789 1214
rect 762 1204 774 1206
rect 170 1176 172 1184
rect 1732 1176 1734 1184
rect 2052 1176 2054 1184
rect 1332 1156 1334 1164
rect 1796 1156 1798 1164
rect 45 1137 60 1143
rect 316 1132 324 1136
rect 3005 1137 3036 1143
rect 844 1132 852 1136
rect 317 1117 355 1123
rect 173 1097 236 1103
rect 349 1097 387 1103
rect 445 1097 499 1103
rect 589 1103 595 1123
rect 676 1117 691 1123
rect 765 1117 851 1123
rect 1453 1117 1475 1123
rect 1556 1116 1564 1124
rect 548 1097 563 1103
rect 589 1097 627 1103
rect 637 1097 652 1103
rect 660 1097 675 1103
rect 52 1077 67 1083
rect 253 1077 284 1083
rect 669 1077 675 1097
rect 1220 1097 1235 1103
rect 1293 1097 1308 1103
rect 1693 1097 1708 1103
rect 2004 1097 2051 1103
rect 2445 1097 2460 1103
rect 2548 1097 2563 1103
rect 2717 1103 2723 1123
rect 2829 1117 2851 1123
rect 2717 1097 2755 1103
rect 2765 1097 2780 1103
rect 2845 1097 2876 1103
rect 1245 1077 1283 1083
rect 1277 1064 1283 1077
rect 2013 1077 2028 1083
rect 2100 1077 2115 1083
rect 2141 1077 2156 1083
rect 2141 1057 2147 1077
rect 2468 1077 2483 1083
rect 2788 1077 2803 1083
rect 2813 1077 2828 1083
rect 836 1037 851 1043
rect 938 1036 940 1044
rect 1844 1036 1848 1044
rect 2628 1036 2632 1044
rect 2708 1036 2710 1044
rect 2266 1014 2278 1016
rect 2251 1006 2253 1014
rect 2261 1006 2263 1014
rect 2271 1006 2273 1014
rect 2281 1006 2283 1014
rect 2291 1006 2293 1014
rect 2266 1004 2278 1006
rect 2602 976 2604 984
rect 205 957 259 963
rect 77 937 124 943
rect 276 937 307 943
rect 173 917 204 923
rect 228 917 243 923
rect 429 923 435 943
rect 717 943 723 963
rect 717 937 812 943
rect 829 937 844 943
rect 900 937 947 943
rect 1149 937 1203 943
rect 1844 937 1875 943
rect 2013 943 2019 956
rect 1940 937 1955 943
rect 1997 937 2019 943
rect 2029 937 2067 943
rect 429 917 451 923
rect 845 917 867 923
rect 1981 917 2012 923
rect 2157 923 2163 936
rect 2205 923 2211 963
rect 2228 937 2243 943
rect 2365 943 2371 963
rect 2749 957 2771 963
rect 2365 937 2396 943
rect 2477 943 2483 956
rect 2477 937 2499 943
rect 2157 917 2179 923
rect 2205 917 2220 923
rect 2324 917 2339 923
rect 2429 917 2444 923
rect 2893 923 2899 943
rect 2868 917 2899 923
rect 532 896 540 904
rect 1684 896 1692 904
rect 1917 897 1955 903
rect 2093 897 2115 903
rect 2932 896 2936 904
rect 1018 876 1020 884
rect 1252 836 1254 844
rect 1316 836 1318 844
rect 1556 836 1558 844
rect 2276 837 2339 843
rect 2516 836 2518 844
rect 762 814 774 816
rect 747 806 749 814
rect 757 806 759 814
rect 767 806 769 814
rect 777 806 779 814
rect 787 806 789 814
rect 762 804 774 806
rect 1060 776 1062 784
rect 1146 776 1148 784
rect 621 737 652 743
rect 1572 736 1574 744
rect 2004 736 2006 744
rect 2202 736 2204 744
rect 45 703 51 723
rect 477 717 499 723
rect 685 717 707 723
rect 1085 717 1107 723
rect 2317 717 2332 723
rect 45 697 60 703
rect 308 697 323 703
rect 333 697 348 703
rect 532 697 547 703
rect 749 697 812 703
rect 1044 697 1059 703
rect 1517 697 1571 703
rect 2301 703 2307 716
rect 2205 697 2307 703
rect 2637 697 2676 703
rect 2717 697 2739 703
rect 2668 692 2676 697
rect 100 677 115 683
rect 525 677 540 683
rect 573 677 604 683
rect 644 677 659 683
rect 1021 677 1043 683
rect 1277 677 1331 683
rect 1757 677 1795 683
rect 1860 677 1891 683
rect 1965 677 1980 683
rect 93 657 99 676
rect 1165 657 1180 663
rect 1908 656 1916 664
rect 1965 657 1971 677
rect 2445 677 2492 683
rect 2525 677 2547 683
rect 2733 677 2739 697
rect 2900 677 2915 683
rect 2132 657 2147 663
rect 2365 657 2380 663
rect 2909 657 2915 677
rect 2948 657 2972 663
rect 506 636 508 644
rect 2061 637 2076 643
rect 2970 636 2972 644
rect 3021 637 3036 643
rect 2266 614 2278 616
rect 2251 606 2253 614
rect 2261 606 2263 614
rect 2271 606 2273 614
rect 2281 606 2283 614
rect 2291 606 2293 614
rect 2266 604 2278 606
rect 186 576 188 584
rect 2013 544 2019 563
rect 2029 557 2044 563
rect 2573 557 2595 563
rect 29 537 51 543
rect 397 537 412 543
rect 612 537 643 543
rect 1028 537 1043 543
rect 1389 537 1404 543
rect 1560 537 1580 543
rect 1693 537 1715 543
rect 1997 537 2012 543
rect 2237 537 2252 543
rect 2605 537 2620 543
rect 61 517 92 523
rect 109 517 131 523
rect 1396 517 1427 523
rect 1917 517 1939 523
rect 2173 523 2179 536
rect 2157 517 2179 523
rect 2412 523 2420 528
rect 2397 517 2420 523
rect 77 497 115 503
rect 212 497 227 503
rect 20 477 35 483
rect 861 483 867 503
rect 1348 496 1358 504
rect 2397 497 2403 517
rect 2621 517 2643 523
rect 861 477 899 483
rect 330 456 332 464
rect 893 457 899 477
rect 948 477 963 483
rect 2372 456 2374 464
rect 138 436 140 444
rect 458 436 460 444
rect 538 436 540 444
rect 1124 436 1126 444
rect 762 414 774 416
rect 747 406 749 414
rect 757 406 759 414
rect 767 406 769 414
rect 777 406 779 414
rect 787 406 789 414
rect 762 404 774 406
rect 714 376 716 384
rect 874 376 876 384
rect 1130 376 1132 384
rect 1210 376 1212 384
rect 1572 376 1574 384
rect 1642 376 1644 384
rect 1690 376 1692 384
rect 1834 376 1836 384
rect 1988 376 1990 384
rect 237 337 252 343
rect 413 317 435 323
rect 301 297 316 303
rect 589 297 611 303
rect 925 297 940 303
rect 1213 297 1228 303
rect 1405 297 1459 303
rect 1517 297 1532 303
rect 1668 297 1683 303
rect 1837 297 1852 303
rect 2004 297 2019 303
rect 2093 297 2124 303
rect 2157 297 2188 303
rect 2461 297 2476 303
rect 2612 297 2627 303
rect 2957 297 2979 303
rect 349 283 355 296
rect 244 277 259 283
rect 349 277 371 283
rect 1364 277 1379 283
rect 1485 277 1500 283
rect 1533 277 1555 283
rect 1613 277 1628 283
rect 1533 264 1539 277
rect 1876 277 1891 283
rect 1901 277 1916 283
rect 1949 277 1971 283
rect 1965 264 1971 277
rect 2797 277 2812 283
rect 3005 277 3036 283
rect 1924 256 1932 264
rect 2260 257 2316 263
rect 2868 237 2883 243
rect 2932 237 2947 243
rect 2266 214 2278 216
rect 2251 206 2253 214
rect 2261 206 2263 214
rect 2271 206 2273 214
rect 2281 206 2283 214
rect 2291 206 2293 214
rect 2266 204 2278 206
rect 68 176 70 184
rect 1082 176 1084 184
rect 1994 176 1996 184
rect 2228 176 2230 184
rect 2420 176 2424 184
rect 989 157 1004 163
rect 548 137 579 143
rect 589 137 611 143
rect 669 137 700 143
rect 932 137 947 143
rect 1309 137 1331 143
rect 1212 124 1220 128
rect 1325 124 1331 137
rect 1565 143 1571 163
rect 1565 137 1587 143
rect 1805 137 1820 143
rect 1940 137 1955 143
rect 2045 137 2060 143
rect 2141 143 2147 163
rect 2141 137 2156 143
rect 2173 137 2211 143
rect 2356 137 2387 143
rect 2628 137 2675 143
rect 2765 143 2771 163
rect 2765 137 2803 143
rect 1580 124 1588 128
rect 141 117 172 123
rect 628 117 659 123
rect 1757 117 1772 123
rect 1789 117 1804 123
rect 1828 117 1843 123
rect 1869 117 1907 123
rect 125 97 147 103
rect 164 97 179 103
rect 333 97 348 103
rect 1757 97 1779 103
rect 1869 97 1875 117
rect 2109 117 2131 123
rect 2525 117 2563 123
rect 2237 97 2323 103
rect 2525 97 2531 117
rect 2701 117 2723 123
rect 2877 117 2915 123
rect 1980 84 1988 88
rect 1316 77 1331 83
rect 3021 77 3036 83
rect 762 14 774 16
rect 747 6 749 14
rect 757 6 759 14
rect 767 6 769 14
rect 777 6 779 14
rect 787 6 789 14
rect 762 4 774 6
<< m2contact >>
rect 739 2006 747 2014
rect 749 2006 757 2014
rect 759 2006 767 2014
rect 769 2006 777 2014
rect 779 2006 787 2014
rect 789 2006 797 2014
rect 796 1976 804 1984
rect 1388 1976 1396 1984
rect 1436 1976 1444 1984
rect 860 1936 868 1944
rect 2060 1936 2068 1944
rect 2412 1936 2420 1944
rect 44 1916 52 1924
rect 76 1916 84 1924
rect 332 1916 340 1924
rect 572 1916 580 1924
rect 844 1916 852 1924
rect 892 1916 900 1924
rect 972 1916 980 1924
rect 1020 1916 1028 1924
rect 1084 1916 1092 1924
rect 1132 1916 1140 1924
rect 1612 1916 1620 1924
rect 1852 1916 1860 1924
rect 2092 1916 2100 1924
rect 2172 1916 2180 1924
rect 188 1896 196 1904
rect 300 1896 308 1904
rect 396 1896 404 1904
rect 508 1896 516 1904
rect 684 1896 692 1904
rect 700 1896 708 1904
rect 1276 1896 1284 1904
rect 1356 1896 1364 1904
rect 1404 1896 1412 1904
rect 1660 1896 1668 1904
rect 1708 1896 1716 1904
rect 1740 1896 1748 1904
rect 1852 1896 1860 1904
rect 1884 1896 1892 1904
rect 1980 1896 1988 1904
rect 2044 1896 2052 1904
rect 2076 1896 2084 1904
rect 2108 1896 2116 1904
rect 2364 1916 2372 1924
rect 2380 1916 2388 1924
rect 2508 1916 2516 1924
rect 2524 1916 2532 1924
rect 2764 1916 2772 1924
rect 2796 1916 2804 1924
rect 2828 1916 2836 1924
rect 44 1876 52 1884
rect 92 1876 100 1884
rect 12 1856 20 1864
rect 124 1856 132 1864
rect 172 1876 180 1884
rect 284 1876 292 1884
rect 364 1876 372 1884
rect 460 1876 468 1884
rect 524 1876 532 1884
rect 604 1876 612 1884
rect 636 1876 644 1884
rect 668 1876 676 1884
rect 892 1876 900 1884
rect 924 1876 932 1884
rect 1004 1876 1012 1884
rect 1052 1876 1060 1884
rect 1100 1876 1108 1884
rect 1180 1876 1188 1884
rect 1260 1876 1268 1884
rect 444 1856 452 1864
rect 556 1856 564 1864
rect 652 1856 660 1864
rect 812 1856 820 1864
rect 956 1856 964 1864
rect 1068 1856 1076 1864
rect 1196 1856 1204 1864
rect 1212 1856 1220 1864
rect 1676 1876 1684 1884
rect 1692 1876 1700 1884
rect 1772 1876 1780 1884
rect 1868 1876 1876 1884
rect 1900 1876 1908 1884
rect 1916 1876 1924 1884
rect 1932 1880 1940 1888
rect 1996 1876 2004 1884
rect 2108 1876 2116 1884
rect 2188 1876 2196 1884
rect 2332 1896 2340 1904
rect 2380 1896 2388 1904
rect 2412 1896 2420 1904
rect 2572 1896 2580 1904
rect 2652 1896 2660 1904
rect 2668 1896 2676 1904
rect 2732 1896 2740 1904
rect 2876 1896 2884 1904
rect 2956 1896 2964 1904
rect 2972 1896 2980 1904
rect 2988 1896 2996 1904
rect 2268 1876 2276 1884
rect 2444 1876 2452 1884
rect 2620 1876 2628 1884
rect 1340 1856 1348 1864
rect 1420 1856 1428 1864
rect 1500 1856 1508 1864
rect 1516 1856 1524 1864
rect 1564 1856 1572 1864
rect 1580 1856 1588 1864
rect 1612 1856 1620 1864
rect 1708 1856 1716 1864
rect 1836 1856 1844 1864
rect 2012 1856 2020 1864
rect 2028 1856 2036 1864
rect 2444 1856 2452 1864
rect 2572 1856 2580 1864
rect 2604 1856 2612 1864
rect 2716 1876 2724 1884
rect 2780 1876 2788 1884
rect 2828 1876 2836 1884
rect 3036 1876 3044 1884
rect 2860 1856 2868 1864
rect 2876 1856 2884 1864
rect 2908 1856 2916 1864
rect 156 1836 164 1844
rect 252 1836 260 1844
rect 332 1836 340 1844
rect 428 1836 436 1844
rect 540 1836 548 1844
rect 588 1836 596 1844
rect 892 1836 900 1844
rect 988 1836 996 1844
rect 1020 1836 1028 1844
rect 1116 1836 1124 1844
rect 1164 1836 1172 1844
rect 1244 1836 1252 1844
rect 1324 1836 1332 1844
rect 1628 1836 1636 1844
rect 1804 1836 1812 1844
rect 1964 1836 1972 1844
rect 2140 1836 2148 1844
rect 2220 1836 2228 1844
rect 2492 1836 2500 1844
rect 2524 1836 2532 1844
rect 2700 1836 2708 1844
rect 2796 1836 2804 1844
rect 2924 1836 2932 1844
rect 2243 1806 2251 1814
rect 2253 1806 2261 1814
rect 2263 1806 2271 1814
rect 2273 1806 2281 1814
rect 2283 1806 2291 1814
rect 2293 1806 2301 1814
rect 236 1776 244 1784
rect 636 1776 644 1784
rect 1852 1776 1860 1784
rect 2460 1776 2468 1784
rect 2940 1776 2948 1784
rect 92 1756 100 1764
rect 252 1756 260 1764
rect 316 1756 324 1764
rect 700 1756 708 1764
rect 108 1736 116 1744
rect 380 1736 388 1744
rect 44 1716 52 1724
rect 60 1716 68 1724
rect 124 1716 132 1724
rect 172 1716 180 1724
rect 220 1716 228 1724
rect 268 1716 276 1724
rect 364 1716 372 1724
rect 572 1736 580 1744
rect 588 1736 596 1744
rect 684 1736 692 1744
rect 812 1756 820 1764
rect 892 1756 900 1764
rect 1100 1756 1108 1764
rect 1244 1756 1252 1764
rect 1340 1756 1348 1764
rect 1420 1756 1428 1764
rect 1532 1756 1540 1764
rect 1564 1756 1572 1764
rect 1628 1756 1636 1764
rect 1836 1756 1844 1764
rect 1900 1756 1908 1764
rect 2236 1756 2244 1764
rect 2348 1756 2356 1764
rect 2444 1756 2452 1764
rect 2700 1756 2708 1764
rect 2812 1756 2820 1764
rect 2988 1756 2996 1764
rect 844 1736 852 1744
rect 940 1736 948 1744
rect 1132 1736 1140 1744
rect 412 1716 420 1724
rect 492 1716 500 1724
rect 556 1716 564 1724
rect 604 1716 612 1724
rect 700 1716 708 1724
rect 892 1716 900 1724
rect 924 1716 932 1724
rect 956 1716 964 1724
rect 1036 1716 1044 1724
rect 1100 1716 1108 1724
rect 1132 1716 1140 1724
rect 1180 1736 1188 1744
rect 1292 1736 1300 1744
rect 1404 1736 1412 1744
rect 1500 1736 1508 1744
rect 1660 1736 1668 1744
rect 1692 1736 1700 1744
rect 1724 1736 1732 1744
rect 1820 1736 1828 1744
rect 2044 1736 2052 1744
rect 2172 1736 2180 1744
rect 2268 1736 2276 1744
rect 2348 1736 2356 1744
rect 2396 1736 2404 1744
rect 2428 1736 2436 1744
rect 2476 1736 2484 1744
rect 2572 1736 2580 1744
rect 2620 1736 2628 1744
rect 2732 1736 2740 1744
rect 2796 1736 2804 1744
rect 2860 1736 2868 1744
rect 2956 1736 2964 1744
rect 1196 1716 1204 1724
rect 332 1696 340 1704
rect 444 1696 452 1704
rect 508 1696 516 1704
rect 524 1696 532 1704
rect 556 1696 564 1704
rect 636 1696 644 1704
rect 652 1696 660 1704
rect 668 1696 676 1704
rect 876 1696 884 1704
rect 988 1696 996 1704
rect 1180 1696 1188 1704
rect 1276 1716 1284 1724
rect 1468 1716 1476 1724
rect 1500 1716 1508 1724
rect 1596 1716 1604 1724
rect 1644 1716 1652 1724
rect 1708 1716 1716 1724
rect 1740 1716 1748 1724
rect 1324 1696 1332 1704
rect 1628 1696 1636 1704
rect 1868 1716 1876 1724
rect 1932 1716 1940 1724
rect 1948 1716 1956 1724
rect 2012 1716 2020 1724
rect 2124 1716 2132 1724
rect 2188 1716 2196 1724
rect 2380 1716 2388 1724
rect 2412 1716 2420 1724
rect 2492 1716 2500 1724
rect 2540 1716 2548 1724
rect 2588 1716 2596 1724
rect 2668 1716 2676 1724
rect 2748 1716 2756 1724
rect 2780 1716 2788 1724
rect 2844 1716 2852 1724
rect 2876 1716 2884 1724
rect 1788 1696 1796 1704
rect 1964 1696 1972 1704
rect 2028 1696 2036 1704
rect 2092 1696 2100 1704
rect 2108 1696 2116 1704
rect 2556 1696 2564 1704
rect 2620 1696 2628 1704
rect 2700 1696 2708 1704
rect 2716 1696 2724 1704
rect 2908 1696 2916 1704
rect 2924 1696 2932 1704
rect 2956 1696 2964 1704
rect 12 1676 20 1684
rect 476 1676 484 1684
rect 844 1676 852 1684
rect 1036 1676 1044 1684
rect 1228 1676 1236 1684
rect 1356 1676 1364 1684
rect 1996 1676 2004 1684
rect 2140 1676 2148 1684
rect 2188 1676 2196 1684
rect 2284 1676 2292 1684
rect 2524 1676 2532 1684
rect 1740 1656 1748 1664
rect 2012 1656 2020 1664
rect 2556 1676 2564 1684
rect 2652 1676 2660 1684
rect 364 1636 372 1644
rect 412 1636 420 1644
rect 492 1636 500 1644
rect 924 1636 932 1644
rect 956 1636 964 1644
rect 1036 1636 1044 1644
rect 1212 1636 1220 1644
rect 1308 1636 1316 1644
rect 1372 1636 1380 1644
rect 1436 1636 1444 1644
rect 1516 1636 1524 1644
rect 1660 1636 1668 1644
rect 2060 1636 2068 1644
rect 2156 1636 2164 1644
rect 2668 1636 2676 1644
rect 2748 1636 2756 1644
rect 2828 1636 2836 1644
rect 2876 1636 2884 1644
rect 739 1606 747 1614
rect 749 1606 757 1614
rect 759 1606 767 1614
rect 769 1606 777 1614
rect 779 1606 787 1614
rect 789 1606 797 1614
rect 396 1576 404 1584
rect 940 1576 948 1584
rect 1916 1556 1924 1564
rect 412 1536 420 1544
rect 668 1536 676 1544
rect 108 1516 116 1524
rect 444 1516 452 1524
rect 524 1516 532 1524
rect 556 1516 564 1524
rect 636 1516 644 1524
rect 700 1516 708 1524
rect 28 1496 36 1504
rect 156 1496 164 1504
rect 172 1496 180 1504
rect 236 1496 244 1504
rect 284 1496 292 1504
rect 316 1496 324 1504
rect 428 1496 436 1504
rect 492 1496 500 1504
rect 524 1496 532 1504
rect 556 1496 564 1504
rect 604 1496 612 1504
rect 652 1496 660 1504
rect 732 1536 740 1544
rect 1116 1536 1124 1544
rect 2668 1536 2676 1544
rect 3036 1536 3044 1544
rect 812 1516 820 1524
rect 1020 1516 1028 1524
rect 1084 1516 1092 1524
rect 1148 1516 1156 1524
rect 1596 1516 1604 1524
rect 1612 1516 1620 1524
rect 2140 1516 2148 1524
rect 2236 1516 2244 1524
rect 2492 1516 2500 1524
rect 2684 1516 2692 1524
rect 764 1496 772 1504
rect 860 1496 868 1504
rect 956 1496 964 1504
rect 988 1496 996 1504
rect 1068 1496 1076 1504
rect 1100 1496 1108 1504
rect 1180 1496 1188 1504
rect 1260 1496 1268 1504
rect 1276 1496 1284 1504
rect 1372 1496 1380 1504
rect 1404 1496 1412 1504
rect 1452 1496 1460 1504
rect 1500 1496 1508 1504
rect 1548 1496 1556 1504
rect 1756 1496 1764 1504
rect 1852 1496 1860 1504
rect 1884 1496 1892 1504
rect 1964 1496 1972 1504
rect 1996 1496 2004 1504
rect 2028 1496 2036 1504
rect 2076 1496 2084 1504
rect 2140 1496 2148 1504
rect 2204 1496 2212 1504
rect 2364 1496 2372 1504
rect 2380 1496 2388 1504
rect 2508 1496 2516 1504
rect 2524 1496 2532 1504
rect 2556 1496 2564 1504
rect 2588 1496 2596 1504
rect 2652 1496 2660 1504
rect 2684 1496 2692 1504
rect 2732 1496 2740 1504
rect 2764 1496 2772 1504
rect 2812 1496 2820 1504
rect 2844 1496 2852 1504
rect 2924 1496 2932 1504
rect 2972 1496 2980 1504
rect 2988 1496 2996 1504
rect 12 1476 20 1484
rect 76 1476 84 1484
rect 620 1476 628 1484
rect 732 1476 740 1484
rect 876 1476 884 1484
rect 956 1476 964 1484
rect 1004 1476 1012 1484
rect 1164 1476 1172 1484
rect 1196 1476 1204 1484
rect 1244 1476 1252 1484
rect 1356 1476 1364 1484
rect 1564 1476 1572 1484
rect 1644 1476 1652 1484
rect 1676 1476 1684 1484
rect 1772 1476 1780 1484
rect 1788 1476 1796 1484
rect 1836 1476 1844 1484
rect 1868 1476 1876 1484
rect 1948 1476 1956 1484
rect 1980 1476 1988 1484
rect 2012 1476 2020 1484
rect 2028 1476 2036 1484
rect 2092 1480 2100 1488
rect 124 1456 132 1464
rect 220 1456 228 1464
rect 332 1456 340 1464
rect 380 1456 388 1464
rect 460 1456 468 1464
rect 892 1456 900 1464
rect 924 1456 932 1464
rect 1036 1456 1044 1464
rect 1212 1456 1220 1464
rect 1276 1456 1284 1464
rect 1308 1456 1316 1464
rect 1324 1456 1332 1464
rect 1372 1456 1380 1464
rect 1452 1456 1460 1464
rect 1500 1456 1508 1464
rect 1516 1456 1524 1464
rect 1660 1456 1668 1464
rect 1724 1456 1732 1464
rect 1820 1456 1828 1464
rect 1932 1456 1940 1464
rect 2172 1476 2180 1484
rect 2188 1476 2196 1484
rect 2220 1476 2228 1484
rect 2364 1476 2372 1484
rect 2540 1476 2548 1484
rect 2572 1476 2580 1484
rect 2748 1476 2756 1484
rect 2780 1476 2788 1484
rect 2860 1476 2868 1484
rect 2908 1476 2916 1484
rect 2940 1476 2948 1484
rect 2316 1456 2324 1464
rect 2412 1456 2420 1464
rect 2444 1456 2452 1464
rect 2460 1456 2468 1464
rect 2604 1456 2612 1464
rect 2780 1456 2788 1464
rect 2844 1456 2852 1464
rect 2876 1456 2884 1464
rect 60 1436 68 1444
rect 108 1436 116 1444
rect 140 1436 148 1444
rect 300 1436 308 1444
rect 908 1436 916 1444
rect 1052 1436 1060 1444
rect 1116 1436 1124 1444
rect 1228 1436 1236 1444
rect 1340 1436 1348 1444
rect 1436 1436 1444 1444
rect 1484 1436 1492 1444
rect 1628 1436 1636 1444
rect 1708 1436 1716 1444
rect 1804 1436 1812 1444
rect 2156 1436 2164 1444
rect 2332 1436 2340 1444
rect 2636 1436 2644 1444
rect 2716 1436 2724 1444
rect 2892 1436 2900 1444
rect 2243 1406 2251 1414
rect 2253 1406 2261 1414
rect 2263 1406 2271 1414
rect 2273 1406 2281 1414
rect 2283 1406 2291 1414
rect 2293 1406 2301 1414
rect 204 1376 212 1384
rect 332 1376 340 1384
rect 588 1376 596 1384
rect 956 1376 964 1384
rect 1580 1376 1588 1384
rect 1820 1376 1828 1384
rect 1948 1376 1956 1384
rect 2108 1376 2116 1384
rect 2572 1376 2580 1384
rect 2940 1376 2948 1384
rect 12 1356 20 1364
rect 76 1356 84 1364
rect 316 1356 324 1364
rect 604 1356 612 1364
rect 620 1356 628 1364
rect 748 1356 756 1364
rect 812 1356 820 1364
rect 972 1356 980 1364
rect 1036 1356 1044 1364
rect 172 1336 180 1344
rect 204 1336 212 1344
rect 284 1336 292 1344
rect 332 1336 340 1344
rect 412 1336 420 1344
rect 460 1336 468 1344
rect 492 1336 500 1344
rect 556 1336 564 1344
rect 652 1336 660 1344
rect 716 1336 724 1344
rect 844 1336 852 1344
rect 924 1336 932 1344
rect 972 1336 980 1344
rect 1084 1336 1092 1344
rect 1212 1356 1220 1364
rect 1324 1356 1332 1364
rect 1500 1356 1508 1364
rect 1644 1356 1652 1364
rect 1676 1356 1684 1364
rect 1708 1356 1716 1364
rect 1740 1356 1748 1364
rect 1836 1356 1844 1364
rect 1980 1356 1988 1364
rect 2028 1356 2036 1364
rect 2124 1356 2132 1364
rect 2220 1356 2228 1364
rect 2332 1356 2340 1364
rect 2396 1356 2404 1364
rect 2412 1356 2420 1364
rect 2444 1356 2452 1364
rect 2476 1356 2484 1364
rect 2668 1356 2676 1364
rect 2844 1356 2852 1364
rect 2972 1356 2980 1364
rect 2988 1356 2996 1364
rect 1244 1336 1252 1344
rect 1260 1336 1268 1344
rect 1756 1336 1764 1344
rect 1804 1336 1812 1344
rect 1932 1336 1940 1344
rect 1964 1336 1972 1344
rect 2156 1336 2164 1344
rect 2364 1336 2372 1344
rect 2460 1336 2468 1344
rect 2492 1336 2500 1344
rect 2556 1336 2564 1344
rect 2604 1336 2612 1344
rect 2636 1336 2644 1344
rect 2796 1336 2804 1344
rect 2908 1336 2916 1344
rect 2924 1336 2932 1344
rect 44 1316 52 1324
rect 172 1316 180 1324
rect 220 1316 228 1324
rect 252 1316 260 1324
rect 316 1316 324 1324
rect 348 1316 356 1324
rect 428 1316 436 1324
rect 476 1316 484 1324
rect 540 1316 548 1324
rect 572 1316 580 1324
rect 668 1316 676 1324
rect 828 1316 836 1324
rect 860 1316 868 1324
rect 908 1316 916 1324
rect 156 1296 164 1304
rect 204 1296 212 1304
rect 508 1296 516 1304
rect 876 1296 884 1304
rect 1020 1296 1028 1304
rect 1068 1316 1076 1324
rect 1116 1316 1124 1324
rect 1132 1316 1140 1324
rect 1164 1316 1172 1324
rect 1212 1316 1220 1324
rect 1244 1316 1252 1324
rect 1276 1316 1284 1324
rect 1324 1316 1332 1324
rect 1356 1316 1364 1324
rect 1388 1316 1396 1324
rect 1452 1316 1460 1324
rect 1532 1316 1540 1324
rect 1612 1316 1620 1324
rect 1708 1316 1716 1324
rect 1772 1316 1780 1324
rect 1788 1316 1796 1324
rect 1868 1316 1876 1324
rect 1916 1316 1924 1324
rect 2012 1316 2020 1324
rect 2172 1316 2180 1324
rect 2284 1316 2292 1324
rect 2348 1316 2356 1324
rect 2508 1316 2516 1324
rect 2524 1316 2532 1324
rect 2540 1316 2548 1324
rect 2620 1316 2628 1324
rect 2716 1316 2724 1324
rect 2780 1316 2788 1324
rect 2812 1316 2820 1324
rect 2876 1316 2884 1324
rect 2908 1316 2916 1324
rect 1148 1296 1156 1304
rect 1308 1296 1316 1304
rect 1372 1296 1380 1304
rect 1436 1296 1444 1304
rect 1852 1296 1860 1304
rect 2284 1296 2292 1304
rect 2572 1296 2580 1304
rect 2748 1296 2756 1304
rect 2860 1296 2868 1304
rect 2972 1296 2980 1304
rect 124 1276 132 1284
rect 1164 1276 1172 1284
rect 1404 1276 1412 1284
rect 1468 1276 1476 1284
rect 1884 1276 1892 1284
rect 2060 1276 2068 1284
rect 1452 1256 1460 1264
rect 2396 1256 2404 1264
rect 60 1236 68 1244
rect 540 1236 548 1244
rect 588 1236 596 1244
rect 620 1236 628 1244
rect 684 1236 692 1244
rect 1356 1236 1364 1244
rect 1388 1236 1396 1244
rect 1516 1236 1524 1244
rect 1868 1236 1876 1244
rect 2076 1236 2084 1244
rect 2140 1236 2148 1244
rect 2716 1236 2724 1244
rect 2812 1236 2820 1244
rect 739 1206 747 1214
rect 749 1206 757 1214
rect 759 1206 767 1214
rect 769 1206 777 1214
rect 779 1206 787 1214
rect 789 1206 797 1214
rect 172 1176 180 1184
rect 1628 1176 1636 1184
rect 1692 1176 1700 1184
rect 1724 1176 1732 1184
rect 1916 1176 1924 1184
rect 2044 1176 2052 1184
rect 444 1156 452 1164
rect 1324 1156 1332 1164
rect 1436 1156 1444 1164
rect 1788 1156 1796 1164
rect 2524 1156 2532 1164
rect 60 1136 68 1144
rect 316 1136 324 1144
rect 844 1136 852 1144
rect 1420 1136 1428 1144
rect 1484 1136 1492 1144
rect 1612 1136 1620 1144
rect 1852 1136 1860 1144
rect 1932 1136 1940 1144
rect 2636 1136 2644 1144
rect 3036 1136 3044 1144
rect 268 1116 276 1124
rect 364 1116 372 1124
rect 524 1116 532 1124
rect 44 1096 52 1104
rect 76 1096 84 1104
rect 140 1096 148 1104
rect 236 1096 244 1104
rect 508 1096 516 1104
rect 540 1096 548 1104
rect 604 1116 612 1124
rect 668 1116 676 1124
rect 700 1116 708 1124
rect 1020 1116 1028 1124
rect 1164 1116 1172 1124
rect 1356 1116 1364 1124
rect 1516 1116 1524 1124
rect 1548 1116 1556 1124
rect 1580 1116 1588 1124
rect 1644 1116 1652 1124
rect 1756 1116 1764 1124
rect 1820 1116 1828 1124
rect 1884 1116 1892 1124
rect 1900 1116 1908 1124
rect 1964 1116 1972 1124
rect 2076 1116 2084 1124
rect 2508 1116 2516 1124
rect 2668 1116 2676 1124
rect 652 1096 660 1104
rect 44 1076 52 1084
rect 124 1076 132 1084
rect 188 1076 196 1084
rect 204 1076 212 1084
rect 236 1076 244 1084
rect 284 1076 292 1084
rect 332 1076 340 1084
rect 396 1076 404 1084
rect 476 1076 484 1084
rect 540 1076 548 1084
rect 620 1076 628 1084
rect 652 1076 660 1084
rect 732 1096 740 1104
rect 892 1096 900 1104
rect 956 1096 964 1104
rect 972 1096 980 1104
rect 1036 1096 1044 1104
rect 1084 1096 1092 1104
rect 1148 1096 1156 1104
rect 1180 1096 1188 1104
rect 1196 1096 1204 1104
rect 1212 1096 1220 1104
rect 1308 1096 1316 1104
rect 1324 1096 1332 1104
rect 1388 1096 1396 1104
rect 1436 1096 1444 1104
rect 1500 1096 1508 1104
rect 1548 1096 1556 1104
rect 1628 1096 1636 1104
rect 1708 1096 1716 1104
rect 1724 1096 1732 1104
rect 1788 1096 1796 1104
rect 1868 1096 1876 1104
rect 1916 1096 1924 1104
rect 1996 1096 2004 1104
rect 2092 1096 2100 1104
rect 2204 1096 2212 1104
rect 2252 1096 2260 1104
rect 2332 1096 2340 1104
rect 2460 1096 2468 1104
rect 2540 1096 2548 1104
rect 2652 1096 2660 1104
rect 2732 1116 2740 1124
rect 2924 1116 2932 1124
rect 2780 1096 2788 1104
rect 2876 1096 2884 1104
rect 2908 1096 2916 1104
rect 2972 1096 2980 1104
rect 716 1076 724 1084
rect 876 1076 884 1084
rect 908 1076 916 1084
rect 940 1076 948 1084
rect 988 1076 996 1084
rect 1052 1076 1060 1084
rect 1132 1076 1140 1084
rect 1212 1076 1220 1084
rect 1308 1076 1316 1084
rect 1532 1076 1540 1084
rect 1708 1076 1716 1084
rect 1772 1076 1780 1084
rect 2028 1076 2036 1084
rect 2092 1076 2100 1084
rect 12 1056 20 1064
rect 428 1056 436 1064
rect 460 1056 468 1064
rect 1020 1056 1028 1064
rect 1084 1056 1092 1064
rect 1100 1056 1108 1064
rect 1260 1056 1268 1064
rect 1276 1056 1284 1064
rect 1372 1056 1380 1064
rect 1660 1056 1668 1064
rect 2156 1076 2164 1084
rect 2188 1076 2196 1084
rect 2348 1076 2356 1084
rect 2412 1076 2420 1084
rect 2460 1076 2468 1084
rect 2492 1076 2500 1084
rect 2540 1076 2548 1084
rect 2572 1076 2580 1084
rect 2684 1076 2692 1084
rect 2780 1076 2788 1084
rect 2828 1076 2836 1084
rect 2956 1076 2964 1084
rect 2156 1056 2164 1064
rect 2220 1056 2228 1064
rect 2380 1056 2388 1064
rect 2396 1056 2404 1064
rect 2604 1056 2612 1064
rect 2860 1056 2868 1064
rect 2876 1056 2884 1064
rect 108 1036 116 1044
rect 316 1036 324 1044
rect 412 1036 420 1044
rect 588 1036 596 1044
rect 828 1036 836 1044
rect 940 1036 948 1044
rect 1116 1036 1124 1044
rect 1836 1036 1844 1044
rect 1964 1036 1972 1044
rect 2124 1036 2132 1044
rect 2172 1036 2180 1044
rect 2236 1036 2244 1044
rect 2364 1036 2372 1044
rect 2588 1036 2596 1044
rect 2620 1036 2628 1044
rect 2700 1036 2708 1044
rect 2892 1036 2900 1044
rect 2924 1036 2932 1044
rect 2243 1006 2251 1014
rect 2253 1006 2261 1014
rect 2263 1006 2271 1014
rect 2273 1006 2281 1014
rect 2283 1006 2291 1014
rect 2293 1006 2301 1014
rect 380 976 388 984
rect 1452 976 1460 984
rect 1516 976 1524 984
rect 1820 976 1828 984
rect 2108 976 2116 984
rect 2188 976 2196 984
rect 2604 976 2612 984
rect 3020 976 3028 984
rect 60 956 68 964
rect 268 956 276 964
rect 284 956 292 964
rect 364 956 372 964
rect 572 956 580 964
rect 124 936 132 944
rect 156 936 164 944
rect 188 936 196 944
rect 268 936 276 944
rect 44 916 52 924
rect 92 916 100 924
rect 204 916 212 924
rect 220 916 228 924
rect 316 916 324 924
rect 332 916 340 924
rect 412 916 420 924
rect 492 936 500 944
rect 508 936 516 944
rect 604 936 612 944
rect 796 956 804 964
rect 908 956 916 964
rect 972 956 980 964
rect 1116 956 1124 964
rect 1468 956 1476 964
rect 1644 956 1652 964
rect 1836 956 1844 964
rect 1900 956 1908 964
rect 1932 956 1940 964
rect 2012 956 2020 964
rect 2092 956 2100 964
rect 812 936 820 944
rect 844 936 852 944
rect 892 936 900 944
rect 1036 936 1044 944
rect 1132 936 1140 944
rect 1212 936 1220 944
rect 1228 936 1236 944
rect 1292 936 1300 944
rect 1436 936 1444 944
rect 1484 936 1492 944
rect 1532 936 1540 944
rect 1612 936 1620 944
rect 1660 936 1668 944
rect 1804 936 1812 944
rect 1836 936 1844 944
rect 1932 936 1940 944
rect 2156 936 2164 944
rect 476 916 484 924
rect 524 916 532 924
rect 572 916 580 924
rect 620 916 628 924
rect 668 916 676 924
rect 924 916 932 924
rect 956 916 964 924
rect 1020 916 1028 924
rect 1068 916 1076 924
rect 1164 916 1172 924
rect 1244 916 1252 924
rect 1308 916 1316 924
rect 1388 916 1396 924
rect 1420 916 1428 924
rect 1548 916 1556 924
rect 1596 916 1604 924
rect 1676 916 1684 924
rect 1756 916 1764 924
rect 1788 916 1796 924
rect 1852 916 1860 924
rect 1884 916 1892 924
rect 2012 916 2020 924
rect 2044 916 2052 924
rect 2140 916 2148 924
rect 2220 936 2228 944
rect 2252 936 2260 944
rect 2380 956 2388 964
rect 2476 956 2484 964
rect 3004 956 3012 964
rect 2396 936 2404 944
rect 2572 936 2580 944
rect 2620 936 2628 944
rect 2700 936 2708 944
rect 2796 936 2804 944
rect 2828 936 2836 944
rect 2876 936 2884 944
rect 2220 916 2228 924
rect 2316 916 2324 924
rect 2444 916 2452 924
rect 2508 916 2516 924
rect 2652 916 2660 924
rect 2716 916 2724 924
rect 2780 916 2788 924
rect 2812 916 2820 924
rect 2860 916 2868 924
rect 2988 936 2996 944
rect 348 896 356 904
rect 380 896 388 904
rect 524 896 532 904
rect 556 896 564 904
rect 684 896 692 904
rect 988 896 996 904
rect 1052 896 1060 904
rect 1180 896 1188 904
rect 1276 896 1284 904
rect 1340 896 1348 904
rect 1404 896 1412 904
rect 1516 896 1524 904
rect 1580 896 1588 904
rect 1676 896 1684 904
rect 1708 896 1716 904
rect 1772 896 1780 904
rect 2220 896 2228 904
rect 2540 896 2548 904
rect 2588 896 2596 904
rect 2636 896 2644 904
rect 2748 896 2756 904
rect 2828 896 2836 904
rect 2924 896 2932 904
rect 12 876 20 884
rect 652 876 660 884
rect 1020 876 1028 884
rect 1084 876 1092 884
rect 1372 876 1380 884
rect 1644 876 1652 884
rect 1740 876 1748 884
rect 2668 876 2676 884
rect 668 836 676 844
rect 700 836 708 844
rect 1100 836 1108 844
rect 1244 836 1252 844
rect 1308 836 1316 844
rect 1356 836 1364 844
rect 1548 836 1556 844
rect 1724 836 1732 844
rect 2268 836 2276 844
rect 2444 836 2452 844
rect 2508 836 2516 844
rect 2556 836 2564 844
rect 2684 836 2692 844
rect 739 806 747 814
rect 749 806 757 814
rect 759 806 767 814
rect 769 806 777 814
rect 779 806 787 814
rect 789 806 797 814
rect 924 776 932 784
rect 1052 776 1060 784
rect 1148 776 1156 784
rect 1628 776 1636 784
rect 1660 776 1668 784
rect 1852 756 1860 764
rect 460 736 468 744
rect 652 736 660 744
rect 908 736 916 744
rect 1564 736 1572 744
rect 1676 736 1684 744
rect 1756 736 1764 744
rect 1996 736 2004 744
rect 2060 736 2068 744
rect 2140 736 2148 744
rect 2204 736 2212 744
rect 2364 736 2372 744
rect 2940 736 2948 744
rect 428 716 436 724
rect 604 716 612 724
rect 828 716 836 724
rect 940 716 948 724
rect 1500 716 1508 724
rect 1596 716 1604 724
rect 1644 716 1652 724
rect 1948 716 1956 724
rect 2028 716 2036 724
rect 2092 716 2100 724
rect 2108 716 2116 724
rect 2172 716 2180 724
rect 2300 716 2308 724
rect 2332 716 2340 724
rect 2396 716 2404 724
rect 2604 716 2612 724
rect 2780 716 2788 724
rect 2844 716 2852 724
rect 2956 716 2964 724
rect 60 696 68 704
rect 124 696 132 704
rect 188 696 196 704
rect 220 696 228 704
rect 268 696 276 704
rect 300 696 308 704
rect 348 696 356 704
rect 412 696 420 704
rect 444 696 452 704
rect 524 696 532 704
rect 588 696 596 704
rect 812 696 820 704
rect 860 696 868 704
rect 924 696 932 704
rect 988 696 996 704
rect 1036 696 1044 704
rect 1132 696 1140 704
rect 1228 696 1236 704
rect 1244 696 1252 704
rect 1308 696 1316 704
rect 1372 696 1380 704
rect 1452 696 1460 704
rect 1660 696 1668 704
rect 1708 696 1716 704
rect 1772 696 1780 704
rect 1852 696 1860 704
rect 1868 696 1876 704
rect 1932 696 1940 704
rect 1996 696 2004 704
rect 2076 696 2084 704
rect 2124 696 2132 704
rect 2380 696 2388 704
rect 2460 696 2468 704
rect 2556 696 2564 704
rect 2620 696 2628 704
rect 12 676 20 684
rect 92 676 100 684
rect 172 676 180 684
rect 204 676 212 684
rect 236 676 244 684
rect 284 676 292 684
rect 396 676 404 684
rect 540 676 548 684
rect 604 676 612 684
rect 636 676 644 684
rect 732 676 740 684
rect 876 676 884 684
rect 1212 676 1220 684
rect 1260 676 1268 684
rect 1388 676 1396 684
rect 1436 676 1444 684
rect 1532 676 1540 684
rect 1548 676 1556 684
rect 1612 676 1620 684
rect 1724 676 1732 684
rect 1852 676 1860 684
rect 1916 676 1924 684
rect 252 656 260 664
rect 348 656 356 664
rect 364 656 372 664
rect 540 656 548 664
rect 700 656 708 664
rect 956 656 964 664
rect 1004 656 1012 664
rect 1116 656 1124 664
rect 1180 656 1188 664
rect 1292 656 1300 664
rect 1340 656 1348 664
rect 1356 656 1364 664
rect 1420 656 1428 664
rect 1804 656 1812 664
rect 1820 656 1828 664
rect 1916 656 1924 664
rect 1980 676 1988 684
rect 2220 676 2228 684
rect 2332 676 2340 684
rect 2492 676 2500 684
rect 2652 676 2660 684
rect 2668 676 2676 684
rect 2684 680 2692 688
rect 2748 696 2756 704
rect 2812 696 2820 704
rect 2828 696 2836 704
rect 2876 696 2884 704
rect 2940 696 2948 704
rect 2860 676 2868 684
rect 2892 676 2900 684
rect 2124 656 2132 664
rect 2380 656 2388 664
rect 2412 656 2420 664
rect 2476 656 2484 664
rect 2796 656 2804 664
rect 2988 676 2996 684
rect 2940 656 2948 664
rect 3004 656 3012 664
rect 44 636 52 644
rect 76 636 84 644
rect 156 636 164 644
rect 380 636 388 644
rect 508 636 516 644
rect 684 636 692 644
rect 828 636 836 644
rect 972 636 980 644
rect 1196 636 1204 644
rect 1404 636 1412 644
rect 1484 636 1492 644
rect 2076 636 2084 644
rect 2428 636 2436 644
rect 2588 636 2596 644
rect 2780 636 2788 644
rect 2972 636 2980 644
rect 3036 636 3044 644
rect 2243 606 2251 614
rect 2253 606 2261 614
rect 2263 606 2271 614
rect 2273 606 2281 614
rect 2283 606 2291 614
rect 2293 606 2301 614
rect 188 576 196 584
rect 588 576 596 584
rect 1164 576 1172 584
rect 1500 576 1508 584
rect 1708 576 1716 584
rect 1756 576 1764 584
rect 1852 576 1860 584
rect 1964 576 1972 584
rect 2140 576 2148 584
rect 2220 576 2228 584
rect 2572 576 2580 584
rect 2636 576 2644 584
rect 2700 576 2708 584
rect 2812 576 2820 584
rect 3020 576 3028 584
rect 12 556 20 564
rect 92 556 100 564
rect 156 556 164 564
rect 364 556 372 564
rect 572 556 580 564
rect 988 556 996 564
rect 1100 556 1108 564
rect 1148 556 1156 564
rect 1196 556 1204 564
rect 1260 556 1268 564
rect 1468 556 1476 564
rect 1484 556 1492 564
rect 1628 556 1636 564
rect 1644 556 1652 564
rect 1740 556 1748 564
rect 1868 556 1876 564
rect 1948 556 1956 564
rect 2044 556 2052 564
rect 2124 556 2132 564
rect 2492 556 2500 564
rect 2556 556 2564 564
rect 2652 556 2660 564
rect 2716 556 2724 564
rect 2796 556 2804 564
rect 204 536 212 544
rect 236 536 244 544
rect 268 536 276 544
rect 284 536 292 544
rect 348 536 356 544
rect 412 536 420 544
rect 476 536 484 544
rect 492 536 500 544
rect 556 536 564 544
rect 604 536 612 544
rect 940 536 948 544
rect 1020 536 1028 544
rect 1084 536 1092 544
rect 1228 536 1236 544
rect 1292 536 1300 544
rect 1324 536 1332 544
rect 1404 536 1412 544
rect 1532 536 1540 544
rect 1580 536 1588 544
rect 1724 536 1732 544
rect 1772 536 1780 544
rect 1804 536 1812 544
rect 1900 536 1908 544
rect 2012 536 2020 544
rect 2060 536 2068 544
rect 2172 536 2180 544
rect 2252 536 2260 544
rect 2316 536 2324 544
rect 2348 536 2356 544
rect 2412 536 2420 544
rect 2444 536 2452 544
rect 2476 536 2484 544
rect 2524 536 2532 544
rect 2620 536 2628 544
rect 2684 536 2692 544
rect 2972 536 2980 544
rect 92 516 100 524
rect 252 516 260 524
rect 300 516 308 524
rect 332 516 340 524
rect 412 516 420 524
rect 460 516 468 524
rect 508 516 516 524
rect 540 516 548 524
rect 620 516 628 524
rect 652 516 660 524
rect 716 516 724 524
rect 844 516 852 524
rect 892 516 900 524
rect 1004 516 1012 524
rect 1020 516 1028 524
rect 1068 516 1076 524
rect 1132 516 1140 524
rect 1180 516 1188 524
rect 1244 516 1252 524
rect 1308 516 1316 524
rect 1340 516 1348 524
rect 1372 516 1380 524
rect 1388 516 1396 524
rect 1436 516 1444 524
rect 1580 516 1588 524
rect 1676 516 1684 524
rect 1788 516 1796 524
rect 1820 516 1828 524
rect 2044 516 2052 524
rect 2076 516 2084 524
rect 2108 516 2116 524
rect 2988 532 2996 540
rect 2188 516 2196 524
rect 2220 516 2228 524
rect 2364 516 2372 524
rect 172 496 180 504
rect 204 496 212 504
rect 428 496 436 504
rect 668 496 676 504
rect 732 496 740 504
rect 12 476 20 484
rect 700 476 708 484
rect 828 476 836 484
rect 876 496 884 504
rect 972 496 980 504
rect 1036 496 1044 504
rect 1340 496 1348 504
rect 1452 496 1460 504
rect 1500 496 1508 504
rect 1596 496 1604 504
rect 1644 496 1652 504
rect 1852 496 1860 504
rect 1868 496 1876 504
rect 1964 496 1972 504
rect 2428 516 2436 524
rect 2460 516 2468 524
rect 2540 516 2548 524
rect 2668 516 2676 524
rect 2748 516 2756 524
rect 2828 516 2836 524
rect 2876 516 2884 524
rect 2924 516 2932 524
rect 2732 496 2740 504
rect 2892 496 2900 504
rect 2908 496 2916 504
rect 332 456 340 464
rect 716 456 724 464
rect 908 476 916 484
rect 940 476 948 484
rect 1564 476 1572 484
rect 2492 476 2500 484
rect 2764 476 2772 484
rect 2860 476 2868 484
rect 2940 476 2948 484
rect 2364 456 2372 464
rect 140 436 148 444
rect 364 436 372 444
rect 460 436 468 444
rect 540 436 548 444
rect 572 436 580 444
rect 844 436 852 444
rect 1116 436 1124 444
rect 1196 436 1204 444
rect 1260 436 1268 444
rect 1612 436 1620 444
rect 2332 436 2340 444
rect 2748 436 2756 444
rect 2828 436 2836 444
rect 2844 436 2852 444
rect 2924 436 2932 444
rect 739 406 747 414
rect 749 406 757 414
rect 759 406 767 414
rect 769 406 777 414
rect 779 406 787 414
rect 789 406 797 414
rect 108 376 116 384
rect 348 376 356 384
rect 716 376 724 384
rect 876 376 884 384
rect 1132 376 1140 384
rect 1212 376 1220 384
rect 1564 376 1572 384
rect 1644 376 1652 384
rect 1692 376 1700 384
rect 1756 376 1764 384
rect 1836 376 1844 384
rect 1980 376 1988 384
rect 2572 376 2580 384
rect 988 356 996 364
rect 252 336 260 344
rect 972 336 980 344
rect 2556 336 2564 344
rect 2876 336 2884 344
rect 2940 336 2948 344
rect 124 316 132 324
rect 188 316 196 324
rect 684 316 692 324
rect 844 316 852 324
rect 1004 316 1012 324
rect 1100 316 1108 324
rect 1244 316 1252 324
rect 1372 316 1380 324
rect 1436 316 1444 324
rect 1804 316 1812 324
rect 1868 316 1876 324
rect 1916 316 1924 324
rect 2172 316 2180 324
rect 2236 316 2244 324
rect 2588 316 2596 324
rect 2604 316 2612 324
rect 2844 316 2852 324
rect 2908 316 2916 324
rect 28 296 36 304
rect 60 296 68 304
rect 156 296 164 304
rect 236 296 244 304
rect 268 296 276 304
rect 316 296 324 304
rect 348 296 356 304
rect 380 296 388 304
rect 476 296 484 304
rect 508 296 516 304
rect 668 296 676 304
rect 716 296 724 304
rect 828 296 836 304
rect 876 296 884 304
rect 908 296 916 304
rect 940 296 948 304
rect 988 296 996 304
rect 1020 296 1028 304
rect 1052 296 1060 304
rect 1084 296 1092 304
rect 1132 296 1140 304
rect 1180 296 1188 304
rect 1228 296 1236 304
rect 1276 296 1284 304
rect 1308 296 1316 304
rect 1468 296 1476 304
rect 1500 296 1508 304
rect 1532 296 1540 304
rect 1564 296 1572 304
rect 1596 296 1604 304
rect 1628 296 1636 304
rect 1660 296 1668 304
rect 1740 296 1748 304
rect 1772 296 1780 304
rect 1852 296 1860 304
rect 1996 296 2004 304
rect 2060 296 2068 304
rect 2124 296 2132 304
rect 2140 296 2148 304
rect 2188 296 2196 304
rect 2204 296 2212 304
rect 2348 296 2356 304
rect 2412 296 2420 304
rect 2476 296 2484 304
rect 2524 296 2532 304
rect 2572 296 2580 304
rect 2604 296 2612 304
rect 2700 296 2708 304
rect 2780 296 2788 304
rect 2860 296 2868 304
rect 2924 296 2932 304
rect 12 276 20 284
rect 76 276 84 284
rect 92 276 100 284
rect 140 276 148 284
rect 236 276 244 284
rect 412 276 420 284
rect 492 276 500 284
rect 732 276 740 284
rect 892 276 900 284
rect 1036 276 1044 284
rect 1068 276 1076 284
rect 1148 276 1156 284
rect 1164 276 1172 284
rect 1228 276 1236 284
rect 1292 276 1300 284
rect 1324 276 1332 284
rect 1356 276 1364 284
rect 1420 276 1428 284
rect 1500 276 1508 284
rect 1628 276 1636 284
rect 1724 276 1732 284
rect 1788 276 1796 284
rect 1852 276 1860 284
rect 1868 276 1876 284
rect 1916 276 1924 284
rect 2044 276 2052 284
rect 2108 276 2116 284
rect 2124 276 2132 284
rect 2188 276 2196 284
rect 2380 276 2388 284
rect 2396 276 2404 284
rect 2492 276 2500 284
rect 2636 276 2644 284
rect 2684 276 2692 284
rect 2812 276 2820 284
rect 3036 276 3044 284
rect 204 256 212 264
rect 316 256 324 264
rect 444 256 452 264
rect 460 256 468 264
rect 540 256 548 264
rect 620 256 628 264
rect 812 256 820 264
rect 940 256 948 264
rect 1340 256 1348 264
rect 1356 256 1364 264
rect 1516 256 1524 264
rect 1532 256 1540 264
rect 1660 256 1668 264
rect 1708 256 1716 264
rect 1916 256 1924 264
rect 1964 256 1972 264
rect 2028 256 2036 264
rect 2236 256 2244 264
rect 2252 256 2260 264
rect 2316 256 2324 264
rect 2364 256 2372 264
rect 2428 256 2436 264
rect 2524 256 2532 264
rect 2652 256 2660 264
rect 2812 256 2820 264
rect 28 236 36 244
rect 188 236 196 244
rect 524 236 532 244
rect 556 236 564 244
rect 636 236 644 244
rect 1244 236 1252 244
rect 2060 236 2068 244
rect 2332 236 2340 244
rect 2444 236 2452 244
rect 2668 236 2676 244
rect 2796 236 2804 244
rect 2860 236 2868 244
rect 2924 236 2932 244
rect 2243 206 2251 214
rect 2253 206 2261 214
rect 2263 206 2271 214
rect 2273 206 2281 214
rect 2283 206 2291 214
rect 2293 206 2301 214
rect 60 176 68 184
rect 124 176 132 184
rect 268 176 276 184
rect 396 176 404 184
rect 444 176 452 184
rect 508 176 516 184
rect 716 176 724 184
rect 812 176 820 184
rect 1052 176 1060 184
rect 1084 176 1092 184
rect 1180 176 1188 184
rect 1260 176 1268 184
rect 1372 176 1380 184
rect 1420 176 1428 184
rect 1484 176 1492 184
rect 1548 176 1556 184
rect 1628 176 1636 184
rect 1868 176 1876 184
rect 1996 176 2004 184
rect 2092 176 2100 184
rect 2188 176 2196 184
rect 2220 176 2228 184
rect 2412 176 2420 184
rect 2524 176 2532 184
rect 2748 176 2756 184
rect 2956 176 2964 184
rect 28 156 36 164
rect 156 156 164 164
rect 188 156 196 164
rect 332 156 340 164
rect 492 156 500 164
rect 620 156 628 164
rect 732 156 740 164
rect 956 156 964 164
rect 1004 156 1012 164
rect 1164 156 1172 164
rect 1356 156 1364 164
rect 1436 156 1444 164
rect 1468 156 1476 164
rect 12 136 20 144
rect 44 136 52 144
rect 92 136 100 144
rect 204 136 212 144
rect 220 136 228 144
rect 284 136 292 144
rect 348 136 356 144
rect 428 136 436 144
rect 460 136 468 144
rect 524 136 532 144
rect 540 136 548 144
rect 700 136 708 144
rect 860 136 868 144
rect 908 136 916 144
rect 924 136 932 144
rect 1020 136 1028 144
rect 1100 136 1108 144
rect 1292 136 1300 144
rect 1404 136 1412 144
rect 1516 136 1524 144
rect 1740 156 1748 164
rect 1964 156 1972 164
rect 2060 156 2068 164
rect 2076 156 2084 164
rect 1820 136 1828 144
rect 1932 136 1940 144
rect 2012 136 2020 144
rect 2060 136 2068 144
rect 2364 156 2372 164
rect 2588 156 2596 164
rect 2652 156 2660 164
rect 2156 136 2164 144
rect 2348 136 2356 144
rect 2476 136 2484 144
rect 2492 136 2500 144
rect 2572 136 2580 144
rect 2620 136 2628 144
rect 2732 136 2740 144
rect 2780 156 2788 164
rect 2892 156 2900 164
rect 2972 156 2980 164
rect 172 116 180 124
rect 236 116 244 124
rect 300 116 308 124
rect 364 116 372 124
rect 412 116 420 124
rect 476 116 484 124
rect 540 116 548 124
rect 620 116 628 124
rect 684 116 692 124
rect 844 116 852 124
rect 924 116 932 124
rect 1148 116 1156 124
rect 1196 116 1204 124
rect 1212 116 1220 124
rect 1228 116 1236 124
rect 1324 116 1332 124
rect 1532 116 1540 124
rect 1580 116 1588 124
rect 1596 116 1604 124
rect 1644 116 1652 124
rect 1692 116 1700 124
rect 1772 116 1780 124
rect 1804 116 1812 124
rect 1820 116 1828 124
rect 76 96 84 104
rect 156 96 164 104
rect 268 96 276 104
rect 348 96 356 104
rect 556 96 564 104
rect 636 96 644 104
rect 812 96 820 104
rect 876 96 884 104
rect 892 96 900 104
rect 972 96 980 104
rect 1068 96 1076 104
rect 1276 96 1284 104
rect 1372 96 1380 104
rect 1452 96 1460 104
rect 1484 96 1492 104
rect 1916 116 1924 124
rect 2028 116 2036 124
rect 1884 96 1892 104
rect 2188 96 2196 104
rect 2604 116 2612 124
rect 2636 116 2644 124
rect 2812 116 2820 124
rect 2860 116 2868 124
rect 2988 116 2996 124
rect 2540 96 2548 104
rect 1308 76 1316 84
rect 1980 76 1988 84
rect 3036 76 3044 84
rect 1116 36 1124 44
rect 1676 36 1684 44
rect 1724 36 1732 44
rect 2844 36 2852 44
rect 2940 36 2948 44
rect 739 6 747 14
rect 749 6 757 14
rect 759 6 767 14
rect 769 6 777 14
rect 779 6 787 14
rect 789 6 797 14
<< metal2 >>
rect 762 2014 774 2016
rect 747 2006 749 2014
rect 757 2006 759 2014
rect 767 2006 769 2014
rect 777 2006 779 2014
rect 787 2006 789 2014
rect 762 2004 774 2006
rect 829 1984 835 2063
rect 189 1904 195 1936
rect 973 1924 979 2063
rect 333 1904 339 1916
rect 509 1904 515 1916
rect 45 1884 51 1896
rect 61 1724 67 1896
rect 125 1864 131 1896
rect 93 1764 99 1856
rect 157 1764 163 1836
rect 13 1684 19 1696
rect 45 1644 51 1716
rect 109 1504 115 1516
rect 173 1504 179 1716
rect 237 1704 243 1776
rect 253 1764 259 1836
rect 269 1684 275 1716
rect 285 1664 291 1876
rect 301 1584 307 1896
rect 461 1884 467 1896
rect 637 1884 643 1916
rect 333 1844 339 1876
rect 365 1864 371 1876
rect 605 1864 611 1876
rect 317 1724 323 1756
rect 333 1704 339 1836
rect 381 1744 387 1776
rect 365 1724 371 1736
rect 429 1723 435 1836
rect 445 1744 451 1856
rect 420 1717 435 1723
rect 493 1704 499 1716
rect 509 1704 515 1796
rect 541 1723 547 1836
rect 557 1784 563 1856
rect 573 1744 579 1756
rect 589 1744 595 1836
rect 637 1784 643 1796
rect 589 1724 595 1736
rect 541 1717 556 1723
rect 605 1704 611 1716
rect 653 1704 659 1836
rect 669 1803 675 1876
rect 685 1844 691 1896
rect 701 1884 707 1896
rect 893 1864 899 1876
rect 813 1804 819 1856
rect 669 1797 684 1803
rect 685 1744 691 1796
rect 445 1684 451 1696
rect 477 1684 483 1696
rect 29 1364 35 1496
rect 61 1384 67 1436
rect 77 1364 83 1476
rect 125 1464 131 1476
rect 45 1304 51 1316
rect 61 1224 67 1236
rect 45 1104 51 1116
rect 13 1064 19 1076
rect 61 984 67 1136
rect 77 1104 83 1116
rect 61 964 67 976
rect 93 924 99 1416
rect 109 1344 115 1436
rect 173 1424 179 1496
rect 205 1384 211 1456
rect 221 1444 227 1456
rect 301 1444 307 1516
rect 317 1504 323 1676
rect 317 1423 323 1496
rect 301 1417 323 1423
rect 125 1084 131 1276
rect 141 1104 147 1356
rect 173 1304 179 1316
rect 205 1304 211 1336
rect 221 1324 227 1336
rect 253 1304 259 1316
rect 189 1084 195 1116
rect 109 924 115 1036
rect 13 884 19 896
rect 45 844 51 916
rect 93 724 99 916
rect 157 884 163 936
rect 205 924 211 936
rect 221 924 227 1136
rect 285 1084 291 1336
rect 301 1144 307 1417
rect 333 1384 339 1456
rect 317 1344 323 1356
rect 333 1344 339 1356
rect 349 1324 355 1576
rect 365 1484 371 1636
rect 397 1584 403 1636
rect 397 1544 403 1576
rect 413 1564 419 1636
rect 413 1524 419 1536
rect 445 1524 451 1596
rect 525 1564 531 1696
rect 637 1684 643 1696
rect 429 1504 435 1516
rect 509 1504 515 1556
rect 557 1524 563 1556
rect 573 1524 579 1596
rect 381 1464 387 1496
rect 461 1464 467 1476
rect 493 1444 499 1496
rect 525 1484 531 1496
rect 557 1484 563 1496
rect 477 1404 483 1436
rect 317 1144 323 1316
rect 365 1124 371 1156
rect 333 1084 339 1096
rect 397 1084 403 1376
rect 285 964 291 1076
rect 413 1063 419 1336
rect 477 1324 483 1396
rect 589 1384 595 1476
rect 605 1464 611 1496
rect 637 1484 643 1516
rect 653 1504 659 1616
rect 669 1504 675 1536
rect 621 1444 627 1476
rect 493 1344 499 1376
rect 573 1324 579 1376
rect 605 1364 611 1396
rect 621 1344 627 1356
rect 653 1344 659 1496
rect 669 1484 675 1496
rect 669 1324 675 1476
rect 701 1384 707 1516
rect 429 1064 435 1316
rect 461 1064 467 1116
rect 509 1104 515 1296
rect 525 1124 531 1176
rect 541 1104 547 1156
rect 397 1057 419 1063
rect 189 704 195 716
rect 221 704 227 916
rect 301 723 307 1056
rect 317 964 323 1036
rect 317 924 323 936
rect 333 924 339 1016
rect 381 984 387 996
rect 397 984 403 1057
rect 365 964 371 976
rect 413 943 419 1036
rect 429 1024 435 1056
rect 413 937 435 943
rect 381 884 387 896
rect 429 864 435 937
rect 477 924 483 956
rect 509 944 515 956
rect 493 924 499 936
rect 461 903 467 916
rect 557 904 563 1076
rect 573 964 579 1316
rect 589 1063 595 1236
rect 605 1224 611 1276
rect 605 1124 611 1216
rect 621 1164 627 1236
rect 685 1204 691 1236
rect 701 1143 707 1376
rect 717 1364 723 1656
rect 813 1624 819 1676
rect 762 1614 774 1616
rect 747 1606 749 1614
rect 757 1606 759 1614
rect 767 1606 769 1614
rect 777 1606 779 1614
rect 787 1606 789 1614
rect 762 1604 774 1606
rect 733 1484 739 1516
rect 749 1364 755 1576
rect 765 1504 771 1536
rect 813 1444 819 1516
rect 717 1344 723 1356
rect 813 1284 819 1356
rect 829 1344 835 1736
rect 861 1504 867 1856
rect 925 1844 931 1876
rect 893 1823 899 1836
rect 877 1817 899 1823
rect 877 1704 883 1817
rect 893 1764 899 1796
rect 925 1724 931 1836
rect 941 1744 947 1856
rect 973 1803 979 1916
rect 1005 1884 1011 2063
rect 1069 1924 1075 2063
rect 1005 1864 1011 1876
rect 1069 1864 1075 1916
rect 1101 1884 1107 2063
rect 1213 2043 1219 2063
rect 1197 2037 1219 2043
rect 964 1797 979 1803
rect 957 1724 963 1796
rect 989 1744 995 1836
rect 1021 1744 1027 1836
rect 893 1544 899 1716
rect 973 1697 988 1703
rect 925 1604 931 1636
rect 941 1584 947 1616
rect 957 1604 963 1636
rect 845 1344 851 1436
rect 877 1424 883 1476
rect 925 1464 931 1496
rect 973 1483 979 1697
rect 1021 1664 1027 1736
rect 1069 1724 1075 1856
rect 1101 1764 1107 1876
rect 1101 1704 1107 1716
rect 1037 1664 1043 1676
rect 989 1504 995 1516
rect 973 1477 995 1483
rect 909 1324 915 1436
rect 957 1424 963 1476
rect 957 1384 963 1416
rect 762 1214 774 1216
rect 747 1206 749 1214
rect 757 1206 759 1214
rect 767 1206 769 1214
rect 777 1206 779 1214
rect 787 1206 789 1214
rect 762 1204 774 1206
rect 685 1137 707 1143
rect 653 1104 659 1116
rect 637 1083 643 1096
rect 637 1077 652 1083
rect 589 1057 611 1063
rect 589 1024 595 1036
rect 605 944 611 1057
rect 621 1044 627 1076
rect 605 924 611 936
rect 621 924 627 936
rect 461 897 524 903
rect 541 897 556 903
rect 461 724 467 736
rect 285 717 307 723
rect 269 704 275 716
rect 13 564 19 676
rect 45 544 51 636
rect 61 564 67 696
rect 285 684 291 717
rect 93 584 99 676
rect 157 644 163 656
rect 173 644 179 676
rect 173 604 179 636
rect 157 564 163 576
rect 13 284 19 476
rect 61 324 67 556
rect 205 544 211 616
rect 237 584 243 676
rect 253 664 259 676
rect 301 664 307 696
rect 237 544 243 556
rect 269 544 275 616
rect 317 544 323 716
rect 413 704 419 716
rect 333 657 348 663
rect 333 604 339 657
rect 365 643 371 656
rect 349 637 371 643
rect 349 544 355 637
rect 253 524 259 536
rect 173 504 179 516
rect 29 304 35 316
rect 93 284 99 476
rect 109 384 115 496
rect 205 484 211 496
rect 141 444 147 456
rect 141 324 147 436
rect 253 344 259 516
rect 349 504 355 536
rect 365 463 371 556
rect 381 504 387 636
rect 397 624 403 676
rect 413 544 419 676
rect 429 624 435 716
rect 445 664 451 696
rect 461 684 467 716
rect 509 624 515 636
rect 445 537 476 543
rect 340 457 371 463
rect 349 384 355 396
rect 29 184 35 236
rect 45 144 51 256
rect 61 184 67 236
rect 77 104 83 276
rect 93 244 99 276
rect 125 184 131 316
rect 141 284 147 296
rect 157 284 163 296
rect 253 284 259 336
rect 381 304 387 416
rect 413 304 419 516
rect 445 504 451 537
rect 493 524 499 536
rect 461 504 467 516
rect 429 444 435 496
rect 381 284 387 296
rect 141 164 147 276
rect 157 164 163 276
rect 237 264 243 276
rect 317 264 323 276
rect 189 204 195 236
rect 93 144 99 156
rect 141 103 147 156
rect 157 144 163 156
rect 221 144 227 256
rect 269 184 275 216
rect 285 144 291 256
rect 429 243 435 376
rect 461 264 467 436
rect 509 424 515 516
rect 525 324 531 696
rect 541 684 547 897
rect 653 884 659 936
rect 685 924 691 1137
rect 701 1104 707 1116
rect 733 1104 739 1116
rect 717 1044 723 1076
rect 829 1064 835 1316
rect 845 1144 851 1196
rect 861 1104 867 1316
rect 877 1304 883 1316
rect 877 1084 883 1256
rect 893 1104 899 1116
rect 909 1084 915 1176
rect 941 1084 947 1356
rect 973 1344 979 1356
rect 957 1104 963 1296
rect 989 1284 995 1477
rect 1037 1483 1043 1636
rect 1021 1477 1043 1483
rect 1005 1264 1011 1476
rect 1021 1444 1027 1477
rect 1053 1463 1059 1636
rect 1069 1504 1075 1556
rect 1085 1524 1091 1696
rect 1117 1564 1123 1836
rect 1165 1824 1171 1836
rect 1181 1803 1187 1876
rect 1197 1864 1203 2037
rect 1261 1884 1267 2063
rect 1373 2057 1395 2063
rect 1389 1984 1395 2057
rect 1437 2057 1459 2063
rect 1437 1984 1443 2057
rect 1165 1797 1187 1803
rect 1165 1704 1171 1797
rect 1197 1784 1203 1856
rect 1245 1804 1251 1836
rect 1245 1764 1251 1776
rect 1277 1724 1283 1896
rect 1517 1864 1523 1896
rect 1428 1857 1443 1863
rect 1325 1763 1331 1836
rect 1325 1757 1340 1763
rect 1229 1664 1235 1676
rect 1101 1504 1107 1536
rect 1117 1524 1123 1536
rect 1149 1524 1155 1596
rect 1117 1484 1123 1516
rect 1165 1504 1171 1596
rect 1044 1457 1059 1463
rect 1053 1323 1059 1436
rect 1069 1324 1075 1416
rect 1085 1344 1091 1396
rect 1117 1344 1123 1436
rect 1133 1324 1139 1456
rect 1037 1317 1059 1323
rect 1021 1304 1027 1316
rect 973 1104 979 1196
rect 1005 1103 1011 1256
rect 1037 1184 1043 1317
rect 1149 1304 1155 1476
rect 1181 1464 1187 1496
rect 1197 1484 1203 1536
rect 1213 1504 1219 1636
rect 1261 1504 1267 1676
rect 1277 1664 1283 1716
rect 1325 1704 1331 1757
rect 1277 1483 1283 1496
rect 1309 1483 1315 1636
rect 1373 1624 1379 1636
rect 1261 1477 1283 1483
rect 1293 1477 1315 1483
rect 1213 1464 1219 1476
rect 1229 1364 1235 1436
rect 1245 1404 1251 1476
rect 1261 1384 1267 1477
rect 1293 1384 1299 1477
rect 1325 1464 1331 1556
rect 1373 1504 1379 1536
rect 1373 1484 1379 1496
rect 1357 1464 1363 1476
rect 1389 1464 1395 1776
rect 1405 1544 1411 1736
rect 1421 1724 1427 1756
rect 1437 1744 1443 1857
rect 1501 1804 1507 1856
rect 1421 1544 1427 1716
rect 1437 1524 1443 1636
rect 1453 1584 1459 1796
rect 1501 1744 1507 1756
rect 1517 1723 1523 1856
rect 1549 1764 1555 2063
rect 1581 1764 1587 1856
rect 1613 1764 1619 1856
rect 1661 1844 1667 1896
rect 1693 1884 1699 1916
rect 1709 1904 1715 2063
rect 1629 1783 1635 1836
rect 1629 1777 1651 1783
rect 1508 1717 1523 1723
rect 1565 1704 1571 1756
rect 1405 1504 1411 1516
rect 1453 1504 1459 1576
rect 1517 1564 1523 1636
rect 1453 1464 1459 1476
rect 1517 1464 1523 1536
rect 1380 1457 1388 1463
rect 1325 1364 1331 1416
rect 1197 1357 1212 1363
rect 989 1097 1011 1103
rect 989 1084 995 1097
rect 1053 1084 1059 1296
rect 1028 1057 1043 1063
rect 797 964 803 996
rect 669 764 675 836
rect 605 724 611 736
rect 541 524 547 636
rect 557 544 563 596
rect 589 584 595 696
rect 605 684 611 716
rect 637 684 643 696
rect 701 644 707 656
rect 573 464 579 556
rect 605 544 611 576
rect 621 524 627 536
rect 637 524 643 596
rect 669 504 675 536
rect 685 483 691 636
rect 717 543 723 916
rect 762 814 774 816
rect 747 806 749 814
rect 757 806 759 814
rect 767 806 769 814
rect 777 806 779 814
rect 787 806 789 814
rect 762 804 774 806
rect 829 743 835 1036
rect 909 964 915 1056
rect 845 924 851 936
rect 893 904 899 936
rect 909 923 915 956
rect 941 924 947 1036
rect 909 917 924 923
rect 957 904 963 916
rect 973 904 979 956
rect 1037 944 1043 1057
rect 1037 924 1043 936
rect 925 784 931 816
rect 813 737 835 743
rect 733 684 739 716
rect 813 704 819 737
rect 909 724 915 736
rect 829 704 835 716
rect 829 644 835 676
rect 717 537 739 543
rect 733 504 739 537
rect 685 477 700 483
rect 541 324 547 436
rect 493 284 499 316
rect 509 284 515 296
rect 541 264 547 316
rect 573 264 579 436
rect 717 384 723 436
rect 762 414 774 416
rect 747 406 749 414
rect 757 406 759 414
rect 767 406 769 414
rect 777 406 779 414
rect 787 406 789 414
rect 762 404 774 406
rect 669 304 675 356
rect 621 284 627 296
rect 621 264 627 276
rect 685 244 691 316
rect 429 237 451 243
rect 349 144 355 196
rect 397 184 403 196
rect 445 184 451 237
rect 509 184 515 216
rect 525 184 531 236
rect 429 144 435 176
rect 349 104 355 136
rect 365 124 371 136
rect 413 124 419 136
rect 477 124 483 176
rect 525 144 531 156
rect 557 123 563 236
rect 621 144 627 156
rect 557 117 579 123
rect 141 97 156 103
rect 573 -23 579 117
rect 637 123 643 236
rect 717 184 723 296
rect 733 284 739 316
rect 813 264 819 636
rect 829 524 835 636
rect 861 604 867 696
rect 877 664 883 676
rect 845 524 851 596
rect 925 504 931 696
rect 941 584 947 716
rect 973 684 979 896
rect 989 884 995 896
rect 1037 824 1043 916
rect 1053 904 1059 936
rect 1069 924 1075 1176
rect 1149 1104 1155 1236
rect 1165 1124 1171 1276
rect 1085 1024 1091 1056
rect 1101 1004 1107 1056
rect 1117 984 1123 1036
rect 1133 1004 1139 1076
rect 1165 1004 1171 1116
rect 1181 1104 1187 1256
rect 1197 1224 1203 1357
rect 1229 1323 1235 1336
rect 1229 1317 1244 1323
rect 1197 1104 1203 1156
rect 1213 1104 1219 1316
rect 1261 1244 1267 1336
rect 1341 1324 1347 1436
rect 1357 1424 1363 1456
rect 1389 1324 1395 1356
rect 1309 1304 1315 1316
rect 1325 1304 1331 1316
rect 1437 1304 1443 1436
rect 1453 1324 1459 1336
rect 1485 1284 1491 1436
rect 1501 1364 1507 1456
rect 1533 1444 1539 1676
rect 1581 1604 1587 1736
rect 1645 1724 1651 1777
rect 1629 1684 1635 1696
rect 1661 1664 1667 1736
rect 1677 1684 1683 1876
rect 1709 1864 1715 1876
rect 1709 1724 1715 1776
rect 1549 1484 1555 1496
rect 1565 1464 1571 1476
rect 1533 1324 1539 1436
rect 1581 1384 1587 1596
rect 1597 1524 1603 1656
rect 1597 1484 1603 1516
rect 1613 1424 1619 1516
rect 1661 1484 1667 1636
rect 1677 1484 1683 1576
rect 1645 1457 1660 1463
rect 1645 1444 1651 1457
rect 1629 1404 1635 1436
rect 1661 1404 1667 1436
rect 1693 1424 1699 1656
rect 1709 1463 1715 1556
rect 1725 1544 1731 1736
rect 1741 1724 1747 1756
rect 1773 1704 1779 1876
rect 1789 1864 1795 1916
rect 1805 1864 1811 2063
rect 1885 2057 1907 2063
rect 1901 1884 1907 2057
rect 1997 1884 2003 1916
rect 1869 1864 1875 1876
rect 1917 1864 1923 1876
rect 1933 1844 1939 1880
rect 1853 1784 1859 1816
rect 1965 1804 1971 1836
rect 1821 1744 1827 1776
rect 1901 1764 1907 1796
rect 1789 1704 1795 1736
rect 1773 1644 1779 1696
rect 1837 1624 1843 1756
rect 1869 1724 1875 1756
rect 1757 1504 1763 1516
rect 1837 1484 1843 1556
rect 1709 1457 1724 1463
rect 1412 1277 1459 1283
rect 1453 1264 1459 1277
rect 1197 964 1203 1096
rect 1213 1024 1219 1076
rect 1053 784 1059 816
rect 1037 704 1043 736
rect 941 544 947 576
rect 829 464 835 476
rect 845 364 851 436
rect 861 384 867 496
rect 916 477 940 483
rect 877 384 883 456
rect 813 184 819 256
rect 845 204 851 316
rect 877 304 883 336
rect 893 324 899 436
rect 957 404 963 656
rect 973 504 979 636
rect 989 604 995 696
rect 989 564 995 576
rect 1021 484 1027 516
rect 893 284 899 316
rect 909 304 915 356
rect 973 284 979 336
rect 989 324 995 356
rect 1005 324 1011 356
rect 1037 344 1043 496
rect 1053 304 1059 716
rect 1085 664 1091 876
rect 1069 524 1075 576
rect 1101 564 1107 836
rect 1117 824 1123 956
rect 1229 944 1235 1216
rect 1149 917 1164 923
rect 1149 784 1155 917
rect 1117 564 1123 656
rect 1165 584 1171 816
rect 1181 764 1187 896
rect 1213 864 1219 936
rect 1229 924 1235 936
rect 1245 924 1251 1096
rect 1261 1064 1267 1236
rect 1357 1124 1363 1236
rect 1389 1123 1395 1236
rect 1469 1224 1475 1276
rect 1421 1144 1427 1156
rect 1373 1117 1395 1123
rect 1309 1064 1315 1076
rect 1325 1064 1331 1096
rect 1373 1064 1379 1117
rect 1396 1097 1436 1103
rect 1245 863 1251 916
rect 1277 904 1283 976
rect 1293 944 1299 1016
rect 1453 984 1459 1056
rect 1469 983 1475 1216
rect 1485 1124 1491 1136
rect 1517 1124 1523 1236
rect 1517 984 1523 1096
rect 1533 1084 1539 1236
rect 1549 1004 1555 1096
rect 1581 1004 1587 1116
rect 1469 977 1491 983
rect 1485 964 1491 977
rect 1309 924 1315 956
rect 1437 944 1443 956
rect 1229 857 1251 863
rect 1213 684 1219 856
rect 1229 783 1235 857
rect 1245 804 1251 836
rect 1229 777 1251 783
rect 1229 704 1235 756
rect 1245 704 1251 777
rect 1277 744 1283 896
rect 1181 624 1187 656
rect 1197 604 1203 636
rect 1245 584 1251 696
rect 1268 677 1283 683
rect 1085 464 1091 536
rect 1133 524 1139 536
rect 1149 444 1155 556
rect 1181 464 1187 516
rect 1117 364 1123 436
rect 1133 384 1139 396
rect 1213 384 1219 556
rect 1229 404 1235 536
rect 1277 484 1283 677
rect 1293 664 1299 896
rect 1309 704 1315 836
rect 1357 724 1363 836
rect 1373 764 1379 876
rect 1389 864 1395 916
rect 1405 863 1411 896
rect 1421 884 1427 916
rect 1469 904 1475 956
rect 1485 944 1491 956
rect 1533 944 1539 956
rect 1597 924 1603 1176
rect 1613 1164 1619 1316
rect 1629 1184 1635 1316
rect 1613 1104 1619 1136
rect 1629 1004 1635 1096
rect 1661 1083 1667 1396
rect 1677 1364 1683 1376
rect 1709 1364 1715 1436
rect 1725 1343 1731 1396
rect 1757 1344 1763 1376
rect 1773 1364 1779 1476
rect 1805 1404 1811 1436
rect 1853 1404 1859 1496
rect 1885 1484 1891 1496
rect 1869 1464 1875 1476
rect 1725 1337 1747 1343
rect 1716 1317 1731 1323
rect 1693 1184 1699 1216
rect 1709 1104 1715 1296
rect 1725 1184 1731 1317
rect 1645 1077 1667 1083
rect 1645 964 1651 1077
rect 1613 944 1619 956
rect 1661 944 1667 1056
rect 1709 1003 1715 1076
rect 1709 997 1731 1003
rect 1517 884 1523 896
rect 1581 884 1587 896
rect 1405 857 1427 863
rect 1373 704 1379 756
rect 1389 704 1395 856
rect 1293 544 1299 576
rect 1309 564 1315 696
rect 1389 684 1395 696
rect 1405 684 1411 736
rect 1357 664 1363 676
rect 1421 664 1427 857
rect 1549 824 1555 836
rect 1629 784 1635 936
rect 1437 684 1443 756
rect 1421 604 1427 656
rect 1549 644 1555 676
rect 1597 644 1603 716
rect 1613 684 1619 776
rect 1645 724 1651 856
rect 1661 784 1667 936
rect 1709 904 1715 916
rect 1725 904 1731 997
rect 1741 923 1747 1337
rect 1757 1124 1763 1336
rect 1837 1324 1843 1356
rect 1789 1224 1795 1316
rect 1853 1304 1859 1356
rect 1869 1324 1875 1336
rect 1885 1264 1891 1276
rect 1853 1144 1859 1156
rect 1805 1117 1820 1123
rect 1789 1084 1795 1096
rect 1789 1044 1795 1076
rect 1741 917 1756 923
rect 1773 904 1779 1016
rect 1805 944 1811 1117
rect 1869 1104 1875 1236
rect 1901 1224 1907 1616
rect 1933 1543 1939 1716
rect 1949 1684 1955 1716
rect 1981 1703 1987 1876
rect 2029 1864 2035 1936
rect 2061 1904 2067 1936
rect 2388 1917 2396 1923
rect 2045 1744 2051 1836
rect 2013 1724 2019 1736
rect 1972 1697 1987 1703
rect 2013 1664 2019 1676
rect 2029 1624 2035 1696
rect 1917 1537 1939 1543
rect 1917 1464 1923 1537
rect 1933 1464 1939 1516
rect 1949 1484 1955 1576
rect 1965 1504 1971 1516
rect 2045 1503 2051 1716
rect 2061 1664 2067 1896
rect 2077 1804 2083 1896
rect 2269 1884 2275 1916
rect 2109 1804 2115 1876
rect 2093 1704 2099 1776
rect 2109 1764 2115 1796
rect 2141 1744 2147 1836
rect 2125 1684 2131 1716
rect 2157 1663 2163 1856
rect 2173 1744 2179 1796
rect 2205 1744 2211 1796
rect 2189 1724 2195 1736
rect 2221 1664 2227 1836
rect 2266 1814 2278 1816
rect 2251 1806 2253 1814
rect 2261 1806 2263 1814
rect 2271 1806 2273 1814
rect 2281 1806 2283 1814
rect 2291 1806 2293 1814
rect 2266 1804 2278 1806
rect 2157 1657 2179 1663
rect 2061 1584 2067 1636
rect 2077 1504 2083 1636
rect 2036 1497 2051 1503
rect 1997 1484 2003 1496
rect 2013 1484 2019 1496
rect 2045 1484 2051 1497
rect 1949 1384 1955 1456
rect 1981 1384 1987 1476
rect 2109 1384 2115 1416
rect 1981 1364 1987 1376
rect 2029 1364 2035 1376
rect 1917 1264 1923 1316
rect 1917 1184 1923 1236
rect 1965 1164 1971 1336
rect 2013 1324 2019 1336
rect 2045 1184 2051 1376
rect 2125 1364 2131 1536
rect 2141 1524 2147 1596
rect 2157 1484 2163 1636
rect 2173 1484 2179 1657
rect 2237 1624 2243 1756
rect 2333 1644 2339 1896
rect 2349 1764 2355 1816
rect 2381 1804 2387 1876
rect 2429 1857 2444 1863
rect 2237 1524 2243 1556
rect 2189 1464 2195 1476
rect 2157 1424 2163 1436
rect 2125 1344 2131 1356
rect 2157 1344 2163 1356
rect 2205 1324 2211 1496
rect 2221 1364 2227 1476
rect 2317 1464 2323 1536
rect 2333 1423 2339 1436
rect 2317 1417 2339 1423
rect 2266 1414 2278 1416
rect 2251 1406 2253 1414
rect 2261 1406 2263 1414
rect 2271 1406 2273 1414
rect 2281 1406 2283 1414
rect 2291 1406 2293 1414
rect 2266 1404 2278 1406
rect 1933 1144 1939 1156
rect 1965 1124 1971 1156
rect 2061 1123 2067 1276
rect 2077 1244 2083 1296
rect 2173 1284 2179 1316
rect 2077 1164 2083 1236
rect 2061 1117 2076 1123
rect 1885 1104 1891 1116
rect 1901 1044 1907 1116
rect 2093 1104 2099 1256
rect 2141 1124 2147 1236
rect 1924 1097 1955 1103
rect 1821 984 1827 1016
rect 1725 724 1731 836
rect 1741 824 1747 876
rect 1789 804 1795 916
rect 1325 544 1331 596
rect 1485 584 1491 636
rect 1501 584 1507 616
rect 1517 577 1555 583
rect 1341 524 1347 556
rect 1405 544 1411 556
rect 1453 543 1459 576
rect 1517 543 1523 577
rect 1549 564 1555 577
rect 1533 544 1539 556
rect 1453 537 1523 543
rect 1588 537 1603 543
rect 1316 517 1331 523
rect 1325 503 1331 517
rect 1325 497 1340 503
rect 1261 323 1267 436
rect 1252 317 1267 323
rect 1021 284 1027 296
rect 1085 284 1091 296
rect 1037 264 1043 276
rect 941 244 947 256
rect 1053 184 1059 276
rect 813 164 819 176
rect 733 144 739 156
rect 861 144 867 176
rect 637 117 659 123
rect 621 104 627 116
rect 637 84 643 96
rect 653 -23 659 117
rect 685 84 691 116
rect 701 104 707 136
rect 845 124 851 136
rect 877 104 883 156
rect 909 124 915 136
rect 957 124 963 156
rect 925 104 931 116
rect 973 104 979 156
rect 1069 144 1075 276
rect 1101 263 1107 316
rect 1277 304 1283 336
rect 1309 304 1315 316
rect 1092 257 1107 263
rect 1085 184 1091 256
rect 1133 224 1139 296
rect 1357 284 1363 336
rect 1373 324 1379 376
rect 1389 284 1395 516
rect 1405 283 1411 536
rect 1428 517 1436 523
rect 1533 484 1539 536
rect 1597 524 1603 537
rect 1565 484 1571 516
rect 1581 504 1587 516
rect 1597 484 1603 496
rect 1501 304 1507 316
rect 1533 304 1539 476
rect 1613 464 1619 676
rect 1709 664 1715 696
rect 1629 564 1635 656
rect 1709 584 1715 596
rect 1757 584 1763 636
rect 1773 604 1779 696
rect 1677 524 1683 576
rect 1805 564 1811 656
rect 1821 644 1827 656
rect 1748 557 1763 563
rect 1693 504 1699 536
rect 1565 384 1571 456
rect 1565 304 1571 316
rect 1405 277 1420 283
rect 1165 264 1171 276
rect 1229 264 1235 276
rect 1293 264 1299 276
rect 1149 204 1155 236
rect 1181 224 1187 256
rect 1101 144 1107 156
rect 1021 124 1027 136
rect 1149 124 1155 196
rect 1181 184 1187 216
rect 1245 204 1251 236
rect 1261 184 1267 236
rect 1213 124 1219 156
rect 1069 104 1075 116
rect 762 14 774 16
rect 747 6 749 14
rect 757 6 759 14
rect 767 6 769 14
rect 777 6 779 14
rect 787 6 789 14
rect 762 4 774 6
rect 1069 -23 1075 96
rect 1117 -17 1123 36
rect 1213 3 1219 116
rect 1277 104 1283 196
rect 1325 184 1331 276
rect 1469 204 1475 296
rect 1421 184 1427 196
rect 1485 184 1491 276
rect 1357 124 1363 156
rect 1405 124 1411 136
rect 1437 124 1443 156
rect 1469 144 1475 156
rect 1501 144 1507 276
rect 1533 224 1539 256
rect 1549 184 1555 256
rect 1565 244 1571 296
rect 1597 264 1603 296
rect 1581 124 1587 136
rect 1613 124 1619 436
rect 1629 304 1635 476
rect 1645 384 1651 496
rect 1693 384 1699 496
rect 1741 344 1747 456
rect 1757 384 1763 557
rect 1773 544 1779 556
rect 1773 464 1779 536
rect 1789 524 1795 536
rect 1805 524 1811 536
rect 1821 524 1827 576
rect 1821 444 1827 496
rect 1837 384 1843 936
rect 1853 924 1859 1036
rect 1901 944 1907 956
rect 1901 903 1907 916
rect 1885 897 1907 903
rect 1853 704 1859 716
rect 1869 684 1875 696
rect 1853 664 1859 676
rect 1869 644 1875 676
rect 1853 584 1859 616
rect 1869 564 1875 576
rect 1853 404 1859 476
rect 1741 304 1747 336
rect 1629 264 1635 276
rect 1661 264 1667 296
rect 1629 184 1635 256
rect 1709 244 1715 256
rect 1789 244 1795 276
rect 1325 104 1331 116
rect 1485 104 1491 116
rect 1213 -3 1235 3
rect 1117 -23 1139 -17
rect 1229 -23 1235 -3
rect 1485 -23 1491 96
rect 1581 3 1587 116
rect 1581 -3 1603 3
rect 1597 -23 1603 -3
rect 1677 -17 1683 36
rect 1725 -17 1731 36
rect 1741 24 1747 156
rect 1805 124 1811 316
rect 1853 304 1859 396
rect 1853 264 1859 276
rect 1885 263 1891 897
rect 1901 584 1907 756
rect 1933 704 1939 816
rect 1949 744 1955 1097
rect 1965 684 1971 1036
rect 1981 784 1987 1096
rect 1997 1084 2003 1096
rect 2157 1084 2163 1156
rect 2205 1104 2211 1236
rect 2253 1104 2259 1156
rect 2013 904 2019 916
rect 1901 524 1907 536
rect 1869 257 1891 263
rect 1869 184 1875 257
rect 1901 164 1907 516
rect 1917 424 1923 636
rect 1965 584 1971 596
rect 1949 544 1955 556
rect 1924 277 1939 283
rect 1933 144 1939 277
rect 1949 144 1955 536
rect 1965 504 1971 516
rect 1981 384 1987 676
rect 1997 664 2003 696
rect 2013 684 2019 896
rect 2029 844 2035 1076
rect 2093 984 2099 1076
rect 2125 1024 2131 1036
rect 2157 984 2163 1056
rect 2173 1004 2179 1036
rect 2189 984 2195 1076
rect 2205 1057 2220 1063
rect 2045 864 2051 916
rect 2093 804 2099 956
rect 2205 904 2211 1057
rect 2221 984 2227 1016
rect 2266 1014 2278 1016
rect 2251 1006 2253 1014
rect 2261 1006 2263 1014
rect 2271 1006 2273 1014
rect 2281 1006 2283 1014
rect 2291 1006 2293 1014
rect 2266 1004 2278 1006
rect 2317 944 2323 1417
rect 2333 1364 2339 1396
rect 2349 1324 2355 1516
rect 2365 1504 2371 1756
rect 2381 1724 2387 1796
rect 2429 1744 2435 1857
rect 2461 1784 2467 1916
rect 2509 1904 2515 1916
rect 2573 1904 2579 2063
rect 2653 2057 2675 2063
rect 2493 1804 2499 1836
rect 2525 1824 2531 1836
rect 2557 1804 2563 1896
rect 2621 1884 2627 1916
rect 2653 1904 2659 2057
rect 2573 1824 2579 1856
rect 2445 1744 2451 1756
rect 2493 1724 2499 1756
rect 2397 1717 2412 1723
rect 2397 1604 2403 1717
rect 2541 1684 2547 1716
rect 2557 1704 2563 1796
rect 2573 1744 2579 1756
rect 2589 1724 2595 1876
rect 2653 1864 2659 1896
rect 2701 1764 2707 1836
rect 2525 1664 2531 1676
rect 2381 1504 2387 1556
rect 2365 1464 2371 1476
rect 2365 1424 2371 1456
rect 2365 1404 2371 1416
rect 2397 1384 2403 1596
rect 2397 1324 2403 1356
rect 2413 1344 2419 1356
rect 2333 1084 2339 1096
rect 2381 1064 2387 1216
rect 2397 1064 2403 1096
rect 2413 1084 2419 1336
rect 2381 1044 2387 1056
rect 2365 1024 2371 1036
rect 2381 944 2387 956
rect 2228 917 2243 923
rect 2093 724 2099 776
rect 2141 744 2147 756
rect 2029 644 2035 716
rect 2077 664 2083 696
rect 1997 384 2003 616
rect 2077 543 2083 636
rect 2093 624 2099 716
rect 2109 604 2115 716
rect 2125 704 2131 716
rect 2173 624 2179 716
rect 2141 584 2147 596
rect 2077 537 2099 543
rect 2093 444 2099 537
rect 2109 524 2115 536
rect 1997 304 2003 316
rect 2045 284 2051 416
rect 2061 304 2067 336
rect 2061 284 2067 296
rect 1965 164 1971 256
rect 2013 144 2019 156
rect 1805 104 1811 116
rect 1661 -23 1683 -17
rect 1709 -23 1731 -17
rect 1773 -23 1779 16
rect 1837 -23 1843 136
rect 1981 84 1987 116
rect 1981 -23 1987 76
rect 2013 -17 2019 136
rect 2029 124 2035 256
rect 2045 184 2051 276
rect 2093 184 2099 376
rect 2125 304 2131 516
rect 2141 504 2147 576
rect 2189 524 2195 556
rect 2205 503 2211 716
rect 2221 704 2227 896
rect 2237 683 2243 917
rect 2253 864 2259 936
rect 2317 924 2323 936
rect 2253 724 2259 856
rect 2269 824 2275 836
rect 2301 724 2307 796
rect 2397 784 2403 896
rect 2365 724 2371 736
rect 2381 704 2387 756
rect 2397 724 2403 776
rect 2228 677 2243 683
rect 2221 584 2227 676
rect 2333 644 2339 676
rect 2266 614 2278 616
rect 2251 606 2253 614
rect 2261 606 2263 614
rect 2271 606 2273 614
rect 2281 606 2283 614
rect 2291 606 2293 614
rect 2266 604 2278 606
rect 2221 524 2227 536
rect 2205 497 2227 503
rect 2141 404 2147 496
rect 2189 344 2195 456
rect 2173 324 2179 336
rect 2189 304 2195 316
rect 2205 304 2211 376
rect 2077 104 2083 156
rect 2109 144 2115 276
rect 2125 264 2131 276
rect 2141 104 2147 296
rect 2205 284 2211 296
rect 2157 144 2163 256
rect 2189 184 2195 276
rect 2221 184 2227 497
rect 2253 264 2259 536
rect 2317 424 2323 536
rect 2333 444 2339 536
rect 2333 303 2339 436
rect 2349 424 2355 536
rect 2365 524 2371 556
rect 2397 523 2403 676
rect 2413 664 2419 1036
rect 2429 944 2435 1576
rect 2509 1504 2515 1636
rect 2541 1504 2547 1676
rect 2445 1464 2451 1496
rect 2525 1484 2531 1496
rect 2445 1404 2451 1456
rect 2445 1084 2451 1316
rect 2477 1124 2483 1356
rect 2493 1344 2499 1416
rect 2541 1384 2547 1476
rect 2557 1463 2563 1496
rect 2573 1484 2579 1516
rect 2589 1504 2595 1716
rect 2605 1464 2611 1656
rect 2621 1624 2627 1696
rect 2653 1684 2659 1736
rect 2669 1684 2675 1716
rect 2717 1704 2723 1796
rect 2733 1744 2739 1816
rect 2749 1724 2755 1736
rect 2765 1724 2771 1916
rect 2893 1904 2899 2063
rect 2941 2024 2947 2063
rect 2781 1884 2787 1896
rect 2829 1884 2835 1896
rect 2909 1864 2915 2016
rect 2973 1904 2979 2016
rect 2989 1884 2995 1896
rect 3037 1884 3043 1896
rect 2797 1784 2803 1836
rect 2877 1823 2883 1856
rect 2861 1817 2883 1823
rect 2797 1744 2803 1756
rect 2813 1744 2819 1756
rect 2781 1724 2787 1736
rect 2845 1724 2851 1756
rect 2861 1744 2867 1817
rect 2925 1764 2931 1836
rect 2941 1784 2947 1876
rect 2621 1524 2627 1616
rect 2669 1544 2675 1636
rect 2685 1524 2691 1556
rect 2557 1457 2579 1463
rect 2573 1384 2579 1457
rect 2509 1324 2515 1376
rect 2557 1344 2563 1356
rect 2621 1324 2627 1396
rect 2541 1144 2547 1316
rect 2573 1284 2579 1296
rect 2637 1204 2643 1336
rect 2669 1324 2675 1356
rect 2548 1137 2563 1143
rect 2468 1097 2492 1103
rect 2509 1084 2515 1116
rect 2461 1064 2467 1076
rect 2445 804 2451 836
rect 2461 804 2467 1056
rect 2477 964 2483 976
rect 2429 604 2435 636
rect 2445 583 2451 776
rect 2468 737 2483 743
rect 2461 704 2467 736
rect 2477 664 2483 737
rect 2493 723 2499 1076
rect 2509 964 2515 1076
rect 2541 1044 2547 1076
rect 2557 943 2563 1137
rect 2637 1124 2643 1136
rect 2573 1024 2579 1076
rect 2605 1064 2611 1096
rect 2589 1004 2595 1036
rect 2621 964 2627 1036
rect 2637 984 2643 1116
rect 2653 1044 2659 1096
rect 2669 1024 2675 1116
rect 2557 937 2572 943
rect 2621 924 2627 936
rect 2653 924 2659 956
rect 2509 764 2515 836
rect 2541 764 2547 896
rect 2557 723 2563 836
rect 2589 744 2595 896
rect 2605 724 2611 796
rect 2493 717 2515 723
rect 2493 684 2499 696
rect 2493 664 2499 676
rect 2461 584 2467 656
rect 2429 577 2451 583
rect 2413 544 2419 576
rect 2429 524 2435 577
rect 2477 544 2483 556
rect 2493 544 2499 556
rect 2397 517 2419 523
rect 2333 297 2348 303
rect 2397 284 2403 336
rect 2413 304 2419 517
rect 2429 384 2435 516
rect 2477 304 2483 496
rect 2266 214 2278 216
rect 2251 206 2253 214
rect 2261 206 2263 214
rect 2271 206 2273 214
rect 2281 206 2283 214
rect 2291 206 2293 214
rect 2266 204 2278 206
rect 2317 144 2323 256
rect 2333 144 2339 236
rect 2413 184 2419 296
rect 2429 264 2435 296
rect 2493 284 2499 296
rect 2509 283 2515 717
rect 2541 717 2563 723
rect 2541 543 2547 717
rect 2557 604 2563 696
rect 2573 584 2579 616
rect 2589 604 2595 636
rect 2637 584 2643 756
rect 2653 684 2659 896
rect 2669 884 2675 956
rect 2685 864 2691 1076
rect 2701 1064 2707 1696
rect 2749 1544 2755 1636
rect 2733 1504 2739 1516
rect 2781 1484 2787 1716
rect 2877 1704 2883 1716
rect 2813 1504 2819 1596
rect 2829 1524 2835 1636
rect 2861 1484 2867 1496
rect 2877 1464 2883 1636
rect 2909 1504 2915 1696
rect 2925 1584 2931 1696
rect 3037 1524 3043 1536
rect 2909 1464 2915 1476
rect 2788 1457 2844 1463
rect 2925 1444 2931 1496
rect 2717 1404 2723 1436
rect 2797 1344 2803 1356
rect 2813 1324 2819 1416
rect 2845 1364 2851 1396
rect 2717 1304 2723 1316
rect 2749 1264 2755 1296
rect 2717 1104 2723 1236
rect 2781 1184 2787 1316
rect 2701 964 2707 1036
rect 2701 924 2707 936
rect 2717 924 2723 936
rect 2701 904 2707 916
rect 2685 724 2691 836
rect 2653 664 2659 676
rect 2669 644 2675 676
rect 2685 664 2691 680
rect 2653 564 2659 636
rect 2701 584 2707 636
rect 2733 584 2739 936
rect 2749 904 2755 916
rect 2532 537 2547 543
rect 2525 384 2531 536
rect 2557 523 2563 556
rect 2548 517 2563 523
rect 2541 504 2547 516
rect 2573 384 2579 496
rect 2525 344 2531 376
rect 2509 277 2531 283
rect 2525 264 2531 277
rect 2445 184 2451 236
rect 2557 224 2563 336
rect 2605 324 2611 516
rect 2612 317 2627 323
rect 2589 303 2595 316
rect 2589 297 2604 303
rect 2525 184 2531 216
rect 2157 24 2163 136
rect 2349 104 2355 136
rect 2013 -23 2035 -17
rect 2189 -23 2195 96
rect 2365 24 2371 156
rect 2493 144 2499 176
rect 2589 164 2595 256
rect 2621 163 2627 317
rect 2637 284 2643 536
rect 2685 284 2691 376
rect 2701 304 2707 556
rect 2717 464 2723 556
rect 2749 484 2755 516
rect 2765 503 2771 1116
rect 2797 1103 2803 1196
rect 2813 1124 2819 1236
rect 2797 1097 2819 1103
rect 2781 964 2787 1076
rect 2797 944 2803 1016
rect 2813 924 2819 1097
rect 2845 944 2851 1276
rect 2877 1144 2883 1316
rect 2893 1304 2899 1436
rect 2909 1344 2915 1376
rect 2925 1344 2931 1436
rect 2989 1404 2995 1496
rect 2973 1344 2979 1356
rect 2909 1184 2915 1316
rect 2973 1304 2979 1336
rect 2861 1064 2867 1076
rect 2829 924 2835 936
rect 2861 924 2867 1056
rect 2893 1024 2899 1036
rect 2877 944 2883 956
rect 2893 944 2899 996
rect 2973 983 2979 1096
rect 3021 984 3027 1496
rect 3037 1124 3043 1136
rect 2973 977 2995 983
rect 2989 964 2995 977
rect 3005 964 3011 976
rect 2877 924 2883 936
rect 2989 924 2995 936
rect 2781 724 2787 916
rect 2797 664 2803 896
rect 2829 824 2835 896
rect 2781 563 2787 636
rect 2813 584 2819 656
rect 2829 644 2835 696
rect 2845 684 2851 716
rect 2781 557 2796 563
rect 2829 524 2835 596
rect 2861 524 2867 676
rect 2877 524 2883 676
rect 2765 497 2787 503
rect 2765 444 2771 476
rect 2653 244 2659 256
rect 2669 164 2675 236
rect 2621 157 2652 163
rect 2477 24 2483 136
rect 2637 124 2643 157
rect 2701 144 2707 296
rect 2749 264 2755 436
rect 2765 243 2771 416
rect 2781 384 2787 497
rect 2781 304 2787 356
rect 2813 284 2819 356
rect 2829 323 2835 436
rect 2845 364 2851 436
rect 2877 424 2883 516
rect 2893 504 2899 576
rect 2909 504 2915 796
rect 2941 723 2947 736
rect 2941 717 2956 723
rect 2941 484 2947 656
rect 2829 317 2844 323
rect 2861 304 2867 376
rect 2749 237 2771 243
rect 2749 184 2755 237
rect 2733 124 2739 136
rect 2813 124 2819 256
rect 2877 244 2883 336
rect 2909 284 2915 316
rect 2925 304 2931 436
rect 2861 124 2867 236
rect 2925 224 2931 236
rect 2893 164 2899 216
rect 2957 184 2963 696
rect 2989 684 2995 856
rect 2973 544 2979 636
rect 3021 584 3027 956
rect 2973 164 2979 516
rect 3037 504 3043 636
rect 2989 124 2995 496
rect 3037 284 3043 296
rect 2637 104 2643 116
rect 3037 84 3043 96
rect 2429 -23 2435 16
rect 2845 -17 2851 36
rect 2941 -17 2947 36
rect 2829 -23 2851 -17
rect 2925 -23 2947 -17
<< m3contact >>
rect 739 2006 747 2014
rect 749 2006 757 2014
rect 759 2006 767 2014
rect 769 2006 777 2014
rect 779 2006 787 2014
rect 789 2006 797 2014
rect 796 1976 804 1984
rect 828 1976 836 1984
rect 188 1936 196 1944
rect 860 1936 868 1944
rect 44 1916 52 1924
rect 76 1916 84 1924
rect 508 1916 516 1924
rect 572 1916 580 1924
rect 636 1916 644 1924
rect 844 1916 852 1924
rect 892 1916 900 1924
rect 44 1896 52 1904
rect 60 1896 68 1904
rect 124 1896 132 1904
rect 332 1896 340 1904
rect 396 1896 404 1904
rect 460 1896 468 1904
rect 12 1856 20 1864
rect 92 1876 100 1884
rect 172 1876 180 1884
rect 92 1856 100 1864
rect 156 1756 164 1764
rect 108 1736 116 1744
rect 124 1716 132 1724
rect 220 1716 228 1724
rect 12 1696 20 1704
rect 44 1636 52 1644
rect 236 1696 244 1704
rect 268 1676 276 1684
rect 284 1656 292 1664
rect 332 1876 340 1884
rect 524 1876 532 1884
rect 364 1856 372 1864
rect 444 1856 452 1864
rect 604 1856 612 1864
rect 652 1856 660 1864
rect 316 1716 324 1724
rect 380 1776 388 1784
rect 364 1736 372 1744
rect 508 1796 516 1804
rect 444 1736 452 1744
rect 652 1836 660 1844
rect 556 1776 564 1784
rect 572 1756 580 1764
rect 636 1796 644 1804
rect 588 1716 596 1724
rect 700 1876 708 1884
rect 860 1856 868 1864
rect 892 1856 900 1864
rect 684 1836 692 1844
rect 684 1796 692 1804
rect 812 1796 820 1804
rect 700 1756 708 1764
rect 812 1756 820 1764
rect 828 1736 836 1744
rect 844 1736 852 1744
rect 700 1716 708 1724
rect 476 1696 484 1704
rect 492 1696 500 1704
rect 556 1696 564 1704
rect 604 1696 612 1704
rect 668 1696 676 1704
rect 316 1676 324 1684
rect 444 1676 452 1684
rect 300 1576 308 1584
rect 300 1516 308 1524
rect 28 1496 36 1504
rect 108 1496 116 1504
rect 156 1496 164 1504
rect 236 1496 244 1504
rect 284 1496 292 1504
rect 12 1476 20 1484
rect 76 1476 84 1484
rect 124 1476 132 1484
rect 60 1376 68 1384
rect 140 1436 148 1444
rect 92 1416 100 1424
rect 12 1356 20 1364
rect 28 1356 36 1364
rect 44 1296 52 1304
rect 60 1216 68 1224
rect 44 1116 52 1124
rect 12 1076 20 1084
rect 44 1076 52 1084
rect 76 1116 84 1124
rect 60 976 68 984
rect 204 1456 212 1464
rect 172 1416 180 1424
rect 396 1636 404 1644
rect 492 1636 500 1644
rect 348 1576 356 1584
rect 220 1436 228 1444
rect 140 1356 148 1364
rect 108 1336 116 1344
rect 172 1336 180 1344
rect 220 1336 228 1344
rect 156 1296 164 1304
rect 172 1296 180 1304
rect 204 1296 212 1304
rect 252 1296 260 1304
rect 172 1176 180 1184
rect 220 1136 228 1144
rect 188 1116 196 1124
rect 204 1076 212 1084
rect 124 936 132 944
rect 188 936 196 944
rect 204 936 212 944
rect 108 916 116 924
rect 12 896 20 904
rect 44 836 52 844
rect 268 1116 276 1124
rect 236 1096 244 1104
rect 332 1356 340 1364
rect 316 1336 324 1344
rect 444 1596 452 1604
rect 412 1556 420 1564
rect 396 1536 404 1544
rect 636 1676 644 1684
rect 812 1676 820 1684
rect 716 1656 724 1664
rect 652 1616 660 1624
rect 572 1596 580 1604
rect 508 1556 516 1564
rect 524 1556 532 1564
rect 556 1556 564 1564
rect 412 1516 420 1524
rect 428 1516 436 1524
rect 524 1516 532 1524
rect 556 1516 564 1524
rect 572 1516 580 1524
rect 380 1496 388 1504
rect 492 1496 500 1504
rect 508 1496 516 1504
rect 364 1476 372 1484
rect 460 1476 468 1484
rect 380 1456 388 1464
rect 460 1456 468 1464
rect 524 1476 532 1484
rect 556 1476 564 1484
rect 588 1476 596 1484
rect 476 1436 484 1444
rect 492 1436 500 1444
rect 476 1396 484 1404
rect 396 1376 404 1384
rect 364 1156 372 1164
rect 300 1136 308 1144
rect 332 1096 340 1104
rect 460 1336 468 1344
rect 236 1076 244 1084
rect 300 1056 308 1064
rect 668 1496 676 1504
rect 636 1476 644 1484
rect 604 1456 612 1464
rect 620 1436 628 1444
rect 604 1396 612 1404
rect 492 1376 500 1384
rect 572 1376 580 1384
rect 556 1336 564 1344
rect 668 1476 676 1484
rect 620 1336 628 1344
rect 700 1376 708 1384
rect 540 1316 548 1324
rect 668 1316 676 1324
rect 444 1156 452 1164
rect 460 1116 468 1124
rect 540 1236 548 1244
rect 524 1176 532 1184
rect 540 1156 548 1164
rect 476 1076 484 1084
rect 540 1076 548 1084
rect 556 1076 564 1084
rect 268 956 276 964
rect 268 936 276 944
rect 156 876 164 884
rect 92 716 100 724
rect 188 716 196 724
rect 268 716 276 724
rect 332 1016 340 1024
rect 316 956 324 964
rect 316 936 324 944
rect 380 996 388 1004
rect 364 976 372 984
rect 396 976 404 984
rect 428 1016 436 1024
rect 476 956 484 964
rect 508 956 516 964
rect 332 916 340 924
rect 412 916 420 924
rect 348 896 356 904
rect 380 876 388 884
rect 460 916 468 924
rect 492 916 500 924
rect 524 916 532 924
rect 604 1276 612 1284
rect 604 1216 612 1224
rect 684 1196 692 1204
rect 620 1156 628 1164
rect 812 1616 820 1624
rect 739 1606 747 1614
rect 749 1606 757 1614
rect 759 1606 767 1614
rect 769 1606 777 1614
rect 779 1606 787 1614
rect 789 1606 797 1614
rect 748 1576 756 1584
rect 732 1536 740 1544
rect 732 1516 740 1524
rect 764 1536 772 1544
rect 812 1436 820 1444
rect 716 1356 724 1364
rect 844 1676 852 1684
rect 940 1856 948 1864
rect 956 1856 964 1864
rect 924 1836 932 1844
rect 892 1796 900 1804
rect 956 1796 964 1804
rect 1020 1916 1028 1924
rect 1068 1916 1076 1924
rect 1084 1916 1092 1924
rect 1052 1876 1060 1884
rect 1132 1916 1140 1924
rect 1100 1876 1108 1884
rect 1004 1856 1012 1864
rect 988 1736 996 1744
rect 1020 1736 1028 1744
rect 940 1616 948 1624
rect 924 1596 932 1604
rect 956 1596 964 1604
rect 892 1536 900 1544
rect 860 1496 868 1504
rect 924 1496 932 1504
rect 956 1496 964 1504
rect 844 1436 852 1444
rect 1036 1716 1044 1724
rect 1068 1716 1076 1724
rect 1084 1696 1092 1704
rect 1100 1696 1108 1704
rect 1020 1656 1028 1664
rect 1036 1656 1044 1664
rect 1052 1636 1060 1644
rect 988 1516 996 1524
rect 1020 1516 1028 1524
rect 892 1456 900 1464
rect 876 1416 884 1424
rect 828 1336 836 1344
rect 956 1416 964 1424
rect 940 1356 948 1364
rect 924 1336 932 1344
rect 876 1316 884 1324
rect 908 1316 916 1324
rect 812 1276 820 1284
rect 739 1206 747 1214
rect 749 1206 757 1214
rect 759 1206 767 1214
rect 769 1206 777 1214
rect 779 1206 787 1214
rect 789 1206 797 1214
rect 652 1116 660 1124
rect 668 1116 676 1124
rect 636 1096 644 1104
rect 588 1016 596 1024
rect 620 1036 628 1044
rect 620 936 628 944
rect 652 936 660 944
rect 572 916 580 924
rect 604 916 612 924
rect 428 856 436 864
rect 60 696 68 704
rect 124 696 132 704
rect 220 696 228 704
rect 12 676 20 684
rect 316 716 324 724
rect 412 716 420 724
rect 460 716 468 724
rect 92 676 100 684
rect 204 676 212 684
rect 252 676 260 684
rect 284 676 292 684
rect 76 636 84 644
rect 156 656 164 664
rect 172 636 180 644
rect 204 616 212 624
rect 172 596 180 604
rect 92 576 100 584
rect 156 576 164 584
rect 188 576 196 584
rect 60 556 68 564
rect 92 556 100 564
rect 44 536 52 544
rect 300 656 308 664
rect 268 616 276 624
rect 236 576 244 584
rect 236 556 244 564
rect 348 696 356 704
rect 412 676 420 684
rect 364 656 372 664
rect 332 596 340 604
rect 204 536 212 544
rect 252 536 260 544
rect 284 536 292 544
rect 316 536 324 544
rect 92 516 100 524
rect 172 516 180 524
rect 300 516 308 524
rect 332 516 340 524
rect 108 496 116 504
rect 92 476 100 484
rect 28 316 36 324
rect 60 316 68 324
rect 60 296 68 304
rect 204 476 212 484
rect 140 456 148 464
rect 348 496 356 504
rect 396 616 404 624
rect 460 676 468 684
rect 444 656 452 664
rect 428 616 436 624
rect 508 616 516 624
rect 412 516 420 524
rect 380 496 388 504
rect 364 436 372 444
rect 380 416 388 424
rect 348 396 356 404
rect 140 316 148 324
rect 188 316 196 324
rect 76 276 84 284
rect 44 256 52 264
rect 28 176 36 184
rect 28 156 36 164
rect 60 236 68 244
rect 12 136 20 144
rect 44 136 52 144
rect 92 236 100 244
rect 140 296 148 304
rect 156 296 164 304
rect 236 296 244 304
rect 492 516 500 524
rect 444 496 452 504
rect 460 496 468 504
rect 428 436 436 444
rect 428 376 436 384
rect 268 296 276 304
rect 316 296 324 304
rect 348 296 356 304
rect 412 296 420 304
rect 156 276 164 284
rect 252 276 260 284
rect 316 276 324 284
rect 380 276 388 284
rect 412 276 420 284
rect 204 256 212 264
rect 220 256 228 264
rect 236 256 244 264
rect 284 256 292 264
rect 188 196 196 204
rect 92 156 100 164
rect 140 156 148 164
rect 188 156 196 164
rect 268 216 276 224
rect 508 416 516 424
rect 732 1116 740 1124
rect 700 1096 708 1104
rect 844 1196 852 1204
rect 876 1256 884 1264
rect 860 1096 868 1104
rect 908 1176 916 1184
rect 892 1116 900 1124
rect 972 1336 980 1344
rect 956 1296 964 1304
rect 988 1276 996 1284
rect 1068 1556 1076 1564
rect 1164 1816 1172 1824
rect 1356 1896 1364 1904
rect 1404 1896 1412 1904
rect 1516 1896 1524 1904
rect 1212 1856 1220 1864
rect 1132 1736 1140 1744
rect 1132 1716 1140 1724
rect 1244 1796 1252 1804
rect 1196 1776 1204 1784
rect 1244 1776 1252 1784
rect 1180 1736 1188 1744
rect 1340 1856 1348 1864
rect 1388 1776 1396 1784
rect 1292 1736 1300 1744
rect 1196 1716 1204 1724
rect 1164 1696 1172 1704
rect 1180 1696 1188 1704
rect 1260 1676 1268 1684
rect 1228 1656 1236 1664
rect 1148 1596 1156 1604
rect 1164 1596 1172 1604
rect 1116 1556 1124 1564
rect 1100 1536 1108 1544
rect 1116 1516 1124 1524
rect 1196 1536 1204 1544
rect 1164 1496 1172 1504
rect 1116 1476 1124 1484
rect 1148 1476 1156 1484
rect 1164 1476 1172 1484
rect 1132 1456 1140 1464
rect 1020 1436 1028 1444
rect 1036 1356 1044 1364
rect 1020 1316 1028 1324
rect 1068 1416 1076 1424
rect 1084 1396 1092 1404
rect 1116 1336 1124 1344
rect 1004 1256 1012 1264
rect 972 1196 980 1204
rect 1116 1316 1124 1324
rect 1356 1676 1364 1684
rect 1276 1656 1284 1664
rect 1212 1496 1220 1504
rect 1276 1496 1284 1504
rect 1212 1476 1220 1484
rect 1372 1616 1380 1624
rect 1324 1556 1332 1564
rect 1180 1456 1188 1464
rect 1244 1396 1252 1404
rect 1276 1456 1284 1464
rect 1372 1536 1380 1544
rect 1372 1476 1380 1484
rect 1452 1796 1460 1804
rect 1500 1796 1508 1804
rect 1436 1736 1444 1744
rect 1420 1716 1428 1724
rect 1404 1536 1412 1544
rect 1420 1536 1428 1544
rect 1500 1756 1508 1764
rect 1468 1716 1476 1724
rect 1500 1716 1508 1724
rect 1612 1916 1620 1924
rect 1692 1916 1700 1924
rect 1564 1856 1572 1864
rect 1788 1916 1796 1924
rect 1708 1896 1716 1904
rect 1740 1896 1748 1904
rect 1676 1876 1684 1884
rect 1708 1876 1716 1884
rect 1772 1876 1780 1884
rect 1660 1836 1668 1844
rect 1532 1756 1540 1764
rect 1548 1756 1556 1764
rect 1580 1756 1588 1764
rect 1612 1756 1620 1764
rect 1628 1756 1636 1764
rect 1580 1736 1588 1744
rect 1564 1696 1572 1704
rect 1532 1676 1540 1684
rect 1452 1576 1460 1584
rect 1404 1516 1412 1524
rect 1436 1516 1444 1524
rect 1516 1556 1524 1564
rect 1516 1536 1524 1544
rect 1500 1496 1508 1504
rect 1452 1476 1460 1484
rect 1308 1456 1316 1464
rect 1356 1456 1364 1464
rect 1388 1456 1396 1464
rect 1324 1416 1332 1424
rect 1260 1376 1268 1384
rect 1292 1376 1300 1384
rect 1164 1316 1172 1324
rect 1052 1296 1060 1304
rect 1148 1296 1156 1304
rect 1036 1176 1044 1184
rect 1020 1116 1028 1124
rect 1036 1096 1044 1104
rect 1148 1236 1156 1244
rect 1068 1176 1076 1184
rect 828 1056 836 1064
rect 908 1056 916 1064
rect 716 1036 724 1044
rect 796 996 804 1004
rect 812 936 820 944
rect 668 916 676 924
rect 684 916 692 924
rect 716 916 724 924
rect 684 896 692 904
rect 700 836 708 844
rect 668 756 676 764
rect 604 736 612 744
rect 652 736 660 744
rect 540 656 548 664
rect 540 636 548 644
rect 556 596 564 604
rect 636 696 644 704
rect 700 636 708 644
rect 636 596 644 604
rect 604 576 612 584
rect 620 536 628 544
rect 668 536 676 544
rect 636 516 644 524
rect 652 516 660 524
rect 739 806 747 814
rect 749 806 757 814
rect 759 806 767 814
rect 769 806 777 814
rect 779 806 787 814
rect 789 806 797 814
rect 844 916 852 924
rect 972 956 980 964
rect 940 916 948 924
rect 1052 936 1060 944
rect 1020 916 1028 924
rect 1036 916 1044 924
rect 892 896 900 904
rect 956 896 964 904
rect 972 896 980 904
rect 924 816 932 824
rect 732 716 740 724
rect 908 716 916 724
rect 828 696 836 704
rect 828 676 836 684
rect 812 636 820 644
rect 716 516 724 524
rect 732 496 740 504
rect 572 456 580 464
rect 716 456 724 464
rect 716 436 724 444
rect 492 316 500 324
rect 524 316 532 324
rect 540 316 548 324
rect 476 296 484 304
rect 508 276 516 284
rect 739 406 747 414
rect 749 406 757 414
rect 759 406 767 414
rect 769 406 777 414
rect 779 406 787 414
rect 789 406 797 414
rect 668 356 676 364
rect 732 316 740 324
rect 620 296 628 304
rect 620 276 628 284
rect 444 256 452 264
rect 572 256 580 264
rect 348 196 356 204
rect 396 196 404 204
rect 332 156 340 164
rect 684 236 692 244
rect 508 216 516 224
rect 428 176 436 184
rect 476 176 484 184
rect 524 176 532 184
rect 156 136 164 144
rect 204 136 212 144
rect 364 136 372 144
rect 412 136 420 144
rect 460 136 468 144
rect 172 116 180 124
rect 236 116 244 124
rect 300 116 308 124
rect 492 156 500 164
rect 524 156 532 164
rect 540 136 548 144
rect 476 116 484 124
rect 540 116 548 124
rect 620 136 628 144
rect 268 96 276 104
rect 556 96 564 104
rect 876 656 884 664
rect 844 596 852 604
rect 860 596 868 604
rect 828 516 836 524
rect 892 516 900 524
rect 988 876 996 884
rect 1020 876 1028 884
rect 1180 1256 1188 1264
rect 1084 1096 1092 1104
rect 1084 1016 1092 1024
rect 1100 996 1108 1004
rect 1228 1356 1236 1364
rect 1228 1336 1236 1344
rect 1244 1336 1252 1344
rect 1212 1316 1220 1324
rect 1196 1216 1204 1224
rect 1196 1156 1204 1164
rect 1356 1416 1364 1424
rect 1388 1356 1396 1364
rect 1276 1316 1284 1324
rect 1308 1316 1316 1324
rect 1340 1316 1348 1324
rect 1356 1316 1364 1324
rect 1452 1336 1460 1344
rect 1324 1296 1332 1304
rect 1372 1296 1380 1304
rect 1596 1716 1604 1724
rect 1628 1676 1636 1684
rect 1708 1776 1716 1784
rect 1692 1736 1700 1744
rect 1740 1756 1748 1764
rect 1676 1676 1684 1684
rect 1596 1656 1604 1664
rect 1660 1656 1668 1664
rect 1692 1656 1700 1664
rect 1580 1596 1588 1604
rect 1548 1476 1556 1484
rect 1564 1456 1572 1464
rect 1532 1436 1540 1444
rect 1596 1476 1604 1484
rect 1676 1576 1684 1584
rect 1644 1476 1652 1484
rect 1660 1476 1668 1484
rect 1644 1436 1652 1444
rect 1660 1436 1668 1444
rect 1612 1416 1620 1424
rect 1708 1556 1716 1564
rect 1852 1916 1860 1924
rect 1852 1896 1860 1904
rect 1884 1896 1892 1904
rect 2028 1936 2036 1944
rect 2412 1936 2420 1944
rect 1996 1916 2004 1924
rect 1980 1896 1988 1904
rect 1900 1876 1908 1884
rect 1788 1856 1796 1864
rect 1804 1856 1812 1864
rect 1836 1856 1844 1864
rect 1868 1856 1876 1864
rect 1916 1856 1924 1864
rect 1980 1876 1988 1884
rect 1804 1836 1812 1844
rect 1932 1836 1940 1844
rect 1852 1816 1860 1824
rect 1900 1796 1908 1804
rect 1964 1796 1972 1804
rect 1820 1776 1828 1784
rect 1868 1756 1876 1764
rect 1788 1736 1796 1744
rect 1772 1696 1780 1704
rect 1788 1696 1796 1704
rect 1740 1656 1748 1664
rect 1772 1636 1780 1644
rect 1836 1616 1844 1624
rect 1900 1616 1908 1624
rect 1836 1556 1844 1564
rect 1724 1536 1732 1544
rect 1756 1516 1764 1524
rect 1852 1496 1860 1504
rect 1788 1476 1796 1484
rect 1692 1416 1700 1424
rect 1628 1396 1636 1404
rect 1660 1396 1668 1404
rect 1644 1356 1652 1364
rect 1532 1316 1540 1324
rect 1628 1316 1636 1324
rect 1484 1276 1492 1284
rect 1260 1236 1268 1244
rect 1228 1216 1236 1224
rect 1132 996 1140 1004
rect 1164 996 1172 1004
rect 1116 976 1124 984
rect 1212 1016 1220 1024
rect 1196 956 1204 964
rect 1036 816 1044 824
rect 1052 816 1060 824
rect 1036 736 1044 744
rect 1052 716 1060 724
rect 1036 696 1044 704
rect 972 676 980 684
rect 956 656 964 664
rect 940 576 948 584
rect 860 496 868 504
rect 876 496 884 504
rect 924 496 932 504
rect 828 456 836 464
rect 876 456 884 464
rect 892 436 900 444
rect 860 376 868 384
rect 844 356 852 364
rect 876 336 884 344
rect 828 296 836 304
rect 1004 656 1012 664
rect 988 596 996 604
rect 988 576 996 584
rect 1020 536 1028 544
rect 1004 516 1012 524
rect 1020 476 1028 484
rect 956 396 964 404
rect 908 356 916 364
rect 1004 356 1012 364
rect 892 316 900 324
rect 876 296 884 304
rect 940 296 948 304
rect 1036 336 1044 344
rect 988 316 996 324
rect 1084 656 1092 664
rect 1068 576 1076 584
rect 1244 1096 1252 1104
rect 1132 936 1140 944
rect 1116 816 1124 824
rect 1164 816 1172 824
rect 1132 696 1140 704
rect 1324 1156 1332 1164
rect 1532 1236 1540 1244
rect 1468 1216 1476 1224
rect 1420 1156 1428 1164
rect 1436 1156 1444 1164
rect 1308 1096 1316 1104
rect 1276 1056 1284 1064
rect 1308 1056 1316 1064
rect 1324 1056 1332 1064
rect 1452 1056 1460 1064
rect 1292 1016 1300 1024
rect 1276 976 1284 984
rect 1228 916 1236 924
rect 1212 856 1220 864
rect 1484 1116 1492 1124
rect 1500 1096 1508 1104
rect 1516 1096 1524 1104
rect 1596 1176 1604 1184
rect 1548 1116 1556 1124
rect 1548 996 1556 1004
rect 1580 996 1588 1004
rect 1308 956 1316 964
rect 1436 956 1444 964
rect 1484 956 1492 964
rect 1532 956 1540 964
rect 1292 896 1300 904
rect 1340 896 1348 904
rect 1180 756 1188 764
rect 1244 796 1252 804
rect 1228 756 1236 764
rect 1276 736 1284 744
rect 1180 616 1188 624
rect 1196 596 1204 604
rect 1244 576 1252 584
rect 1116 556 1124 564
rect 1196 556 1204 564
rect 1212 556 1220 564
rect 1260 556 1268 564
rect 1132 536 1140 544
rect 1084 456 1092 464
rect 1180 456 1188 464
rect 1148 436 1156 444
rect 1196 436 1204 444
rect 1132 396 1140 404
rect 1244 516 1252 524
rect 1404 896 1412 904
rect 1388 856 1396 864
rect 1612 1156 1620 1164
rect 1644 1116 1652 1124
rect 1612 1096 1620 1104
rect 1676 1376 1684 1384
rect 1724 1396 1732 1404
rect 1756 1376 1764 1384
rect 1740 1356 1748 1364
rect 1820 1456 1828 1464
rect 1884 1476 1892 1484
rect 1868 1456 1876 1464
rect 1804 1396 1812 1404
rect 1852 1396 1860 1404
rect 1820 1376 1828 1384
rect 1772 1356 1780 1364
rect 1852 1356 1860 1364
rect 1708 1296 1716 1304
rect 1692 1216 1700 1224
rect 1724 1096 1732 1104
rect 1628 996 1636 1004
rect 1612 956 1620 964
rect 1628 936 1636 944
rect 1548 916 1556 924
rect 1596 916 1604 924
rect 1468 896 1476 904
rect 1420 876 1428 884
rect 1516 876 1524 884
rect 1580 876 1588 884
rect 1372 756 1380 764
rect 1356 716 1364 724
rect 1404 736 1412 744
rect 1388 696 1396 704
rect 1292 576 1300 584
rect 1356 676 1364 684
rect 1404 676 1412 684
rect 1548 816 1556 824
rect 1644 876 1652 884
rect 1644 856 1652 864
rect 1612 776 1620 784
rect 1436 756 1444 764
rect 1564 736 1572 744
rect 1500 716 1508 724
rect 1452 696 1460 704
rect 1532 676 1540 684
rect 1340 656 1348 664
rect 1404 636 1412 644
rect 1676 916 1684 924
rect 1708 916 1716 924
rect 1804 1336 1812 1344
rect 1772 1316 1780 1324
rect 1836 1316 1844 1324
rect 1868 1336 1876 1344
rect 1884 1256 1892 1264
rect 1788 1216 1796 1224
rect 1788 1156 1796 1164
rect 1852 1156 1860 1164
rect 1772 1076 1780 1084
rect 1788 1076 1796 1084
rect 1788 1036 1796 1044
rect 1772 1016 1780 1024
rect 1820 1116 1828 1124
rect 1916 1556 1924 1564
rect 2092 1916 2100 1924
rect 2172 1916 2180 1924
rect 2268 1916 2276 1924
rect 2364 1916 2372 1924
rect 2396 1916 2404 1924
rect 2460 1916 2468 1924
rect 2524 1916 2532 1924
rect 2044 1896 2052 1904
rect 2060 1896 2068 1904
rect 2108 1896 2116 1904
rect 2012 1856 2020 1864
rect 2044 1836 2052 1844
rect 2012 1736 2020 1744
rect 2044 1736 2052 1744
rect 2044 1716 2052 1724
rect 1948 1676 1956 1684
rect 1996 1676 2004 1684
rect 2012 1676 2020 1684
rect 2028 1616 2036 1624
rect 1948 1576 1956 1584
rect 1932 1516 1940 1524
rect 1964 1516 1972 1524
rect 2012 1496 2020 1504
rect 2380 1896 2388 1904
rect 2412 1896 2420 1904
rect 2188 1876 2196 1884
rect 2156 1856 2164 1864
rect 2076 1796 2084 1804
rect 2108 1796 2116 1804
rect 2092 1776 2100 1784
rect 2108 1756 2116 1764
rect 2140 1736 2148 1744
rect 2108 1696 2116 1704
rect 2124 1676 2132 1684
rect 2140 1676 2148 1684
rect 2060 1656 2068 1664
rect 2172 1796 2180 1804
rect 2204 1796 2212 1804
rect 2188 1736 2196 1744
rect 2204 1736 2212 1744
rect 2188 1676 2196 1684
rect 2243 1806 2251 1814
rect 2253 1806 2261 1814
rect 2263 1806 2271 1814
rect 2273 1806 2281 1814
rect 2283 1806 2291 1814
rect 2293 1806 2301 1814
rect 2076 1636 2084 1644
rect 2060 1576 2068 1584
rect 2140 1596 2148 1604
rect 2124 1536 2132 1544
rect 1996 1476 2004 1484
rect 2028 1476 2036 1484
rect 2044 1476 2052 1484
rect 2092 1480 2100 1484
rect 2092 1476 2100 1480
rect 1916 1456 1924 1464
rect 1948 1456 1956 1464
rect 2108 1416 2116 1424
rect 1980 1376 1988 1384
rect 2028 1376 2036 1384
rect 2044 1376 2052 1384
rect 1932 1336 1940 1344
rect 2012 1336 2020 1344
rect 1916 1256 1924 1264
rect 1916 1236 1924 1244
rect 1900 1216 1908 1224
rect 2140 1496 2148 1504
rect 2220 1656 2228 1664
rect 2268 1736 2276 1744
rect 2284 1676 2292 1684
rect 2380 1876 2388 1884
rect 2444 1876 2452 1884
rect 2348 1816 2356 1824
rect 2380 1796 2388 1804
rect 2364 1756 2372 1764
rect 2348 1736 2356 1744
rect 2332 1636 2340 1644
rect 2236 1616 2244 1624
rect 2236 1556 2244 1564
rect 2316 1536 2324 1544
rect 2204 1496 2212 1504
rect 2156 1476 2164 1484
rect 2188 1456 2196 1464
rect 2156 1416 2164 1424
rect 2156 1356 2164 1364
rect 2124 1336 2132 1344
rect 2348 1516 2356 1524
rect 2243 1406 2251 1414
rect 2253 1406 2261 1414
rect 2263 1406 2271 1414
rect 2273 1406 2281 1414
rect 2283 1406 2291 1414
rect 2293 1406 2301 1414
rect 2172 1316 2180 1324
rect 2204 1316 2212 1324
rect 2284 1316 2292 1324
rect 2076 1296 2084 1304
rect 1932 1156 1940 1164
rect 1964 1156 1972 1164
rect 2284 1296 2292 1304
rect 2172 1276 2180 1284
rect 2092 1256 2100 1264
rect 2076 1156 2084 1164
rect 1884 1096 1892 1104
rect 2204 1236 2212 1244
rect 2156 1156 2164 1164
rect 2140 1116 2148 1124
rect 1836 1036 1844 1044
rect 1852 1036 1860 1044
rect 1900 1036 1908 1044
rect 1820 1016 1828 1024
rect 1836 956 1844 964
rect 1804 936 1812 944
rect 1676 896 1684 904
rect 1724 896 1732 904
rect 1676 736 1684 744
rect 1740 816 1748 824
rect 1788 796 1796 804
rect 1756 736 1764 744
rect 1724 716 1732 724
rect 1660 696 1668 704
rect 1548 636 1556 644
rect 1596 636 1604 644
rect 1324 596 1332 604
rect 1420 596 1428 604
rect 1308 556 1316 564
rect 1500 616 1508 624
rect 1452 576 1460 584
rect 1484 576 1492 584
rect 1340 556 1348 564
rect 1404 556 1412 564
rect 1468 556 1476 564
rect 1484 556 1492 564
rect 1532 556 1540 564
rect 1548 556 1556 564
rect 1372 516 1380 524
rect 1276 476 1284 484
rect 1228 396 1236 404
rect 1116 356 1124 364
rect 1372 376 1380 384
rect 1276 336 1284 344
rect 1356 336 1364 344
rect 988 296 996 304
rect 972 276 980 284
rect 1020 276 1028 284
rect 1052 276 1060 284
rect 1084 276 1092 284
rect 1036 256 1044 264
rect 940 236 948 244
rect 844 196 852 204
rect 860 176 868 184
rect 812 156 820 164
rect 876 156 884 164
rect 972 156 980 164
rect 1004 156 1012 164
rect 732 136 740 144
rect 844 136 852 144
rect 620 96 628 104
rect 636 76 644 84
rect 924 136 932 144
rect 908 116 916 124
rect 956 116 964 124
rect 1084 256 1092 264
rect 1308 316 1316 324
rect 1180 296 1188 304
rect 1228 296 1236 304
rect 1148 276 1156 284
rect 1388 276 1396 284
rect 1420 516 1428 524
rect 1452 496 1460 504
rect 1500 496 1508 504
rect 1564 516 1572 524
rect 1596 516 1604 524
rect 1580 496 1588 504
rect 1532 476 1540 484
rect 1596 476 1604 484
rect 1436 316 1444 324
rect 1500 316 1508 324
rect 1724 676 1732 684
rect 1628 656 1636 664
rect 1708 656 1716 664
rect 1756 636 1764 644
rect 1708 596 1716 604
rect 1772 596 1780 604
rect 1676 576 1684 584
rect 1644 556 1652 564
rect 1820 636 1828 644
rect 1820 576 1828 584
rect 1692 536 1700 544
rect 1724 536 1732 544
rect 1692 496 1700 504
rect 1628 476 1636 484
rect 1564 456 1572 464
rect 1612 456 1620 464
rect 1564 316 1572 324
rect 1164 256 1172 264
rect 1180 256 1188 264
rect 1228 256 1236 264
rect 1292 256 1300 264
rect 1148 236 1156 244
rect 1132 216 1140 224
rect 1260 236 1268 244
rect 1180 216 1188 224
rect 1148 196 1156 204
rect 1100 156 1108 164
rect 1068 136 1076 144
rect 1244 196 1252 204
rect 1276 196 1284 204
rect 1164 156 1172 164
rect 1212 156 1220 164
rect 1020 116 1028 124
rect 1068 116 1076 124
rect 1196 116 1204 124
rect 1228 116 1236 124
rect 700 96 708 104
rect 812 96 820 104
rect 892 96 900 104
rect 924 96 932 104
rect 972 96 980 104
rect 684 76 692 84
rect 739 6 747 14
rect 749 6 757 14
rect 759 6 767 14
rect 769 6 777 14
rect 779 6 787 14
rect 789 6 797 14
rect 1340 256 1348 264
rect 1356 256 1364 264
rect 1484 276 1492 284
rect 1420 196 1428 204
rect 1468 196 1476 204
rect 1324 176 1332 184
rect 1372 176 1380 184
rect 1292 136 1300 144
rect 1516 256 1524 264
rect 1548 256 1556 264
rect 1532 216 1540 224
rect 1596 256 1604 264
rect 1564 236 1572 244
rect 1468 136 1476 144
rect 1500 136 1508 144
rect 1516 136 1524 144
rect 1580 136 1588 144
rect 1740 456 1748 464
rect 1772 556 1780 564
rect 1804 556 1812 564
rect 1788 536 1796 544
rect 1804 516 1812 524
rect 1820 496 1828 504
rect 1772 456 1780 464
rect 1820 436 1828 444
rect 1932 956 1940 964
rect 1900 936 1908 944
rect 1932 936 1940 944
rect 1884 916 1892 924
rect 1900 916 1908 924
rect 1852 756 1860 764
rect 1852 716 1860 724
rect 1868 676 1876 684
rect 1852 656 1860 664
rect 1868 636 1876 644
rect 1852 616 1860 624
rect 1868 576 1876 584
rect 1852 496 1860 504
rect 1868 496 1876 504
rect 1852 476 1860 484
rect 1852 396 1860 404
rect 1740 336 1748 344
rect 1772 296 1780 304
rect 1724 276 1732 284
rect 1628 256 1636 264
rect 1660 256 1668 264
rect 1708 236 1716 244
rect 1788 236 1796 244
rect 1740 156 1748 164
rect 1356 116 1364 124
rect 1404 116 1412 124
rect 1436 116 1444 124
rect 1484 116 1492 124
rect 1532 116 1540 124
rect 1596 116 1604 124
rect 1612 116 1620 124
rect 1644 116 1652 124
rect 1692 116 1700 124
rect 1324 96 1332 104
rect 1372 96 1380 104
rect 1452 96 1460 104
rect 1308 76 1316 84
rect 1868 316 1876 324
rect 1868 276 1876 284
rect 1852 256 1860 264
rect 1932 816 1940 824
rect 1900 756 1908 764
rect 1980 1096 1988 1104
rect 1948 736 1956 744
rect 1948 716 1956 724
rect 2252 1156 2260 1164
rect 1996 1076 2004 1084
rect 2012 956 2020 964
rect 2012 896 2020 904
rect 1980 776 1988 784
rect 1996 736 2004 744
rect 1916 676 1924 684
rect 1964 676 1972 684
rect 1916 656 1924 664
rect 1916 636 1924 644
rect 1900 576 1908 584
rect 1900 516 1908 524
rect 1964 596 1972 604
rect 1964 576 1972 584
rect 1948 536 1956 544
rect 1916 416 1924 424
rect 1916 316 1924 324
rect 1916 256 1924 264
rect 1900 156 1908 164
rect 1964 516 1972 524
rect 2124 1016 2132 1024
rect 2172 996 2180 1004
rect 2092 976 2100 984
rect 2108 976 2116 984
rect 2156 976 2164 984
rect 2044 856 2052 864
rect 2028 836 2036 844
rect 2156 936 2164 944
rect 2140 916 2148 924
rect 2236 1036 2244 1044
rect 2220 1016 2228 1024
rect 2243 1006 2251 1014
rect 2253 1006 2261 1014
rect 2263 1006 2271 1014
rect 2273 1006 2281 1014
rect 2283 1006 2291 1014
rect 2293 1006 2301 1014
rect 2220 976 2228 984
rect 2332 1396 2340 1404
rect 2444 1856 2452 1864
rect 2620 1916 2628 1924
rect 2508 1896 2516 1904
rect 2556 1896 2564 1904
rect 2572 1896 2580 1904
rect 2524 1816 2532 1824
rect 2796 1916 2804 1924
rect 2828 1916 2836 1924
rect 2668 1896 2676 1904
rect 2732 1896 2740 1904
rect 2588 1876 2596 1884
rect 2620 1876 2628 1884
rect 2572 1856 2580 1864
rect 2572 1816 2580 1824
rect 2492 1796 2500 1804
rect 2556 1796 2564 1804
rect 2492 1756 2500 1764
rect 2396 1736 2404 1744
rect 2444 1736 2452 1744
rect 2476 1736 2484 1744
rect 2572 1756 2580 1764
rect 2716 1876 2724 1884
rect 2604 1856 2612 1864
rect 2652 1856 2660 1864
rect 2732 1816 2740 1824
rect 2716 1796 2724 1804
rect 2700 1756 2708 1764
rect 2620 1736 2628 1744
rect 2652 1736 2660 1744
rect 2540 1676 2548 1684
rect 2556 1676 2564 1684
rect 2524 1656 2532 1664
rect 2508 1636 2516 1644
rect 2396 1596 2404 1604
rect 2380 1556 2388 1564
rect 2364 1456 2372 1464
rect 2364 1416 2372 1424
rect 2364 1396 2372 1404
rect 2428 1576 2436 1584
rect 2412 1456 2420 1464
rect 2396 1376 2404 1384
rect 2396 1356 2404 1364
rect 2364 1336 2372 1344
rect 2412 1336 2420 1344
rect 2396 1316 2404 1324
rect 2396 1256 2404 1264
rect 2380 1216 2388 1224
rect 2332 1096 2340 1104
rect 2332 1076 2340 1084
rect 2348 1076 2356 1084
rect 2396 1096 2404 1104
rect 2412 1076 2420 1084
rect 2380 1036 2388 1044
rect 2412 1036 2420 1044
rect 2364 1016 2372 1024
rect 2220 936 2228 944
rect 2316 936 2324 944
rect 2380 936 2388 944
rect 2396 936 2404 944
rect 2204 896 2212 904
rect 2092 796 2100 804
rect 2092 776 2100 784
rect 2060 736 2068 744
rect 2140 756 2148 764
rect 2204 736 2212 744
rect 2124 716 2132 724
rect 2204 716 2212 724
rect 2012 676 2020 684
rect 1996 656 2004 664
rect 2076 656 2084 664
rect 2028 636 2036 644
rect 1996 616 2004 624
rect 2044 556 2052 564
rect 2012 536 2020 544
rect 2060 536 2068 544
rect 2092 616 2100 624
rect 2124 656 2132 664
rect 2172 616 2180 624
rect 2108 596 2116 604
rect 2140 596 2148 604
rect 2124 556 2132 564
rect 2044 516 2052 524
rect 2076 516 2084 524
rect 2108 536 2116 544
rect 2124 516 2132 524
rect 2092 436 2100 444
rect 2044 416 2052 424
rect 1996 376 2004 384
rect 1996 316 2004 324
rect 2092 376 2100 384
rect 2060 336 2068 344
rect 2060 276 2068 284
rect 1996 176 2004 184
rect 1964 156 1972 164
rect 2012 156 2020 164
rect 1820 136 1828 144
rect 1836 136 1844 144
rect 1948 136 1956 144
rect 1772 116 1780 124
rect 1820 116 1828 124
rect 1804 96 1812 104
rect 1740 16 1748 24
rect 1772 16 1780 24
rect 1916 116 1924 124
rect 1980 116 1988 124
rect 1884 96 1892 104
rect 2060 236 2068 244
rect 2188 556 2196 564
rect 2172 536 2180 544
rect 2140 496 2148 504
rect 2220 696 2228 704
rect 2396 896 2404 904
rect 2252 856 2260 864
rect 2268 816 2276 824
rect 2300 796 2308 804
rect 2396 776 2404 784
rect 2380 756 2388 764
rect 2252 716 2260 724
rect 2332 716 2340 724
rect 2364 716 2372 724
rect 2396 676 2404 684
rect 2380 656 2388 664
rect 2332 636 2340 644
rect 2243 606 2251 614
rect 2253 606 2261 614
rect 2263 606 2271 614
rect 2273 606 2281 614
rect 2283 606 2291 614
rect 2293 606 2301 614
rect 2364 556 2372 564
rect 2220 536 2228 544
rect 2332 536 2340 544
rect 2188 456 2196 464
rect 2140 396 2148 404
rect 2204 376 2212 384
rect 2172 336 2180 344
rect 2188 336 2196 344
rect 2188 316 2196 324
rect 2124 296 2132 304
rect 2044 176 2052 184
rect 2060 156 2068 164
rect 2060 136 2068 144
rect 2028 116 2036 124
rect 2124 256 2132 264
rect 2108 136 2116 144
rect 2204 276 2212 284
rect 2156 256 2164 264
rect 2236 316 2244 324
rect 2316 416 2324 424
rect 2492 1516 2500 1524
rect 2572 1516 2580 1524
rect 2444 1496 2452 1504
rect 2540 1496 2548 1504
rect 2524 1476 2532 1484
rect 2460 1456 2468 1464
rect 2492 1416 2500 1424
rect 2444 1396 2452 1404
rect 2444 1356 2452 1364
rect 2460 1336 2468 1344
rect 2444 1316 2452 1324
rect 2604 1656 2612 1664
rect 2748 1736 2756 1744
rect 2908 2016 2916 2024
rect 2940 2016 2948 2024
rect 2972 2016 2980 2024
rect 2780 1896 2788 1904
rect 2828 1896 2836 1904
rect 2876 1896 2884 1904
rect 2892 1896 2900 1904
rect 2956 1896 2964 1904
rect 3036 1896 3044 1904
rect 2940 1876 2948 1884
rect 2988 1876 2996 1884
rect 2860 1856 2868 1864
rect 2908 1856 2916 1864
rect 2796 1776 2804 1784
rect 2796 1756 2804 1764
rect 2844 1756 2852 1764
rect 2780 1736 2788 1744
rect 2812 1736 2820 1744
rect 2924 1756 2932 1764
rect 2988 1756 2996 1764
rect 2860 1736 2868 1744
rect 2956 1736 2964 1744
rect 2764 1716 2772 1724
rect 2700 1696 2708 1704
rect 2716 1696 2724 1704
rect 2668 1676 2676 1684
rect 2620 1616 2628 1624
rect 2684 1556 2692 1564
rect 2620 1516 2628 1524
rect 2652 1496 2660 1504
rect 2684 1496 2692 1504
rect 2636 1436 2644 1444
rect 2620 1396 2628 1404
rect 2508 1376 2516 1384
rect 2540 1376 2548 1384
rect 2556 1356 2564 1364
rect 2604 1336 2612 1344
rect 2524 1316 2532 1324
rect 2524 1156 2532 1164
rect 2572 1276 2580 1284
rect 2668 1316 2676 1324
rect 2636 1196 2644 1204
rect 2540 1136 2548 1144
rect 2476 1116 2484 1124
rect 2492 1096 2500 1104
rect 2540 1096 2548 1104
rect 2444 1076 2452 1084
rect 2492 1076 2500 1084
rect 2508 1076 2516 1084
rect 2460 1056 2468 1064
rect 2428 936 2436 944
rect 2444 916 2452 924
rect 2476 976 2484 984
rect 2444 796 2452 804
rect 2460 796 2468 804
rect 2444 776 2452 784
rect 2428 596 2436 604
rect 2412 576 2420 584
rect 2460 736 2468 744
rect 2540 1036 2548 1044
rect 2508 956 2516 964
rect 2636 1116 2644 1124
rect 2604 1096 2612 1104
rect 2572 1016 2580 1024
rect 2588 996 2596 1004
rect 2604 976 2612 984
rect 2652 1036 2660 1044
rect 2668 1016 2676 1024
rect 2636 976 2644 984
rect 2620 956 2628 964
rect 2652 956 2660 964
rect 2668 956 2676 964
rect 2572 936 2580 944
rect 2508 916 2516 924
rect 2620 916 2628 924
rect 2636 896 2644 904
rect 2652 896 2660 904
rect 2556 836 2564 844
rect 2508 756 2516 764
rect 2540 756 2548 764
rect 2604 796 2612 804
rect 2588 736 2596 744
rect 2636 756 2644 764
rect 2492 696 2500 704
rect 2460 656 2468 664
rect 2492 656 2500 664
rect 2460 576 2468 584
rect 2476 556 2484 564
rect 2444 536 2452 544
rect 2492 536 2500 544
rect 2364 456 2372 464
rect 2348 416 2356 424
rect 2396 336 2404 344
rect 2348 296 2356 304
rect 2460 516 2468 524
rect 2476 496 2484 504
rect 2428 376 2436 384
rect 2492 476 2500 484
rect 2428 296 2436 304
rect 2492 296 2500 304
rect 2380 276 2388 284
rect 2236 256 2244 264
rect 2364 256 2372 264
rect 2243 206 2251 214
rect 2253 206 2261 214
rect 2263 206 2271 214
rect 2273 206 2281 214
rect 2283 206 2291 214
rect 2293 206 2301 214
rect 2620 696 2628 704
rect 2572 616 2580 624
rect 2556 596 2564 604
rect 2588 596 2596 604
rect 2748 1536 2756 1544
rect 2732 1516 2740 1524
rect 2764 1496 2772 1504
rect 2876 1696 2884 1704
rect 2908 1696 2916 1704
rect 2956 1696 2964 1704
rect 2812 1596 2820 1604
rect 2828 1516 2836 1524
rect 2844 1496 2852 1504
rect 2860 1496 2868 1504
rect 2748 1476 2756 1484
rect 2924 1576 2932 1584
rect 3036 1516 3044 1524
rect 2908 1496 2916 1504
rect 2972 1496 2980 1504
rect 3020 1496 3028 1504
rect 2908 1456 2916 1464
rect 2940 1476 2948 1484
rect 2924 1436 2932 1444
rect 2812 1416 2820 1424
rect 2716 1396 2724 1404
rect 2796 1356 2804 1364
rect 2844 1396 2852 1404
rect 2716 1296 2724 1304
rect 2748 1256 2756 1264
rect 2860 1296 2868 1304
rect 2844 1276 2852 1284
rect 2796 1196 2804 1204
rect 2780 1176 2788 1184
rect 2732 1116 2740 1124
rect 2764 1116 2772 1124
rect 2716 1096 2724 1104
rect 2700 1056 2708 1064
rect 2700 956 2708 964
rect 2716 936 2724 944
rect 2732 936 2740 944
rect 2700 916 2708 924
rect 2700 896 2708 904
rect 2684 856 2692 864
rect 2684 716 2692 724
rect 2652 656 2660 664
rect 2684 656 2692 664
rect 2652 636 2660 644
rect 2668 636 2676 644
rect 2700 636 2708 644
rect 2748 916 2756 924
rect 2748 696 2756 704
rect 2732 576 2740 584
rect 2652 556 2660 564
rect 2700 556 2708 564
rect 2620 536 2628 544
rect 2636 536 2644 544
rect 2684 536 2692 544
rect 2604 516 2612 524
rect 2540 496 2548 504
rect 2572 496 2580 504
rect 2524 376 2532 384
rect 2524 336 2532 344
rect 2524 296 2532 304
rect 2524 256 2532 264
rect 2572 296 2580 304
rect 2588 256 2596 264
rect 2524 216 2532 224
rect 2556 216 2564 224
rect 2444 176 2452 184
rect 2492 176 2500 184
rect 2316 136 2324 144
rect 2332 136 2340 144
rect 2076 96 2084 104
rect 2140 96 2148 104
rect 2188 96 2196 104
rect 2348 96 2356 104
rect 2156 16 2164 24
rect 2668 516 2676 524
rect 2684 376 2692 384
rect 2732 496 2740 504
rect 2780 1096 2788 1104
rect 2812 1116 2820 1124
rect 2796 1016 2804 1024
rect 2780 956 2788 964
rect 2828 1076 2836 1084
rect 2908 1376 2916 1384
rect 2988 1396 2996 1404
rect 2940 1376 2948 1384
rect 2988 1356 2996 1364
rect 2972 1336 2980 1344
rect 2892 1296 2900 1304
rect 2908 1176 2916 1184
rect 2876 1136 2884 1144
rect 2924 1116 2932 1124
rect 2876 1096 2884 1104
rect 2908 1096 2916 1104
rect 2860 1076 2868 1084
rect 2956 1076 2964 1084
rect 2876 1056 2884 1064
rect 2844 936 2852 944
rect 2924 1036 2932 1044
rect 2892 1016 2900 1024
rect 2892 996 2900 1004
rect 2876 956 2884 964
rect 3036 1116 3044 1124
rect 3004 976 3012 984
rect 2988 956 2996 964
rect 3020 956 3028 964
rect 2892 936 2900 944
rect 2828 916 2836 924
rect 2876 916 2884 924
rect 2988 916 2996 924
rect 2796 896 2804 904
rect 2924 896 2932 904
rect 2988 856 2996 864
rect 2828 816 2836 824
rect 2908 796 2916 804
rect 2812 696 2820 704
rect 2812 656 2820 664
rect 2876 696 2884 704
rect 2844 676 2852 684
rect 2876 676 2884 684
rect 2892 676 2900 684
rect 2828 636 2836 644
rect 2828 596 2836 604
rect 2892 576 2900 584
rect 2860 516 2868 524
rect 2748 476 2756 484
rect 2716 456 2724 464
rect 2764 436 2772 444
rect 2652 236 2660 244
rect 2572 136 2580 144
rect 2620 136 2628 144
rect 2668 156 2676 164
rect 2764 416 2772 424
rect 2748 256 2756 264
rect 2860 476 2868 484
rect 2780 376 2788 384
rect 2780 356 2788 364
rect 2812 356 2820 364
rect 2940 696 2948 704
rect 2956 696 2964 704
rect 2924 516 2932 524
rect 2876 416 2884 424
rect 2860 376 2868 384
rect 2844 356 2852 364
rect 2812 256 2820 264
rect 2796 236 2804 244
rect 2780 156 2788 164
rect 2700 136 2708 144
rect 2940 336 2948 344
rect 2908 276 2916 284
rect 2876 236 2884 244
rect 2892 216 2900 224
rect 2924 216 2932 224
rect 3004 656 3012 664
rect 2988 540 2996 544
rect 2988 536 2996 540
rect 2972 516 2980 524
rect 2988 496 2996 504
rect 3036 496 3044 504
rect 3036 296 3044 304
rect 2604 116 2612 124
rect 2732 116 2740 124
rect 2540 96 2548 104
rect 2636 96 2644 104
rect 3036 96 3044 104
rect 2364 16 2372 24
rect 2428 16 2436 24
rect 2476 16 2484 24
<< metal3 >>
rect 2916 2017 2940 2023
rect 2948 2017 2972 2023
rect 738 2014 798 2016
rect 738 2006 739 2014
rect 748 2006 749 2014
rect 787 2006 788 2014
rect 797 2006 798 2014
rect 738 2004 798 2006
rect 804 1977 828 1983
rect 196 1937 860 1943
rect 2036 1937 2412 1943
rect 52 1917 76 1923
rect 516 1917 572 1923
rect 580 1917 636 1923
rect 852 1917 892 1923
rect 1028 1917 1068 1923
rect 1092 1917 1132 1923
rect 1620 1917 1692 1923
rect 1796 1917 1852 1923
rect 1876 1917 1996 1923
rect 2100 1917 2172 1923
rect 2180 1917 2268 1923
rect 2372 1917 2380 1923
rect 2404 1917 2460 1923
rect 2532 1917 2620 1923
rect 2804 1917 2828 1923
rect -35 1897 44 1903
rect 52 1897 60 1903
rect 68 1897 124 1903
rect 132 1897 332 1903
rect 340 1897 396 1903
rect 404 1897 460 1903
rect 468 1897 876 1903
rect 1364 1897 1404 1903
rect 1524 1897 1708 1903
rect 1748 1897 1852 1903
rect 1860 1897 1884 1903
rect 1988 1897 2044 1903
rect 2068 1897 2108 1903
rect 2388 1897 2412 1903
rect 2516 1897 2556 1903
rect 2580 1897 2668 1903
rect 2676 1897 2732 1903
rect 2788 1897 2828 1903
rect 2836 1897 2876 1903
rect 2884 1897 2892 1903
rect 2900 1897 2956 1903
rect 3044 1897 3075 1903
rect 100 1877 172 1883
rect 180 1877 268 1883
rect 340 1877 524 1883
rect 596 1877 700 1883
rect 1060 1877 1100 1883
rect 1684 1877 1708 1883
rect 1780 1877 1900 1883
rect 1988 1877 2188 1883
rect 2196 1877 2380 1883
rect 2452 1877 2588 1883
rect 2628 1877 2716 1883
rect 2948 1877 2988 1883
rect -35 1857 12 1863
rect 20 1857 92 1863
rect 100 1857 364 1863
rect 372 1857 444 1863
rect 525 1863 531 1876
rect 525 1857 604 1863
rect 660 1857 860 1863
rect 900 1857 940 1863
rect 948 1857 956 1863
rect 964 1857 1004 1863
rect 1220 1857 1340 1863
rect 1572 1857 1740 1863
rect 1748 1857 1788 1863
rect 1812 1857 1836 1863
rect 1876 1857 1916 1863
rect 1940 1857 2012 1863
rect 2020 1857 2156 1863
rect 2452 1857 2572 1863
rect 2612 1857 2652 1863
rect 2868 1857 2908 1863
rect 660 1837 684 1843
rect 692 1837 924 1843
rect 1668 1837 1804 1843
rect 1812 1837 1932 1843
rect 2052 1837 2355 1843
rect 2349 1824 2355 1837
rect 1172 1817 1292 1823
rect 1860 1817 1868 1823
rect 1885 1817 1932 1823
rect 516 1797 636 1803
rect 692 1797 812 1803
rect 820 1797 892 1803
rect 900 1797 956 1803
rect 1252 1797 1452 1803
rect 1885 1803 1891 1817
rect 2356 1817 2524 1823
rect 2580 1817 2732 1823
rect 2242 1814 2302 1816
rect 2242 1806 2243 1814
rect 2252 1806 2253 1814
rect 2291 1806 2292 1814
rect 2301 1806 2302 1814
rect 2242 1804 2302 1806
rect 1508 1797 1891 1803
rect 1908 1797 1964 1803
rect 1972 1797 2076 1803
rect 2084 1797 2108 1803
rect 2180 1797 2204 1803
rect 2388 1797 2492 1803
rect 2500 1797 2540 1803
rect 2564 1797 2716 1803
rect 388 1777 556 1783
rect 564 1777 819 1783
rect 813 1764 819 1777
rect 1204 1777 1244 1783
rect 1252 1777 1388 1783
rect 1716 1777 1820 1783
rect 1828 1777 2092 1783
rect 2100 1777 2796 1783
rect 164 1757 524 1763
rect 580 1757 700 1763
rect 820 1757 851 1763
rect 845 1744 851 1757
rect 1508 1757 1532 1763
rect 1540 1757 1548 1763
rect 1556 1757 1580 1763
rect 1588 1757 1612 1763
rect 1636 1757 1740 1763
rect 1876 1757 2067 1763
rect 116 1737 364 1743
rect 452 1737 828 1743
rect 852 1737 988 1743
rect 1028 1737 1100 1743
rect 1140 1737 1180 1743
rect 1188 1737 1292 1743
rect 1444 1737 1580 1743
rect 1700 1737 1788 1743
rect 2020 1737 2044 1743
rect 2061 1743 2067 1757
rect 2116 1757 2364 1763
rect 2500 1757 2572 1763
rect 2580 1757 2700 1763
rect 2804 1757 2844 1763
rect 2852 1757 2924 1763
rect 2932 1757 2988 1763
rect 2061 1737 2140 1743
rect 2148 1737 2188 1743
rect 2212 1737 2268 1743
rect 2404 1737 2444 1743
rect 2628 1737 2652 1743
rect 2701 1743 2707 1756
rect 2701 1737 2748 1743
rect 2788 1737 2812 1743
rect 2820 1737 2860 1743
rect 132 1717 220 1723
rect 324 1717 588 1723
rect 596 1717 700 1723
rect 1044 1717 1068 1723
rect 1076 1717 1132 1723
rect 1204 1717 1420 1723
rect 1476 1717 1500 1723
rect 1604 1717 1804 1723
rect 1812 1717 2044 1723
rect 2061 1717 2764 1723
rect -35 1697 12 1703
rect 244 1697 476 1703
rect 500 1697 556 1703
rect 612 1697 668 1703
rect 701 1703 707 1716
rect 701 1697 1084 1703
rect 1108 1697 1164 1703
rect 1172 1697 1180 1703
rect 1572 1697 1772 1703
rect 2061 1703 2067 1717
rect 1796 1697 2067 1703
rect 2100 1697 2108 1703
rect 2388 1697 2700 1703
rect 2724 1697 2876 1703
rect 2916 1697 2956 1703
rect 276 1677 316 1683
rect 605 1683 611 1696
rect 452 1677 611 1683
rect 644 1677 812 1683
rect 852 1677 1260 1683
rect 1364 1677 1532 1683
rect 1636 1677 1676 1683
rect 1956 1677 1996 1683
rect 2020 1677 2124 1683
rect 2148 1677 2188 1683
rect 2292 1677 2540 1683
rect 2564 1677 2668 1683
rect 292 1657 716 1663
rect 724 1657 1020 1663
rect 1044 1657 1228 1663
rect 1284 1657 1596 1663
rect 1668 1657 1692 1663
rect 1748 1657 2028 1663
rect 2228 1657 2524 1663
rect 2548 1657 2604 1663
rect 52 1637 396 1643
rect 500 1637 588 1643
rect 596 1637 1052 1643
rect 1780 1637 2076 1643
rect 2340 1637 2508 1643
rect 276 1617 652 1623
rect 820 1617 940 1623
rect 1380 1617 1836 1623
rect 1844 1617 1900 1623
rect 2036 1617 2236 1623
rect 2244 1617 2620 1623
rect 738 1614 798 1616
rect 738 1606 739 1614
rect 748 1606 749 1614
rect 787 1606 788 1614
rect 797 1606 798 1614
rect 738 1604 798 1606
rect 452 1597 572 1603
rect 916 1597 924 1603
rect 964 1597 1148 1603
rect 1373 1603 1379 1616
rect 1172 1597 1379 1603
rect 1588 1597 2140 1603
rect 2404 1597 2812 1603
rect 308 1577 348 1583
rect 356 1577 748 1583
rect 756 1577 1452 1583
rect 1501 1577 1676 1583
rect 420 1557 508 1563
rect 532 1557 556 1563
rect 685 1557 1068 1563
rect 685 1543 691 1557
rect 1124 1557 1324 1563
rect 1501 1563 1507 1577
rect 1837 1577 1948 1583
rect 1837 1564 1843 1577
rect 2068 1577 2428 1583
rect 1332 1557 1507 1563
rect 1524 1557 1708 1563
rect 1716 1557 1836 1563
rect 1924 1557 2236 1563
rect 2244 1557 2380 1563
rect 2516 1557 2684 1563
rect 404 1537 691 1543
rect 740 1537 764 1543
rect 900 1537 1100 1543
rect 1108 1537 1196 1543
rect 1380 1537 1404 1543
rect 1428 1537 1516 1543
rect 1732 1537 2124 1543
rect 2132 1537 2316 1543
rect 2324 1537 2748 1543
rect 308 1517 412 1523
rect 436 1517 524 1523
rect 580 1517 732 1523
rect 925 1517 988 1523
rect 925 1504 931 1517
rect 1028 1517 1116 1523
rect 1300 1517 1404 1523
rect 1444 1517 1756 1523
rect 1764 1517 1932 1523
rect 1940 1517 1964 1523
rect 1972 1517 2348 1523
rect 2500 1517 2572 1523
rect 2628 1517 2732 1523
rect 2740 1517 2828 1523
rect 3044 1517 3075 1523
rect 36 1497 108 1503
rect 116 1497 156 1503
rect 244 1497 284 1503
rect 388 1497 492 1503
rect 516 1497 668 1503
rect 868 1497 924 1503
rect 964 1497 972 1503
rect 980 1497 1164 1503
rect 1220 1497 1228 1503
rect 1284 1497 1500 1503
rect 1524 1497 1852 1503
rect 2020 1497 2140 1503
rect 2148 1497 2204 1503
rect 2212 1497 2444 1503
rect 2548 1497 2652 1503
rect 2692 1497 2764 1503
rect 2836 1497 2844 1503
rect 2868 1497 2908 1503
rect 2980 1497 3020 1503
rect -35 1477 12 1483
rect 20 1477 76 1483
rect 84 1477 124 1483
rect 372 1477 460 1483
rect 532 1477 556 1483
rect 596 1477 636 1483
rect 676 1477 1027 1483
rect 212 1457 380 1463
rect 468 1457 588 1463
rect 596 1457 604 1463
rect 884 1457 892 1463
rect 1021 1463 1027 1477
rect 1124 1477 1148 1483
rect 1172 1477 1212 1483
rect 1380 1477 1452 1483
rect 1460 1477 1548 1483
rect 1604 1477 1644 1483
rect 1668 1477 1676 1483
rect 1780 1477 1788 1483
rect 1892 1477 1900 1483
rect 2004 1477 2028 1483
rect 2052 1477 2092 1483
rect 2164 1477 2508 1483
rect 2532 1477 2540 1483
rect 2740 1477 2748 1483
rect 2948 1477 3075 1483
rect 1021 1457 1132 1463
rect 1188 1457 1276 1463
rect 1316 1457 1356 1463
rect 1396 1457 1564 1463
rect 1828 1457 1868 1463
rect 1924 1457 1948 1463
rect 2029 1463 2035 1476
rect 2029 1457 2188 1463
rect 2196 1457 2364 1463
rect 2420 1457 2460 1463
rect 2468 1457 2908 1463
rect 148 1437 220 1443
rect 228 1437 476 1443
rect 500 1437 620 1443
rect 628 1437 812 1443
rect 820 1437 844 1443
rect 861 1437 1020 1443
rect 100 1417 172 1423
rect 861 1423 867 1437
rect 1028 1437 1516 1443
rect 1540 1437 1644 1443
rect 1668 1437 2188 1443
rect 2221 1437 2627 1443
rect 180 1417 867 1423
rect 884 1417 956 1423
rect 964 1417 1068 1423
rect 1108 1417 1324 1423
rect 1364 1417 1612 1423
rect 1700 1417 2108 1423
rect 2221 1423 2227 1437
rect 2164 1417 2227 1423
rect 2372 1417 2492 1423
rect 2621 1423 2627 1437
rect 2644 1437 2924 1443
rect 2621 1417 2812 1423
rect 2242 1414 2302 1416
rect 2242 1406 2243 1414
rect 2252 1406 2253 1414
rect 2291 1406 2292 1414
rect 2301 1406 2302 1414
rect 2242 1404 2302 1406
rect 484 1397 604 1403
rect 916 1397 1084 1403
rect 1252 1397 1420 1403
rect 1636 1397 1660 1403
rect 1732 1397 1804 1403
rect 1860 1397 2227 1403
rect 68 1377 396 1383
rect 404 1377 492 1383
rect 500 1377 572 1383
rect 708 1377 1260 1383
rect 1300 1377 1676 1383
rect 1764 1377 1820 1383
rect 1988 1377 2028 1383
rect 2052 1377 2060 1383
rect 2221 1383 2227 1397
rect 2340 1397 2364 1403
rect 2452 1397 2620 1403
rect 2724 1397 2844 1403
rect 2852 1397 2988 1403
rect 2221 1377 2396 1383
rect 2404 1377 2444 1383
rect 2452 1377 2508 1383
rect 2548 1377 2803 1383
rect 2797 1364 2803 1377
rect 2916 1377 2940 1383
rect -35 1357 12 1363
rect 20 1357 28 1363
rect 36 1357 140 1363
rect 340 1357 716 1363
rect 948 1357 1036 1363
rect 1236 1357 1388 1363
rect 1652 1357 1740 1363
rect 1780 1357 1852 1363
rect 1860 1357 2156 1363
rect 2196 1357 2396 1363
rect 2452 1357 2556 1363
rect 2804 1357 2988 1363
rect 116 1337 172 1343
rect 180 1337 220 1343
rect 228 1337 316 1343
rect 468 1337 556 1343
rect 564 1337 620 1343
rect 836 1337 924 1343
rect 932 1337 972 1343
rect 1124 1337 1228 1343
rect 1252 1337 1452 1343
rect 1460 1337 1804 1343
rect 1876 1337 1932 1343
rect 2020 1337 2124 1343
rect 2372 1337 2412 1343
rect 2468 1337 2604 1343
rect 2612 1337 2972 1343
rect 532 1317 540 1323
rect 676 1317 876 1323
rect 916 1317 1020 1323
rect 1124 1317 1164 1323
rect 1220 1317 1276 1323
rect 1316 1317 1340 1323
rect 1364 1317 1532 1323
rect 1636 1317 1772 1323
rect 1844 1317 1964 1323
rect 2132 1317 2172 1323
rect 2212 1317 2284 1323
rect 2404 1317 2444 1323
rect 2532 1317 2668 1323
rect 2868 1317 2924 1323
rect 52 1297 156 1303
rect 180 1297 204 1303
rect 260 1297 956 1303
rect 964 1297 1052 1303
rect 1060 1297 1148 1303
rect 1332 1297 1372 1303
rect 1716 1297 2076 1303
rect 2292 1297 2716 1303
rect 2868 1297 2892 1303
rect 612 1277 812 1283
rect 996 1277 1484 1283
rect 1492 1277 2156 1283
rect 2180 1277 2572 1283
rect 2852 1277 2956 1283
rect 884 1257 1004 1263
rect 1188 1257 1884 1263
rect 1892 1257 1916 1263
rect 1924 1257 2092 1263
rect 2404 1257 2748 1263
rect 548 1237 1148 1243
rect 1268 1237 1532 1243
rect 1540 1237 1916 1243
rect 2036 1237 2204 1243
rect 68 1217 604 1223
rect 1204 1217 1228 1223
rect 1476 1217 1692 1223
rect 1700 1217 1788 1223
rect 1908 1217 2380 1223
rect 738 1214 798 1216
rect 738 1206 739 1214
rect 748 1206 749 1214
rect 787 1206 788 1214
rect 797 1206 798 1214
rect 738 1204 798 1206
rect 468 1197 684 1203
rect 852 1197 972 1203
rect 1428 1197 2476 1203
rect 2484 1197 2636 1203
rect 2644 1197 2796 1203
rect 180 1177 524 1183
rect 532 1177 908 1183
rect 1044 1177 1068 1183
rect 1604 1177 2540 1183
rect 2548 1177 2780 1183
rect 2788 1177 2908 1183
rect 372 1157 444 1163
rect 452 1157 540 1163
rect 628 1157 1196 1163
rect 1332 1157 1420 1163
rect 1444 1157 1612 1163
rect 1796 1157 1852 1163
rect 1940 1157 1964 1163
rect 2084 1157 2156 1163
rect 2260 1157 2524 1163
rect 228 1137 300 1143
rect 308 1137 1228 1143
rect 1236 1137 1356 1143
rect 1364 1137 2348 1143
rect 2356 1137 2540 1143
rect 2644 1137 2876 1143
rect -35 1117 44 1123
rect 52 1117 76 1123
rect 84 1117 188 1123
rect 196 1117 268 1123
rect 276 1117 460 1123
rect 468 1117 652 1123
rect 676 1117 732 1123
rect 740 1117 892 1123
rect 1028 1117 1452 1123
rect 1492 1117 1548 1123
rect 1556 1117 1635 1123
rect 244 1097 332 1103
rect 340 1097 636 1103
rect 644 1097 700 1103
rect 868 1097 1036 1103
rect 1092 1097 1244 1103
rect 1316 1097 1500 1103
rect 1524 1097 1612 1103
rect 1629 1103 1635 1117
rect 1828 1117 2140 1123
rect 2148 1117 2476 1123
rect 2644 1117 2732 1123
rect 2772 1117 2812 1123
rect 2932 1117 2956 1123
rect 3044 1117 3075 1123
rect 1629 1097 1724 1103
rect 1892 1097 1980 1103
rect 1988 1097 2092 1103
rect 2340 1097 2396 1103
rect 2452 1097 2476 1103
rect 2500 1097 2540 1103
rect 2612 1097 2716 1103
rect 2788 1097 2876 1103
rect 2884 1097 2908 1103
rect -35 1077 12 1083
rect 20 1077 44 1083
rect 52 1077 204 1083
rect 212 1077 236 1083
rect 244 1077 476 1083
rect 484 1077 540 1083
rect 564 1077 876 1083
rect 884 1077 1555 1083
rect 1549 1064 1555 1077
rect 1716 1077 1772 1083
rect 1796 1077 1996 1083
rect 2036 1077 2332 1083
rect 2356 1077 2412 1083
rect 2452 1077 2492 1083
rect 2516 1077 2828 1083
rect 2868 1077 2956 1083
rect 2964 1077 3075 1083
rect 308 1057 771 1063
rect 628 1037 716 1043
rect 765 1043 771 1057
rect 836 1057 908 1063
rect 1284 1057 1308 1063
rect 1332 1057 1452 1063
rect 1556 1057 2460 1063
rect 2468 1057 2700 1063
rect 2884 1057 2956 1063
rect 765 1037 1420 1043
rect 1460 1037 1788 1043
rect 1805 1037 1836 1043
rect 340 1017 428 1023
rect 596 1017 1084 1023
rect 1092 1017 1212 1023
rect 1220 1017 1292 1023
rect 1805 1023 1811 1037
rect 1860 1037 1900 1043
rect 1908 1037 2236 1043
rect 2388 1037 2412 1043
rect 2548 1037 2652 1043
rect 2660 1037 2924 1043
rect 1780 1017 1811 1023
rect 1828 1017 2028 1023
rect 2132 1017 2220 1023
rect 2372 1017 2572 1023
rect 2804 1017 2892 1023
rect 2242 1014 2302 1016
rect 2242 1006 2243 1014
rect 2252 1006 2253 1014
rect 2291 1006 2292 1014
rect 2301 1006 2302 1014
rect 2242 1004 2302 1006
rect 388 997 796 1003
rect 948 997 1100 1003
rect 1140 997 1164 1003
rect 1261 997 1548 1003
rect 68 977 364 983
rect 372 977 396 983
rect 1261 983 1267 997
rect 1588 997 1628 1003
rect 1636 997 2172 1003
rect 2596 997 2851 1003
rect 1124 977 1267 983
rect 1284 977 1932 983
rect 1940 977 2092 983
rect 2116 977 2156 983
rect 2228 977 2476 983
rect 2612 977 2636 983
rect 2845 983 2851 997
rect 2868 997 2892 1003
rect 2804 977 3004 983
rect 276 957 316 963
rect 324 957 476 963
rect 484 957 508 963
rect 1204 957 1308 963
rect 1444 957 1484 963
rect 1540 957 1612 963
rect 1620 957 1651 963
rect 132 937 188 943
rect 212 937 268 943
rect 324 937 460 943
rect 596 937 620 943
rect 628 937 652 943
rect 820 937 1052 943
rect 1140 937 1411 943
rect 116 917 332 923
rect 420 917 460 923
rect 500 917 524 923
rect 532 917 572 923
rect 612 917 668 923
rect 692 917 716 923
rect 852 917 915 923
rect -35 897 12 903
rect 356 897 684 903
rect 692 897 892 903
rect 909 903 915 917
rect 948 917 1020 923
rect 1044 917 1228 923
rect 1405 923 1411 937
rect 1428 937 1628 943
rect 1645 943 1651 957
rect 1748 957 1836 963
rect 1940 957 1964 963
rect 2020 957 2508 963
rect 2628 957 2652 963
rect 2676 957 2700 963
rect 2788 957 2876 963
rect 2996 957 3020 963
rect 1645 937 1804 943
rect 1908 937 1932 943
rect 2164 937 2220 943
rect 2324 937 2380 943
rect 2404 937 2428 943
rect 2580 937 2716 943
rect 2740 937 2844 943
rect 2868 937 2892 943
rect 1405 917 1548 923
rect 1556 917 1596 923
rect 1716 917 1884 923
rect 1908 917 2140 923
rect 2452 917 2508 923
rect 2628 917 2700 923
rect 2756 917 2828 923
rect 2884 917 2988 923
rect 2996 917 3020 923
rect 3028 917 3075 923
rect 909 897 956 903
rect 980 897 1292 903
rect 1348 897 1404 903
rect 1476 897 1676 903
rect 1732 897 2012 903
rect 2020 897 2204 903
rect 2404 897 2636 903
rect 2660 897 2700 903
rect 2708 897 2796 903
rect 2804 897 2924 903
rect 164 877 380 883
rect 660 877 988 883
rect 1028 877 1420 883
rect 1428 877 1516 883
rect 1588 877 1644 883
rect 1940 877 2124 883
rect 436 857 1212 863
rect 1220 857 1388 863
rect 1652 857 2044 863
rect 2052 857 2252 863
rect 2260 857 2684 863
rect 2692 857 2988 863
rect 52 837 700 843
rect 980 837 1708 843
rect 1716 837 2028 843
rect 2164 837 2547 843
rect 932 817 1036 823
rect 1060 817 1116 823
rect 1140 817 1164 823
rect 1556 817 1740 823
rect 1940 817 2268 823
rect 2541 823 2547 837
rect 2564 837 2732 843
rect 2541 817 2828 823
rect 738 814 798 816
rect 738 806 739 814
rect 748 806 749 814
rect 787 806 788 814
rect 797 806 798 814
rect 738 804 798 806
rect 1252 797 1788 803
rect 1972 797 2028 803
rect 2036 797 2092 803
rect 2308 797 2444 803
rect 2468 797 2604 803
rect 2612 797 2908 803
rect 692 777 1164 783
rect 1172 777 1612 783
rect 1620 777 1900 783
rect 1988 777 2092 783
rect 2100 777 2396 783
rect 2452 777 2828 783
rect 676 757 1180 763
rect 1188 757 1228 763
rect 1236 757 1372 763
rect 1380 757 1436 763
rect 1860 757 1900 763
rect 2148 757 2380 763
rect 2388 757 2508 763
rect 2548 757 2636 763
rect 468 737 604 743
rect 660 737 1036 743
rect 1108 737 1276 743
rect 1412 737 1564 743
rect 1684 737 1756 743
rect 1764 737 1948 743
rect 2004 737 2060 743
rect 2212 737 2460 743
rect 2468 737 2588 743
rect 100 717 188 723
rect 196 717 236 723
rect 276 717 316 723
rect 420 717 460 723
rect 740 717 908 723
rect 916 717 1052 723
rect 1364 717 1500 723
rect 1684 717 1724 723
rect 1860 717 1948 723
rect 1956 717 2124 723
rect 2212 717 2252 723
rect 2340 717 2364 723
rect 2692 717 2700 723
rect 68 697 124 703
rect 228 697 332 703
rect 356 697 636 703
rect 644 697 828 703
rect 1044 697 1132 703
rect 1396 697 1452 703
rect 1668 697 2220 703
rect 2228 697 2492 703
rect 2628 697 2748 703
rect 2820 697 2876 703
rect 2884 697 2940 703
rect -35 677 12 683
rect 20 677 92 683
rect 212 677 252 683
rect 292 677 412 683
rect 468 677 828 683
rect 845 677 972 683
rect 164 657 300 663
rect 372 657 444 663
rect 845 663 851 677
rect 1364 677 1404 683
rect 1460 677 1532 683
rect 1540 677 1548 683
rect 1732 677 1868 683
rect 1924 677 1964 683
rect 2020 677 2396 683
rect 2404 677 2668 683
rect 2676 677 2844 683
rect 2868 677 2876 683
rect 548 657 851 663
rect 884 657 956 663
rect 964 657 1004 663
rect 1092 657 1340 663
rect 1348 657 1628 663
rect 1716 657 1804 663
rect 1812 657 1852 663
rect 1924 657 1996 663
rect 2084 657 2124 663
rect 2388 657 2460 663
rect 2500 657 2652 663
rect 2660 657 2684 663
rect 2820 657 3004 663
rect 84 637 172 643
rect 301 643 307 656
rect 301 637 540 643
rect 708 637 812 643
rect 1412 637 1548 643
rect 1604 637 1756 643
rect 1828 637 1836 643
rect 1876 637 1916 643
rect 2036 637 2323 643
rect 212 617 268 623
rect 276 617 396 623
rect 404 617 428 623
rect 516 617 524 623
rect 1188 617 1500 623
rect 1860 617 1932 623
rect 2004 617 2092 623
rect 2132 617 2172 623
rect 2317 623 2323 637
rect 2340 637 2652 643
rect 2676 637 2700 643
rect 2708 637 2828 643
rect 2317 617 2572 623
rect 2242 614 2302 616
rect 2242 606 2243 614
rect 2252 606 2253 614
rect 2291 606 2292 614
rect 2301 606 2302 614
rect 2242 604 2302 606
rect 180 597 332 603
rect 340 597 556 603
rect 644 597 844 603
rect 868 597 988 603
rect 996 597 1196 603
rect 1204 597 1324 603
rect 1428 597 1708 603
rect 1780 597 1964 603
rect 2116 597 2140 603
rect 2436 597 2556 603
rect 2596 597 2828 603
rect 100 577 156 583
rect 196 577 236 583
rect 244 577 604 583
rect 612 577 940 583
rect 948 577 988 583
rect 1076 577 1244 583
rect 1300 577 1452 583
rect 1492 577 1676 583
rect 1684 577 1820 583
rect 1876 577 1900 583
rect 1972 577 2412 583
rect 2468 577 2732 583
rect 2740 577 2892 583
rect 68 557 92 563
rect 244 557 1116 563
rect 1124 557 1196 563
rect 1220 557 1260 563
rect 1316 557 1324 563
rect 1348 557 1388 563
rect 1412 557 1468 563
rect 1492 557 1532 563
rect 1556 557 1644 563
rect 1812 557 2044 563
rect 2052 557 2124 563
rect 2132 557 2188 563
rect 2196 557 2364 563
rect 2372 557 2476 563
rect 2660 557 2700 563
rect 52 537 204 543
rect 260 537 284 543
rect 324 537 611 543
rect 100 517 172 523
rect 244 517 300 523
rect 420 517 492 523
rect 605 523 611 537
rect 628 537 668 543
rect 676 537 1020 543
rect 1140 537 1676 543
rect 1700 537 1724 543
rect 1732 537 1788 543
rect 1956 537 2012 543
rect 2020 537 2060 543
rect 2116 537 2172 543
rect 2228 537 2332 543
rect 2452 537 2492 543
rect 2628 537 2636 543
rect 2644 537 2684 543
rect 2925 537 2988 543
rect 2925 524 2931 537
rect 605 517 636 523
rect 660 517 716 523
rect 836 517 892 523
rect 1012 517 1244 523
rect 1364 517 1372 523
rect 1396 517 1420 523
rect 1437 517 1564 523
rect 116 497 348 503
rect 388 497 444 503
rect 468 497 524 503
rect 740 497 860 503
rect 1245 503 1251 516
rect 1437 503 1443 517
rect 1604 517 1804 523
rect 1908 517 1964 523
rect 1972 517 2044 523
rect 2052 517 2076 523
rect 2132 517 2460 523
rect 2468 517 2476 523
rect 2612 517 2636 523
rect 2644 517 2668 523
rect 2868 517 2924 523
rect 2980 517 3020 523
rect 1245 497 1443 503
rect 1508 497 1580 503
rect 1588 497 1692 503
rect 1828 497 1852 503
rect 1876 497 2124 503
rect 2148 497 2476 503
rect 2484 497 2540 503
rect 2580 497 2732 503
rect 2996 497 3036 503
rect 100 477 204 483
rect 349 483 355 496
rect 925 483 931 496
rect 349 477 1020 483
rect 1501 483 1507 496
rect 1284 477 1507 483
rect 1540 477 1596 483
rect 1604 477 1628 483
rect 1844 477 1852 483
rect 2500 477 2748 483
rect 2804 477 2860 483
rect 148 457 572 463
rect 724 457 828 463
rect 884 457 972 463
rect 1092 457 1180 463
rect 1188 457 1564 463
rect 1620 457 1740 463
rect 1780 457 2188 463
rect 2372 457 2716 463
rect 372 437 428 443
rect 724 437 883 443
rect 388 417 508 423
rect 877 423 883 437
rect 900 437 1148 443
rect 1204 437 1820 443
rect 2100 437 2764 443
rect 877 417 940 423
rect 1924 417 2044 423
rect 2052 417 2316 423
rect 2324 417 2348 423
rect 2772 417 2876 423
rect 738 414 798 416
rect 738 406 739 414
rect 748 406 749 414
rect 787 406 788 414
rect 797 406 798 414
rect 738 404 798 406
rect 356 397 460 403
rect 964 397 1132 403
rect 1140 397 1228 403
rect 1860 397 2140 403
rect 436 377 652 383
rect 868 377 1372 383
rect 1380 377 1996 383
rect 2036 377 2092 383
rect 2212 377 2428 383
rect 2532 377 2684 383
rect 2788 377 2860 383
rect 676 357 844 363
rect 852 357 908 363
rect 1012 357 1116 363
rect 1300 357 2780 363
rect 2820 357 2844 363
rect 884 337 1036 343
rect 1284 337 1356 343
rect 1748 337 2060 343
rect 2164 337 2172 343
rect 2196 337 2396 343
rect 2404 337 2524 343
rect 2708 337 2940 343
rect -35 317 28 323
rect 36 317 60 323
rect 148 317 188 323
rect 500 317 524 323
rect 548 317 732 323
rect 740 317 892 323
rect 996 317 1292 323
rect 1316 317 1324 323
rect 1332 317 1436 323
rect 1508 317 1564 323
rect 1876 317 1916 323
rect 1924 317 1996 323
rect 2196 317 2236 323
rect 68 297 140 303
rect 164 297 236 303
rect 244 297 268 303
rect 324 297 348 303
rect 356 297 412 303
rect 484 297 620 303
rect 836 297 876 303
rect 948 297 988 303
rect 1172 297 1180 303
rect 1236 297 1772 303
rect 1780 297 2124 303
rect 2356 297 2428 303
rect 2436 297 2492 303
rect 2532 297 2572 303
rect 3044 297 3075 303
rect -35 277 76 283
rect 84 277 156 283
rect 260 277 316 283
rect 324 277 380 283
rect 420 277 508 283
rect 628 277 972 283
rect 1028 277 1052 283
rect 1092 277 1148 283
rect 1156 277 1388 283
rect 1396 277 1484 283
rect 1492 277 1724 283
rect 1812 277 1868 283
rect 2068 277 2204 283
rect 2388 277 2908 283
rect 52 257 204 263
rect 212 257 220 263
rect 228 257 236 263
rect 244 257 284 263
rect 452 257 572 263
rect 1044 257 1084 263
rect 1092 257 1164 263
rect 1188 257 1228 263
rect 1300 257 1340 263
rect 1364 257 1516 263
rect 1556 257 1596 263
rect 1636 257 1660 263
rect 1860 257 1916 263
rect 2132 257 2156 263
rect 2244 257 2364 263
rect 2532 257 2588 263
rect 2756 257 2812 263
rect 68 237 92 243
rect 493 237 684 243
rect 493 223 499 237
rect 948 237 1148 243
rect 1268 237 1564 243
rect 1597 243 1603 256
rect 1597 237 1708 243
rect 1716 237 1788 243
rect 2068 237 2652 243
rect 2804 237 2876 243
rect 276 217 499 223
rect 516 217 1100 223
rect 1140 217 1180 223
rect 1188 217 1532 223
rect 2532 217 2556 223
rect 2900 217 2924 223
rect 2242 214 2302 216
rect 2242 206 2243 214
rect 2252 206 2253 214
rect 2291 206 2292 214
rect 2301 206 2302 214
rect 2242 204 2302 206
rect 196 197 348 203
rect 404 197 844 203
rect 1156 197 1244 203
rect 1284 197 1420 203
rect 1428 197 1468 203
rect 36 177 268 183
rect 276 177 428 183
rect 484 177 524 183
rect 868 177 1324 183
rect 1332 177 1372 183
rect 2004 177 2044 183
rect 2452 177 2492 183
rect 36 157 92 163
rect 100 157 140 163
rect 196 157 243 163
rect -35 137 12 143
rect 20 137 44 143
rect 164 137 204 143
rect 237 143 243 157
rect 340 157 492 163
rect 532 157 812 163
rect 884 157 972 163
rect 1012 157 1100 163
rect 1108 157 1164 163
rect 1172 157 1212 163
rect 1748 157 1900 163
rect 1972 157 2012 163
rect 2020 157 2060 163
rect 2676 157 2780 163
rect 237 137 364 143
rect 372 137 412 143
rect 468 137 540 143
rect 628 137 732 143
rect 740 137 844 143
rect 852 137 924 143
rect 1076 137 1292 143
rect 1476 137 1500 143
rect 1508 137 1516 143
rect 1524 137 1580 143
rect 1828 137 1836 143
rect 1844 137 1948 143
rect 2068 137 2108 143
rect 2116 137 2316 143
rect 2340 137 2572 143
rect 2580 137 2620 143
rect 2628 137 2700 143
rect 180 117 236 123
rect 244 117 300 123
rect 484 117 540 123
rect 916 117 956 123
rect 964 117 1020 123
rect 1028 117 1068 123
rect 1076 117 1196 123
rect 1204 117 1228 123
rect 1364 117 1404 123
rect 1412 117 1436 123
rect 1444 117 1484 123
rect 1492 117 1532 123
rect 1540 117 1596 123
rect 1620 117 1644 123
rect 1684 117 1692 123
rect 1780 117 1820 123
rect 1924 117 1980 123
rect 1988 117 2028 123
rect 2612 117 2732 123
rect 564 97 620 103
rect 708 97 812 103
rect 820 97 892 103
rect 932 97 972 103
rect 1332 97 1372 103
rect 1380 97 1452 103
rect 1812 97 1884 103
rect 2084 97 2140 103
rect 2148 97 2188 103
rect 2196 97 2348 103
rect 2548 97 2636 103
rect 3044 97 3075 103
rect 644 77 684 83
rect 692 77 1308 83
rect 1748 17 1772 23
rect 2164 17 2364 23
rect 2372 17 2428 23
rect 2436 17 2476 23
rect 738 14 798 16
rect 738 6 739 14
rect 748 6 749 14
rect 787 6 788 14
rect 797 6 798 14
rect 738 4 798 6
<< m4contact >>
rect 740 2006 747 2014
rect 747 2006 748 2014
rect 752 2006 757 2014
rect 757 2006 759 2014
rect 759 2006 760 2014
rect 764 2006 767 2014
rect 767 2006 769 2014
rect 769 2006 772 2014
rect 776 2006 777 2014
rect 777 2006 779 2014
rect 779 2006 784 2014
rect 788 2006 789 2014
rect 789 2006 796 2014
rect 1868 1916 1876 1924
rect 2380 1916 2388 1924
rect 876 1896 884 1904
rect 268 1876 276 1884
rect 588 1876 596 1884
rect 1740 1856 1748 1864
rect 1804 1856 1812 1864
rect 1932 1856 1940 1864
rect 1292 1816 1300 1824
rect 1868 1816 1876 1824
rect 1932 1816 1940 1824
rect 2244 1806 2251 1814
rect 2251 1806 2252 1814
rect 2256 1806 2261 1814
rect 2261 1806 2263 1814
rect 2263 1806 2264 1814
rect 2268 1806 2271 1814
rect 2271 1806 2273 1814
rect 2273 1806 2276 1814
rect 2280 1806 2281 1814
rect 2281 1806 2283 1814
rect 2283 1806 2288 1814
rect 2292 1806 2293 1814
rect 2293 1806 2300 1814
rect 2540 1796 2548 1804
rect 524 1756 532 1764
rect 1100 1736 1108 1744
rect 2348 1736 2356 1744
rect 2476 1736 2484 1744
rect 2956 1736 2964 1744
rect 1804 1716 1812 1724
rect 2092 1696 2100 1704
rect 2380 1696 2388 1704
rect 2028 1656 2036 1664
rect 2060 1656 2068 1664
rect 2540 1656 2548 1664
rect 588 1636 596 1644
rect 268 1616 276 1624
rect 740 1606 747 1614
rect 747 1606 748 1614
rect 752 1606 757 1614
rect 757 1606 759 1614
rect 759 1606 760 1614
rect 764 1606 767 1614
rect 767 1606 769 1614
rect 769 1606 772 1614
rect 776 1606 777 1614
rect 777 1606 779 1614
rect 779 1606 784 1614
rect 788 1606 789 1614
rect 789 1606 796 1614
rect 908 1596 916 1604
rect 2924 1576 2932 1584
rect 2508 1556 2516 1564
rect 556 1516 564 1524
rect 1292 1516 1300 1524
rect 972 1496 980 1504
rect 1228 1496 1236 1504
rect 1516 1496 1524 1504
rect 2828 1496 2836 1504
rect 588 1456 596 1464
rect 876 1456 884 1464
rect 1676 1476 1684 1484
rect 1772 1476 1780 1484
rect 1900 1476 1908 1484
rect 2508 1476 2516 1484
rect 2540 1476 2548 1484
rect 2732 1476 2740 1484
rect 1516 1436 1524 1444
rect 2188 1436 2196 1444
rect 1100 1416 1108 1424
rect 2244 1406 2251 1414
rect 2251 1406 2252 1414
rect 2256 1406 2261 1414
rect 2261 1406 2263 1414
rect 2263 1406 2264 1414
rect 2268 1406 2271 1414
rect 2271 1406 2273 1414
rect 2273 1406 2276 1414
rect 2280 1406 2281 1414
rect 2281 1406 2283 1414
rect 2283 1406 2288 1414
rect 2292 1406 2293 1414
rect 2293 1406 2300 1414
rect 908 1396 916 1404
rect 1420 1396 1428 1404
rect 2060 1376 2068 1384
rect 2444 1376 2452 1384
rect 2188 1356 2196 1364
rect 1932 1336 1940 1344
rect 524 1316 532 1324
rect 1964 1316 1972 1324
rect 2124 1316 2132 1324
rect 2860 1316 2868 1324
rect 2924 1316 2932 1324
rect 2156 1276 2164 1284
rect 2956 1276 2964 1284
rect 2028 1236 2036 1244
rect 740 1206 747 1214
rect 747 1206 748 1214
rect 752 1206 757 1214
rect 757 1206 759 1214
rect 759 1206 760 1214
rect 764 1206 767 1214
rect 767 1206 769 1214
rect 769 1206 772 1214
rect 776 1206 777 1214
rect 777 1206 779 1214
rect 779 1206 784 1214
rect 788 1206 789 1214
rect 789 1206 796 1214
rect 460 1196 468 1204
rect 684 1196 692 1204
rect 1420 1196 1428 1204
rect 2476 1196 2484 1204
rect 2540 1176 2548 1184
rect 1228 1136 1236 1144
rect 1356 1136 1364 1144
rect 2348 1136 2356 1144
rect 2636 1136 2644 1144
rect 1452 1116 1460 1124
rect 1644 1116 1652 1124
rect 2956 1116 2964 1124
rect 2092 1096 2100 1104
rect 2444 1096 2452 1104
rect 2476 1096 2484 1104
rect 556 1076 564 1084
rect 876 1076 884 1084
rect 1708 1076 1716 1084
rect 2028 1076 2036 1084
rect 1548 1056 1556 1064
rect 2956 1056 2964 1064
rect 1420 1036 1428 1044
rect 1452 1036 1460 1044
rect 2028 1016 2036 1024
rect 2668 1016 2676 1024
rect 2892 1016 2900 1024
rect 2244 1006 2251 1014
rect 2251 1006 2252 1014
rect 2256 1006 2261 1014
rect 2261 1006 2263 1014
rect 2263 1006 2264 1014
rect 2268 1006 2271 1014
rect 2271 1006 2273 1014
rect 2273 1006 2276 1014
rect 2280 1006 2281 1014
rect 2281 1006 2283 1014
rect 2283 1006 2288 1014
rect 2292 1006 2293 1014
rect 2293 1006 2300 1014
rect 940 996 948 1004
rect 1132 996 1140 1004
rect 1932 976 1940 984
rect 2796 976 2804 984
rect 2860 996 2868 1004
rect 972 956 980 964
rect 460 936 468 944
rect 588 936 596 944
rect 1420 936 1428 944
rect 1740 956 1748 964
rect 1964 956 1972 964
rect 2860 936 2868 944
rect 1676 916 1684 924
rect 3020 916 3028 924
rect 652 876 660 884
rect 1932 876 1940 884
rect 2124 876 2132 884
rect 1644 856 1652 864
rect 972 836 980 844
rect 1708 836 1716 844
rect 2156 836 2164 844
rect 1132 816 1140 824
rect 2732 836 2740 844
rect 740 806 747 814
rect 747 806 748 814
rect 752 806 757 814
rect 757 806 759 814
rect 759 806 760 814
rect 764 806 767 814
rect 767 806 769 814
rect 769 806 772 814
rect 776 806 777 814
rect 777 806 779 814
rect 779 806 784 814
rect 788 806 789 814
rect 789 806 796 814
rect 1964 796 1972 804
rect 2028 796 2036 804
rect 684 776 692 784
rect 1164 776 1172 784
rect 1900 776 1908 784
rect 2828 776 2836 784
rect 460 736 468 744
rect 1100 736 1108 744
rect 236 716 244 724
rect 1676 716 1684 724
rect 2700 716 2708 724
rect 332 696 340 704
rect 2956 696 2964 704
rect 1452 676 1460 684
rect 1548 676 1556 684
rect 2668 676 2676 684
rect 2860 676 2868 684
rect 2892 676 2900 684
rect 1804 656 1812 664
rect 1836 636 1844 644
rect 524 616 532 624
rect 1932 616 1940 624
rect 2124 616 2132 624
rect 2244 606 2251 614
rect 2251 606 2252 614
rect 2256 606 2261 614
rect 2261 606 2263 614
rect 2263 606 2264 614
rect 2268 606 2271 614
rect 2271 606 2273 614
rect 2273 606 2276 614
rect 2280 606 2281 614
rect 2281 606 2283 614
rect 2283 606 2288 614
rect 2292 606 2293 614
rect 2293 606 2300 614
rect 1324 556 1332 564
rect 1388 556 1396 564
rect 1772 556 1780 564
rect 236 516 244 524
rect 332 516 340 524
rect 1676 536 1684 544
rect 1356 516 1364 524
rect 1388 516 1396 524
rect 524 496 532 504
rect 876 496 884 504
rect 2476 516 2484 524
rect 2636 516 2644 524
rect 3020 516 3028 524
rect 1452 496 1460 504
rect 2124 496 2132 504
rect 1836 476 1844 484
rect 2796 476 2804 484
rect 972 456 980 464
rect 940 416 948 424
rect 740 406 747 414
rect 747 406 748 414
rect 752 406 757 414
rect 757 406 759 414
rect 759 406 760 414
rect 764 406 767 414
rect 767 406 769 414
rect 769 406 772 414
rect 776 406 777 414
rect 777 406 779 414
rect 779 406 784 414
rect 788 406 789 414
rect 789 406 796 414
rect 460 396 468 404
rect 652 376 660 384
rect 2028 376 2036 384
rect 1292 356 1300 364
rect 2156 336 2164 344
rect 2700 336 2708 344
rect 1292 316 1300 324
rect 1324 316 1332 324
rect 1164 296 1172 304
rect 1804 276 1812 284
rect 1100 216 1108 224
rect 2244 206 2251 214
rect 2251 206 2252 214
rect 2256 206 2261 214
rect 2261 206 2263 214
rect 2263 206 2264 214
rect 2268 206 2271 214
rect 2271 206 2273 214
rect 2273 206 2276 214
rect 2280 206 2281 214
rect 2281 206 2283 214
rect 2283 206 2288 214
rect 2292 206 2293 214
rect 2293 206 2300 214
rect 268 176 276 184
rect 1676 116 1684 124
rect 268 96 276 104
rect 740 6 747 14
rect 747 6 748 14
rect 752 6 757 14
rect 757 6 759 14
rect 759 6 760 14
rect 764 6 767 14
rect 767 6 769 14
rect 769 6 772 14
rect 776 6 777 14
rect 777 6 779 14
rect 779 6 784 14
rect 788 6 789 14
rect 789 6 796 14
<< metal4 >>
rect 736 2014 800 2016
rect 736 2006 740 2014
rect 748 2006 752 2014
rect 760 2006 764 2014
rect 772 2006 776 2014
rect 784 2006 788 2014
rect 796 2006 800 2014
rect 266 1884 278 1886
rect 266 1876 268 1884
rect 276 1876 278 1884
rect 266 1624 278 1876
rect 586 1884 598 1886
rect 586 1876 588 1884
rect 596 1876 598 1884
rect 266 1616 268 1624
rect 276 1616 278 1624
rect 266 1614 278 1616
rect 522 1764 534 1766
rect 522 1756 524 1764
rect 532 1756 534 1764
rect 522 1324 534 1756
rect 586 1644 598 1876
rect 586 1636 588 1644
rect 596 1636 598 1644
rect 586 1634 598 1636
rect 736 1614 800 2006
rect 1866 1924 1878 1926
rect 1866 1916 1868 1924
rect 1876 1916 1878 1924
rect 736 1606 740 1614
rect 748 1606 752 1614
rect 760 1606 764 1614
rect 772 1606 776 1614
rect 784 1606 788 1614
rect 796 1606 800 1614
rect 522 1316 524 1324
rect 532 1316 534 1324
rect 522 1314 534 1316
rect 554 1524 566 1526
rect 554 1516 556 1524
rect 564 1516 566 1524
rect 458 1204 470 1206
rect 458 1196 460 1204
rect 468 1196 470 1204
rect 458 944 470 1196
rect 554 1084 566 1516
rect 554 1076 556 1084
rect 564 1076 566 1084
rect 554 1074 566 1076
rect 586 1464 598 1466
rect 586 1456 588 1464
rect 596 1456 598 1464
rect 458 936 460 944
rect 468 936 470 944
rect 458 934 470 936
rect 586 944 598 1456
rect 736 1214 800 1606
rect 874 1904 886 1906
rect 874 1896 876 1904
rect 884 1896 886 1904
rect 874 1464 886 1896
rect 1738 1864 1750 1866
rect 1738 1856 1740 1864
rect 1748 1856 1750 1864
rect 1290 1824 1302 1826
rect 1290 1816 1292 1824
rect 1300 1816 1302 1824
rect 1098 1744 1110 1746
rect 1098 1736 1100 1744
rect 1108 1736 1110 1744
rect 874 1456 876 1464
rect 884 1456 886 1464
rect 874 1454 886 1456
rect 906 1604 918 1606
rect 906 1596 908 1604
rect 916 1596 918 1604
rect 906 1404 918 1596
rect 906 1396 908 1404
rect 916 1396 918 1404
rect 906 1394 918 1396
rect 970 1504 982 1506
rect 970 1496 972 1504
rect 980 1496 982 1504
rect 736 1206 740 1214
rect 748 1206 752 1214
rect 760 1206 764 1214
rect 772 1206 776 1214
rect 784 1206 788 1214
rect 796 1206 800 1214
rect 586 936 588 944
rect 596 936 598 944
rect 586 934 598 936
rect 682 1204 694 1206
rect 682 1196 684 1204
rect 692 1196 694 1204
rect 650 884 662 886
rect 650 876 652 884
rect 660 876 662 884
rect 458 744 470 746
rect 458 736 460 744
rect 468 736 470 744
rect 234 724 246 726
rect 234 716 236 724
rect 244 716 246 724
rect 234 524 246 716
rect 234 516 236 524
rect 244 516 246 524
rect 234 514 246 516
rect 330 704 342 706
rect 330 696 332 704
rect 340 696 342 704
rect 330 524 342 696
rect 330 516 332 524
rect 340 516 342 524
rect 330 514 342 516
rect 458 404 470 736
rect 522 624 534 626
rect 522 616 524 624
rect 532 616 534 624
rect 522 504 534 616
rect 522 496 524 504
rect 532 496 534 504
rect 522 494 534 496
rect 458 396 460 404
rect 468 396 470 404
rect 458 394 470 396
rect 650 384 662 876
rect 682 784 694 1196
rect 682 776 684 784
rect 692 776 694 784
rect 682 774 694 776
rect 736 814 800 1206
rect 736 806 740 814
rect 748 806 752 814
rect 760 806 764 814
rect 772 806 776 814
rect 784 806 788 814
rect 796 806 800 814
rect 650 376 652 384
rect 660 376 662 384
rect 650 374 662 376
rect 736 414 800 806
rect 874 1084 886 1086
rect 874 1076 876 1084
rect 884 1076 886 1084
rect 874 504 886 1076
rect 874 496 876 504
rect 884 496 886 504
rect 874 494 886 496
rect 938 1004 950 1006
rect 938 996 940 1004
rect 948 996 950 1004
rect 938 424 950 996
rect 970 964 982 1496
rect 1098 1424 1110 1736
rect 1290 1524 1302 1816
rect 1290 1516 1292 1524
rect 1300 1516 1302 1524
rect 1290 1514 1302 1516
rect 1098 1416 1100 1424
rect 1108 1416 1110 1424
rect 1098 1414 1110 1416
rect 1226 1504 1238 1506
rect 1226 1496 1228 1504
rect 1236 1496 1238 1504
rect 1226 1144 1238 1496
rect 1514 1504 1526 1506
rect 1514 1496 1516 1504
rect 1524 1496 1526 1504
rect 1514 1444 1526 1496
rect 1514 1436 1516 1444
rect 1524 1436 1526 1444
rect 1514 1434 1526 1436
rect 1674 1484 1686 1486
rect 1674 1476 1676 1484
rect 1684 1476 1686 1484
rect 1418 1404 1430 1406
rect 1418 1396 1420 1404
rect 1428 1396 1430 1404
rect 1418 1204 1430 1396
rect 1418 1196 1420 1204
rect 1428 1196 1430 1204
rect 1226 1136 1228 1144
rect 1236 1136 1238 1144
rect 1226 1134 1238 1136
rect 1354 1144 1366 1146
rect 1354 1136 1356 1144
rect 1364 1136 1366 1144
rect 970 956 972 964
rect 980 956 982 964
rect 970 954 982 956
rect 1130 1004 1142 1006
rect 1130 996 1132 1004
rect 1140 996 1142 1004
rect 970 844 982 846
rect 970 836 972 844
rect 980 836 982 844
rect 970 464 982 836
rect 1130 824 1142 996
rect 1130 816 1132 824
rect 1140 816 1142 824
rect 1130 814 1142 816
rect 1162 784 1174 786
rect 1162 776 1164 784
rect 1172 776 1174 784
rect 970 456 972 464
rect 980 456 982 464
rect 970 454 982 456
rect 1098 744 1110 746
rect 1098 736 1100 744
rect 1108 736 1110 744
rect 938 416 940 424
rect 948 416 950 424
rect 938 414 950 416
rect 736 406 740 414
rect 748 406 752 414
rect 760 406 764 414
rect 772 406 776 414
rect 784 406 788 414
rect 796 406 800 414
rect 266 184 278 186
rect 266 176 268 184
rect 276 176 278 184
rect 266 104 278 176
rect 266 96 268 104
rect 276 96 278 104
rect 266 94 278 96
rect 736 14 800 406
rect 1098 224 1110 736
rect 1162 304 1174 776
rect 1322 564 1334 566
rect 1322 556 1324 564
rect 1332 556 1334 564
rect 1290 364 1302 366
rect 1290 356 1292 364
rect 1300 356 1302 364
rect 1290 324 1302 356
rect 1290 316 1292 324
rect 1300 316 1302 324
rect 1290 314 1302 316
rect 1322 324 1334 556
rect 1354 524 1366 1136
rect 1418 1044 1430 1196
rect 1418 1036 1420 1044
rect 1428 1036 1430 1044
rect 1418 944 1430 1036
rect 1450 1124 1462 1126
rect 1450 1116 1452 1124
rect 1460 1116 1462 1124
rect 1450 1044 1462 1116
rect 1642 1124 1654 1126
rect 1642 1116 1644 1124
rect 1652 1116 1654 1124
rect 1450 1036 1452 1044
rect 1460 1036 1462 1044
rect 1450 1034 1462 1036
rect 1546 1064 1558 1066
rect 1546 1056 1548 1064
rect 1556 1056 1558 1064
rect 1418 936 1420 944
rect 1428 936 1430 944
rect 1418 934 1430 936
rect 1450 684 1462 686
rect 1450 676 1452 684
rect 1460 676 1462 684
rect 1354 516 1356 524
rect 1364 516 1366 524
rect 1354 514 1366 516
rect 1386 564 1398 566
rect 1386 556 1388 564
rect 1396 556 1398 564
rect 1386 524 1398 556
rect 1386 516 1388 524
rect 1396 516 1398 524
rect 1386 514 1398 516
rect 1450 504 1462 676
rect 1546 684 1558 1056
rect 1642 864 1654 1116
rect 1674 924 1686 1476
rect 1674 916 1676 924
rect 1684 916 1686 924
rect 1674 914 1686 916
rect 1706 1084 1718 1086
rect 1706 1076 1708 1084
rect 1716 1076 1718 1084
rect 1642 856 1644 864
rect 1652 856 1654 864
rect 1642 854 1654 856
rect 1706 844 1718 1076
rect 1738 964 1750 1856
rect 1802 1864 1814 1866
rect 1802 1856 1804 1864
rect 1812 1856 1814 1864
rect 1802 1724 1814 1856
rect 1866 1824 1878 1916
rect 1866 1816 1868 1824
rect 1876 1816 1878 1824
rect 1866 1814 1878 1816
rect 1930 1864 1942 1866
rect 1930 1856 1932 1864
rect 1940 1856 1942 1864
rect 1930 1824 1942 1856
rect 1930 1816 1932 1824
rect 1940 1816 1942 1824
rect 1930 1814 1942 1816
rect 2240 1814 2304 2016
rect 1802 1716 1804 1724
rect 1812 1716 1814 1724
rect 1802 1714 1814 1716
rect 2240 1806 2244 1814
rect 2252 1806 2256 1814
rect 2264 1806 2268 1814
rect 2276 1806 2280 1814
rect 2288 1806 2292 1814
rect 2300 1806 2304 1814
rect 2090 1704 2102 1706
rect 2090 1696 2092 1704
rect 2100 1696 2102 1704
rect 2026 1664 2038 1666
rect 2026 1656 2028 1664
rect 2036 1656 2038 1664
rect 1738 956 1740 964
rect 1748 956 1750 964
rect 1738 954 1750 956
rect 1770 1484 1782 1486
rect 1770 1476 1772 1484
rect 1780 1476 1782 1484
rect 1706 836 1708 844
rect 1716 836 1718 844
rect 1706 834 1718 836
rect 1546 676 1548 684
rect 1556 676 1558 684
rect 1546 674 1558 676
rect 1674 724 1686 726
rect 1674 716 1676 724
rect 1684 716 1686 724
rect 1450 496 1452 504
rect 1460 496 1462 504
rect 1450 494 1462 496
rect 1674 544 1686 716
rect 1770 564 1782 1476
rect 1898 1484 1910 1486
rect 1898 1476 1900 1484
rect 1908 1476 1910 1484
rect 1898 784 1910 1476
rect 1930 1344 1942 1346
rect 1930 1336 1932 1344
rect 1940 1336 1942 1344
rect 1930 984 1942 1336
rect 1930 976 1932 984
rect 1940 976 1942 984
rect 1930 974 1942 976
rect 1962 1324 1974 1326
rect 1962 1316 1964 1324
rect 1972 1316 1974 1324
rect 1962 964 1974 1316
rect 2026 1244 2038 1656
rect 2058 1664 2070 1666
rect 2058 1656 2060 1664
rect 2068 1656 2070 1664
rect 2058 1384 2070 1656
rect 2058 1376 2060 1384
rect 2068 1376 2070 1384
rect 2058 1374 2070 1376
rect 2026 1236 2028 1244
rect 2036 1236 2038 1244
rect 2026 1234 2038 1236
rect 2090 1104 2102 1696
rect 2186 1444 2198 1446
rect 2186 1436 2188 1444
rect 2196 1436 2198 1444
rect 2186 1364 2198 1436
rect 2186 1356 2188 1364
rect 2196 1356 2198 1364
rect 2186 1354 2198 1356
rect 2240 1414 2304 1806
rect 2378 1924 2390 1926
rect 2378 1916 2380 1924
rect 2388 1916 2390 1924
rect 2240 1406 2244 1414
rect 2252 1406 2256 1414
rect 2264 1406 2268 1414
rect 2276 1406 2280 1414
rect 2288 1406 2292 1414
rect 2300 1406 2304 1414
rect 2090 1096 2092 1104
rect 2100 1096 2102 1104
rect 2090 1094 2102 1096
rect 2122 1324 2134 1326
rect 2122 1316 2124 1324
rect 2132 1316 2134 1324
rect 2026 1084 2038 1086
rect 2026 1076 2028 1084
rect 2036 1076 2038 1084
rect 2026 1024 2038 1076
rect 2026 1016 2028 1024
rect 2036 1016 2038 1024
rect 2026 1014 2038 1016
rect 1962 956 1964 964
rect 1972 956 1974 964
rect 1898 776 1900 784
rect 1908 776 1910 784
rect 1898 774 1910 776
rect 1930 884 1942 886
rect 1930 876 1932 884
rect 1940 876 1942 884
rect 1770 556 1772 564
rect 1780 556 1782 564
rect 1770 554 1782 556
rect 1802 664 1814 666
rect 1802 656 1804 664
rect 1812 656 1814 664
rect 1674 536 1676 544
rect 1684 536 1686 544
rect 1322 316 1324 324
rect 1332 316 1334 324
rect 1322 314 1334 316
rect 1162 296 1164 304
rect 1172 296 1174 304
rect 1162 294 1174 296
rect 1098 216 1100 224
rect 1108 216 1110 224
rect 1098 214 1110 216
rect 1674 124 1686 536
rect 1802 284 1814 656
rect 1834 644 1846 646
rect 1834 636 1836 644
rect 1844 636 1846 644
rect 1834 484 1846 636
rect 1930 624 1942 876
rect 1962 804 1974 956
rect 2122 884 2134 1316
rect 2122 876 2124 884
rect 2132 876 2134 884
rect 2122 874 2134 876
rect 2154 1284 2166 1286
rect 2154 1276 2156 1284
rect 2164 1276 2166 1284
rect 2154 844 2166 1276
rect 2154 836 2156 844
rect 2164 836 2166 844
rect 1962 796 1964 804
rect 1972 796 1974 804
rect 1962 794 1974 796
rect 2026 804 2038 806
rect 2026 796 2028 804
rect 2036 796 2038 804
rect 1930 616 1932 624
rect 1940 616 1942 624
rect 1930 614 1942 616
rect 1834 476 1836 484
rect 1844 476 1846 484
rect 1834 474 1846 476
rect 2026 384 2038 796
rect 2122 624 2134 626
rect 2122 616 2124 624
rect 2132 616 2134 624
rect 2122 504 2134 616
rect 2122 496 2124 504
rect 2132 496 2134 504
rect 2122 494 2134 496
rect 2026 376 2028 384
rect 2036 376 2038 384
rect 2026 374 2038 376
rect 2154 344 2166 836
rect 2154 336 2156 344
rect 2164 336 2166 344
rect 2154 334 2166 336
rect 2240 1014 2304 1406
rect 2346 1744 2358 1746
rect 2346 1736 2348 1744
rect 2356 1736 2358 1744
rect 2346 1144 2358 1736
rect 2378 1704 2390 1916
rect 2538 1804 2550 1806
rect 2538 1796 2540 1804
rect 2548 1796 2550 1804
rect 2378 1696 2380 1704
rect 2388 1696 2390 1704
rect 2378 1694 2390 1696
rect 2474 1744 2486 1746
rect 2474 1736 2476 1744
rect 2484 1736 2486 1744
rect 2346 1136 2348 1144
rect 2356 1136 2358 1144
rect 2346 1134 2358 1136
rect 2442 1384 2454 1386
rect 2442 1376 2444 1384
rect 2452 1376 2454 1384
rect 2442 1104 2454 1376
rect 2474 1204 2486 1736
rect 2538 1664 2550 1796
rect 2538 1656 2540 1664
rect 2548 1656 2550 1664
rect 2538 1654 2550 1656
rect 2954 1744 2966 1746
rect 2954 1736 2956 1744
rect 2964 1736 2966 1744
rect 2922 1584 2934 1586
rect 2922 1576 2924 1584
rect 2932 1576 2934 1584
rect 2506 1564 2518 1566
rect 2506 1556 2508 1564
rect 2516 1556 2518 1564
rect 2506 1484 2518 1556
rect 2826 1504 2838 1506
rect 2826 1496 2828 1504
rect 2836 1496 2838 1504
rect 2506 1476 2508 1484
rect 2516 1476 2518 1484
rect 2506 1474 2518 1476
rect 2538 1484 2550 1486
rect 2538 1476 2540 1484
rect 2548 1476 2550 1484
rect 2474 1196 2476 1204
rect 2484 1196 2486 1204
rect 2474 1194 2486 1196
rect 2538 1184 2550 1476
rect 2538 1176 2540 1184
rect 2548 1176 2550 1184
rect 2538 1174 2550 1176
rect 2730 1484 2742 1486
rect 2730 1476 2732 1484
rect 2740 1476 2742 1484
rect 2634 1144 2646 1146
rect 2634 1136 2636 1144
rect 2644 1136 2646 1144
rect 2442 1096 2444 1104
rect 2452 1096 2454 1104
rect 2442 1094 2454 1096
rect 2474 1104 2486 1106
rect 2474 1096 2476 1104
rect 2484 1096 2486 1104
rect 2240 1006 2244 1014
rect 2252 1006 2256 1014
rect 2264 1006 2268 1014
rect 2276 1006 2280 1014
rect 2288 1006 2292 1014
rect 2300 1006 2304 1014
rect 2240 614 2304 1006
rect 2240 606 2244 614
rect 2252 606 2256 614
rect 2264 606 2268 614
rect 2276 606 2280 614
rect 2288 606 2292 614
rect 2300 606 2304 614
rect 1802 276 1804 284
rect 1812 276 1814 284
rect 1802 274 1814 276
rect 1674 116 1676 124
rect 1684 116 1686 124
rect 1674 114 1686 116
rect 2240 214 2304 606
rect 2474 524 2486 1096
rect 2474 516 2476 524
rect 2484 516 2486 524
rect 2474 514 2486 516
rect 2634 524 2646 1136
rect 2666 1024 2678 1026
rect 2666 1016 2668 1024
rect 2676 1016 2678 1024
rect 2666 684 2678 1016
rect 2730 844 2742 1476
rect 2730 836 2732 844
rect 2740 836 2742 844
rect 2730 834 2742 836
rect 2794 984 2806 986
rect 2794 976 2796 984
rect 2804 976 2806 984
rect 2666 676 2668 684
rect 2676 676 2678 684
rect 2666 674 2678 676
rect 2698 724 2710 726
rect 2698 716 2700 724
rect 2708 716 2710 724
rect 2634 516 2636 524
rect 2644 516 2646 524
rect 2634 514 2646 516
rect 2698 344 2710 716
rect 2794 484 2806 976
rect 2826 784 2838 1496
rect 2858 1324 2870 1326
rect 2858 1316 2860 1324
rect 2868 1316 2870 1324
rect 2858 1004 2870 1316
rect 2922 1324 2934 1576
rect 2922 1316 2924 1324
rect 2932 1316 2934 1324
rect 2922 1314 2934 1316
rect 2954 1284 2966 1736
rect 2954 1276 2956 1284
rect 2964 1276 2966 1284
rect 2954 1274 2966 1276
rect 2954 1124 2966 1126
rect 2954 1116 2956 1124
rect 2964 1116 2966 1124
rect 2954 1064 2966 1116
rect 2954 1056 2956 1064
rect 2964 1056 2966 1064
rect 2858 996 2860 1004
rect 2868 996 2870 1004
rect 2858 994 2870 996
rect 2890 1024 2902 1026
rect 2890 1016 2892 1024
rect 2900 1016 2902 1024
rect 2826 776 2828 784
rect 2836 776 2838 784
rect 2826 774 2838 776
rect 2858 944 2870 946
rect 2858 936 2860 944
rect 2868 936 2870 944
rect 2858 684 2870 936
rect 2858 676 2860 684
rect 2868 676 2870 684
rect 2858 674 2870 676
rect 2890 684 2902 1016
rect 2954 704 2966 1056
rect 2954 696 2956 704
rect 2964 696 2966 704
rect 2954 694 2966 696
rect 3018 924 3030 926
rect 3018 916 3020 924
rect 3028 916 3030 924
rect 2890 676 2892 684
rect 2900 676 2902 684
rect 2890 674 2902 676
rect 3018 524 3030 916
rect 3018 516 3020 524
rect 3028 516 3030 524
rect 3018 514 3030 516
rect 2794 476 2796 484
rect 2804 476 2806 484
rect 2794 474 2806 476
rect 2698 336 2700 344
rect 2708 336 2710 344
rect 2698 334 2710 336
rect 2240 206 2244 214
rect 2252 206 2256 214
rect 2264 206 2268 214
rect 2276 206 2280 214
rect 2288 206 2292 214
rect 2300 206 2304 214
rect 736 6 740 14
rect 748 6 752 14
rect 760 6 764 14
rect 772 6 776 14
rect 784 6 788 14
rect 796 6 800 14
rect 736 -10 800 6
rect 2240 -10 2304 206
use INVX2  _556_
timestamp 1589549099
transform 1 0 8 0 -1 210
box -4 -6 36 206
use NAND2X1  _595_
timestamp 1589549099
transform 1 0 40 0 -1 210
box -4 -6 52 206
use NAND2X1  _596_
timestamp 1589549099
transform 1 0 88 0 -1 210
box -4 -6 52 206
use INVX1  _555_
timestamp 1589549099
transform -1 0 168 0 -1 210
box -4 -6 36 206
use OAI22X1  _558_
timestamp 1589549099
transform -1 0 88 0 1 210
box -4 -6 84 206
use NAND2X1  _597_
timestamp 1589549099
transform 1 0 88 0 1 210
box -4 -6 52 206
use OAI21X1  _826_
timestamp 1589549099
transform 1 0 136 0 1 210
box -4 -6 68 206
use NAND2X1  _629_
timestamp 1589549099
transform -1 0 216 0 -1 210
box -4 -6 52 206
use OAI21X1  _559_
timestamp 1589549099
transform 1 0 216 0 -1 210
box -4 -6 68 206
use OAI21X1  _827_
timestamp 1589549099
transform 1 0 280 0 -1 210
box -4 -6 68 206
use NOR2X1  _547_
timestamp 1589549099
transform 1 0 200 0 1 210
box -4 -6 52 206
use AND2X2  _546_
timestamp 1589549099
transform 1 0 248 0 1 210
box -4 -6 68 206
use AND2X2  _831_
timestamp 1589549099
transform 1 0 344 0 -1 210
box -4 -6 68 206
use AOI22X1  _633_
timestamp 1589549099
transform 1 0 408 0 -1 210
box -4 -6 84 206
use NOR2X1  _803_
timestamp 1589549099
transform 1 0 312 0 1 210
box -4 -6 52 206
use OAI21X1  _802_
timestamp 1589549099
transform 1 0 360 0 1 210
box -4 -6 68 206
use AOI21X1  _828_
timestamp 1589549099
transform -1 0 552 0 -1 210
box -4 -6 68 206
use NAND2X1  _632_
timestamp 1589549099
transform -1 0 600 0 -1 210
box -4 -6 52 206
use INVX1  _801_
timestamp 1589549099
transform -1 0 456 0 1 210
box -4 -6 36 206
use AOI21X1  _811_
timestamp 1589549099
transform -1 0 520 0 1 210
box -4 -6 68 206
use INVX1  _628_
timestamp 1589549099
transform -1 0 552 0 1 210
box -4 -6 36 206
use BUFX2  _994_
timestamp 1589549099
transform -1 0 600 0 1 210
box -4 -6 52 206
use INVX1  _630_
timestamp 1589549099
transform -1 0 632 0 -1 210
box -4 -6 36 206
use NAND2X1  _631_
timestamp 1589549099
transform -1 0 680 0 -1 210
box -4 -6 52 206
use AOI21X1  _565_
timestamp 1589549099
transform 1 0 680 0 -1 210
box -4 -6 68 206
use INVX1  _812_
timestamp 1589549099
transform -1 0 632 0 1 210
box -4 -6 36 206
use BUFX2  _993_
timestamp 1589549099
transform -1 0 680 0 1 210
box -4 -6 52 206
use OAI21X1  _566_
timestamp 1589549099
transform -1 0 744 0 1 210
box -4 -6 68 206
use FILL  SFILL7440x2100
timestamp 1589549099
transform 1 0 744 0 1 210
box -4 -6 20 206
use FILL  SFILL7440x100
timestamp 1589549099
transform -1 0 760 0 -1 210
box -4 -6 20 206
use FILL  SFILL7920x2100
timestamp 1589549099
transform 1 0 792 0 1 210
box -4 -6 20 206
use FILL  SFILL7760x2100
timestamp 1589549099
transform 1 0 776 0 1 210
box -4 -6 20 206
use FILL  SFILL7600x2100
timestamp 1589549099
transform 1 0 760 0 1 210
box -4 -6 20 206
use FILL  SFILL7920x100
timestamp 1589549099
transform -1 0 808 0 -1 210
box -4 -6 20 206
use FILL  SFILL7760x100
timestamp 1589549099
transform -1 0 792 0 -1 210
box -4 -6 20 206
use FILL  SFILL7600x100
timestamp 1589549099
transform -1 0 776 0 -1 210
box -4 -6 20 206
use INVX1  _792_
timestamp 1589549099
transform 1 0 808 0 1 210
box -4 -6 36 206
use OAI21X1  _789_
timestamp 1589549099
transform -1 0 872 0 -1 210
box -4 -6 68 206
use NAND2X1  _564_
timestamp 1589549099
transform -1 0 920 0 -1 210
box -4 -6 52 206
use NOR2X1  _561_
timestamp 1589549099
transform -1 0 968 0 -1 210
box -4 -6 52 206
use OAI21X1  _832_
timestamp 1589549099
transform -1 0 904 0 1 210
box -4 -6 68 206
use NOR2X1  _979_
timestamp 1589549099
transform -1 0 952 0 1 210
box -4 -6 52 206
use NAND3X1  _980_
timestamp 1589549099
transform -1 0 1016 0 1 210
box -4 -6 68 206
use INVX1  _560_
timestamp 1589549099
transform -1 0 1000 0 -1 210
box -4 -6 36 206
use OR2X2  _599_
timestamp 1589549099
transform 1 0 1000 0 -1 210
box -4 -6 68 206
use NAND2X1  _598_
timestamp 1589549099
transform -1 0 1112 0 -1 210
box -4 -6 52 206
use AOI22X1  _603_
timestamp 1589549099
transform 1 0 1016 0 1 210
box -4 -6 84 206
use OAI21X1  _781_
timestamp 1589549099
transform -1 0 1160 0 1 210
box -4 -6 68 206
use BUFX2  _992_
timestamp 1589549099
transform -1 0 1160 0 -1 210
box -4 -6 52 206
use NOR2X1  _550_
timestamp 1589549099
transform 1 0 1160 0 -1 210
box -4 -6 52 206
use AND2X2  _549_
timestamp 1589549099
transform 1 0 1208 0 -1 210
box -4 -6 68 206
use OAI22X1  _770_
timestamp 1589549099
transform -1 0 1240 0 1 210
box -4 -6 84 206
use NAND2X1  _602_
timestamp 1589549099
transform -1 0 1320 0 -1 210
box -4 -6 52 206
use NOR2X1  _563_
timestamp 1589549099
transform -1 0 1368 0 -1 210
box -4 -6 52 206
use NAND2X1  _765_
timestamp 1589549099
transform -1 0 1416 0 -1 210
box -4 -6 52 206
use OAI21X1  _779_
timestamp 1589549099
transform -1 0 1304 0 1 210
box -4 -6 68 206
use AOI21X1  _766_
timestamp 1589549099
transform 1 0 1304 0 1 210
box -4 -6 68 206
use OAI21X1  _769_
timestamp 1589549099
transform -1 0 1432 0 1 210
box -4 -6 68 206
use INVX1  _601_
timestamp 1589549099
transform -1 0 1448 0 -1 210
box -4 -6 36 206
use INVX1  _562_
timestamp 1589549099
transform -1 0 1480 0 -1 210
box -4 -6 36 206
use NAND2X1  _600_
timestamp 1589549099
transform -1 0 1528 0 -1 210
box -4 -6 52 206
use OAI21X1  _768_
timestamp 1589549099
transform -1 0 1496 0 1 210
box -4 -6 68 206
use NOR2X1  _764_
timestamp 1589549099
transform -1 0 1544 0 1 210
box -4 -6 52 206
use NOR2X1  _552_
timestamp 1589549099
transform -1 0 1576 0 -1 210
box -4 -6 52 206
use AND2X2  _551_
timestamp 1589549099
transform 1 0 1576 0 -1 210
box -4 -6 68 206
use BUFX2  _991_
timestamp 1589549099
transform 1 0 1640 0 -1 210
box -4 -6 52 206
use OAI22X1  _553_
timestamp 1589549099
transform 1 0 1544 0 1 210
box -4 -6 84 206
use NOR2X1  _772_
timestamp 1589549099
transform -1 0 1672 0 1 210
box -4 -6 52 206
use BUFX2  _995_
timestamp 1589549099
transform 1 0 1688 0 -1 210
box -4 -6 52 206
use INVX1  _534_
timestamp 1589549099
transform 1 0 1736 0 -1 210
box -4 -6 36 206
use NAND2X1  _535_
timestamp 1589549099
transform -1 0 1816 0 -1 210
box -4 -6 52 206
use NOR2X1  _745_
timestamp 1589549099
transform -1 0 1720 0 1 210
box -4 -6 52 206
use OAI22X1  _759_
timestamp 1589549099
transform -1 0 1800 0 1 210
box -4 -6 84 206
use OAI21X1  _537_
timestamp 1589549099
transform 1 0 1816 0 -1 210
box -4 -6 68 206
use OAI21X1  _536_
timestamp 1589549099
transform -1 0 1944 0 -1 210
box -4 -6 68 206
use OAI21X1  _666_
timestamp 1589549099
transform -1 0 1864 0 1 210
box -4 -6 68 206
use NAND2X1  _507_
timestamp 1589549099
transform -1 0 1912 0 1 210
box -4 -6 52 206
use NAND2X1  _665_
timestamp 1589549099
transform -1 0 1960 0 1 210
box -4 -6 52 206
use INVX1  _505_
timestamp 1589549099
transform -1 0 1976 0 -1 210
box -4 -6 36 206
use NAND2X1  _504_
timestamp 1589549099
transform -1 0 2024 0 -1 210
box -4 -6 52 206
use NOR2X1  _519_
timestamp 1589549099
transform -1 0 2072 0 -1 210
box -4 -6 52 206
use NOR2X1  _935_
timestamp 1589549099
transform 1 0 1960 0 1 210
box -4 -6 52 206
use INVX1  _506_
timestamp 1589549099
transform -1 0 2040 0 1 210
box -4 -6 36 206
use OAI22X1  _919_
timestamp 1589549099
transform -1 0 2120 0 1 210
box -4 -6 84 206
use NOR2X1  _540_
timestamp 1589549099
transform 1 0 2072 0 -1 210
box -4 -6 52 206
use INVX1  _539_
timestamp 1589549099
transform -1 0 2152 0 -1 210
box -4 -6 36 206
use NAND2X1  _513_
timestamp 1589549099
transform 1 0 2152 0 -1 210
box -4 -6 52 206
use OAI21X1  _972_
timestamp 1589549099
transform 1 0 2120 0 1 210
box -4 -6 68 206
use OAI21X1  _973_
timestamp 1589549099
transform 1 0 2184 0 1 210
box -4 -6 68 206
use FILL  SFILL22480x2100
timestamp 1589549099
transform 1 0 2248 0 1 210
box -4 -6 20 206
use FILL  SFILL22480x100
timestamp 1589549099
transform -1 0 2264 0 -1 210
box -4 -6 20 206
use NAND2X1  _515_
timestamp 1589549099
transform 1 0 2200 0 -1 210
box -4 -6 52 206
use FILL  SFILL22960x2100
timestamp 1589549099
transform 1 0 2296 0 1 210
box -4 -6 20 206
use FILL  SFILL22800x2100
timestamp 1589549099
transform 1 0 2280 0 1 210
box -4 -6 20 206
use FILL  SFILL22640x2100
timestamp 1589549099
transform 1 0 2264 0 1 210
box -4 -6 20 206
use FILL  SFILL22960x100
timestamp 1589549099
transform -1 0 2312 0 -1 210
box -4 -6 20 206
use FILL  SFILL22800x100
timestamp 1589549099
transform -1 0 2296 0 -1 210
box -4 -6 20 206
use FILL  SFILL22640x100
timestamp 1589549099
transform -1 0 2280 0 -1 210
box -4 -6 20 206
use NOR2X1  _902_
timestamp 1589549099
transform 1 0 2312 0 1 210
box -4 -6 52 206
use OR2X2  _514_
timestamp 1589549099
transform -1 0 2376 0 -1 210
box -4 -6 68 206
use XOR2X1  _486_
timestamp 1589549099
transform -1 0 2488 0 -1 210
box -4 -6 116 206
use AOI21X1  _974_
timestamp 1589549099
transform -1 0 2424 0 1 210
box -4 -6 68 206
use NOR2X1  _928_
timestamp 1589549099
transform 1 0 2424 0 1 210
box -4 -6 52 206
use NAND2X1  _929_
timestamp 1589549099
transform 1 0 2488 0 -1 210
box -4 -6 52 206
use NAND2X1  _927_
timestamp 1589549099
transform -1 0 2584 0 -1 210
box -4 -6 52 206
use AOI21X1  _918_
timestamp 1589549099
transform -1 0 2648 0 -1 210
box -4 -6 68 206
use AOI21X1  _930_
timestamp 1589549099
transform 1 0 2472 0 1 210
box -4 -6 68 206
use NAND3X1  _931_
timestamp 1589549099
transform -1 0 2600 0 1 210
box -4 -6 68 206
use NAND2X1  _926_
timestamp 1589549099
transform -1 0 2648 0 1 210
box -4 -6 52 206
use OR2X2  _917_
timestamp 1589549099
transform 1 0 2648 0 -1 210
box -4 -6 68 206
use AOI21X1  _922_
timestamp 1589549099
transform 1 0 2712 0 -1 210
box -4 -6 68 206
use AOI21X1  _920_
timestamp 1589549099
transform -1 0 2712 0 1 210
box -4 -6 68 206
use NOR3X1  _982_
timestamp 1589549099
transform -1 0 2840 0 1 210
box -4 -6 132 206
use INVX1  _921_
timestamp 1589549099
transform 1 0 2776 0 -1 210
box -4 -6 36 206
use BUFX2  _1000_
timestamp 1589549099
transform 1 0 2808 0 -1 210
box -4 -6 52 206
use NOR2X1  _986_
timestamp 1589549099
transform -1 0 2904 0 -1 210
box -4 -6 52 206
use NAND3X1  _985_
timestamp 1589549099
transform 1 0 2840 0 1 210
box -4 -6 68 206
use BUFX2  _1004_
timestamp 1589549099
transform 1 0 2904 0 -1 210
box -4 -6 52 206
use INVX1  _498_
timestamp 1589549099
transform -1 0 2984 0 -1 210
box -4 -6 36 206
use BUFX2  _1001_
timestamp 1589549099
transform 1 0 2984 0 -1 210
box -4 -6 52 206
use NAND3X1  _975_
timestamp 1589549099
transform 1 0 2904 0 1 210
box -4 -6 68 206
use BUFX2  _1002_
timestamp 1589549099
transform 1 0 2968 0 1 210
box -4 -6 52 206
use FILL  FILL28880x2100
timestamp 1589549099
transform 1 0 3016 0 1 210
box -4 -6 20 206
use INVX1  _557_
timestamp 1589549099
transform 1 0 8 0 -1 610
box -4 -6 36 206
use NAND2X1  _593_
timestamp 1589549099
transform 1 0 40 0 -1 610
box -4 -6 52 206
use INVX1  _592_
timestamp 1589549099
transform 1 0 88 0 -1 610
box -4 -6 36 206
use NOR2X1  _799_
timestamp 1589549099
transform -1 0 168 0 -1 610
box -4 -6 52 206
use NAND2X1  _594_
timestamp 1589549099
transform -1 0 216 0 -1 610
box -4 -6 52 206
use OAI21X1  _819_
timestamp 1589549099
transform -1 0 280 0 -1 610
box -4 -6 68 206
use OAI22X1  _808_
timestamp 1589549099
transform -1 0 360 0 -1 610
box -4 -6 84 206
use AOI21X1  _809_
timestamp 1589549099
transform -1 0 424 0 -1 610
box -4 -6 68 206
use OAI21X1  _810_
timestamp 1589549099
transform -1 0 488 0 -1 610
box -4 -6 68 206
use OAI22X1  _548_
timestamp 1589549099
transform -1 0 568 0 -1 610
box -4 -6 84 206
use AOI21X1  _800_
timestamp 1589549099
transform -1 0 632 0 -1 610
box -4 -6 68 206
use NAND2X1  _794_
timestamp 1589549099
transform 1 0 632 0 -1 610
box -4 -6 52 206
use NAND3X1  _795_
timestamp 1589549099
transform -1 0 744 0 -1 610
box -4 -6 68 206
use NAND3X1  _798_
timestamp 1589549099
transform -1 0 872 0 -1 610
box -4 -6 68 206
use FILL  SFILL7440x4100
timestamp 1589549099
transform -1 0 760 0 -1 610
box -4 -6 20 206
use FILL  SFILL7600x4100
timestamp 1589549099
transform -1 0 776 0 -1 610
box -4 -6 20 206
use FILL  SFILL7760x4100
timestamp 1589549099
transform -1 0 792 0 -1 610
box -4 -6 20 206
use FILL  SFILL7920x4100
timestamp 1589549099
transform -1 0 808 0 -1 610
box -4 -6 20 206
use NAND3X1  _785_
timestamp 1589549099
transform 1 0 872 0 -1 610
box -4 -6 68 206
use NAND2X1  _784_
timestamp 1589549099
transform 1 0 936 0 -1 610
box -4 -6 52 206
use NOR2X1  _846_
timestamp 1589549099
transform 1 0 984 0 -1 610
box -4 -6 52 206
use OAI21X1  _793_
timestamp 1589549099
transform -1 0 1096 0 -1 610
box -4 -6 68 206
use NOR2X1  _978_
timestamp 1589549099
transform 1 0 1096 0 -1 610
box -4 -6 52 206
use NOR2X1  _554_
timestamp 1589549099
transform 1 0 1144 0 -1 610
box -4 -6 52 206
use AOI21X1  _848_
timestamp 1589549099
transform -1 0 1256 0 -1 610
box -4 -6 68 206
use AOI21X1  _778_
timestamp 1589549099
transform -1 0 1320 0 -1 610
box -4 -6 68 206
use OAI22X1  _777_
timestamp 1589549099
transform -1 0 1400 0 -1 610
box -4 -6 84 206
use OAI21X1  _776_
timestamp 1589549099
transform 1 0 1400 0 -1 610
box -4 -6 68 206
use INVX1  _767_
timestamp 1589549099
transform -1 0 1496 0 -1 610
box -4 -6 36 206
use NAND2X1  _774_
timestamp 1589549099
transform -1 0 1544 0 -1 610
box -4 -6 52 206
use NAND3X1  _847_
timestamp 1589549099
transform -1 0 1608 0 -1 610
box -4 -6 68 206
use INVX1  _763_
timestamp 1589549099
transform -1 0 1640 0 -1 610
box -4 -6 36 206
use OAI21X1  _773_
timestamp 1589549099
transform -1 0 1704 0 -1 610
box -4 -6 68 206
use INVX2  _746_
timestamp 1589549099
transform -1 0 1736 0 -1 610
box -4 -6 36 206
use AOI21X1  _760_
timestamp 1589549099
transform -1 0 1800 0 -1 610
box -4 -6 68 206
use OAI21X1  _849_
timestamp 1589549099
transform 1 0 1800 0 -1 610
box -4 -6 68 206
use AOI21X1  _945_
timestamp 1589549099
transform -1 0 1928 0 -1 610
box -4 -6 68 206
use INVX1  _943_
timestamp 1589549099
transform -1 0 1960 0 -1 610
box -4 -6 36 206
use NAND2X1  _508_
timestamp 1589549099
transform -1 0 2008 0 -1 610
box -4 -6 52 206
use NOR2X1  _509_
timestamp 1589549099
transform 1 0 2008 0 -1 610
box -4 -6 52 206
use AND2X2  _520_
timestamp 1589549099
transform 1 0 2056 0 -1 610
box -4 -6 68 206
use NOR2X1  _664_
timestamp 1589549099
transform 1 0 2120 0 -1 610
box -4 -6 52 206
use OAI22X1  _521_
timestamp 1589549099
transform 1 0 2168 0 -1 610
box -4 -6 84 206
use INVX2  _518_
timestamp 1589549099
transform 1 0 2312 0 -1 610
box -4 -6 36 206
use FILL  SFILL22480x4100
timestamp 1589549099
transform -1 0 2264 0 -1 610
box -4 -6 20 206
use FILL  SFILL22640x4100
timestamp 1589549099
transform -1 0 2280 0 -1 610
box -4 -6 20 206
use FILL  SFILL22800x4100
timestamp 1589549099
transform -1 0 2296 0 -1 610
box -4 -6 20 206
use FILL  SFILL22960x4100
timestamp 1589549099
transform -1 0 2312 0 -1 610
box -4 -6 20 206
use OAI21X1  _950_
timestamp 1589549099
transform 1 0 2344 0 -1 610
box -4 -6 68 206
use OAI22X1  _940_
timestamp 1589549099
transform -1 0 2488 0 -1 610
box -4 -6 84 206
use AOI21X1  _941_
timestamp 1589549099
transform -1 0 2552 0 -1 610
box -4 -6 68 206
use INVX1  _924_
timestamp 1589549099
transform 1 0 2552 0 -1 610
box -4 -6 36 206
use NOR2X1  _925_
timestamp 1589549099
transform 1 0 2584 0 -1 610
box -4 -6 52 206
use INVX1  _909_
timestamp 1589549099
transform -1 0 2664 0 -1 610
box -4 -6 36 206
use AOI21X1  _951_
timestamp 1589549099
transform 1 0 2664 0 -1 610
box -4 -6 68 206
use NAND3X1  _942_
timestamp 1589549099
transform 1 0 2728 0 -1 610
box -4 -6 68 206
use NOR2X1  _959_
timestamp 1589549099
transform 1 0 2792 0 -1 610
box -4 -6 52 206
use NAND3X1  _981_
timestamp 1589549099
transform -1 0 2904 0 -1 610
box -4 -6 68 206
use NAND3X1  _966_
timestamp 1589549099
transform 1 0 2904 0 -1 610
box -4 -6 68 206
use AND2X2  _965_
timestamp 1589549099
transform 1 0 2968 0 -1 610
box -4 -6 68 206
use NAND2X1  _591_
timestamp 1589549099
transform 1 0 8 0 1 610
box -4 -6 52 206
use NOR2X1  _545_
timestamp 1589549099
transform -1 0 104 0 1 610
box -4 -6 52 206
use AND2X2  _544_
timestamp 1589549099
transform 1 0 104 0 1 610
box -4 -6 68 206
use OAI22X1  _796_
timestamp 1589549099
transform -1 0 248 0 1 610
box -4 -6 84 206
use AOI21X1  _797_
timestamp 1589549099
transform -1 0 312 0 1 610
box -4 -6 68 206
use NOR2X1  _780_
timestamp 1589549099
transform -1 0 360 0 1 610
box -4 -6 52 206
use AOI21X1  _805_
timestamp 1589549099
transform -1 0 424 0 1 610
box -4 -6 68 206
use NAND3X1  _806_
timestamp 1589549099
transform 1 0 424 0 1 610
box -4 -6 68 206
use NAND2X1  _807_
timestamp 1589549099
transform -1 0 536 0 1 610
box -4 -6 52 206
use AOI21X1  _804_
timestamp 1589549099
transform -1 0 600 0 1 610
box -4 -6 68 206
use NAND2X1  _816_
timestamp 1589549099
transform -1 0 648 0 1 610
box -4 -6 52 206
use NAND2X1  _791_
timestamp 1589549099
transform 1 0 648 0 1 610
box -4 -6 52 206
use AOI21X1  _790_
timestamp 1589549099
transform -1 0 760 0 1 610
box -4 -6 68 206
use OAI21X1  _782_
timestamp 1589549099
transform -1 0 888 0 1 610
box -4 -6 68 206
use FILL  SFILL7600x6100
timestamp 1589549099
transform 1 0 760 0 1 610
box -4 -6 20 206
use FILL  SFILL7760x6100
timestamp 1589549099
transform 1 0 776 0 1 610
box -4 -6 20 206
use FILL  SFILL7920x6100
timestamp 1589549099
transform 1 0 792 0 1 610
box -4 -6 20 206
use FILL  SFILL8080x6100
timestamp 1589549099
transform 1 0 808 0 1 610
box -4 -6 20 206
use NAND3X1  _604_
timestamp 1589549099
transform -1 0 952 0 1 610
box -4 -6 68 206
use NOR2X1  _783_
timestamp 1589549099
transform 1 0 952 0 1 610
box -4 -6 52 206
use INVX1  _818_
timestamp 1589549099
transform 1 0 1000 0 1 610
box -4 -6 36 206
use OAI21X1  _821_
timestamp 1589549099
transform 1 0 1032 0 1 610
box -4 -6 68 206
use INVX1  _820_
timestamp 1589549099
transform -1 0 1128 0 1 610
box -4 -6 36 206
use NOR2X1  _817_
timestamp 1589549099
transform -1 0 1176 0 1 610
box -4 -6 52 206
use AOI21X1  _775_
timestamp 1589549099
transform -1 0 1240 0 1 610
box -4 -6 68 206
use AOI21X1  _752_
timestamp 1589549099
transform 1 0 1240 0 1 610
box -4 -6 68 206
use AOI21X1  _762_
timestamp 1589549099
transform 1 0 1304 0 1 610
box -4 -6 68 206
use AOI21X1  _755_
timestamp 1589549099
transform 1 0 1368 0 1 610
box -4 -6 68 206
use AND2X2  _771_
timestamp 1589549099
transform 1 0 1432 0 1 610
box -4 -6 68 206
use NAND2X1  _757_
timestamp 1589549099
transform -1 0 1544 0 1 610
box -4 -6 52 206
use OAI21X1  _761_
timestamp 1589549099
transform 1 0 1544 0 1 610
box -4 -6 68 206
use INVX2  _678_
timestamp 1589549099
transform 1 0 1608 0 1 610
box -4 -6 36 206
use NAND3X1  _589_
timestamp 1589549099
transform 1 0 1640 0 1 610
box -4 -6 68 206
use AOI22X1  _511_
timestamp 1589549099
transform 1 0 1704 0 1 610
box -4 -6 84 206
use INVX1  _510_
timestamp 1589549099
transform -1 0 1816 0 1 610
box -4 -6 36 206
use NOR2X1  _944_
timestamp 1589549099
transform 1 0 1816 0 1 610
box -4 -6 52 206
use AOI22X1  _934_
timestamp 1589549099
transform 1 0 1864 0 1 610
box -4 -6 84 206
use INVX1  _937_
timestamp 1589549099
transform -1 0 1976 0 1 610
box -4 -6 36 206
use OAI21X1  _936_
timestamp 1589549099
transform 1 0 1976 0 1 610
box -4 -6 68 206
use NAND3X1  _939_
timestamp 1589549099
transform -1 0 2104 0 1 610
box -4 -6 68 206
use NAND3X1  _938_
timestamp 1589549099
transform 1 0 2104 0 1 610
box -4 -6 68 206
use OAI21X1  _946_
timestamp 1589549099
transform -1 0 2232 0 1 610
box -4 -6 68 206
use NAND2X1  _908_
timestamp 1589549099
transform -1 0 2344 0 1 610
box -4 -6 52 206
use FILL  SFILL22320x6100
timestamp 1589549099
transform 1 0 2232 0 1 610
box -4 -6 20 206
use FILL  SFILL22480x6100
timestamp 1589549099
transform 1 0 2248 0 1 610
box -4 -6 20 206
use FILL  SFILL22640x6100
timestamp 1589549099
transform 1 0 2264 0 1 610
box -4 -6 20 206
use FILL  SFILL22800x6100
timestamp 1589549099
transform 1 0 2280 0 1 610
box -4 -6 20 206
use NAND3X1  _911_
timestamp 1589549099
transform -1 0 2408 0 1 610
box -4 -6 68 206
use AOI21X1  _948_
timestamp 1589549099
transform -1 0 2472 0 1 610
box -4 -6 68 206
use OR2X2  _947_
timestamp 1589549099
transform 1 0 2472 0 1 610
box -4 -6 68 206
use AND2X2  _949_
timestamp 1589549099
transform 1 0 2536 0 1 610
box -4 -6 68 206
use OAI21X1  _953_
timestamp 1589549099
transform -1 0 2664 0 1 610
box -4 -6 68 206
use AND2X2  _952_
timestamp 1589549099
transform 1 0 2664 0 1 610
box -4 -6 68 206
use OAI21X1  _958_
timestamp 1589549099
transform 1 0 2728 0 1 610
box -4 -6 68 206
use NOR2X1  _961_
timestamp 1589549099
transform 1 0 2792 0 1 610
box -4 -6 52 206
use OAI21X1  _964_
timestamp 1589549099
transform -1 0 2904 0 1 610
box -4 -6 68 206
use NOR2X1  _962_
timestamp 1589549099
transform 1 0 2904 0 1 610
box -4 -6 52 206
use NAND2X1  _963_
timestamp 1589549099
transform -1 0 3000 0 1 610
box -4 -6 52 206
use INVX1  _960_
timestamp 1589549099
transform 1 0 3000 0 1 610
box -4 -6 36 206
use BUFX2  _990_
timestamp 1589549099
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use NOR2X1  _740_
timestamp 1589549099
transform 1 0 56 0 -1 1010
box -4 -6 52 206
use NOR3X1  _741_
timestamp 1589549099
transform -1 0 232 0 -1 1010
box -4 -6 132 206
use NOR2X1  _738_
timestamp 1589549099
transform -1 0 280 0 -1 1010
box -4 -6 52 206
use NOR2X1  _739_
timestamp 1589549099
transform 1 0 280 0 -1 1010
box -4 -6 52 206
use NOR2X1  _728_
timestamp 1589549099
transform -1 0 376 0 -1 1010
box -4 -6 52 206
use OAI21X1  _742_
timestamp 1589549099
transform -1 0 440 0 -1 1010
box -4 -6 68 206
use AND2X2  _736_
timestamp 1589549099
transform -1 0 504 0 -1 1010
box -4 -6 68 206
use OAI21X1  _737_
timestamp 1589549099
transform 1 0 504 0 -1 1010
box -4 -6 68 206
use AOI21X1  _735_
timestamp 1589549099
transform -1 0 632 0 -1 1010
box -4 -6 68 206
use NAND3X1  _754_
timestamp 1589549099
transform -1 0 696 0 -1 1010
box -4 -6 68 206
use INVX1  _744_
timestamp 1589549099
transform -1 0 728 0 -1 1010
box -4 -6 36 206
use AOI21X1  _743_
timestamp 1589549099
transform -1 0 856 0 -1 1010
box -4 -6 68 206
use FILL  SFILL7280x8100
timestamp 1589549099
transform -1 0 744 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7440x8100
timestamp 1589549099
transform -1 0 760 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7600x8100
timestamp 1589549099
transform -1 0 776 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7760x8100
timestamp 1589549099
transform -1 0 792 0 -1 1010
box -4 -6 20 206
use OR2X2  _732_
timestamp 1589549099
transform -1 0 920 0 -1 1010
box -4 -6 68 206
use AOI21X1  _733_
timestamp 1589549099
transform 1 0 920 0 -1 1010
box -4 -6 68 206
use OAI21X1  _641_
timestamp 1589549099
transform -1 0 1048 0 -1 1010
box -4 -6 68 206
use NAND3X1  _977_
timestamp 1589549099
transform 1 0 1048 0 -1 1010
box -4 -6 68 206
use AOI21X1  _822_
timestamp 1589549099
transform -1 0 1176 0 -1 1010
box -4 -6 68 206
use NAND2X1  _815_
timestamp 1589549099
transform -1 0 1224 0 -1 1010
box -4 -6 52 206
use OAI21X1  _840_
timestamp 1589549099
transform 1 0 1224 0 -1 1010
box -4 -6 68 206
use OAI21X1  _750_
timestamp 1589549099
transform 1 0 1288 0 -1 1010
box -4 -6 68 206
use NAND3X1  _756_
timestamp 1589549099
transform -1 0 1416 0 -1 1010
box -4 -6 68 206
use AOI21X1  _671_
timestamp 1589549099
transform 1 0 1416 0 -1 1010
box -4 -6 68 206
use NAND2X1  _642_
timestamp 1589549099
transform 1 0 1480 0 -1 1010
box -4 -6 52 206
use OAI21X1  _824_
timestamp 1589549099
transform 1 0 1528 0 -1 1010
box -4 -6 68 206
use AOI21X1  _823_
timestamp 1589549099
transform 1 0 1592 0 -1 1010
box -4 -6 68 206
use OAI21X1  _670_
timestamp 1589549099
transform 1 0 1656 0 -1 1010
box -4 -6 68 206
use NAND3X1  _838_
timestamp 1589549099
transform -1 0 1784 0 -1 1010
box -4 -6 68 206
use AOI21X1  _843_
timestamp 1589549099
transform 1 0 1784 0 -1 1010
box -4 -6 68 206
use AOI21X1  _669_
timestamp 1589549099
transform 1 0 1848 0 -1 1010
box -4 -6 68 206
use INVX1  _667_
timestamp 1589549099
transform -1 0 1944 0 -1 1010
box -4 -6 36 206
use OAI21X1  _668_
timestamp 1589549099
transform -1 0 2008 0 -1 1010
box -4 -6 68 206
use INVX1  _538_
timestamp 1589549099
transform 1 0 2008 0 -1 1010
box -4 -6 36 206
use AOI21X1  _541_
timestamp 1589549099
transform 1 0 2040 0 -1 1010
box -4 -6 68 206
use OAI21X1  _542_
timestamp 1589549099
transform -1 0 2168 0 -1 1010
box -4 -6 68 206
use NOR2X1  _522_
timestamp 1589549099
transform -1 0 2216 0 -1 1010
box -4 -6 52 206
use NAND2X1  _517_
timestamp 1589549099
transform -1 0 2264 0 -1 1010
box -4 -6 52 206
use NOR2X1  _933_
timestamp 1589549099
transform -1 0 2376 0 -1 1010
box -4 -6 52 206
use FILL  SFILL22640x8100
timestamp 1589549099
transform -1 0 2280 0 -1 1010
box -4 -6 20 206
use FILL  SFILL22800x8100
timestamp 1589549099
transform -1 0 2296 0 -1 1010
box -4 -6 20 206
use FILL  SFILL22960x8100
timestamp 1589549099
transform -1 0 2312 0 -1 1010
box -4 -6 20 206
use FILL  SFILL23120x8100
timestamp 1589549099
transform -1 0 2328 0 -1 1010
box -4 -6 20 206
use OR2X2  _906_
timestamp 1589549099
transform 1 0 2376 0 -1 1010
box -4 -6 68 206
use NOR2X1  _907_
timestamp 1589549099
transform -1 0 2488 0 -1 1010
box -4 -6 52 206
use OAI21X1  _910_
timestamp 1589549099
transform 1 0 2488 0 -1 1010
box -4 -6 68 206
use INVX2  _758_
timestamp 1589549099
transform -1 0 2584 0 -1 1010
box -4 -6 36 206
use NAND2X1  _967_
timestamp 1589549099
transform -1 0 2632 0 -1 1010
box -4 -6 52 206
use NAND3X1  _971_
timestamp 1589549099
transform 1 0 2632 0 -1 1010
box -4 -6 68 206
use OAI21X1  _956_
timestamp 1589549099
transform 1 0 2696 0 -1 1010
box -4 -6 68 206
use AOI21X1  _957_
timestamp 1589549099
transform -1 0 2824 0 -1 1010
box -4 -6 68 206
use OAI21X1  _955_
timestamp 1589549099
transform -1 0 2888 0 -1 1010
box -4 -6 68 206
use XNOR2X1  _516_
timestamp 1589549099
transform -1 0 3000 0 -1 1010
box -4 -6 116 206
use INVX1  _861_
timestamp 1589549099
transform 1 0 3000 0 -1 1010
box -4 -6 36 206
use NOR2X1  _568_
timestamp 1589549099
transform 1 0 8 0 1 1010
box -4 -6 52 206
use AND2X2  _567_
timestamp 1589549099
transform 1 0 56 0 1 1010
box -4 -6 68 206
use OAI22X1  _581_
timestamp 1589549099
transform -1 0 200 0 1 1010
box -4 -6 84 206
use INVX2  _579_
timestamp 1589549099
transform 1 0 200 0 1 1010
box -4 -6 36 206
use NAND2X1  _605_
timestamp 1589549099
transform 1 0 232 0 1 1010
box -4 -6 52 206
use NAND2X1  _734_
timestamp 1589549099
transform 1 0 280 0 1 1010
box -4 -6 52 206
use NAND2X1  _606_
timestamp 1589549099
transform 1 0 328 0 1 1010
box -4 -6 52 206
use AOI21X1  _753_
timestamp 1589549099
transform 1 0 376 0 1 1010
box -4 -6 68 206
use INVX1  _578_
timestamp 1589549099
transform -1 0 472 0 1 1010
box -4 -6 36 206
use OAI21X1  _582_
timestamp 1589549099
transform 1 0 472 0 1 1010
box -4 -6 68 206
use OAI21X1  _749_
timestamp 1589549099
transform 1 0 536 0 1 1010
box -4 -6 68 206
use OAI21X1  _748_
timestamp 1589549099
transform -1 0 664 0 1 1010
box -4 -6 68 206
use NAND2X1  _639_
timestamp 1589549099
transform 1 0 664 0 1 1010
box -4 -6 52 206
use AND2X2  _787_
timestamp 1589549099
transform 1 0 712 0 1 1010
box -4 -6 68 206
use FILL  SFILL7760x10100
timestamp 1589549099
transform 1 0 776 0 1 1010
box -4 -6 20 206
use FILL  SFILL7920x10100
timestamp 1589549099
transform 1 0 792 0 1 1010
box -4 -6 20 206
use FILL  SFILL8080x10100
timestamp 1589549099
transform 1 0 808 0 1 1010
box -4 -6 20 206
use FILL  SFILL8240x10100
timestamp 1589549099
transform 1 0 824 0 1 1010
box -4 -6 20 206
use NAND2X1  _788_
timestamp 1589549099
transform -1 0 888 0 1 1010
box -4 -6 52 206
use AOI22X1  _640_
timestamp 1589549099
transform 1 0 888 0 1 1010
box -4 -6 84 206
use AOI21X1  _830_
timestamp 1589549099
transform 1 0 968 0 1 1010
box -4 -6 68 206
use AOI21X1  _751_
timestamp 1589549099
transform 1 0 1032 0 1 1010
box -4 -6 68 206
use AOI21X1  _584_
timestamp 1589549099
transform -1 0 1160 0 1 1010
box -4 -6 68 206
use OAI21X1  _825_
timestamp 1589549099
transform -1 0 1224 0 1 1010
box -4 -6 68 206
use NOR2X1  _655_
timestamp 1589549099
transform -1 0 1272 0 1 1010
box -4 -6 52 206
use INVX1  _656_
timestamp 1589549099
transform 1 0 1272 0 1 1010
box -4 -6 36 206
use OAI21X1  _674_
timestamp 1589549099
transform 1 0 1304 0 1 1010
box -4 -6 68 206
use INVX1  _693_
timestamp 1589549099
transform 1 0 1368 0 1 1010
box -4 -6 36 206
use NAND3X1  _694_
timestamp 1589549099
transform -1 0 1464 0 1 1010
box -4 -6 68 206
use NAND3X1  _660_
timestamp 1589549099
transform -1 0 1528 0 1 1010
box -4 -6 68 206
use OAI21X1  _585_
timestamp 1589549099
transform 1 0 1528 0 1 1010
box -4 -6 68 206
use NAND3X1  _643_
timestamp 1589549099
transform -1 0 1656 0 1 1010
box -4 -6 68 206
use NOR2X1  _590_
timestamp 1589549099
transform 1 0 1656 0 1 1010
box -4 -6 52 206
use OAI21X1  _621_
timestamp 1589549099
transform 1 0 1704 0 1 1010
box -4 -6 68 206
use OAI21X1  _833_
timestamp 1589549099
transform 1 0 1768 0 1 1010
box -4 -6 68 206
use NAND3X1  _834_
timestamp 1589549099
transform -1 0 1896 0 1 1010
box -4 -6 68 206
use NAND3X1  _512_
timestamp 1589549099
transform 1 0 1896 0 1 1010
box -4 -6 68 206
use OAI21X1  _932_
timestamp 1589549099
transform -1 0 2024 0 1 1010
box -4 -6 68 206
use OAI21X1  _866_
timestamp 1589549099
transform 1 0 2024 0 1 1010
box -4 -6 68 206
use AOI21X1  _903_
timestamp 1589549099
transform 1 0 2088 0 1 1010
box -4 -6 68 206
use AOI21X1  _543_
timestamp 1589549099
transform -1 0 2216 0 1 1010
box -4 -6 68 206
use NOR2X1  _503_
timestamp 1589549099
transform 1 0 2216 0 1 1010
box -4 -6 52 206
use AOI21X1  _845_
timestamp 1589549099
transform 1 0 2328 0 1 1010
box -4 -6 68 206
use FILL  SFILL22640x10100
timestamp 1589549099
transform 1 0 2264 0 1 1010
box -4 -6 20 206
use FILL  SFILL22800x10100
timestamp 1589549099
transform 1 0 2280 0 1 1010
box -4 -6 20 206
use FILL  SFILL22960x10100
timestamp 1589549099
transform 1 0 2296 0 1 1010
box -4 -6 20 206
use FILL  SFILL23120x10100
timestamp 1589549099
transform 1 0 2312 0 1 1010
box -4 -6 20 206
use OR2X2  _844_
timestamp 1589549099
transform 1 0 2392 0 1 1010
box -4 -6 68 206
use INVX4  _698_
timestamp 1589549099
transform -1 0 2504 0 1 1010
box -4 -6 52 206
use NAND2X1  _502_
timestamp 1589549099
transform -1 0 2552 0 1 1010
box -4 -6 52 206
use AOI21X1  _860_
timestamp 1589549099
transform 1 0 2552 0 1 1010
box -4 -6 68 206
use NAND3X1  _970_
timestamp 1589549099
transform -1 0 2680 0 1 1010
box -4 -6 68 206
use NAND2X1  _969_
timestamp 1589549099
transform 1 0 2680 0 1 1010
box -4 -6 52 206
use OAI21X1  _968_
timestamp 1589549099
transform -1 0 2792 0 1 1010
box -4 -6 68 206
use NAND2X1  _501_
timestamp 1589549099
transform 1 0 2792 0 1 1010
box -4 -6 52 206
use INVX1  _500_
timestamp 1589549099
transform -1 0 2872 0 1 1010
box -4 -6 36 206
use NOR2X1  _954_
timestamp 1589549099
transform 1 0 2872 0 1 1010
box -4 -6 52 206
use NAND2X1  _499_
timestamp 1589549099
transform -1 0 2968 0 1 1010
box -4 -6 52 206
use BUFX2  _1003_
timestamp 1589549099
transform 1 0 2968 0 1 1010
box -4 -6 52 206
use FILL  FILL28880x10100
timestamp 1589549099
transform 1 0 3016 0 1 1010
box -4 -6 20 206
use INVX1  _608_
timestamp 1589549099
transform 1 0 8 0 -1 1410
box -4 -6 36 206
use NOR2X1  _730_
timestamp 1589549099
transform -1 0 88 0 -1 1410
box -4 -6 52 206
use INVX1  _580_
timestamp 1589549099
transform 1 0 88 0 -1 1410
box -4 -6 36 206
use NAND2X1  _609_
timestamp 1589549099
transform 1 0 120 0 -1 1410
box -4 -6 52 206
use NAND2X1  _714_
timestamp 1589549099
transform 1 0 168 0 -1 1410
box -4 -6 52 206
use AOI22X1  _610_
timestamp 1589549099
transform -1 0 296 0 -1 1410
box -4 -6 84 206
use NOR3X1  _724_
timestamp 1589549099
transform 1 0 296 0 -1 1410
box -4 -6 132 206
use OAI22X1  _571_
timestamp 1589549099
transform 1 0 424 0 -1 1410
box -4 -6 84 206
use OAI21X1  _583_
timestamp 1589549099
transform -1 0 568 0 -1 1410
box -4 -6 68 206
use NOR2X1  _716_
timestamp 1589549099
transform -1 0 616 0 -1 1410
box -4 -6 52 206
use AOI21X1  _747_
timestamp 1589549099
transform -1 0 680 0 -1 1410
box -4 -6 68 206
use OR2X2  _677_
timestamp 1589549099
transform -1 0 744 0 -1 1410
box -4 -6 68 206
use AOI21X1  _731_
timestamp 1589549099
transform -1 0 872 0 -1 1410
box -4 -6 68 206
use FILL  SFILL7440x12100
timestamp 1589549099
transform -1 0 760 0 -1 1410
box -4 -6 20 206
use FILL  SFILL7600x12100
timestamp 1589549099
transform -1 0 776 0 -1 1410
box -4 -6 20 206
use FILL  SFILL7760x12100
timestamp 1589549099
transform -1 0 792 0 -1 1410
box -4 -6 20 206
use FILL  SFILL7920x12100
timestamp 1589549099
transform -1 0 808 0 -1 1410
box -4 -6 20 206
use OAI21X1  _729_
timestamp 1589549099
transform -1 0 936 0 -1 1410
box -4 -6 68 206
use NOR2X1  _637_
timestamp 1589549099
transform -1 0 984 0 -1 1410
box -4 -6 52 206
use NAND2X1  _635_
timestamp 1589549099
transform 1 0 984 0 -1 1410
box -4 -6 52 206
use OAI21X1  _638_
timestamp 1589549099
transform -1 0 1096 0 -1 1410
box -4 -6 68 206
use NOR2X1  _653_
timestamp 1589549099
transform 1 0 1096 0 -1 1410
box -4 -6 52 206
use NAND3X1  _654_
timestamp 1589549099
transform 1 0 1144 0 -1 1410
box -4 -6 68 206
use NOR2X1  _619_
timestamp 1589549099
transform 1 0 1208 0 -1 1410
box -4 -6 52 206
use OAI21X1  _689_
timestamp 1589549099
transform 1 0 1256 0 -1 1410
box -4 -6 68 206
use NOR2X1  _673_
timestamp 1589549099
transform 1 0 1320 0 -1 1410
box -4 -6 52 206
use NAND3X1  _692_
timestamp 1589549099
transform 1 0 1368 0 -1 1410
box -4 -6 68 206
use NAND3X1  _691_
timestamp 1589549099
transform 1 0 1432 0 -1 1410
box -4 -6 68 206
use NOR2X1  _659_
timestamp 1589549099
transform 1 0 1496 0 -1 1410
box -4 -6 52 206
use NOR3X1  _695_
timestamp 1589549099
transform -1 0 1672 0 -1 1410
box -4 -6 132 206
use NOR2X1  _627_
timestamp 1589549099
transform 1 0 1672 0 -1 1410
box -4 -6 52 206
use AOI21X1  _648_
timestamp 1589549099
transform -1 0 1784 0 -1 1410
box -4 -6 68 206
use AOI21X1  _620_
timestamp 1589549099
transform 1 0 1784 0 -1 1410
box -4 -6 68 206
use NAND3X1  _829_
timestamp 1589549099
transform 1 0 1848 0 -1 1410
box -4 -6 68 206
use AOI21X1  _893_
timestamp 1589549099
transform 1 0 1912 0 -1 1410
box -4 -6 68 206
use NOR2X1  _497_
timestamp 1589549099
transform 1 0 1976 0 -1 1410
box -4 -6 52 206
use INVX1  _586_
timestamp 1589549099
transform 1 0 2024 0 -1 1410
box -4 -6 36 206
use NAND2X1  _588_
timestamp 1589549099
transform 1 0 2056 0 -1 1410
box -4 -6 52 206
use INVX1  _587_
timestamp 1589549099
transform -1 0 2136 0 -1 1410
box -4 -6 36 206
use INVX2  _814_
timestamp 1589549099
transform -1 0 2168 0 -1 1410
box -4 -6 36 206
use AOI21X1  _851_
timestamp 1589549099
transform 1 0 2168 0 -1 1410
box -4 -6 68 206
use NOR2X1  _839_
timestamp 1589549099
transform -1 0 2344 0 -1 1410
box -4 -6 52 206
use FILL  SFILL22320x12100
timestamp 1589549099
transform -1 0 2248 0 -1 1410
box -4 -6 20 206
use FILL  SFILL22480x12100
timestamp 1589549099
transform -1 0 2264 0 -1 1410
box -4 -6 20 206
use FILL  SFILL22640x12100
timestamp 1589549099
transform -1 0 2280 0 -1 1410
box -4 -6 20 206
use FILL  SFILL22800x12100
timestamp 1589549099
transform -1 0 2296 0 -1 1410
box -4 -6 20 206
use AOI21X1  _855_
timestamp 1589549099
transform 1 0 2344 0 -1 1410
box -4 -6 68 206
use INVX1  _852_
timestamp 1589549099
transform 1 0 2408 0 -1 1410
box -4 -6 36 206
use NOR2X1  _853_
timestamp 1589549099
transform -1 0 2488 0 -1 1410
box -4 -6 52 206
use OAI22X1  _857_
timestamp 1589549099
transform -1 0 2568 0 -1 1410
box -4 -6 84 206
use NAND2X1  _872_
timestamp 1589549099
transform -1 0 2616 0 -1 1410
box -4 -6 52 206
use AOI21X1  _858_
timestamp 1589549099
transform 1 0 2616 0 -1 1410
box -4 -6 68 206
use OAI21X1  _859_
timestamp 1589549099
transform -1 0 2744 0 -1 1410
box -4 -6 68 206
use OAI21X1  _856_
timestamp 1589549099
transform -1 0 2808 0 -1 1410
box -4 -6 68 206
use NOR2X1  _984_
timestamp 1589549099
transform -1 0 2856 0 -1 1410
box -4 -6 52 206
use OAI21X1  _916_
timestamp 1589549099
transform -1 0 2920 0 -1 1410
box -4 -6 68 206
use NAND2X1  _913_
timestamp 1589549099
transform 1 0 2920 0 -1 1410
box -4 -6 52 206
use INVX1  _854_
timestamp 1589549099
transform 1 0 2968 0 -1 1410
box -4 -6 36 206
use FILL  FILL28720x12100
timestamp 1589549099
transform -1 0 3016 0 -1 1410
box -4 -6 20 206
use FILL  FILL28880x12100
timestamp 1589549099
transform -1 0 3032 0 -1 1410
box -4 -6 20 206
use AND2X2  _569_
timestamp 1589549099
transform 1 0 8 0 1 1410
box -4 -6 68 206
use NAND2X1  _607_
timestamp 1589549099
transform 1 0 72 0 1 1410
box -4 -6 52 206
use NOR2X1  _570_
timestamp 1589549099
transform 1 0 120 0 1 1410
box -4 -6 52 206
use NOR2X1  _725_
timestamp 1589549099
transform -1 0 216 0 1 1410
box -4 -6 52 206
use NOR3X1  _726_
timestamp 1589549099
transform -1 0 344 0 1 1410
box -4 -6 132 206
use NOR2X1  _723_
timestamp 1589549099
transform -1 0 392 0 1 1410
box -4 -6 52 206
use NAND3X1  _727_
timestamp 1589549099
transform -1 0 456 0 1 1410
box -4 -6 68 206
use NOR2X1  _720_
timestamp 1589549099
transform 1 0 456 0 1 1410
box -4 -6 52 206
use OAI21X1  _722_
timestamp 1589549099
transform 1 0 504 0 1 1410
box -4 -6 68 206
use AND2X2  _721_
timestamp 1589549099
transform -1 0 632 0 1 1410
box -4 -6 68 206
use NAND3X1  _717_
timestamp 1589549099
transform 1 0 632 0 1 1410
box -4 -6 68 206
use NAND3X1  _718_
timestamp 1589549099
transform 1 0 696 0 1 1410
box -4 -6 68 206
use OAI21X1  _715_
timestamp 1589549099
transform -1 0 888 0 1 1410
box -4 -6 68 206
use FILL  SFILL7600x14100
timestamp 1589549099
transform 1 0 760 0 1 1410
box -4 -6 20 206
use FILL  SFILL7760x14100
timestamp 1589549099
transform 1 0 776 0 1 1410
box -4 -6 20 206
use FILL  SFILL7920x14100
timestamp 1589549099
transform 1 0 792 0 1 1410
box -4 -6 20 206
use FILL  SFILL8080x14100
timestamp 1589549099
transform 1 0 808 0 1 1410
box -4 -6 20 206
use INVX1  _634_
timestamp 1589549099
transform 1 0 888 0 1 1410
box -4 -6 36 206
use NOR2X1  _704_
timestamp 1589549099
transform 1 0 920 0 1 1410
box -4 -6 52 206
use OAI21X1  _786_
timestamp 1589549099
transform 1 0 968 0 1 1410
box -4 -6 68 206
use NOR2X1  _976_
timestamp 1589549099
transform 1 0 1032 0 1 1410
box -4 -6 52 206
use NAND3X1  _618_
timestamp 1589549099
transform 1 0 1080 0 1 1410
box -4 -6 68 206
use OAI21X1  _686_
timestamp 1589549099
transform -1 0 1208 0 1 1410
box -4 -6 68 206
use AOI21X1  _687_
timestamp 1589549099
transform -1 0 1272 0 1 1410
box -4 -6 68 206
use NOR2X1  _683_
timestamp 1589549099
transform -1 0 1320 0 1 1410
box -4 -6 52 206
use NOR2X1  _688_
timestamp 1589549099
transform 1 0 1320 0 1 1410
box -4 -6 52 206
use NOR2X1  _680_
timestamp 1589549099
transform 1 0 1368 0 1 1410
box -4 -6 52 206
use NOR2X1  _690_
timestamp 1589549099
transform -1 0 1464 0 1 1410
box -4 -6 52 206
use NOR2X1  _684_
timestamp 1589549099
transform -1 0 1512 0 1 1410
box -4 -6 52 206
use NOR2X1  _682_
timestamp 1589549099
transform 1 0 1512 0 1 1410
box -4 -6 52 206
use NAND2X1  _681_
timestamp 1589549099
transform 1 0 1560 0 1 1410
box -4 -6 52 206
use NAND2X1  _697_
timestamp 1589549099
transform -1 0 1656 0 1 1410
box -4 -6 52 206
use OR2X2  _647_
timestamp 1589549099
transform 1 0 1656 0 1 1410
box -4 -6 68 206
use NOR2X1  _813_
timestamp 1589549099
transform 1 0 1720 0 1 1410
box -4 -6 52 206
use AOI21X1  _837_
timestamp 1589549099
transform 1 0 1768 0 1 1410
box -4 -6 68 206
use OAI22X1  _836_
timestamp 1589549099
transform 1 0 1832 0 1 1410
box -4 -6 84 206
use INVX1  _835_
timestamp 1589549099
transform -1 0 1944 0 1 1410
box -4 -6 36 206
use OAI22X1  _491_
timestamp 1589549099
transform 1 0 1944 0 1 1410
box -4 -6 84 206
use NOR2X1  _490_
timestamp 1589549099
transform -1 0 2072 0 1 1410
box -4 -6 52 206
use AND2X2  _489_
timestamp 1589549099
transform 1 0 2072 0 1 1410
box -4 -6 68 206
use NAND2X1  _983_
timestamp 1589549099
transform -1 0 2184 0 1 1410
box -4 -6 52 206
use OAI21X1  _850_
timestamp 1589549099
transform 1 0 2184 0 1 1410
box -4 -6 68 206
use NOR2X1  _904_
timestamp 1589549099
transform 1 0 2312 0 1 1410
box -4 -6 52 206
use FILL  SFILL22480x14100
timestamp 1589549099
transform 1 0 2248 0 1 1410
box -4 -6 20 206
use FILL  SFILL22640x14100
timestamp 1589549099
transform 1 0 2264 0 1 1410
box -4 -6 20 206
use FILL  SFILL22800x14100
timestamp 1589549099
transform 1 0 2280 0 1 1410
box -4 -6 20 206
use FILL  SFILL22960x14100
timestamp 1589549099
transform 1 0 2296 0 1 1410
box -4 -6 20 206
use OAI21X1  _874_
timestamp 1589549099
transform 1 0 2360 0 1 1410
box -4 -6 68 206
use INVX1  _873_
timestamp 1589549099
transform -1 0 2456 0 1 1410
box -4 -6 36 206
use INVX1  _875_
timestamp 1589549099
transform 1 0 2456 0 1 1410
box -4 -6 36 206
use OAI21X1  _877_
timestamp 1589549099
transform -1 0 2552 0 1 1410
box -4 -6 68 206
use AOI21X1  _876_
timestamp 1589549099
transform 1 0 2552 0 1 1410
box -4 -6 68 206
use NOR2X1  _912_
timestamp 1589549099
transform 1 0 2616 0 1 1410
box -4 -6 52 206
use NAND3X1  _901_
timestamp 1589549099
transform 1 0 2664 0 1 1410
box -4 -6 68 206
use AOI21X1  _900_
timestamp 1589549099
transform 1 0 2728 0 1 1410
box -4 -6 68 206
use OAI22X1  _899_
timestamp 1589549099
transform 1 0 2792 0 1 1410
box -4 -6 84 206
use AOI21X1  _915_
timestamp 1589549099
transform -1 0 2936 0 1 1410
box -4 -6 68 206
use BUFX2  _996_
timestamp 1589549099
transform -1 0 2984 0 1 1410
box -4 -6 52 206
use BUFX2  _998_
timestamp 1589549099
transform 1 0 2984 0 1 1410
box -4 -6 52 206
use BUFX2  _989_
timestamp 1589549099
transform -1 0 56 0 -1 1810
box -4 -6 52 206
use NOR2X1  _650_
timestamp 1589549099
transform -1 0 104 0 -1 1810
box -4 -6 52 206
use NOR2X1  _711_
timestamp 1589549099
transform 1 0 104 0 -1 1810
box -4 -6 52 206
use NOR3X1  _712_
timestamp 1589549099
transform -1 0 280 0 -1 1810
box -4 -6 132 206
use NOR2X1  _708_
timestamp 1589549099
transform -1 0 328 0 -1 1810
box -4 -6 52 206
use OAI21X1  _719_
timestamp 1589549099
transform -1 0 392 0 -1 1810
box -4 -6 68 206
use OAI21X1  _652_
timestamp 1589549099
transform 1 0 392 0 -1 1810
box -4 -6 68 206
use NAND3X1  _713_
timestamp 1589549099
transform -1 0 520 0 -1 1810
box -4 -6 68 206
use OAI21X1  _701_
timestamp 1589549099
transform -1 0 584 0 -1 1810
box -4 -6 68 206
use OAI21X1  _705_
timestamp 1589549099
transform 1 0 584 0 -1 1810
box -4 -6 68 206
use NAND2X1  _651_
timestamp 1589549099
transform -1 0 696 0 -1 1810
box -4 -6 52 206
use NOR2X1  _699_
timestamp 1589549099
transform -1 0 744 0 -1 1810
box -4 -6 52 206
use INVX1  _675_
timestamp 1589549099
transform 1 0 808 0 -1 1810
box -4 -6 36 206
use FILL  SFILL7440x16100
timestamp 1589549099
transform -1 0 760 0 -1 1810
box -4 -6 20 206
use FILL  SFILL7600x16100
timestamp 1589549099
transform -1 0 776 0 -1 1810
box -4 -6 20 206
use FILL  SFILL7760x16100
timestamp 1589549099
transform -1 0 792 0 -1 1810
box -4 -6 20 206
use FILL  SFILL7920x16100
timestamp 1589549099
transform -1 0 808 0 -1 1810
box -4 -6 20 206
use NAND2X1  _617_
timestamp 1589549099
transform 1 0 840 0 -1 1810
box -4 -6 52 206
use NOR2X1  _636_
timestamp 1589549099
transform 1 0 888 0 -1 1810
box -4 -6 52 206
use OAI21X1  _685_
timestamp 1589549099
transform 1 0 936 0 -1 1810
box -4 -6 68 206
use NAND3X1  _710_
timestamp 1589549099
transform -1 0 1064 0 -1 1810
box -4 -6 68 206
use INVX1  _657_
timestamp 1589549099
transform -1 0 1096 0 -1 1810
box -4 -6 36 206
use NOR2X1  _622_
timestamp 1589549099
transform 1 0 1096 0 -1 1810
box -4 -6 52 206
use NAND2X1  _658_
timestamp 1589549099
transform 1 0 1144 0 -1 1810
box -4 -6 52 206
use NAND2X1  _707_
timestamp 1589549099
transform 1 0 1192 0 -1 1810
box -4 -6 52 206
use NOR2X1  _706_
timestamp 1589549099
transform 1 0 1240 0 -1 1810
box -4 -6 52 206
use NAND2X1  _626_
timestamp 1589549099
transform 1 0 1288 0 -1 1810
box -4 -6 52 206
use INVX1  _644_
timestamp 1589549099
transform 1 0 1336 0 -1 1810
box -4 -6 36 206
use OR2X2  _703_
timestamp 1589549099
transform -1 0 1432 0 -1 1810
box -4 -6 68 206
use AND2X2  _487_
timestamp 1589549099
transform -1 0 1496 0 -1 1810
box -4 -6 68 206
use NOR2X1  _488_
timestamp 1589549099
transform -1 0 1544 0 -1 1810
box -4 -6 52 206
use INVX1  _523_
timestamp 1589549099
transform -1 0 1576 0 -1 1810
box -4 -6 36 206
use OAI21X1  _527_
timestamp 1589549099
transform 1 0 1576 0 -1 1810
box -4 -6 68 206
use AOI22X1  _663_
timestamp 1589549099
transform -1 0 1720 0 -1 1810
box -4 -6 84 206
use OAI21X1  _533_
timestamp 1589549099
transform 1 0 1720 0 -1 1810
box -4 -6 68 206
use NAND2X1  _532_
timestamp 1589549099
transform -1 0 1832 0 -1 1810
box -4 -6 52 206
use NOR2X1  _871_
timestamp 1589549099
transform 1 0 1832 0 -1 1810
box -4 -6 52 206
use INVX1  _894_
timestamp 1589549099
transform -1 0 1912 0 -1 1810
box -4 -6 36 206
use OAI21X1  _895_
timestamp 1589549099
transform 1 0 1912 0 -1 1810
box -4 -6 68 206
use NAND3X1  _896_
timestamp 1589549099
transform -1 0 2040 0 -1 1810
box -4 -6 68 206
use OAI21X1  _905_
timestamp 1589549099
transform 1 0 2040 0 -1 1810
box -4 -6 68 206
use NAND3X1  _897_
timestamp 1589549099
transform 1 0 2104 0 -1 1810
box -4 -6 68 206
use OAI21X1  _892_
timestamp 1589549099
transform 1 0 2168 0 -1 1810
box -4 -6 68 206
use INVX1  _885_
timestamp 1589549099
transform 1 0 2232 0 -1 1810
box -4 -6 36 206
use INVX1  _891_
timestamp 1589549099
transform -1 0 2360 0 -1 1810
box -4 -6 36 206
use FILL  SFILL22640x16100
timestamp 1589549099
transform -1 0 2280 0 -1 1810
box -4 -6 20 206
use FILL  SFILL22800x16100
timestamp 1589549099
transform -1 0 2296 0 -1 1810
box -4 -6 20 206
use FILL  SFILL22960x16100
timestamp 1589549099
transform -1 0 2312 0 -1 1810
box -4 -6 20 206
use FILL  SFILL23120x16100
timestamp 1589549099
transform -1 0 2328 0 -1 1810
box -4 -6 20 206
use OAI22X1  _879_
timestamp 1589549099
transform -1 0 2440 0 -1 1810
box -4 -6 84 206
use AOI21X1  _880_
timestamp 1589549099
transform -1 0 2504 0 -1 1810
box -4 -6 68 206
use NAND3X1  _887_
timestamp 1589549099
transform -1 0 2568 0 -1 1810
box -4 -6 68 206
use OAI21X1  _888_
timestamp 1589549099
transform 1 0 2568 0 -1 1810
box -4 -6 68 206
use NAND3X1  _889_
timestamp 1589549099
transform -1 0 2696 0 -1 1810
box -4 -6 68 206
use INVX1  _862_
timestamp 1589549099
transform 1 0 2696 0 -1 1810
box -4 -6 36 206
use OAI22X1  _496_
timestamp 1589549099
transform 1 0 2728 0 -1 1810
box -4 -6 84 206
use NOR2X1  _884_
timestamp 1589549099
transform 1 0 2808 0 -1 1810
box -4 -6 52 206
use OAI21X1  _914_
timestamp 1589549099
transform 1 0 2856 0 -1 1810
box -4 -6 68 206
use NAND2X1  _923_
timestamp 1589549099
transform -1 0 2968 0 -1 1810
box -4 -6 52 206
use INVX1  _898_
timestamp 1589549099
transform -1 0 3000 0 -1 1810
box -4 -6 36 206
use FILL  FILL28720x16100
timestamp 1589549099
transform -1 0 3016 0 -1 1810
box -4 -6 20 206
use FILL  FILL28880x16100
timestamp 1589549099
transform -1 0 3032 0 -1 1810
box -4 -6 20 206
use INVX1  _572_
timestamp 1589549099
transform 1 0 8 0 1 1810
box -4 -6 36 206
use NAND2X1  _576_
timestamp 1589549099
transform 1 0 40 0 1 1810
box -4 -6 52 206
use NOR2X1  _573_
timestamp 1589549099
transform -1 0 136 0 1 1810
box -4 -6 52 206
use AOI21X1  _577_
timestamp 1589549099
transform -1 0 200 0 1 1810
box -4 -6 68 206
use NOR3X1  _709_
timestamp 1589549099
transform -1 0 328 0 1 1810
box -4 -6 132 206
use NAND2X1  _611_
timestamp 1589549099
transform -1 0 376 0 1 1810
box -4 -6 52 206
use AND2X2  _649_
timestamp 1589549099
transform 1 0 376 0 1 1810
box -4 -6 68 206
use OR2X2  _612_
timestamp 1589549099
transform 1 0 440 0 1 1810
box -4 -6 68 206
use AOI21X1  _700_
timestamp 1589549099
transform 1 0 504 0 1 1810
box -4 -6 68 206
use NAND2X1  _613_
timestamp 1589549099
transform -1 0 616 0 1 1810
box -4 -6 52 206
use AOI22X1  _702_
timestamp 1589549099
transform -1 0 696 0 1 1810
box -4 -6 84 206
use BUFX2  _988_
timestamp 1589549099
transform 1 0 696 0 1 1810
box -4 -6 52 206
use INVX1  _574_
timestamp 1589549099
transform 1 0 808 0 1 1810
box -4 -6 36 206
use FILL  SFILL7440x18100
timestamp 1589549099
transform 1 0 744 0 1 1810
box -4 -6 20 206
use FILL  SFILL7600x18100
timestamp 1589549099
transform 1 0 760 0 1 1810
box -4 -6 20 206
use FILL  SFILL7760x18100
timestamp 1589549099
transform 1 0 776 0 1 1810
box -4 -6 20 206
use FILL  SFILL7920x18100
timestamp 1589549099
transform 1 0 792 0 1 1810
box -4 -6 20 206
use NAND2X1  _575_
timestamp 1589549099
transform -1 0 888 0 1 1810
box -4 -6 52 206
use NAND2X1  _616_
timestamp 1589549099
transform -1 0 936 0 1 1810
box -4 -6 52 206
use INVX1  _615_
timestamp 1589549099
transform -1 0 968 0 1 1810
box -4 -6 36 206
use NAND2X1  _614_
timestamp 1589549099
transform -1 0 1016 0 1 1810
box -4 -6 52 206
use NAND2X1  _672_
timestamp 1589549099
transform -1 0 1064 0 1 1810
box -4 -6 52 206
use INVX1  _645_
timestamp 1589549099
transform 1 0 1064 0 1 1810
box -4 -6 36 206
use NAND2X1  _646_
timestamp 1589549099
transform 1 0 1096 0 1 1810
box -4 -6 52 206
use NAND2X1  _679_
timestamp 1589549099
transform -1 0 1192 0 1 1810
box -4 -6 52 206
use INVX1  _623_
timestamp 1589549099
transform 1 0 1192 0 1 1810
box -4 -6 36 206
use NAND2X1  _676_
timestamp 1589549099
transform -1 0 1272 0 1 1810
box -4 -6 52 206
use INVX1  _624_
timestamp 1589549099
transform 1 0 1272 0 1 1810
box -4 -6 36 206
use NOR2X1  _625_
timestamp 1589549099
transform -1 0 1352 0 1 1810
box -4 -6 52 206
use BUFX2  _987_
timestamp 1589549099
transform 1 0 1352 0 1 1810
box -4 -6 52 206
use INVX1  _696_
timestamp 1589549099
transform -1 0 1432 0 1 1810
box -4 -6 36 206
use BUFX2  _997_
timestamp 1589549099
transform -1 0 1480 0 1 1810
box -4 -6 52 206
use INVX1  _883_
timestamp 1589549099
transform -1 0 1512 0 1 1810
box -4 -6 36 206
use INVX1  _841_
timestamp 1589549099
transform 1 0 1512 0 1 1810
box -4 -6 36 206
use NOR2X1  _842_
timestamp 1589549099
transform -1 0 1592 0 1 1810
box -4 -6 52 206
use INVX1  _525_
timestamp 1589549099
transform -1 0 1624 0 1 1810
box -4 -6 36 206
use AND2X2  _662_
timestamp 1589549099
transform -1 0 1688 0 1 1810
box -4 -6 68 206
use OAI22X1  _526_
timestamp 1589549099
transform -1 0 1768 0 1 1810
box -4 -6 84 206
use NAND2X1  _661_
timestamp 1589549099
transform 1 0 1768 0 1 1810
box -4 -6 52 206
use INVX1  _524_
timestamp 1589549099
transform -1 0 1848 0 1 1810
box -4 -6 36 206
use OAI21X1  _867_
timestamp 1589549099
transform -1 0 1912 0 1 1810
box -4 -6 68 206
use AND2X2  _868_
timestamp 1589549099
transform 1 0 1912 0 1 1810
box -4 -6 68 206
use AOI21X1  _882_
timestamp 1589549099
transform 1 0 1976 0 1 1810
box -4 -6 68 206
use NAND3X1  _869_
timestamp 1589549099
transform -1 0 2104 0 1 1810
box -4 -6 68 206
use AOI21X1  _870_
timestamp 1589549099
transform 1 0 2104 0 1 1810
box -4 -6 68 206
use INVX2  _865_
timestamp 1589549099
transform -1 0 2200 0 1 1810
box -4 -6 36 206
use NAND2X1  _886_
timestamp 1589549099
transform 1 0 2200 0 1 1810
box -4 -6 52 206
use OAI21X1  _878_
timestamp 1589549099
transform 1 0 2312 0 1 1810
box -4 -6 68 206
use FILL  SFILL22480x18100
timestamp 1589549099
transform 1 0 2248 0 1 1810
box -4 -6 20 206
use FILL  SFILL22640x18100
timestamp 1589549099
transform 1 0 2264 0 1 1810
box -4 -6 20 206
use FILL  SFILL22800x18100
timestamp 1589549099
transform 1 0 2280 0 1 1810
box -4 -6 20 206
use FILL  SFILL22960x18100
timestamp 1589549099
transform 1 0 2296 0 1 1810
box -4 -6 20 206
use OAI21X1  _881_
timestamp 1589549099
transform -1 0 2440 0 1 1810
box -4 -6 68 206
use INVX1  _863_
timestamp 1589549099
transform 1 0 2440 0 1 1810
box -4 -6 36 206
use NAND2X1  _864_
timestamp 1589549099
transform 1 0 2472 0 1 1810
box -4 -6 52 206
use NAND2X1  _890_
timestamp 1589549099
transform -1 0 2568 0 1 1810
box -4 -6 52 206
use NOR2X1  _493_
timestamp 1589549099
transform -1 0 2616 0 1 1810
box -4 -6 52 206
use INVX1  _530_
timestamp 1589549099
transform -1 0 2648 0 1 1810
box -4 -6 36 206
use AND2X2  _492_
timestamp 1589549099
transform 1 0 2648 0 1 1810
box -4 -6 68 206
use OAI22X1  _531_
timestamp 1589549099
transform -1 0 2792 0 1 1810
box -4 -6 84 206
use NAND2X1  _529_
timestamp 1589549099
transform -1 0 2840 0 1 1810
box -4 -6 52 206
use INVX1  _528_
timestamp 1589549099
transform -1 0 2872 0 1 1810
box -4 -6 36 206
use NOR2X1  _495_
timestamp 1589549099
transform -1 0 2920 0 1 1810
box -4 -6 52 206
use AND2X2  _494_
timestamp 1589549099
transform -1 0 2984 0 1 1810
box -4 -6 68 206
use BUFX2  _999_
timestamp 1589549099
transform 1 0 2984 0 1 1810
box -4 -6 52 206
<< labels >>
flabel metal4 s 2240 -10 2304 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 736 -10 800 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 2189 -23 2195 -17 7 FreeSans 24 270 0 0 a[15]
port 2 nsew
flabel metal3 s 3069 1077 3075 1083 3 FreeSans 24 0 0 0 a[14]
port 3 nsew
flabel metal2 s 1773 -23 1779 -17 7 FreeSans 24 270 0 0 a[13]
port 4 nsew
flabel metal2 s 1981 -23 1987 -17 7 FreeSans 24 270 0 0 a[12]
port 5 nsew
flabel metal2 s 2893 2057 2899 2063 3 FreeSans 24 90 0 0 a[11]
port 6 nsew
flabel metal2 s 2573 2057 2579 2063 3 FreeSans 24 90 0 0 a[10]
port 7 nsew
flabel metal2 s 1885 2057 1891 2063 3 FreeSans 24 90 0 0 a[9]
port 8 nsew
flabel metal2 s 1709 2057 1715 2063 3 FreeSans 24 90 0 0 a[8]
port 9 nsew
flabel metal3 s -35 277 -29 283 7 FreeSans 24 0 0 0 a[7]
port 10 nsew
flabel metal3 s -35 317 -29 323 7 FreeSans 24 0 0 0 a[6]
port 11 nsew
flabel metal2 s 1069 -23 1075 -17 7 FreeSans 24 270 0 0 a[5]
port 12 nsew
flabel metal2 s 1485 -23 1491 -17 7 FreeSans 24 270 0 0 a[4]
port 13 nsew
flabel metal3 s -35 1117 -29 1123 7 FreeSans 24 0 0 0 a[3]
port 14 nsew
flabel metal3 s -35 1357 -29 1363 7 FreeSans 24 0 0 0 a[2]
port 15 nsew
flabel metal3 s -35 1897 -29 1903 7 FreeSans 24 0 0 0 a[1]
port 16 nsew
flabel metal2 s 1005 2057 1011 2063 3 FreeSans 24 90 0 0 a[0]
port 17 nsew
flabel metal3 s 3069 297 3075 303 3 FreeSans 24 0 0 0 alu_output[15]
port 18 nsew
flabel metal3 s 3069 97 3075 103 3 FreeSans 24 0 0 0 alu_output[14]
port 19 nsew
flabel metal2 s 2829 -23 2835 -17 7 FreeSans 24 270 0 0 alu_output[13]
port 20 nsew
flabel metal3 s 3069 1897 3075 1903 3 FreeSans 24 0 0 0 alu_output[12]
port 21 nsew
flabel metal3 s 3069 1517 3075 1523 3 FreeSans 24 0 0 0 alu_output[11]
port 22 nsew
flabel metal2 s 1453 2057 1459 2063 3 FreeSans 24 90 0 0 alu_output[10]
port 23 nsew
flabel metal3 s 3069 1477 3075 1483 3 FreeSans 24 0 0 0 alu_output[9]
port 24 nsew
flabel metal2 s 1709 -23 1715 -17 7 FreeSans 24 270 0 0 alu_output[8]
port 25 nsew
flabel metal2 s 573 -23 579 -17 7 FreeSans 24 270 0 0 alu_output[7]
port 26 nsew
flabel metal2 s 653 -23 659 -17 7 FreeSans 24 270 0 0 alu_output[6]
port 27 nsew
flabel metal2 s 1133 -23 1139 -17 7 FreeSans 24 270 0 0 alu_output[5]
port 28 nsew
flabel metal2 s 1661 -23 1667 -17 7 FreeSans 24 270 0 0 alu_output[4]
port 29 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 alu_output[3]
port 30 nsew
flabel metal3 s -35 1697 -29 1703 7 FreeSans 24 0 0 0 alu_output[2]
port 31 nsew
flabel metal2 s 829 2057 835 2063 3 FreeSans 24 90 0 0 alu_output[1]
port 32 nsew
flabel metal2 s 1373 2057 1379 2063 3 FreeSans 24 90 0 0 alu_output[0]
port 33 nsew
flabel metal2 s 2429 -23 2435 -17 7 FreeSans 24 270 0 0 b[15]
port 34 nsew
flabel metal3 s 3069 917 3075 923 3 FreeSans 24 0 0 0 b[14]
port 35 nsew
flabel metal2 s 1837 -23 1843 -17 7 FreeSans 24 270 0 0 b[13]
port 36 nsew
flabel metal2 s 2029 -23 2035 -17 7 FreeSans 24 270 0 0 b[12]
port 37 nsew
flabel metal2 s 2941 2057 2947 2063 3 FreeSans 24 90 0 0 b[11]
port 38 nsew
flabel metal2 s 2669 2057 2675 2063 3 FreeSans 24 90 0 0 b[10]
port 39 nsew
flabel metal2 s 1805 2057 1811 2063 3 FreeSans 24 90 0 0 b[9]
port 40 nsew
flabel metal2 s 1549 2057 1555 2063 3 FreeSans 24 90 0 0 b[8]
port 41 nsew
flabel metal3 s -35 137 -29 143 7 FreeSans 24 0 0 0 b[7]
port 42 nsew
flabel metal3 s -35 677 -29 683 7 FreeSans 24 0 0 0 b[6]
port 43 nsew
flabel metal2 s 1229 -23 1235 -17 7 FreeSans 24 270 0 0 b[5]
port 44 nsew
flabel metal2 s 1597 -23 1603 -17 7 FreeSans 24 270 0 0 b[4]
port 45 nsew
flabel metal3 s -35 1077 -29 1083 7 FreeSans 24 0 0 0 b[3]
port 46 nsew
flabel metal3 s -35 1477 -29 1483 7 FreeSans 24 0 0 0 b[2]
port 47 nsew
flabel metal3 s -35 1857 -29 1863 7 FreeSans 24 0 0 0 b[1]
port 48 nsew
flabel metal2 s 973 2057 979 2063 3 FreeSans 24 90 0 0 b[0]
port 49 nsew
flabel metal3 s 3069 1117 3075 1123 3 FreeSans 24 0 0 0 carryout
port 50 nsew
flabel metal2 s 1213 2057 1219 2063 3 FreeSans 24 90 0 0 op_code[3]
port 51 nsew
flabel metal2 s 1261 2057 1267 2063 3 FreeSans 24 90 0 0 op_code[2]
port 52 nsew
flabel metal2 s 1069 2057 1075 2063 3 FreeSans 24 90 0 0 op_code[1]
port 53 nsew
flabel metal2 s 1101 2057 1107 2063 3 FreeSans 24 90 0 0 op_code[0]
port 54 nsew
flabel metal2 s 2925 -23 2931 -17 7 FreeSans 24 270 0 0 zero_flag
port 55 nsew
<< end >>
