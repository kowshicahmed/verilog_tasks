magic
tech scmos
magscale 1 2
timestamp 1597059762
<< metal1 >>
rect 762 5214 774 5216
rect 3770 5214 3782 5216
rect 6778 5214 6790 5216
rect 747 5206 749 5214
rect 757 5206 759 5214
rect 767 5206 769 5214
rect 777 5206 779 5214
rect 787 5206 789 5214
rect 3755 5206 3757 5214
rect 3765 5206 3767 5214
rect 3775 5206 3777 5214
rect 3785 5206 3787 5214
rect 3795 5206 3797 5214
rect 6763 5206 6765 5214
rect 6773 5206 6775 5214
rect 6783 5206 6785 5214
rect 6793 5206 6795 5214
rect 6803 5206 6805 5214
rect 762 5204 774 5206
rect 3770 5204 3782 5206
rect 6778 5204 6790 5206
rect 5261 5177 5324 5183
rect 4909 5137 4924 5143
rect 1012 5116 1020 5124
rect 4717 5117 4732 5123
rect 5076 5117 5091 5123
rect 5188 5117 5203 5123
rect 5501 5117 5523 5123
rect 5757 5117 5779 5123
rect 6228 5117 6243 5123
rect 6340 5117 6355 5123
rect 7357 5117 7379 5123
rect 5516 5104 5524 5108
rect 852 5097 883 5103
rect 2093 5097 2108 5103
rect 2244 5097 2275 5103
rect 2845 5097 2860 5103
rect 4861 5097 4876 5103
rect 6061 5097 6076 5103
rect 6733 5097 6819 5103
rect 6893 5097 6915 5103
rect 7053 5103 7059 5116
rect 7037 5097 7059 5103
rect 7117 5097 7132 5103
rect 7204 5097 7219 5103
rect 7364 5097 7379 5103
rect 7549 5097 7564 5103
rect 333 5077 371 5083
rect 253 5057 291 5063
rect 365 5057 371 5077
rect 532 5076 534 5084
rect 925 5077 963 5083
rect 925 5057 931 5077
rect 1757 5077 1772 5083
rect 2093 5077 2131 5083
rect 1453 5057 1491 5063
rect 2093 5057 2099 5077
rect 2332 5077 2348 5083
rect 2429 5077 2467 5083
rect 2461 5057 2467 5077
rect 2749 5077 2764 5083
rect 3148 5077 3172 5083
rect 3373 5077 3411 5083
rect 3405 5057 3411 5077
rect 4012 5077 4036 5083
rect 4797 5077 4812 5083
rect 4884 5077 4899 5083
rect 3709 5057 3747 5063
rect 3764 5057 3827 5063
rect 3821 5043 3827 5057
rect 4893 5057 4899 5077
rect 5021 5077 5059 5083
rect 5597 5077 5635 5083
rect 5821 5077 5843 5083
rect 5949 5077 5964 5083
rect 5156 5056 5164 5064
rect 5924 5057 5939 5063
rect 5949 5057 5955 5077
rect 6989 5077 7027 5083
rect 6308 5056 6316 5064
rect 6845 5057 6860 5063
rect 6989 5057 6995 5077
rect 7044 5077 7075 5083
rect 7149 5077 7164 5083
rect 7261 5077 7299 5083
rect 7261 5057 7267 5077
rect 3821 5037 3843 5043
rect 5604 5036 5606 5044
rect 5688 5036 5692 5044
rect 2266 5014 2278 5016
rect 5274 5014 5286 5016
rect 2251 5006 2253 5014
rect 2261 5006 2263 5014
rect 2271 5006 2273 5014
rect 2281 5006 2283 5014
rect 2291 5006 2293 5014
rect 5259 5006 5261 5014
rect 5269 5006 5271 5014
rect 5279 5006 5281 5014
rect 5289 5006 5291 5014
rect 5299 5006 5301 5014
rect 2266 5004 2278 5006
rect 5274 5004 5286 5006
rect 6618 4976 6620 4984
rect 7348 4976 7352 4984
rect 253 4943 259 4963
rect 1732 4957 1747 4963
rect 2653 4957 2691 4963
rect 2957 4957 2995 4963
rect 3069 4957 3107 4963
rect 3533 4957 3571 4963
rect 3981 4957 4003 4963
rect 4109 4957 4131 4963
rect 5181 4957 5203 4963
rect 5549 4957 5564 4963
rect 6244 4957 6259 4963
rect 253 4937 291 4943
rect 941 4937 963 4943
rect 324 4917 339 4923
rect 397 4917 412 4923
rect 941 4923 947 4937
rect 1188 4937 1203 4943
rect 1709 4937 1724 4943
rect 2916 4937 2931 4943
rect 4829 4943 4835 4956
rect 4813 4937 4835 4943
rect 5037 4943 5043 4956
rect 5037 4937 5059 4943
rect 5204 4937 5219 4943
rect 5789 4937 5827 4943
rect 932 4917 947 4923
rect 989 4917 1020 4923
rect 989 4897 995 4917
rect 1053 4917 1091 4923
rect 1053 4897 1059 4917
rect 1156 4917 1187 4923
rect 1181 4897 1187 4917
rect 1404 4917 1443 4923
rect 1404 4914 1412 4917
rect 1725 4917 1731 4936
rect 2029 4917 2044 4923
rect 2429 4917 2444 4923
rect 3428 4917 3443 4923
rect 3860 4917 3891 4923
rect 4157 4917 4172 4923
rect 4989 4923 4995 4936
rect 6205 4937 6227 4943
rect 6269 4937 6307 4943
rect 6445 4943 6451 4963
rect 6461 4957 6483 4963
rect 6685 4957 6707 4963
rect 6436 4937 6451 4943
rect 6692 4937 6707 4943
rect 6989 4937 7004 4943
rect 7156 4937 7171 4943
rect 5324 4923 5332 4928
rect 6204 4924 6212 4928
rect 4989 4917 5011 4923
rect 5245 4917 5332 4923
rect 5581 4917 5596 4923
rect 6372 4917 6387 4923
rect 6740 4917 6819 4923
rect 7053 4917 7068 4923
rect 7085 4917 7116 4923
rect 6525 4897 6547 4903
rect 2854 4876 2860 4884
rect 6548 4877 6579 4883
rect 5892 4856 5896 4864
rect 362 4836 364 4844
rect 458 4836 460 4844
rect 1466 4836 1468 4844
rect 1562 4836 1564 4844
rect 2004 4836 2006 4844
rect 2554 4836 2556 4844
rect 4794 4836 4796 4844
rect 4932 4836 4936 4844
rect 5092 4836 5096 4844
rect 5448 4836 5452 4844
rect 6004 4836 6008 4844
rect 6324 4836 6326 4844
rect 7524 4836 7526 4844
rect 762 4814 774 4816
rect 3770 4814 3782 4816
rect 6778 4814 6790 4816
rect 747 4806 749 4814
rect 757 4806 759 4814
rect 767 4806 769 4814
rect 777 4806 779 4814
rect 787 4806 789 4814
rect 3755 4806 3757 4814
rect 3765 4806 3767 4814
rect 3775 4806 3777 4814
rect 3785 4806 3787 4814
rect 3795 4806 3797 4814
rect 6763 4806 6765 4814
rect 6773 4806 6775 4814
rect 6783 4806 6785 4814
rect 6793 4806 6795 4814
rect 6803 4806 6805 4814
rect 762 4804 774 4806
rect 3770 4804 3782 4806
rect 6778 4804 6790 4806
rect 820 4776 822 4784
rect 2090 4776 2092 4784
rect 5261 4777 5308 4783
rect 7549 4777 7564 4783
rect 490 4756 492 4764
rect 1898 4736 1900 4744
rect 2682 4736 2684 4744
rect 3757 4737 3820 4743
rect 4342 4736 4348 4744
rect 5021 4737 5036 4743
rect 557 4697 572 4703
rect 845 4703 851 4723
rect 845 4697 883 4703
rect 1236 4697 1251 4703
rect 1341 4703 1347 4723
rect 1341 4697 1379 4703
rect 1837 4703 1843 4723
rect 1837 4697 1860 4703
rect 1852 4692 1860 4697
rect 2541 4697 2595 4703
rect 2653 4703 2659 4723
rect 4925 4717 4947 4723
rect 5933 4717 5955 4723
rect 2636 4697 2659 4703
rect 2636 4692 2644 4697
rect 3037 4697 3052 4703
rect 3076 4697 3091 4703
rect 4980 4697 4995 4703
rect 5540 4697 5555 4703
rect 5645 4697 5660 4703
rect 5677 4697 5699 4703
rect 6269 4703 6275 4723
rect 7101 4717 7116 4723
rect 7309 4717 7347 4723
rect 6269 4697 6323 4703
rect 6429 4697 6460 4703
rect 6781 4697 6867 4703
rect 6964 4697 6979 4703
rect 7357 4703 7363 4716
rect 7357 4697 7379 4703
rect 7389 4697 7404 4703
rect 509 4677 531 4683
rect 580 4677 595 4683
rect 637 4677 659 4683
rect 740 4677 803 4683
rect 1053 4677 1075 4683
rect 1341 4677 1356 4683
rect 3261 4677 3283 4683
rect 4893 4677 4908 4683
rect 5197 4683 5203 4696
rect 5181 4677 5203 4683
rect 5373 4677 5388 4683
rect 5476 4677 5507 4683
rect 5517 4677 5548 4683
rect 5565 4677 5603 4683
rect 2877 4657 2915 4663
rect 3501 4657 3523 4663
rect 3629 4657 3651 4663
rect 3757 4657 3843 4663
rect 5597 4657 5603 4677
rect 5700 4677 5715 4683
rect 5908 4677 5923 4683
rect 5917 4657 5923 4677
rect 7005 4677 7020 4683
rect 7005 4657 7011 4677
rect 7341 4677 7372 4683
rect 7501 4677 7532 4683
rect 7524 4657 7539 4663
rect 4676 4636 4680 4644
rect 4954 4636 4956 4644
rect 5962 4636 5964 4644
rect 6184 4636 6188 4644
rect 6260 4636 6262 4644
rect 7092 4636 7094 4644
rect 2266 4614 2278 4616
rect 5274 4614 5286 4616
rect 2251 4606 2253 4614
rect 2261 4606 2263 4614
rect 2271 4606 2273 4614
rect 2281 4606 2283 4614
rect 2291 4606 2293 4614
rect 5259 4606 5261 4614
rect 5269 4606 5271 4614
rect 5279 4606 5281 4614
rect 5289 4606 5291 4614
rect 5299 4606 5301 4614
rect 2266 4604 2278 4606
rect 5274 4604 5286 4606
rect 29 4557 67 4563
rect 269 4557 307 4563
rect 100 4537 131 4543
rect 205 4537 220 4543
rect 317 4543 323 4563
rect 477 4557 492 4563
rect 893 4557 908 4563
rect 1597 4557 1635 4563
rect 317 4537 332 4543
rect 701 4537 787 4543
rect 868 4537 883 4543
rect 2125 4543 2131 4556
rect 2084 4537 2115 4543
rect 2125 4537 2147 4543
rect 2237 4537 2252 4543
rect 2653 4537 2668 4543
rect 2860 4543 2868 4548
rect 2781 4537 2803 4543
rect 2845 4537 2868 4543
rect 3261 4537 3283 4543
rect 3549 4543 3555 4563
rect 4253 4557 4275 4563
rect 5044 4557 5059 4563
rect 3517 4537 3555 4543
rect 4797 4537 4819 4543
rect 5044 4537 5075 4543
rect 5325 4543 5331 4563
rect 5469 4557 5491 4563
rect 5988 4557 6003 4563
rect 6109 4557 6140 4563
rect 7229 4557 7251 4563
rect 5252 4537 5331 4543
rect 5469 4537 5484 4543
rect 5597 4537 5635 4543
rect 5965 4537 5996 4543
rect 6061 4537 6099 4543
rect 6317 4537 6332 4543
rect 6916 4537 6931 4543
rect 7316 4537 7331 4543
rect 7364 4537 7395 4543
rect 7460 4537 7475 4543
rect 1796 4517 1811 4523
rect 2077 4517 2092 4523
rect 2157 4517 2195 4523
rect 1197 4497 1235 4503
rect 1924 4496 1932 4504
rect 2189 4497 2195 4517
rect 2221 4517 2236 4523
rect 2557 4517 2595 4523
rect 2557 4497 2563 4517
rect 2829 4517 2844 4523
rect 2948 4517 2979 4523
rect 3060 4517 3075 4523
rect 3101 4517 3139 4523
rect 3076 4496 3084 4504
rect 3101 4497 3107 4517
rect 3156 4517 3171 4523
rect 3420 4523 3428 4528
rect 3420 4517 3443 4523
rect 3437 4497 3443 4517
rect 4253 4517 4268 4523
rect 4397 4517 4412 4523
rect 4845 4517 4876 4523
rect 5268 4517 5347 4523
rect 5524 4517 5539 4523
rect 5725 4517 5747 4523
rect 5821 4517 5843 4523
rect 5917 4517 5948 4523
rect 6141 4517 6156 4523
rect 6461 4517 6499 4523
rect 6493 4504 6499 4517
rect 6893 4517 6924 4523
rect 7181 4517 7212 4523
rect 7469 4523 7475 4537
rect 7469 4517 7507 4523
rect 4861 4497 4899 4503
rect 4909 4497 4931 4503
rect 6116 4497 6131 4503
rect 6733 4497 6796 4503
rect 6813 4497 6828 4503
rect 7432 4498 7436 4506
rect 1172 4476 1174 4484
rect 2356 4476 2362 4484
rect 2900 4476 2906 4484
rect 6804 4477 6851 4483
rect 356 4436 358 4444
rect 1450 4436 1452 4444
rect 2762 4436 2764 4444
rect 3322 4436 3324 4444
rect 4708 4436 4712 4444
rect 5140 4436 5142 4444
rect 7178 4436 7180 4444
rect 7508 4436 7510 4444
rect 762 4414 774 4416
rect 3770 4414 3782 4416
rect 6778 4414 6790 4416
rect 747 4406 749 4414
rect 757 4406 759 4414
rect 767 4406 769 4414
rect 777 4406 779 4414
rect 787 4406 789 4414
rect 3755 4406 3757 4414
rect 3765 4406 3767 4414
rect 3775 4406 3777 4414
rect 3785 4406 3787 4414
rect 3795 4406 3797 4414
rect 6763 4406 6765 4414
rect 6773 4406 6775 4414
rect 6783 4406 6785 4414
rect 6793 4406 6795 4414
rect 6803 4406 6805 4414
rect 762 4404 774 4406
rect 3770 4404 3782 4406
rect 6778 4404 6790 4406
rect 554 4376 556 4384
rect 842 4376 844 4384
rect 1018 4376 1020 4384
rect 1834 4376 1836 4384
rect 2221 4377 2268 4383
rect 3130 4376 3132 4384
rect 3444 4376 3446 4384
rect 4026 4376 4028 4384
rect 4282 4376 4284 4384
rect 7412 4376 7414 4384
rect 1188 4336 1190 4344
rect 1514 4336 1516 4344
rect 3188 4336 3190 4344
rect 4916 4337 4931 4343
rect 5544 4336 5548 4344
rect 557 4297 572 4303
rect 701 4297 732 4303
rect 845 4297 899 4303
rect 980 4297 995 4303
rect 1085 4297 1100 4303
rect 1325 4297 1340 4303
rect 1453 4303 1459 4323
rect 3700 4316 3708 4324
rect 5805 4317 5820 4323
rect 5917 4317 5939 4323
rect 6013 4317 6028 4323
rect 6301 4317 6323 4323
rect 6333 4317 6348 4323
rect 6733 4317 6764 4323
rect 1412 4297 1427 4303
rect 1453 4297 1476 4303
rect 1468 4292 1476 4297
rect 1517 4297 1571 4303
rect 2381 4297 2396 4303
rect 2532 4297 2547 4303
rect 3277 4297 3308 4303
rect 3709 4297 3724 4303
rect 4236 4303 4244 4306
rect 4236 4297 4252 4303
rect 4733 4297 4748 4303
rect 4868 4297 4883 4303
rect 5629 4297 5667 4303
rect 5773 4297 5811 4303
rect 6381 4297 6403 4303
rect 6461 4297 6499 4303
rect 6701 4297 6739 4303
rect 7092 4297 7139 4303
rect 7325 4297 7340 4303
rect 7517 4297 7564 4303
rect 253 4277 291 4283
rect 253 4257 259 4277
rect 701 4277 780 4283
rect 1396 4277 1411 4283
rect 2125 4277 2163 4283
rect 362 4256 364 4264
rect 2125 4257 2131 4277
rect 2580 4277 2611 4283
rect 2781 4277 2796 4283
rect 2909 4277 2924 4283
rect 3085 4277 3116 4283
rect 3588 4277 3603 4283
rect 4788 4277 4808 4283
rect 4893 4277 4915 4283
rect 4909 4264 4915 4277
rect 5165 4277 5203 4283
rect 5261 4277 5363 4283
rect 5709 4277 5763 4283
rect 5860 4277 5891 4283
rect 6045 4277 6099 4283
rect 6356 4277 6364 4283
rect 6685 4277 6716 4283
rect 6932 4277 6947 4283
rect 6996 4277 7011 4283
rect 7044 4277 7075 4283
rect 7213 4277 7228 4283
rect 7357 4277 7395 4283
rect 2813 4257 2828 4263
rect 3156 4257 3171 4263
rect 5613 4257 5628 4263
rect 6125 4257 6163 4263
rect 6365 4257 6371 4276
rect 6964 4256 6972 4264
rect 7140 4257 7155 4263
rect 6836 4236 6838 4244
rect 7028 4236 7030 4244
rect 2266 4214 2278 4216
rect 5274 4214 5286 4216
rect 2251 4206 2253 4214
rect 2261 4206 2263 4214
rect 2271 4206 2273 4214
rect 2281 4206 2283 4214
rect 2291 4206 2293 4214
rect 5259 4206 5261 4214
rect 5269 4206 5271 4214
rect 5279 4206 5281 4214
rect 5289 4206 5291 4214
rect 5299 4206 5301 4214
rect 2266 4204 2278 4206
rect 5274 4204 5286 4206
rect 6088 4176 6092 4184
rect 6538 4176 6540 4184
rect 6632 4176 6636 4184
rect 6765 4177 6828 4183
rect 253 4143 259 4163
rect 820 4157 835 4163
rect 3325 4157 3363 4163
rect 3949 4157 3971 4163
rect 4541 4157 4579 4163
rect 4612 4157 4627 4163
rect 4637 4157 4675 4163
rect 253 4137 291 4143
rect 733 4137 796 4143
rect 1476 4137 1491 4143
rect 3140 4137 3155 4143
rect 3261 4137 3283 4143
rect 605 4117 643 4123
rect 580 4096 588 4104
rect 605 4097 611 4117
rect 1309 4117 1347 4123
rect 1309 4097 1315 4117
rect 1645 4117 1699 4123
rect 1740 4123 1748 4128
rect 1740 4117 1763 4123
rect 1757 4097 1763 4117
rect 2077 4117 2115 4123
rect 2109 4097 2115 4117
rect 2493 4117 2531 4123
rect 2525 4097 2531 4117
rect 2893 4117 2908 4123
rect 3277 4124 3283 4137
rect 3533 4137 3548 4143
rect 4733 4143 4739 4163
rect 6292 4157 6307 4163
rect 6957 4157 6979 4163
rect 4733 4137 4771 4143
rect 4845 4137 4860 4143
rect 4957 4137 4979 4143
rect 5469 4137 5484 4143
rect 5645 4137 5660 4143
rect 6269 4137 6300 4143
rect 3028 4117 3043 4123
rect 3069 4117 3107 4123
rect 3117 4117 3148 4123
rect 3044 4096 3052 4104
rect 3069 4097 3075 4117
rect 3156 4117 3171 4123
rect 3181 4117 3219 4123
rect 3213 4097 3219 4117
rect 3533 4117 3571 4123
rect 3533 4097 3539 4117
rect 4605 4117 4620 4123
rect 4717 4117 4748 4123
rect 4781 4117 4803 4123
rect 5316 4117 5347 4123
rect 5565 4117 5603 4123
rect 5661 4117 5708 4123
rect 6573 4123 6579 4143
rect 7053 4137 7075 4143
rect 7316 4137 7331 4143
rect 6564 4117 6579 4123
rect 6877 4117 6892 4123
rect 7197 4117 7212 4123
rect 7533 4117 7548 4123
rect 5732 4096 5740 4104
rect 6461 4097 6492 4103
rect 6509 4097 6531 4103
rect 7197 4097 7219 4103
rect 7437 4097 7452 4103
rect 922 4076 924 4084
rect 2554 4076 2556 4084
rect 7229 4077 7244 4083
rect 330 4036 332 4044
rect 3242 4036 3244 4044
rect 4692 4036 4694 4044
rect 7128 4036 7132 4044
rect 7290 4036 7292 4044
rect 762 4014 774 4016
rect 3770 4014 3782 4016
rect 6778 4014 6790 4016
rect 747 4006 749 4014
rect 757 4006 759 4014
rect 767 4006 769 4014
rect 777 4006 779 4014
rect 787 4006 789 4014
rect 3755 4006 3757 4014
rect 3765 4006 3767 4014
rect 3775 4006 3777 4014
rect 3785 4006 3787 4014
rect 3795 4006 3797 4014
rect 6763 4006 6765 4014
rect 6773 4006 6775 4014
rect 6783 4006 6785 4014
rect 6793 4006 6795 4014
rect 6803 4006 6805 4014
rect 762 4004 774 4006
rect 3770 4004 3782 4006
rect 6778 4004 6790 4006
rect 189 3937 204 3943
rect 454 3936 460 3944
rect 749 3937 764 3943
rect 1556 3936 1558 3944
rect 7108 3936 7110 3944
rect 253 3903 259 3923
rect 221 3897 259 3903
rect 2333 3903 2339 3923
rect 2356 3916 2364 3924
rect 2237 3897 2339 3903
rect 2733 3903 2739 3923
rect 4813 3917 4828 3923
rect 5444 3917 5459 3923
rect 7133 3917 7155 3923
rect 7341 3917 7356 3923
rect 2701 3897 2739 3903
rect 2765 3897 2780 3903
rect 2996 3897 3011 3903
rect 3293 3897 3308 3903
rect 3428 3897 3443 3903
rect 3828 3897 3859 3903
rect 4317 3897 4339 3903
rect 4589 3897 4611 3903
rect 5565 3897 5587 3903
rect 5836 3903 5844 3908
rect 5836 3897 5859 3903
rect 772 3877 828 3883
rect 1037 3877 1052 3883
rect 1844 3877 1859 3883
rect 4253 3877 4268 3883
rect 4381 3877 4396 3883
rect 5236 3877 5299 3883
rect 5444 3877 5475 3883
rect 5853 3877 5859 3897
rect 5997 3897 6051 3903
rect 6109 3897 6124 3903
rect 5869 3877 5907 3883
rect 5997 3877 6003 3897
rect 6109 3884 6115 3897
rect 6141 3897 6163 3903
rect 6196 3897 6211 3903
rect 6301 3897 6339 3903
rect 6541 3897 6563 3903
rect 6621 3897 6643 3903
rect 6756 3897 6819 3903
rect 7276 3903 7284 3908
rect 7276 3897 7299 3903
rect 6173 3877 6211 3883
rect 6237 3877 6291 3883
rect 6365 3877 6380 3883
rect 6205 3864 6211 3877
rect 6605 3877 6620 3883
rect 6692 3877 6707 3883
rect 7069 3877 7091 3883
rect 7293 3877 7299 3897
rect 7485 3877 7500 3883
rect 7549 3877 7564 3883
rect 7021 3857 7052 3863
rect 852 3836 854 3844
rect 4436 3836 4438 3844
rect 5213 3837 5228 3843
rect 5428 3836 5430 3844
rect 5626 3836 5628 3844
rect 7380 3836 7382 3844
rect 2266 3814 2278 3816
rect 5274 3814 5286 3816
rect 2251 3806 2253 3814
rect 2261 3806 2263 3814
rect 2271 3806 2273 3814
rect 2281 3806 2283 3814
rect 2291 3806 2293 3814
rect 5259 3806 5261 3814
rect 5269 3806 5271 3814
rect 5279 3806 5281 3814
rect 5289 3806 5291 3814
rect 5299 3806 5301 3814
rect 2266 3804 2278 3806
rect 5274 3804 5286 3806
rect 5832 3776 5836 3784
rect 221 3757 259 3763
rect 477 3737 492 3743
rect 845 3737 867 3743
rect 1181 3737 1196 3743
rect 1981 3737 1996 3743
rect 3197 3737 3212 3743
rect 3437 3743 3443 3763
rect 3437 3737 3475 3743
rect 3788 3737 3852 3743
rect 4189 3743 4195 3763
rect 4452 3756 4460 3764
rect 5485 3757 5507 3763
rect 6884 3757 6899 3763
rect 6909 3757 6947 3763
rect 4157 3737 4195 3743
rect 4365 3743 4371 3756
rect 4349 3737 4371 3743
rect 4484 3737 4531 3743
rect 4829 3737 4844 3743
rect 5197 3737 5235 3743
rect 5677 3737 5715 3743
rect 6196 3737 6211 3743
rect 6413 3743 6419 3756
rect 6308 3737 6323 3743
rect 6413 3737 6435 3743
rect 7149 3737 7171 3743
rect 436 3717 451 3723
rect 477 3717 515 3723
rect 477 3697 483 3717
rect 1140 3717 1155 3723
rect 1181 3717 1219 3723
rect 1181 3697 1187 3717
rect 1853 3717 1891 3723
rect 1460 3696 1468 3704
rect 1885 3697 1891 3717
rect 2061 3717 2076 3723
rect 2397 3717 2435 3723
rect 2636 3717 2675 3723
rect 2397 3697 2403 3717
rect 2636 3714 2644 3717
rect 2756 3717 2771 3723
rect 7165 3724 7171 3737
rect 7220 3737 7235 3743
rect 7533 3737 7564 3743
rect 3268 3717 3283 3723
rect 3485 3717 3500 3723
rect 3517 3717 3555 3723
rect 2861 3697 2899 3703
rect 3549 3697 3555 3717
rect 4180 3717 4211 3723
rect 4221 3717 4243 3723
rect 4413 3717 4435 3723
rect 4573 3717 4595 3723
rect 4765 3717 4787 3723
rect 5005 3717 5027 3723
rect 5117 3717 5132 3723
rect 5277 3717 5363 3723
rect 5533 3717 5555 3723
rect 6013 3717 6028 3723
rect 6173 3717 6204 3723
rect 6253 3717 6291 3723
rect 3572 3696 3580 3704
rect 6141 3697 6156 3703
rect 6253 3697 6259 3717
rect 6349 3717 6387 3723
rect 6612 3717 6627 3723
rect 6772 3717 6835 3723
rect 7181 3717 7212 3723
rect 1821 3677 1836 3683
rect 3094 3676 3100 3684
rect 3652 3676 3658 3684
rect 4653 3677 4668 3683
rect 6084 3677 6099 3683
rect 964 3636 966 3644
rect 2020 3636 2022 3644
rect 2794 3636 2796 3644
rect 3306 3636 3308 3644
rect 5944 3636 5948 3644
rect 6052 3636 6054 3644
rect 6394 3636 6396 3644
rect 6964 3636 6966 3644
rect 7112 3636 7116 3644
rect 7316 3636 7320 3644
rect 762 3614 774 3616
rect 3770 3614 3782 3616
rect 6778 3614 6790 3616
rect 747 3606 749 3614
rect 757 3606 759 3614
rect 767 3606 769 3614
rect 777 3606 779 3614
rect 787 3606 789 3614
rect 3755 3606 3757 3614
rect 3765 3606 3767 3614
rect 3775 3606 3777 3614
rect 3785 3606 3787 3614
rect 3795 3606 3797 3614
rect 6763 3606 6765 3614
rect 6773 3606 6775 3614
rect 6783 3606 6785 3614
rect 6793 3606 6795 3614
rect 6803 3606 6805 3614
rect 762 3604 774 3606
rect 3770 3604 3782 3606
rect 6778 3604 6790 3606
rect 602 3576 604 3584
rect 1444 3576 1446 3584
rect 1818 3576 1820 3584
rect 3821 3577 3884 3583
rect 6484 3576 6486 3584
rect 733 3557 796 3563
rect 1622 3536 1628 3544
rect 6285 3537 6316 3543
rect 6900 3537 6915 3543
rect 850 3516 860 3524
rect 452 3497 467 3503
rect 532 3497 579 3503
rect 1021 3497 1036 3503
rect 1357 3503 1363 3523
rect 1325 3497 1363 3503
rect 1748 3497 1795 3503
rect 2061 3497 2076 3503
rect 2429 3503 2435 3523
rect 2429 3497 2467 3503
rect 2781 3497 2835 3503
rect 3181 3497 3212 3503
rect 3325 3503 3331 3523
rect 4900 3517 4915 3523
rect 3325 3497 3363 3503
rect 4637 3497 4684 3503
rect 5101 3497 5139 3503
rect 5252 3497 5315 3503
rect 5421 3497 5459 3503
rect 5965 3497 5980 3503
rect 6061 3497 6099 3503
rect 6221 3503 6227 3523
rect 6189 3497 6227 3503
rect 6372 3497 6387 3503
rect 6509 3503 6515 3523
rect 7460 3516 7468 3524
rect 6468 3497 6483 3503
rect 6509 3497 6547 3503
rect 6660 3497 6675 3503
rect 7140 3497 7155 3503
rect 7341 3497 7356 3503
rect 7444 3497 7459 3503
rect 1101 3477 1124 3483
rect 1116 3472 1124 3477
rect 2077 3477 2099 3483
rect 2429 3477 2444 3483
rect 2941 3477 2956 3483
rect 3588 3477 3603 3483
rect 4077 3477 4115 3483
rect 4173 3477 4195 3483
rect 1644 3472 1652 3476
rect 397 3457 435 3463
rect 2205 3457 2243 3463
rect 3997 3457 4035 3463
rect 4109 3457 4115 3477
rect 4733 3477 4755 3483
rect 4957 3477 4979 3483
rect 5181 3477 5196 3483
rect 5236 3477 5331 3483
rect 5373 3477 5395 3483
rect 5565 3477 5587 3483
rect 5805 3477 5843 3483
rect 6036 3477 6051 3483
rect 6445 3477 6467 3483
rect 6605 3477 6643 3483
rect 6733 3483 6739 3496
rect 6733 3477 6819 3483
rect 6852 3477 6883 3483
rect 6989 3477 7036 3483
rect 7197 3477 7235 3483
rect 4141 3457 4163 3463
rect 4141 3437 4147 3457
rect 4820 3456 4828 3464
rect 5021 3457 5036 3463
rect 5204 3457 5219 3463
rect 7229 3457 7235 3477
rect 7277 3477 7292 3483
rect 7357 3477 7372 3483
rect 4394 3436 4396 3444
rect 5652 3436 5656 3444
rect 5876 3436 5880 3444
rect 6692 3436 6694 3444
rect 7172 3436 7174 3444
rect 2266 3414 2278 3416
rect 5274 3414 5286 3416
rect 2251 3406 2253 3414
rect 2261 3406 2263 3414
rect 2271 3406 2273 3414
rect 2281 3406 2283 3414
rect 2291 3406 2293 3414
rect 5259 3406 5261 3414
rect 5269 3406 5271 3414
rect 5279 3406 5281 3414
rect 5289 3406 5291 3414
rect 5299 3406 5301 3414
rect 2266 3404 2278 3406
rect 5274 3404 5286 3406
rect 5060 3376 5062 3384
rect 5188 3376 5190 3384
rect 7373 3377 7388 3383
rect 205 3343 211 3363
rect 1661 3357 1699 3363
rect 1965 3357 2003 3363
rect 2932 3357 2964 3363
rect 2956 3348 2964 3357
rect 3981 3357 4003 3363
rect 4468 3357 4483 3363
rect 173 3337 211 3343
rect 1076 3337 1091 3343
rect 333 3317 364 3323
rect 852 3317 867 3323
rect 925 3317 940 3323
rect 1005 3317 1036 3323
rect 1149 3323 1155 3343
rect 3421 3337 3443 3343
rect 4125 3337 4163 3343
rect 4381 3337 4403 3343
rect 4500 3337 4531 3343
rect 4621 3343 4627 3363
rect 5284 3357 5356 3363
rect 5412 3356 5420 3364
rect 4621 3337 4636 3343
rect 4653 3337 4675 3343
rect 4964 3337 4979 3343
rect 5092 3337 5107 3343
rect 5261 3337 5292 3343
rect 5437 3337 5475 3343
rect 5588 3337 5603 3343
rect 5645 3343 5651 3363
rect 5645 3337 5683 3343
rect 5725 3343 5731 3363
rect 5837 3357 5875 3363
rect 6861 3357 6892 3363
rect 6948 3356 6956 3364
rect 5725 3337 5763 3343
rect 5972 3337 5987 3343
rect 1140 3317 1155 3323
rect 1197 3317 1235 3323
rect 1069 3297 1075 3316
rect 1197 3297 1203 3317
rect 1517 3317 1532 3323
rect 1540 3317 1571 3323
rect 2781 3317 2796 3323
rect 2916 3317 2931 3323
rect 3117 3317 3171 3323
rect 3293 3317 3308 3323
rect 3428 3317 3459 3323
rect 3581 3317 3596 3323
rect 4029 3317 4060 3323
rect 4429 3317 4467 3323
rect 4740 3317 4755 3323
rect 4765 3317 4780 3323
rect 5901 3317 5923 3323
rect 6040 3317 6076 3323
rect 6365 3323 6371 3343
rect 6429 3337 6451 3343
rect 6973 3337 6988 3343
rect 6996 3337 7027 3343
rect 7220 3337 7235 3343
rect 7476 3337 7507 3343
rect 6164 3317 6200 3323
rect 6365 3317 6387 3323
rect 6669 3317 6691 3323
rect 6996 3317 7011 3323
rect 3186 3296 3196 3304
rect 406 3276 412 3284
rect 1796 3276 1802 3284
rect 2602 3276 2604 3284
rect 4180 3277 4195 3283
rect 6308 3276 6312 3284
rect 1492 3236 1494 3244
rect 3044 3236 3046 3244
rect 3556 3236 3558 3244
rect 4330 3236 4332 3244
rect 4714 3236 4716 3244
rect 5892 3236 5894 3244
rect 6772 3237 6835 3243
rect 762 3214 774 3216
rect 3770 3214 3782 3216
rect 6778 3214 6790 3216
rect 747 3206 749 3214
rect 757 3206 759 3214
rect 767 3206 769 3214
rect 777 3206 779 3214
rect 787 3206 789 3214
rect 3755 3206 3757 3214
rect 3765 3206 3767 3214
rect 3775 3206 3777 3214
rect 3785 3206 3787 3214
rect 3795 3206 3797 3214
rect 6763 3206 6765 3214
rect 6773 3206 6775 3214
rect 6783 3206 6785 3214
rect 6793 3206 6795 3214
rect 6803 3206 6805 3214
rect 762 3204 774 3206
rect 3770 3204 3782 3206
rect 6778 3204 6790 3206
rect 2106 3176 2108 3184
rect 2740 3176 2742 3184
rect 4874 3176 4876 3184
rect 4996 3176 4998 3184
rect 7284 3156 7288 3164
rect 644 3136 646 3144
rect 3030 3136 3036 3144
rect 3108 3136 3110 3144
rect 4266 3136 4268 3144
rect 6426 3136 6428 3144
rect 580 3116 588 3124
rect 1261 3103 1267 3123
rect 1229 3097 1267 3103
rect 1437 3097 1468 3103
rect 1917 3097 1932 3103
rect 2068 3097 2083 3103
rect 2596 3097 2611 3103
rect 3133 3103 3139 3123
rect 4756 3116 4764 3124
rect 4813 3117 4851 3123
rect 3133 3097 3171 3103
rect 3188 3097 3235 3103
rect 3396 3097 3411 3103
rect 3661 3097 3708 3103
rect 3844 3097 3859 3103
rect 4029 3097 4044 3103
rect 4404 3097 4435 3103
rect 5021 3103 5027 3123
rect 5021 3097 5059 3103
rect 5229 3097 5331 3103
rect 5405 3097 5420 3103
rect 5517 3103 5523 3123
rect 5508 3097 5523 3103
rect 5661 3103 5667 3123
rect 5629 3097 5667 3103
rect 5805 3103 5811 3123
rect 7133 3117 7155 3123
rect 5805 3097 5843 3103
rect 6077 3097 6092 3103
rect 6132 3097 6147 3103
rect 6717 3097 6732 3103
rect 6868 3097 6931 3103
rect 7140 3097 7155 3103
rect 7444 3097 7459 3103
rect 100 3077 131 3083
rect 733 3077 835 3083
rect 925 3077 963 3083
rect 29 3057 67 3063
rect 733 3057 739 3077
rect 756 3057 819 3063
rect 957 3057 963 3077
rect 1933 3077 1948 3083
rect 1933 3057 1939 3077
rect 2173 3077 2211 3083
rect 2205 3057 2211 3077
rect 2508 3077 2531 3083
rect 2573 3077 2595 3083
rect 2508 3072 2516 3077
rect 2701 3077 2716 3083
rect 3204 3077 3219 3083
rect 3492 3077 3507 3083
rect 3916 3077 3932 3083
rect 3965 3077 3980 3083
rect 4157 3077 4179 3083
rect 4372 3077 4387 3083
rect 4717 3077 4739 3083
rect 4893 3077 4915 3083
rect 4957 3077 4979 3083
rect 5421 3077 5443 3083
rect 5565 3077 5603 3083
rect 5709 3077 5731 3083
rect 5917 3077 5939 3083
rect 6020 3077 6035 3083
rect 6061 3077 6076 3083
rect 6324 3077 6339 3083
rect 6493 3077 6515 3083
rect 6564 3077 6595 3083
rect 6637 3077 6675 3083
rect 6701 3077 6716 3083
rect 2861 3057 2876 3063
rect 3645 3057 3692 3063
rect 3981 3057 4003 3063
rect 4612 3057 4627 3063
rect 4660 3057 4675 3063
rect 5124 3056 5132 3064
rect 5268 3057 5347 3063
rect 6637 3057 6643 3077
rect 7005 3077 7020 3083
rect 7117 3077 7132 3083
rect 7172 3077 7203 3083
rect 5492 3036 5494 3044
rect 6212 3037 6227 3043
rect 6836 3036 6840 3044
rect 7380 3036 7382 3044
rect 7498 3036 7500 3044
rect 2266 3014 2278 3016
rect 5274 3014 5286 3016
rect 2251 3006 2253 3014
rect 2261 3006 2263 3014
rect 2271 3006 2273 3014
rect 2281 3006 2283 3014
rect 2291 3006 2293 3014
rect 5259 3006 5261 3014
rect 5269 3006 5271 3014
rect 5279 3006 5281 3014
rect 5289 3006 5291 3014
rect 5299 3006 5301 3014
rect 2266 3004 2278 3006
rect 5274 3004 5286 3006
rect 733 2977 748 2983
rect 1290 2976 1292 2984
rect 5508 2976 5510 2984
rect 253 2957 291 2963
rect 804 2957 819 2963
rect 1021 2957 1036 2963
rect 1453 2957 1491 2963
rect 308 2937 323 2943
rect 1437 2937 1468 2943
rect 1757 2943 1763 2963
rect 2109 2957 2147 2963
rect 1725 2937 1763 2943
rect 2541 2937 2572 2943
rect 2781 2937 2803 2943
rect 3597 2937 3619 2943
rect 3996 2937 4020 2943
rect 4340 2937 4355 2943
rect 4381 2937 4403 2943
rect 4653 2937 4691 2943
rect 4788 2937 4819 2943
rect 5021 2943 5027 2963
rect 4909 2937 4931 2943
rect 5021 2937 5036 2943
rect 5053 2937 5075 2943
rect 100 2917 131 2923
rect 349 2917 364 2923
rect 621 2917 636 2923
rect 909 2917 924 2923
rect 1252 2917 1267 2923
rect 1508 2917 1523 2923
rect 1588 2917 1635 2923
rect 1956 2917 1987 2923
rect 2564 2917 2579 2923
rect 2829 2917 2844 2923
rect 3076 2917 3091 2923
rect 3620 2917 3635 2923
rect 3741 2917 3804 2923
rect 3924 2917 3939 2923
rect 4532 2917 4563 2923
rect 1196 2904 1204 2914
rect 3636 2896 3644 2904
rect 2205 2877 2268 2883
rect 4621 2883 4627 2923
rect 4932 2917 4947 2923
rect 4980 2917 4995 2923
rect 5373 2923 5379 2963
rect 5613 2957 5619 2983
rect 5658 2976 5660 2984
rect 6692 2976 6694 2984
rect 6932 2977 6974 2983
rect 5716 2956 5724 2964
rect 6109 2957 6140 2963
rect 6189 2957 6227 2963
rect 6237 2957 6252 2963
rect 6285 2957 6300 2963
rect 6580 2957 6595 2963
rect 5597 2937 5635 2943
rect 5741 2937 5756 2943
rect 6077 2937 6099 2943
rect 7005 2937 7036 2943
rect 7108 2937 7139 2943
rect 5373 2917 5388 2923
rect 6429 2917 6451 2923
rect 6541 2917 6579 2923
rect 6756 2917 6819 2923
rect 7373 2923 7379 2943
rect 7492 2937 7507 2943
rect 7293 2917 7347 2923
rect 7373 2917 7432 2923
rect 4733 2897 4771 2903
rect 5570 2896 5580 2904
rect 4621 2877 4636 2883
rect 5821 2883 5827 2903
rect 7101 2897 7123 2903
rect 7341 2897 7347 2917
rect 6556 2884 6564 2888
rect 5805 2877 5827 2883
rect 2762 2856 2764 2864
rect 3498 2856 3500 2864
rect 410 2836 412 2844
rect 506 2836 508 2844
rect 1364 2836 1366 2844
rect 1658 2836 1660 2844
rect 4858 2836 4860 2844
rect 4948 2836 4950 2844
rect 762 2814 774 2816
rect 3770 2814 3782 2816
rect 6778 2814 6790 2816
rect 747 2806 749 2814
rect 757 2806 759 2814
rect 767 2806 769 2814
rect 777 2806 779 2814
rect 787 2806 789 2814
rect 3755 2806 3757 2814
rect 3765 2806 3767 2814
rect 3775 2806 3777 2814
rect 3785 2806 3787 2814
rect 3795 2806 3797 2814
rect 6763 2806 6765 2814
rect 6773 2806 6775 2814
rect 6783 2806 6785 2814
rect 6793 2806 6795 2814
rect 6803 2806 6805 2814
rect 762 2804 774 2806
rect 3770 2804 3782 2806
rect 6778 2804 6790 2806
rect 458 2776 460 2784
rect 554 2776 556 2784
rect 922 2776 924 2784
rect 1876 2776 1878 2784
rect 3540 2776 3542 2784
rect 1914 2736 1916 2744
rect 4045 2737 4068 2743
rect 4957 2737 4979 2743
rect 493 2697 508 2703
rect 964 2697 979 2703
rect 989 2697 1020 2703
rect 1316 2697 1331 2703
rect 1508 2697 1523 2703
rect 1668 2697 1683 2703
rect 1997 2697 2012 2703
rect 285 2677 316 2683
rect 941 2683 947 2696
rect 2781 2703 2787 2723
rect 4973 2717 4979 2737
rect 5837 2737 5852 2743
rect 6596 2737 6611 2743
rect 2781 2697 2804 2703
rect 2796 2692 2804 2697
rect 2845 2697 2860 2703
rect 2884 2697 2899 2703
rect 3037 2697 3052 2703
rect 3213 2697 3228 2703
rect 3588 2697 3603 2703
rect 4724 2697 4755 2703
rect 4845 2697 4860 2703
rect 4893 2697 4924 2703
rect 5309 2703 5315 2723
rect 5956 2716 5964 2724
rect 6669 2717 6691 2723
rect 7188 2716 7196 2724
rect 5213 2697 5315 2703
rect 5341 2697 5356 2703
rect 5868 2703 5876 2708
rect 5868 2697 5907 2703
rect 5917 2697 5932 2703
rect 6132 2697 6147 2703
rect 6189 2697 6204 2703
rect 6909 2697 6931 2703
rect 6989 2697 7011 2703
rect 7197 2697 7212 2703
rect 7485 2697 7507 2703
rect 941 2677 956 2683
rect 1245 2677 1260 2683
rect 1300 2677 1315 2683
rect 1773 2677 1795 2683
rect 2476 2677 2500 2683
rect 3060 2677 3075 2683
rect 3380 2677 3411 2683
rect 3661 2677 3676 2683
rect 4685 2677 4707 2683
rect 5044 2677 5059 2683
rect 5284 2677 5315 2683
rect 5357 2677 5395 2683
rect 5924 2677 5939 2683
rect 6269 2677 6307 2683
rect 6365 2677 6403 2683
rect 6477 2677 6499 2683
rect 7213 2677 7235 2683
rect 349 2657 387 2663
rect 1277 2657 1292 2663
rect 3357 2657 3395 2663
rect 3741 2657 3756 2663
rect 5812 2657 5832 2663
rect 5476 2636 5478 2644
rect 5672 2636 5676 2644
rect 5748 2636 5750 2644
rect 6948 2636 6950 2644
rect 2266 2614 2278 2616
rect 5274 2614 5286 2616
rect 2251 2606 2253 2614
rect 2261 2606 2263 2614
rect 2271 2606 2273 2614
rect 2281 2606 2283 2614
rect 2291 2606 2293 2614
rect 5259 2606 5261 2614
rect 5269 2606 5271 2614
rect 5279 2606 5281 2614
rect 5289 2606 5291 2614
rect 5299 2606 5301 2614
rect 2266 2604 2278 2606
rect 5274 2604 5286 2606
rect 5896 2576 5900 2584
rect 6692 2576 6694 2584
rect 6836 2577 6910 2583
rect 317 2557 355 2563
rect 621 2557 659 2563
rect 669 2557 716 2563
rect 957 2557 995 2563
rect 3533 2557 3555 2563
rect 4125 2557 4147 2563
rect 4669 2557 4691 2563
rect 4701 2557 4739 2563
rect 996 2537 1011 2543
rect 1421 2537 1443 2543
rect 2493 2537 2508 2543
rect 2749 2537 2764 2543
rect 3101 2537 3116 2543
rect 253 2517 268 2523
rect 1053 2523 1059 2536
rect 1037 2517 1059 2523
rect 1085 2517 1116 2523
rect 1629 2517 1644 2523
rect 2077 2517 2115 2523
rect 1901 2497 1939 2503
rect 2109 2497 2115 2517
rect 2148 2517 2195 2523
rect 2221 2517 2323 2523
rect 2221 2497 2227 2517
rect 2452 2517 2467 2523
rect 2749 2517 2787 2523
rect 2749 2497 2755 2517
rect 3012 2517 3027 2523
rect 3053 2517 3091 2523
rect 3053 2497 3059 2517
rect 3165 2523 3171 2543
rect 4068 2537 4092 2543
rect 4445 2537 4467 2543
rect 4509 2537 4531 2543
rect 4669 2537 4684 2543
rect 4916 2537 4931 2543
rect 5181 2543 5187 2563
rect 5725 2557 5763 2563
rect 5773 2557 5811 2563
rect 5149 2537 5187 2543
rect 5220 2537 5315 2543
rect 5325 2537 5340 2543
rect 5453 2537 5475 2543
rect 5517 2537 5539 2543
rect 5613 2537 5635 2543
rect 5693 2537 5715 2543
rect 5933 2537 5948 2543
rect 6045 2537 6067 2543
rect 6189 2537 6243 2543
rect 6317 2537 6355 2543
rect 6596 2537 6611 2543
rect 6724 2537 6739 2543
rect 6765 2537 6780 2543
rect 6941 2537 6995 2543
rect 7460 2537 7475 2543
rect 3108 2517 3171 2523
rect 3213 2517 3251 2523
rect 3213 2497 3219 2517
rect 3533 2517 3548 2523
rect 3604 2517 3619 2523
rect 4308 2517 4323 2523
rect 4573 2517 4611 2523
rect 3684 2497 3699 2503
rect 4573 2497 4579 2517
rect 4765 2517 4787 2523
rect 4973 2517 5011 2523
rect 5069 2517 5084 2523
rect 5373 2517 5411 2523
rect 4861 2497 4876 2503
rect 5069 2497 5091 2503
rect 5101 2497 5116 2503
rect 5341 2497 5356 2503
rect 5405 2497 5411 2517
rect 5965 2517 6003 2523
rect 6509 2517 6547 2523
rect 6580 2517 6595 2523
rect 6948 2517 6972 2523
rect 7021 2517 7052 2523
rect 7108 2517 7123 2523
rect 7149 2517 7187 2523
rect 5581 2497 5596 2503
rect 6018 2496 6028 2504
rect 6061 2497 6099 2503
rect 6109 2497 6147 2503
rect 7149 2497 7155 2517
rect 7277 2517 7299 2523
rect 7501 2517 7516 2523
rect 7517 2497 7532 2503
rect 1140 2476 1142 2484
rect 1876 2476 1878 2484
rect 3636 2477 3651 2483
rect 3910 2476 3916 2484
rect 5434 2476 5436 2484
rect 7396 2476 7400 2484
rect 7124 2456 7126 2464
rect 1482 2436 1484 2444
rect 1604 2436 1606 2444
rect 3188 2436 3190 2444
rect 5012 2436 5014 2444
rect 5652 2436 5654 2444
rect 6260 2436 6262 2444
rect 762 2414 774 2416
rect 3770 2414 3782 2416
rect 6778 2414 6790 2416
rect 747 2406 749 2414
rect 757 2406 759 2414
rect 767 2406 769 2414
rect 777 2406 779 2414
rect 787 2406 789 2414
rect 3755 2406 3757 2414
rect 3765 2406 3767 2414
rect 3775 2406 3777 2414
rect 3785 2406 3787 2414
rect 3795 2406 3797 2414
rect 6763 2406 6765 2414
rect 6773 2406 6775 2414
rect 6783 2406 6785 2414
rect 6793 2406 6795 2414
rect 6803 2406 6805 2414
rect 762 2404 774 2406
rect 3770 2404 3782 2406
rect 6778 2404 6790 2406
rect 1572 2376 1574 2384
rect 5194 2376 5196 2384
rect 3174 2336 3180 2344
rect 3340 2337 3363 2343
rect 4973 2337 5004 2343
rect 5716 2337 5731 2343
rect 5978 2336 5980 2344
rect 6733 2337 6796 2343
rect 1332 2316 1340 2324
rect 365 2297 387 2303
rect 493 2297 508 2303
rect 621 2297 636 2303
rect 845 2297 860 2303
rect 1357 2303 1363 2323
rect 1357 2297 1395 2303
rect 1533 2303 1539 2323
rect 1492 2297 1507 2303
rect 1533 2297 1556 2303
rect 1548 2292 1556 2297
rect 1597 2297 1651 2303
rect 1661 2297 1676 2303
rect 1796 2297 1811 2303
rect 2100 2297 2115 2303
rect 2445 2303 2451 2323
rect 2413 2297 2451 2303
rect 3101 2297 3116 2303
rect 3300 2297 3315 2303
rect 3700 2297 3715 2303
rect 3773 2297 3859 2303
rect 3869 2297 3884 2303
rect 173 2277 188 2283
rect 1421 2277 1436 2283
rect 1773 2277 1795 2283
rect 3020 2277 3044 2283
rect 3693 2277 3708 2283
rect 445 2257 467 2263
rect 1668 2257 1683 2263
rect 3453 2257 3475 2263
rect 3773 2263 3779 2297
rect 4269 2303 4275 2323
rect 6980 2316 6984 2324
rect 4269 2297 4307 2303
rect 4381 2297 4403 2303
rect 4580 2297 4595 2303
rect 4205 2277 4227 2283
rect 4429 2277 4467 2283
rect 3757 2257 3779 2263
rect 4429 2257 4435 2277
rect 4532 2277 4547 2283
rect 4516 2256 4524 2264
rect 4541 2257 4547 2277
rect 4669 2283 4675 2303
rect 4861 2297 4915 2303
rect 4669 2277 4739 2283
rect 4557 2257 4572 2263
rect 4733 2257 4739 2277
rect 4909 2277 4915 2297
rect 5124 2297 5139 2303
rect 5149 2297 5187 2303
rect 5261 2297 5324 2303
rect 5805 2297 5820 2303
rect 5837 2297 5875 2303
rect 5956 2297 5971 2303
rect 6285 2297 6307 2303
rect 6365 2297 6387 2303
rect 6484 2297 6499 2303
rect 6653 2297 6668 2303
rect 7204 2297 7235 2303
rect 7252 2297 7299 2303
rect 7309 2297 7363 2303
rect 7421 2297 7436 2303
rect 5053 2277 5084 2283
rect 5101 2277 5123 2283
rect 5581 2277 5619 2283
rect 5645 2277 5676 2283
rect 6045 2277 6060 2283
rect 6077 2277 6131 2283
rect 6413 2277 6444 2283
rect 7309 2277 7315 2297
rect 7421 2277 7427 2297
rect 7492 2297 7507 2303
rect 7469 2277 7484 2283
rect 5949 2257 5964 2263
rect 6221 2257 6236 2263
rect 5300 2237 5324 2243
rect 6154 2236 6156 2244
rect 2266 2214 2278 2216
rect 5274 2214 5286 2216
rect 2251 2206 2253 2214
rect 2261 2206 2263 2214
rect 2271 2206 2273 2214
rect 2281 2206 2283 2214
rect 2291 2206 2293 2214
rect 5259 2206 5261 2214
rect 5269 2206 5271 2214
rect 5279 2206 5281 2214
rect 5289 2206 5291 2214
rect 5299 2206 5301 2214
rect 2266 2204 2278 2206
rect 5274 2204 5286 2206
rect 458 2176 460 2184
rect 554 2176 556 2184
rect 125 2157 147 2163
rect 1117 2157 1155 2163
rect 3101 2157 3139 2163
rect 3725 2157 3811 2163
rect 4557 2163 4563 2183
rect 5866 2176 5868 2184
rect 7476 2176 7480 2184
rect 4557 2157 4579 2163
rect 4765 2157 4803 2163
rect 5156 2156 5164 2164
rect 6436 2156 6444 2164
rect 7053 2157 7068 2163
rect 29 2137 44 2143
rect 484 2137 499 2143
rect 1101 2143 1107 2156
rect 1021 2137 1043 2143
rect 1085 2137 1107 2143
rect 1388 2143 1396 2148
rect 1388 2137 1411 2143
rect 2925 2137 2956 2143
rect 132 2117 147 2123
rect 509 2117 540 2123
rect 637 2117 675 2123
rect 429 2097 444 2103
rect 637 2097 643 2117
rect 692 2117 707 2123
rect 1917 2117 1955 2123
rect 1684 2096 1692 2104
rect 1949 2097 1955 2117
rect 2237 2117 2300 2123
rect 2525 2117 2563 2123
rect 1972 2096 1980 2104
rect 2557 2097 2563 2117
rect 2797 2117 2835 2123
rect 2829 2097 2835 2117
rect 2925 2117 2931 2137
rect 2996 2137 3011 2143
rect 3661 2137 3676 2143
rect 4557 2137 4572 2143
rect 3668 2117 3683 2123
rect 4557 2117 4563 2137
rect 4589 2137 4611 2143
rect 4788 2137 4819 2143
rect 5085 2137 5123 2143
rect 5533 2137 5555 2143
rect 5805 2137 5827 2143
rect 6109 2137 6131 2143
rect 6301 2137 6323 2143
rect 6788 2137 6851 2143
rect 7181 2143 7187 2163
rect 7181 2137 7219 2143
rect 4941 2117 4956 2123
rect 5220 2117 5331 2123
rect 5421 2117 5475 2123
rect 5597 2117 5635 2123
rect 5725 2117 5763 2123
rect 3725 2097 3772 2103
rect 3796 2097 3811 2103
rect 4708 2097 4723 2103
rect 5037 2097 5059 2103
rect 5597 2097 5603 2117
rect 5757 2097 5763 2117
rect 6189 2117 6243 2123
rect 6237 2097 6243 2117
rect 6365 2117 6403 2123
rect 6557 2117 6572 2123
rect 7261 2117 7283 2123
rect 7293 2117 7331 2123
rect 6548 2096 6556 2104
rect 6605 2097 6620 2103
rect 106 2076 108 2084
rect 3302 2076 3308 2084
rect 4006 2076 4012 2084
rect 6637 2077 6652 2083
rect 2858 2036 2860 2044
rect 5476 2036 5478 2044
rect 5786 2036 5788 2044
rect 762 2014 774 2016
rect 3770 2014 3782 2016
rect 6778 2014 6790 2016
rect 747 2006 749 2014
rect 757 2006 759 2014
rect 767 2006 769 2014
rect 777 2006 779 2014
rect 787 2006 789 2014
rect 3755 2006 3757 2014
rect 3765 2006 3767 2014
rect 3775 2006 3777 2014
rect 3785 2006 3787 2014
rect 3795 2006 3797 2014
rect 6763 2006 6765 2014
rect 6773 2006 6775 2014
rect 6783 2006 6785 2014
rect 6793 2006 6795 2014
rect 6803 2006 6805 2014
rect 762 2004 774 2006
rect 3770 2004 3782 2006
rect 6778 2004 6790 2006
rect 1524 1976 1526 1984
rect 3588 1976 3590 1984
rect 4532 1976 4534 1984
rect 5156 1976 5160 1984
rect 5962 1976 5964 1984
rect 6324 1976 6326 1984
rect 650 1956 652 1964
rect 4102 1936 4108 1944
rect 4644 1937 4659 1943
rect 253 1903 259 1923
rect 1005 1917 1043 1923
rect 1284 1916 1292 1924
rect 1924 1916 1932 1924
rect 253 1897 291 1903
rect 381 1897 396 1903
rect 580 1897 627 1903
rect 1325 1903 1331 1916
rect 1293 1897 1331 1903
rect 1949 1903 1955 1923
rect 1908 1897 1923 1903
rect 1949 1897 1987 1903
rect 2276 1897 2387 1903
rect 2445 1897 2460 1903
rect 2813 1903 2819 1923
rect 3332 1916 3340 1924
rect 3652 1916 3660 1924
rect 4397 1917 4412 1923
rect 4477 1917 4492 1923
rect 4589 1917 4636 1923
rect 5620 1917 5635 1923
rect 6372 1916 6380 1924
rect 2781 1897 2819 1903
rect 3172 1897 3187 1903
rect 3300 1897 3331 1903
rect 5005 1897 5043 1903
rect 5421 1897 5459 1903
rect 6285 1897 6300 1903
rect 6333 1897 6348 1903
rect 1613 1877 1651 1883
rect 460 1864 468 1872
rect 1492 1857 1507 1863
rect 1645 1857 1651 1877
rect 2356 1877 2387 1883
rect 4596 1877 4611 1883
rect 2477 1857 2515 1863
rect 4372 1857 4387 1863
rect 4605 1857 4611 1877
rect 4925 1877 4947 1883
rect 5069 1877 5107 1883
rect 5245 1877 5331 1883
rect 5485 1877 5507 1883
rect 5524 1877 5555 1883
rect 5773 1877 5795 1883
rect 5773 1864 5779 1877
rect 5981 1877 6019 1883
rect 6029 1877 6044 1883
rect 5373 1857 5395 1863
rect 6029 1857 6035 1877
rect 6205 1877 6220 1883
rect 6756 1877 6835 1883
rect 6861 1877 6876 1883
rect 7012 1877 7027 1883
rect 7181 1877 7212 1883
rect 7252 1877 7283 1883
rect 7412 1877 7427 1883
rect 7293 1857 7331 1863
rect 7421 1857 7427 1877
rect 7437 1857 7452 1863
rect 2244 1836 2246 1844
rect 4580 1836 4582 1844
rect 4660 1836 4662 1844
rect 4820 1836 4822 1844
rect 5604 1836 5606 1844
rect 6132 1836 6134 1844
rect 7124 1836 7128 1844
rect 2266 1814 2278 1816
rect 5274 1814 5286 1816
rect 2251 1806 2253 1814
rect 2261 1806 2263 1814
rect 2271 1806 2273 1814
rect 2281 1806 2283 1814
rect 2291 1806 2293 1814
rect 5259 1806 5261 1814
rect 5269 1806 5271 1814
rect 5279 1806 5281 1814
rect 5289 1806 5291 1814
rect 5299 1806 5301 1814
rect 2266 1804 2278 1806
rect 5274 1804 5286 1806
rect 2676 1776 2678 1784
rect 2890 1776 2892 1784
rect 3178 1776 3180 1784
rect 3226 1776 3228 1784
rect 4138 1776 4140 1784
rect 4525 1777 4540 1783
rect 4730 1776 4732 1784
rect 6468 1776 6470 1784
rect 6996 1776 6998 1784
rect 253 1757 291 1763
rect 413 1757 451 1763
rect 1236 1757 1251 1763
rect 1261 1757 1276 1763
rect 1364 1757 1379 1763
rect 3757 1757 3843 1763
rect 4269 1757 4284 1763
rect 4445 1757 4467 1763
rect 349 1737 380 1743
rect 893 1737 915 1743
rect 1037 1737 1059 1743
rect 1268 1737 1299 1743
rect 2093 1737 2115 1743
rect 2253 1737 2316 1743
rect 493 1717 531 1723
rect 525 1697 531 1717
rect 820 1717 867 1723
rect 916 1717 931 1723
rect 1309 1717 1324 1723
rect 1677 1717 1708 1723
rect 1821 1717 1875 1723
rect 2013 1717 2044 1723
rect 2116 1717 2131 1723
rect 2925 1723 2931 1743
rect 4045 1737 4115 1743
rect 4157 1737 4188 1743
rect 4445 1743 4451 1757
rect 4548 1757 4563 1763
rect 6148 1756 6156 1764
rect 6836 1756 6844 1764
rect 6932 1756 6940 1764
rect 4413 1737 4451 1743
rect 4909 1737 4931 1743
rect 5069 1737 5107 1743
rect 5197 1737 5219 1743
rect 5700 1737 5715 1743
rect 5764 1737 5779 1743
rect 5837 1737 5875 1743
rect 6260 1737 6307 1743
rect 6356 1737 6387 1743
rect 6541 1737 6556 1743
rect 6884 1737 6915 1743
rect 7028 1737 7043 1743
rect 2916 1717 2931 1723
rect 4253 1717 4284 1723
rect 4573 1723 4579 1736
rect 4525 1717 4579 1723
rect 932 1696 940 1704
rect 2146 1696 2156 1704
rect 2685 1697 2707 1703
rect 2797 1697 2819 1703
rect 2957 1697 2979 1703
rect 3092 1697 3107 1703
rect 3149 1697 3171 1703
rect 3828 1697 3843 1703
rect 4109 1697 4131 1703
rect 4525 1697 4531 1717
rect 4829 1717 4867 1723
rect 4861 1697 4867 1717
rect 4989 1717 5004 1723
rect 5741 1717 5763 1723
rect 5917 1717 5955 1723
rect 6045 1717 6083 1723
rect 5028 1696 5036 1704
rect 5204 1697 5219 1703
rect 5444 1696 5452 1704
rect 5917 1697 5923 1717
rect 6669 1717 6707 1723
rect 7012 1717 7027 1723
rect 7149 1717 7164 1723
rect 7437 1717 7475 1723
rect 1876 1676 1878 1684
rect 3494 1676 3500 1684
rect 5386 1676 5388 1684
rect 7204 1676 7208 1684
rect 1466 1656 1468 1664
rect 1754 1636 1756 1644
rect 762 1614 774 1616
rect 3770 1614 3782 1616
rect 6778 1614 6790 1616
rect 747 1606 749 1614
rect 757 1606 759 1614
rect 767 1606 769 1614
rect 777 1606 779 1614
rect 787 1606 789 1614
rect 3755 1606 3757 1614
rect 3765 1606 3767 1614
rect 3775 1606 3777 1614
rect 3785 1606 3787 1614
rect 3795 1606 3797 1614
rect 6763 1606 6765 1614
rect 6773 1606 6775 1614
rect 6783 1606 6785 1614
rect 6793 1606 6795 1614
rect 6803 1606 6805 1614
rect 762 1604 774 1606
rect 3770 1604 3782 1606
rect 6778 1604 6790 1606
rect 1060 1576 1062 1584
rect 1156 1576 1158 1584
rect 2253 1577 2300 1583
rect 4164 1576 4166 1584
rect 4922 1576 4924 1584
rect 7396 1576 7400 1584
rect 1994 1536 1996 1544
rect 2180 1537 2211 1543
rect 173 1517 211 1523
rect 109 1497 131 1503
rect 125 1484 131 1497
rect 340 1497 355 1503
rect 893 1497 908 1503
rect 1325 1497 1340 1503
rect 1421 1497 1436 1503
rect 1485 1503 1491 1523
rect 2205 1517 2211 1537
rect 2388 1537 2403 1543
rect 2413 1537 2428 1543
rect 2452 1537 2467 1543
rect 2964 1536 2966 1544
rect 3284 1537 3299 1543
rect 4093 1537 4124 1543
rect 4506 1536 4508 1544
rect 7220 1536 7224 1544
rect 2349 1517 2371 1523
rect 3092 1516 3100 1524
rect 3197 1517 3219 1523
rect 3252 1517 3267 1523
rect 3757 1517 3804 1523
rect 3812 1517 3843 1523
rect 3988 1514 3992 1522
rect 4116 1517 4131 1523
rect 4708 1517 4723 1523
rect 4980 1517 4995 1523
rect 5428 1517 5443 1523
rect 5508 1516 5518 1524
rect 5684 1516 5692 1524
rect 1485 1497 1516 1503
rect 1668 1497 1683 1503
rect 1965 1497 1987 1503
rect 2797 1497 2844 1503
rect 3220 1497 3235 1503
rect 3508 1497 3523 1503
rect 3876 1497 3891 1503
rect 4013 1497 4028 1503
rect 4589 1497 4620 1503
rect 4884 1497 4899 1503
rect 5021 1497 5036 1503
rect 5101 1497 5116 1503
rect 5693 1497 5708 1503
rect 5821 1497 5836 1503
rect 5869 1497 5891 1503
rect 6045 1497 6067 1503
rect 6157 1497 6195 1503
rect 6340 1497 6355 1503
rect 6580 1497 6595 1503
rect 6781 1497 6860 1503
rect 7165 1497 7180 1503
rect 93 1477 108 1483
rect 532 1477 563 1483
rect 685 1477 700 1483
rect 1204 1477 1235 1483
rect 2813 1477 2828 1483
rect 3892 1477 3907 1483
rect 3917 1477 3948 1483
rect 4029 1477 4044 1483
rect 4205 1477 4243 1483
rect 4308 1477 4323 1483
rect 4445 1477 4467 1483
rect 4525 1477 4563 1483
rect 4669 1477 4691 1483
rect 4861 1477 4883 1483
rect 4941 1477 4963 1483
rect 5037 1477 5059 1483
rect 5197 1477 5219 1483
rect 5469 1477 5491 1483
rect 5613 1477 5651 1483
rect 5709 1477 5731 1483
rect 5748 1477 5763 1483
rect 5828 1477 5859 1483
rect 5933 1477 5948 1483
rect 6068 1477 6083 1483
rect 6429 1477 6444 1483
rect 6557 1477 6572 1483
rect 6580 1477 6611 1483
rect 6765 1477 6780 1483
rect 6868 1477 6883 1483
rect 6925 1477 6963 1483
rect 29 1457 67 1463
rect 477 1457 515 1463
rect 589 1457 627 1463
rect 701 1457 739 1463
rect 1476 1456 1484 1464
rect 3933 1457 3964 1463
rect 4020 1457 4035 1463
rect 4349 1457 4371 1463
rect 4605 1457 4627 1463
rect 4701 1457 4723 1463
rect 5261 1457 5347 1463
rect 5437 1457 5459 1463
rect 5805 1457 5843 1463
rect 6221 1457 6236 1463
rect 6532 1456 6540 1464
rect 6628 1456 6636 1464
rect 6925 1457 6931 1477
rect 7165 1477 7171 1497
rect 7300 1477 7315 1483
rect 7453 1477 7468 1483
rect 7549 1477 7564 1483
rect 5396 1436 5400 1444
rect 6692 1436 6694 1444
rect 7060 1436 7064 1444
rect 2266 1414 2278 1416
rect 5274 1414 5286 1416
rect 2251 1406 2253 1414
rect 2261 1406 2263 1414
rect 2271 1406 2273 1414
rect 2281 1406 2283 1414
rect 2291 1406 2293 1414
rect 5259 1406 5261 1414
rect 5269 1406 5271 1414
rect 5279 1406 5281 1414
rect 5289 1406 5291 1414
rect 5299 1406 5301 1414
rect 2266 1404 2278 1406
rect 5274 1404 5286 1406
rect 2388 1376 2390 1384
rect 2660 1376 2662 1384
rect 2708 1376 2710 1384
rect 2906 1376 2908 1384
rect 2964 1376 2966 1384
rect 3172 1376 3174 1384
rect 3258 1376 3260 1384
rect 4157 1377 4172 1383
rect 4242 1377 4268 1383
rect 4292 1377 4307 1383
rect 5930 1376 5932 1384
rect 6740 1376 6744 1384
rect 1085 1357 1123 1363
rect 2548 1356 2556 1364
rect 4717 1357 4755 1363
rect 4868 1357 4883 1363
rect 188 1337 212 1343
rect 2221 1337 2284 1343
rect 2573 1337 2611 1343
rect 2628 1337 2643 1343
rect 2932 1337 2947 1343
rect 3085 1337 3123 1343
rect 3140 1337 3155 1343
rect 3229 1337 3244 1343
rect 4164 1337 4211 1343
rect 4893 1343 4899 1363
rect 4893 1337 4931 1343
rect 5053 1337 5075 1343
rect 5229 1337 5315 1343
rect 5460 1337 5475 1343
rect 5549 1337 5571 1343
rect 5645 1337 5667 1343
rect 5789 1337 5827 1343
rect 6125 1343 6131 1356
rect 6125 1337 6147 1343
rect 6269 1337 6307 1343
rect 6541 1343 6547 1363
rect 6628 1357 6652 1363
rect 6516 1337 6547 1343
rect 6685 1343 6691 1356
rect 6877 1343 6883 1356
rect 6685 1337 6707 1343
rect 6797 1337 6883 1343
rect 6989 1337 7027 1343
rect 100 1317 131 1323
rect 692 1317 707 1323
rect 765 1317 812 1323
rect 1197 1317 1251 1323
rect 1284 1317 1299 1323
rect 2205 1317 2220 1323
rect 3476 1317 3507 1323
rect 3540 1317 3555 1323
rect 3844 1317 3859 1323
rect 4340 1317 4355 1323
rect 4413 1317 4428 1323
rect 4493 1317 4515 1323
rect 4781 1317 4803 1323
rect 4989 1317 5027 1323
rect 5588 1317 5619 1323
rect 5725 1317 5763 1323
rect 5949 1317 5971 1323
rect 6109 1317 6124 1323
rect 6381 1317 6403 1323
rect 6461 1317 6483 1323
rect 6893 1317 6931 1323
rect 7021 1317 7027 1337
rect 7277 1337 7315 1343
rect 7309 1324 7315 1337
rect 7421 1343 7427 1363
rect 7412 1337 7427 1343
rect 7188 1317 7219 1323
rect 7348 1317 7363 1323
rect 1508 1296 1516 1304
rect 1668 1296 1676 1304
rect 2397 1297 2419 1303
rect 3444 1296 3452 1304
rect 3508 1296 3516 1304
rect 3604 1297 3619 1303
rect 4109 1297 4124 1303
rect 5332 1296 5342 1304
rect 5588 1297 5603 1303
rect 2588 1284 2596 1288
rect 634 1276 636 1284
rect 2668 1284 2676 1288
rect 2716 1283 2724 1288
rect 2764 1284 2772 1288
rect 2716 1277 2732 1283
rect 2892 1283 2900 1288
rect 2884 1277 2900 1283
rect 2972 1284 2980 1288
rect 3100 1284 3108 1288
rect 3180 1284 3188 1288
rect 3196 1284 3204 1288
rect 3380 1276 3382 1284
rect 7236 1277 7251 1283
rect 7533 1277 7564 1283
rect 1322 1256 1324 1264
rect 1802 1256 1804 1264
rect 3316 1256 3318 1264
rect 4410 1256 4412 1264
rect 1194 1236 1196 1244
rect 762 1214 774 1216
rect 3770 1214 3782 1216
rect 6778 1214 6790 1216
rect 747 1206 749 1214
rect 757 1206 759 1214
rect 767 1206 769 1214
rect 777 1206 779 1214
rect 787 1206 789 1214
rect 3755 1206 3757 1214
rect 3765 1206 3767 1214
rect 3775 1206 3777 1214
rect 3785 1206 3787 1214
rect 3795 1206 3797 1214
rect 6763 1206 6765 1214
rect 6773 1206 6775 1214
rect 6783 1206 6785 1214
rect 6793 1206 6795 1214
rect 6803 1206 6805 1214
rect 762 1204 774 1206
rect 3770 1204 3782 1206
rect 6778 1204 6790 1206
rect 1188 1176 1190 1184
rect 2221 1177 2268 1183
rect 4984 1176 4988 1184
rect 5348 1176 5352 1184
rect 6424 1176 6428 1184
rect 6733 1177 6796 1183
rect 7050 1176 7052 1184
rect 717 1137 780 1143
rect 2093 1137 2124 1143
rect 2372 1137 2387 1143
rect 5485 1137 5500 1143
rect 6301 1137 6316 1143
rect 6596 1137 6611 1143
rect 2813 1117 2828 1123
rect 3261 1117 3276 1123
rect 3453 1117 3491 1123
rect 3757 1117 3859 1123
rect 5949 1117 5971 1123
rect 6052 1116 6056 1124
rect 477 1097 492 1103
rect 1133 1097 1164 1103
rect 1485 1097 1500 1103
rect 1693 1097 1708 1103
rect 1949 1097 1964 1103
rect 2244 1097 2323 1103
rect 2909 1097 2931 1103
rect 3780 1097 3820 1103
rect 4365 1097 4380 1103
rect 4413 1097 4428 1103
rect 5229 1097 5244 1103
rect 5501 1097 5560 1103
rect 644 1077 659 1083
rect 1085 1077 1100 1083
rect 1037 1057 1075 1063
rect 1085 1057 1091 1077
rect 2573 1077 2595 1083
rect 3053 1077 3075 1083
rect 3149 1077 3164 1083
rect 3053 1064 3059 1077
rect 3316 1077 3331 1083
rect 3645 1077 3660 1083
rect 3828 1077 3843 1083
rect 3988 1077 4019 1083
rect 4077 1077 4092 1083
rect 4909 1077 4924 1083
rect 5181 1077 5203 1083
rect 5300 1077 5315 1083
rect 5405 1077 5420 1083
rect 5437 1077 5468 1083
rect 5501 1077 5507 1097
rect 5620 1097 5635 1103
rect 6468 1097 6499 1103
rect 6756 1097 6835 1103
rect 7021 1097 7043 1103
rect 7261 1097 7292 1103
rect 7309 1097 7331 1103
rect 7501 1097 7548 1103
rect 5661 1077 5683 1083
rect 5821 1077 5836 1083
rect 5917 1077 5932 1083
rect 5997 1077 6012 1083
rect 6301 1077 6323 1083
rect 6525 1077 6547 1083
rect 6557 1077 6595 1083
rect 6541 1064 6547 1077
rect 6628 1077 6659 1083
rect 7357 1077 7372 1083
rect 1533 1057 1571 1063
rect 2957 1057 2979 1063
rect 3204 1057 3219 1063
rect 4093 1057 4115 1063
rect 4365 1057 4387 1063
rect 5917 1057 5939 1063
rect 6852 1057 6867 1063
rect 7357 1057 7363 1077
rect 628 1036 630 1044
rect 3530 1036 3532 1044
rect 3684 1036 3686 1044
rect 5716 1036 5720 1044
rect 5802 1036 5804 1044
rect 5860 1036 5862 1044
rect 7412 1036 7416 1044
rect 2266 1014 2278 1016
rect 5274 1014 5286 1016
rect 2251 1006 2253 1014
rect 2261 1006 2263 1014
rect 2271 1006 2273 1014
rect 2281 1006 2283 1014
rect 2291 1006 2293 1014
rect 5259 1006 5261 1014
rect 5269 1006 5271 1014
rect 5279 1006 5281 1014
rect 5289 1006 5291 1014
rect 5299 1006 5301 1014
rect 2266 1004 2278 1006
rect 5274 1004 5286 1006
rect 452 976 454 984
rect 2056 976 2060 984
rect 2442 976 2444 984
rect 5604 976 5606 984
rect 5738 976 5740 984
rect 5924 976 5926 984
rect 6196 976 6200 984
rect 6504 976 6508 984
rect 685 957 700 963
rect 260 937 291 943
rect 573 937 588 943
rect 621 937 636 943
rect 1165 937 1180 943
rect 1380 937 1395 943
rect 1469 937 1484 943
rect 2205 937 2220 943
rect 2557 943 2563 963
rect 4356 956 4364 964
rect 4772 956 4780 964
rect 5252 957 5284 963
rect 5276 948 5284 957
rect 5508 957 5540 963
rect 5532 948 5540 957
rect 7117 957 7155 963
rect 2468 937 2483 943
rect 2557 937 2572 943
rect 2797 937 2812 943
rect 3053 937 3084 943
rect 3581 937 3603 943
rect 3748 937 3827 943
rect 3924 937 3939 943
rect 4029 937 4051 943
rect 4324 937 4339 943
rect 4660 937 4675 943
rect 4724 937 4755 943
rect 5661 937 5699 943
rect 5997 937 6012 943
rect 6637 937 6668 943
rect 173 917 211 923
rect 333 917 371 923
rect 525 917 563 923
rect 605 917 643 923
rect 685 917 748 923
rect 1188 917 1203 923
rect 1332 917 1347 923
rect 1469 917 1507 923
rect 580 897 595 903
rect 1469 897 1475 917
rect 2084 917 2099 923
rect 2109 917 2124 923
rect 2237 917 2316 923
rect 2653 917 2675 923
rect 2957 917 2995 923
rect 3028 917 3043 923
rect 3133 917 3148 923
rect 3213 917 3228 923
rect 3245 917 3260 923
rect 3405 917 3443 923
rect 3453 917 3484 923
rect 3725 917 3820 923
rect 3869 917 3907 923
rect 2925 897 2940 903
rect 3469 897 3507 903
rect 3741 897 3772 903
rect 3869 897 3875 917
rect 4148 917 4179 923
rect 4237 917 4275 923
rect 5981 917 6028 923
rect 6061 917 6099 923
rect 6061 904 6067 917
rect 6116 917 6131 923
rect 6749 923 6755 943
rect 7101 943 7107 956
rect 7085 937 7107 943
rect 7140 937 7171 943
rect 7245 937 7267 943
rect 7261 924 7267 937
rect 7501 943 7507 963
rect 7469 937 7507 943
rect 6749 917 6851 923
rect 7437 917 7459 923
rect 4093 897 4131 903
rect 6701 897 6723 903
rect 2172 884 2180 888
rect 2220 884 2228 888
rect 2428 884 2436 888
rect 3341 877 3356 883
rect 5309 837 5324 843
rect 762 814 774 816
rect 3770 814 3782 816
rect 6778 814 6790 816
rect 747 806 749 814
rect 757 806 759 814
rect 767 806 769 814
rect 777 806 779 814
rect 787 806 789 814
rect 3755 806 3757 814
rect 3765 806 3767 814
rect 3775 806 3777 814
rect 3785 806 3787 814
rect 3795 806 3797 814
rect 6763 806 6765 814
rect 6773 806 6775 814
rect 6783 806 6785 814
rect 6793 806 6795 814
rect 6803 806 6805 814
rect 762 804 774 806
rect 3770 804 3782 806
rect 6778 804 6790 806
rect 5588 776 5592 784
rect 5700 776 5708 784
rect 5940 776 5942 784
rect 7140 776 7142 784
rect 7188 776 7190 784
rect 7496 776 7500 784
rect 2212 737 2227 743
rect 3956 737 3971 743
rect 4566 736 4572 744
rect 4676 737 4691 743
rect 4868 736 4870 744
rect 4948 737 4979 743
rect 4996 737 5052 743
rect 2173 717 2195 723
rect 2276 717 2323 723
rect 3981 717 3996 723
rect 4749 717 4787 723
rect 6301 717 6323 723
rect 6333 717 6348 723
rect 420 697 451 703
rect 637 697 652 703
rect 669 697 707 703
rect 1565 697 1603 703
rect 1709 697 1724 703
rect 2541 697 2572 703
rect 3028 697 3043 703
rect 3133 697 3155 703
rect 4836 697 4851 703
rect 1524 677 1539 683
rect 1549 677 1580 683
rect 2925 677 2940 683
rect 3661 677 3676 683
rect 3940 677 3955 683
rect 4845 677 4851 697
rect 5821 683 5827 703
rect 6084 697 6115 703
rect 6301 697 6316 703
rect 6381 697 6412 703
rect 6669 697 6691 703
rect 6973 697 7011 703
rect 7156 697 7187 703
rect 7373 697 7388 703
rect 5789 677 5827 683
rect 5885 677 5923 683
rect 6036 677 6051 683
rect 6605 677 6620 683
rect 6740 677 6851 683
rect 7037 677 7052 683
rect 7261 677 7276 683
rect 7357 677 7411 683
rect 7428 677 7443 683
rect 749 657 764 663
rect 4604 663 4612 666
rect 4604 657 4627 663
rect 5812 657 5843 663
rect 6909 657 6924 663
rect 7261 657 7283 663
rect 7293 657 7331 663
rect 842 636 844 644
rect 3642 636 3644 644
rect 3690 636 3692 644
rect 3741 637 3804 643
rect 4010 636 4012 644
rect 4740 636 4742 644
rect 5380 636 5382 644
rect 5418 636 5420 644
rect 5466 636 5468 644
rect 5514 636 5516 644
rect 5720 636 5724 644
rect 2266 614 2278 616
rect 5274 614 5286 616
rect 2251 606 2253 614
rect 2261 606 2263 614
rect 2271 606 2273 614
rect 2281 606 2283 614
rect 2291 606 2293 614
rect 5259 606 5261 614
rect 5269 606 5271 614
rect 5279 606 5281 614
rect 5289 606 5291 614
rect 5299 606 5301 614
rect 2266 604 2278 606
rect 5274 604 5286 606
rect 1588 576 1590 584
rect 3898 576 3900 584
rect 5172 577 5187 583
rect 5796 576 5800 584
rect 5908 576 5912 584
rect 6580 576 6582 584
rect 6840 576 6844 584
rect 6964 576 6966 584
rect 1636 556 1644 564
rect 2212 557 2227 563
rect 2988 557 3011 563
rect 2988 554 2996 557
rect 3165 557 3180 563
rect 4388 556 4396 564
rect 4724 556 4732 564
rect 5460 557 5475 563
rect 7405 557 7427 563
rect 1757 537 1772 543
rect 2237 537 2300 543
rect 3124 537 3171 543
rect 269 517 284 523
rect 1453 517 1491 523
rect 1709 517 1747 523
rect 1949 517 1996 523
rect 2349 517 2364 523
rect 2445 517 2476 523
rect 3101 517 3148 523
rect 3172 517 3187 523
rect 3389 523 3395 543
rect 3485 537 3500 543
rect 3565 537 3619 543
rect 4356 537 4371 543
rect 4420 537 4451 543
rect 4692 537 4707 543
rect 4756 537 4787 543
rect 5037 537 5059 543
rect 5965 537 5980 543
rect 6093 537 6108 543
rect 6333 537 6355 543
rect 6445 537 6499 543
rect 6548 537 6563 543
rect 6676 537 6691 543
rect 7172 537 7203 543
rect 3372 517 3395 523
rect 3421 517 3459 523
rect 3372 512 3380 517
rect 717 497 732 503
rect 2749 497 2787 503
rect 3021 497 3036 503
rect 3421 497 3427 517
rect 3492 517 3523 523
rect 3773 517 3820 523
rect 3917 517 3932 523
rect 3949 517 3987 523
rect 5229 517 5331 523
rect 5485 517 5500 523
rect 6013 517 6035 523
rect 6397 517 6412 523
rect 6541 517 6556 523
rect 7005 517 7027 523
rect 7117 517 7139 523
rect 7236 517 7251 523
rect 7453 517 7475 523
rect 3556 497 3571 503
rect 6589 497 6611 503
rect 6637 497 6675 503
rect 6973 497 7011 503
rect 7300 497 7315 503
rect 5140 477 5187 483
rect 5437 477 5468 483
rect 7277 477 7292 483
rect 6442 436 6444 444
rect 7517 437 7532 443
rect 762 414 774 416
rect 3770 414 3782 416
rect 6778 414 6790 416
rect 747 406 749 414
rect 757 406 759 414
rect 767 406 769 414
rect 777 406 779 414
rect 787 406 789 414
rect 3755 406 3757 414
rect 3765 406 3767 414
rect 3775 406 3777 414
rect 3785 406 3787 414
rect 3795 406 3797 414
rect 6763 406 6765 414
rect 6773 406 6775 414
rect 6783 406 6785 414
rect 6793 406 6795 414
rect 6803 406 6805 414
rect 762 404 774 406
rect 3770 404 3782 406
rect 6778 404 6790 406
rect 2164 376 2166 384
rect 2484 376 2486 384
rect 4276 376 4278 384
rect 6340 376 6344 384
rect 7460 376 7462 384
rect 1286 336 1292 344
rect 4634 336 4636 344
rect 4685 337 4700 343
rect 4717 337 4771 343
rect 7172 337 7187 343
rect 989 317 1004 323
rect 605 297 643 303
rect 749 297 764 303
rect 941 297 979 303
rect 1012 297 1027 303
rect 1597 297 1635 303
rect 2125 297 2156 303
rect 308 276 310 284
rect 380 277 403 283
rect 380 272 388 277
rect 884 277 915 283
rect 2125 277 2131 297
rect 2189 303 2195 323
rect 2308 317 2323 323
rect 2381 317 2419 323
rect 2749 317 2787 323
rect 3101 317 3116 323
rect 2189 297 2227 303
rect 2349 297 2364 303
rect 2429 297 2483 303
rect 2788 297 2803 303
rect 3309 303 3315 323
rect 4301 317 4323 323
rect 4424 314 4428 322
rect 4813 317 4835 323
rect 5348 317 5363 323
rect 6472 316 6476 324
rect 6701 317 6716 323
rect 3309 297 3347 303
rect 3364 297 3379 303
rect 3517 297 3548 303
rect 3565 297 3603 303
rect 4100 297 4115 303
rect 4708 297 4723 303
rect 4836 297 4851 303
rect 4861 297 4892 303
rect 4900 297 4947 303
rect 6733 297 6819 303
rect 6884 297 6899 303
rect 7112 297 7171 303
rect 2941 277 2956 283
rect 3076 276 3080 284
rect 3245 277 3260 283
rect 4029 277 4051 283
rect 4237 277 4252 283
rect 4653 277 4691 283
rect 4877 277 4908 283
rect 5092 277 5107 283
rect 5252 277 5272 283
rect 5300 277 5363 283
rect 5556 277 5587 283
rect 5869 277 5884 283
rect 5924 277 5955 283
rect 5972 277 6003 283
rect 6292 277 6307 283
rect 6884 277 6915 283
rect 7165 277 7171 297
rect 7245 277 7267 283
rect 7277 277 7331 283
rect 7357 277 7411 283
rect 1804 266 1812 276
rect 820 257 835 263
rect 2932 256 2940 264
rect 1114 236 1116 244
rect 3748 237 3811 243
rect 6106 236 6108 244
rect 2266 214 2278 216
rect 5274 214 5286 216
rect 2251 206 2253 214
rect 2261 206 2263 214
rect 2271 206 2273 214
rect 2281 206 2283 214
rect 2291 206 2293 214
rect 5259 206 5261 214
rect 5269 206 5271 214
rect 5279 206 5281 214
rect 5289 206 5291 214
rect 5299 206 5301 214
rect 2266 204 2278 206
rect 5274 204 5286 206
rect 3844 177 3859 183
rect 1476 157 1491 163
rect 2436 157 2451 163
rect 3853 163 3859 177
rect 6536 176 6540 184
rect 7396 176 7400 184
rect 3853 157 3923 163
rect 244 137 259 143
rect 2292 137 2355 143
rect 4308 137 4323 143
rect 4372 137 4403 143
rect 4653 143 4659 163
rect 4788 157 4803 163
rect 4980 156 4988 164
rect 6765 157 6780 163
rect 4589 137 4659 143
rect 4740 137 4771 143
rect 4948 137 4963 143
rect 5036 143 5044 144
rect 5036 137 5052 143
rect 6708 137 6739 143
rect 7284 137 7299 143
rect 7341 143 7347 163
rect 7341 137 7356 143
rect 84 117 99 123
rect 173 117 211 123
rect 541 117 572 123
rect 701 117 764 123
rect 845 117 876 123
rect 1581 117 1619 123
rect 2308 117 2371 123
rect 2765 117 2819 123
rect 2973 117 3004 123
rect 3149 117 3187 123
rect 3197 117 3235 123
rect 3725 117 3740 123
rect 3933 117 3971 123
rect 4573 117 4588 123
rect 4884 117 4899 123
rect 5869 117 5907 123
rect 6093 117 6131 123
rect 6253 117 6291 123
rect 6788 117 6860 123
rect 6877 117 6915 123
rect 6989 117 7004 123
rect 7085 117 7100 123
rect 2125 97 2140 103
rect 2269 97 2332 103
rect 2397 97 2419 103
rect 2589 97 2611 103
rect 6653 97 6668 103
rect 6989 97 7011 103
rect 7021 97 7059 103
rect 7316 97 7331 103
rect 4570 76 4572 84
rect 762 14 774 16
rect 3770 14 3782 16
rect 6778 14 6790 16
rect 747 6 749 14
rect 757 6 759 14
rect 767 6 769 14
rect 777 6 779 14
rect 787 6 789 14
rect 3755 6 3757 14
rect 3765 6 3767 14
rect 3775 6 3777 14
rect 3785 6 3787 14
rect 3795 6 3797 14
rect 6763 6 6765 14
rect 6773 6 6775 14
rect 6783 6 6785 14
rect 6793 6 6795 14
rect 6803 6 6805 14
rect 762 4 774 6
rect 3770 4 3782 6
rect 6778 4 6790 6
<< m2contact >>
rect 739 5206 747 5214
rect 749 5206 757 5214
rect 759 5206 767 5214
rect 769 5206 777 5214
rect 779 5206 787 5214
rect 789 5206 797 5214
rect 3747 5206 3755 5214
rect 3757 5206 3765 5214
rect 3767 5206 3775 5214
rect 3777 5206 3785 5214
rect 3787 5206 3795 5214
rect 3797 5206 3805 5214
rect 6755 5206 6763 5214
rect 6765 5206 6773 5214
rect 6775 5206 6783 5214
rect 6785 5206 6793 5214
rect 6795 5206 6803 5214
rect 6805 5206 6813 5214
rect 4220 5176 4228 5184
rect 4460 5176 4468 5184
rect 4508 5176 4516 5184
rect 4684 5176 4692 5184
rect 5324 5176 5332 5184
rect 7468 5176 7476 5184
rect 4204 5156 4212 5164
rect 5532 5156 5540 5164
rect 6156 5156 6164 5164
rect 4444 5136 4452 5144
rect 4924 5136 4932 5144
rect 5548 5136 5556 5144
rect 988 5116 996 5124
rect 1020 5116 1028 5124
rect 4732 5116 4740 5124
rect 4828 5116 4836 5124
rect 4956 5116 4964 5124
rect 4972 5116 4980 5124
rect 5036 5116 5044 5124
rect 5068 5116 5076 5124
rect 5148 5116 5156 5124
rect 5180 5116 5188 5124
rect 5372 5116 5380 5124
rect 5436 5116 5444 5124
rect 5612 5116 5620 5124
rect 6012 5116 6020 5124
rect 6028 5116 6036 5124
rect 6188 5116 6196 5124
rect 6220 5116 6228 5124
rect 6300 5116 6308 5124
rect 6332 5116 6340 5124
rect 7052 5116 7060 5124
rect 7180 5116 7188 5124
rect 76 5096 84 5104
rect 124 5096 132 5104
rect 204 5096 212 5104
rect 268 5096 276 5104
rect 316 5096 324 5104
rect 380 5096 388 5104
rect 412 5096 420 5104
rect 476 5094 484 5102
rect 684 5096 692 5104
rect 748 5094 756 5102
rect 844 5096 852 5104
rect 972 5096 980 5104
rect 1020 5096 1028 5104
rect 1100 5094 1108 5102
rect 1292 5094 1300 5102
rect 1468 5096 1476 5104
rect 1532 5096 1540 5104
rect 1660 5096 1668 5104
rect 1740 5096 1748 5104
rect 1788 5096 1796 5104
rect 1836 5096 1844 5104
rect 1964 5096 1972 5104
rect 2044 5096 2052 5104
rect 2108 5096 2116 5104
rect 2140 5096 2148 5104
rect 2236 5096 2244 5104
rect 2412 5096 2420 5104
rect 2508 5096 2516 5104
rect 2572 5094 2580 5102
rect 2732 5096 2740 5104
rect 2764 5096 2772 5104
rect 2860 5096 2868 5104
rect 2892 5096 2900 5104
rect 3036 5096 3044 5104
rect 3084 5096 3092 5104
rect 3212 5094 3220 5102
rect 3276 5096 3284 5104
rect 3356 5096 3364 5104
rect 3420 5096 3428 5104
rect 3452 5096 3460 5104
rect 3532 5096 3540 5104
rect 3580 5096 3588 5104
rect 3660 5096 3668 5104
rect 3708 5096 3716 5104
rect 3724 5096 3732 5104
rect 3948 5096 3956 5104
rect 4076 5094 4084 5102
rect 4140 5096 4148 5104
rect 4252 5096 4260 5104
rect 4316 5094 4324 5102
rect 4492 5096 4500 5104
rect 4540 5096 4548 5104
rect 4588 5096 4596 5104
rect 4636 5096 4644 5104
rect 4652 5096 4660 5104
rect 4780 5096 4788 5104
rect 4876 5096 4884 5104
rect 5004 5096 5012 5104
rect 5228 5096 5236 5104
rect 5404 5096 5412 5104
rect 5516 5096 5524 5104
rect 5532 5096 5540 5104
rect 5804 5096 5812 5104
rect 5900 5096 5908 5104
rect 5916 5096 5924 5104
rect 5980 5096 5988 5104
rect 6076 5096 6084 5104
rect 6092 5096 6100 5104
rect 6412 5096 6420 5104
rect 6604 5096 6612 5104
rect 6700 5096 6708 5104
rect 6828 5096 6836 5104
rect 6876 5096 6884 5104
rect 6940 5096 6948 5104
rect 7132 5096 7140 5104
rect 7164 5096 7172 5104
rect 7196 5096 7204 5104
rect 7308 5096 7316 5104
rect 7356 5096 7364 5104
rect 7452 5096 7460 5104
rect 7500 5096 7508 5104
rect 7564 5096 7572 5104
rect 220 5076 228 5084
rect 300 5056 308 5064
rect 348 5056 356 5064
rect 396 5076 404 5084
rect 444 5076 452 5084
rect 524 5076 532 5084
rect 892 5076 900 5084
rect 1036 5076 1044 5084
rect 1068 5076 1076 5084
rect 1500 5076 1508 5084
rect 1516 5076 1524 5084
rect 1708 5076 1716 5084
rect 1772 5076 1780 5084
rect 1804 5076 1812 5084
rect 2012 5076 2020 5084
rect 2060 5076 2068 5084
rect 940 5056 948 5064
rect 1292 5056 1300 5064
rect 1436 5056 1444 5064
rect 1772 5056 1780 5064
rect 1836 5056 1844 5064
rect 2252 5076 2260 5084
rect 2348 5076 2356 5084
rect 2108 5056 2116 5064
rect 2444 5056 2452 5064
rect 2476 5076 2484 5084
rect 2492 5076 2500 5084
rect 2540 5076 2548 5084
rect 2764 5076 2772 5084
rect 3068 5076 3076 5084
rect 2716 5056 2724 5064
rect 3388 5056 3396 5064
rect 3436 5076 3444 5084
rect 3676 5076 3684 5084
rect 3900 5076 3908 5084
rect 4348 5076 4356 5084
rect 4556 5076 4564 5084
rect 4604 5076 4612 5084
rect 4748 5076 4756 5084
rect 4764 5076 4772 5084
rect 4812 5076 4820 5084
rect 4876 5076 4884 5084
rect 3756 5056 3764 5064
rect 188 5036 196 5044
rect 236 5036 244 5044
rect 604 5036 612 5044
rect 620 5036 628 5044
rect 908 5036 916 5044
rect 1228 5036 1236 5044
rect 1420 5036 1428 5044
rect 1548 5036 1556 5044
rect 1852 5036 1860 5044
rect 2156 5036 2164 5044
rect 2700 5036 2708 5044
rect 2780 5036 2788 5044
rect 2972 5036 2980 5044
rect 3340 5036 3348 5044
rect 3468 5036 3476 5044
rect 4700 5056 4708 5064
rect 4812 5056 4820 5064
rect 4924 5076 4932 5084
rect 5068 5076 5076 5084
rect 5116 5076 5124 5084
rect 5180 5076 5188 5084
rect 5340 5076 5348 5084
rect 5356 5076 5364 5084
rect 5388 5076 5396 5084
rect 5468 5076 5476 5084
rect 5580 5076 5588 5084
rect 5724 5076 5732 5084
rect 5772 5076 5780 5084
rect 5132 5056 5140 5064
rect 5148 5056 5156 5064
rect 5212 5056 5220 5064
rect 5452 5056 5460 5064
rect 5740 5056 5748 5064
rect 5852 5056 5860 5064
rect 5916 5056 5924 5064
rect 5964 5076 5972 5084
rect 6076 5076 6084 5084
rect 6124 5076 6132 5084
rect 6220 5076 6228 5084
rect 6268 5076 6276 5084
rect 6332 5076 6340 5084
rect 6460 5080 6468 5088
rect 6476 5076 6484 5084
rect 6492 5076 6500 5084
rect 6588 5076 6596 5084
rect 6620 5076 6628 5084
rect 6956 5076 6964 5084
rect 6140 5056 6148 5064
rect 6172 5056 6180 5064
rect 6284 5056 6292 5064
rect 6300 5056 6308 5064
rect 6364 5056 6372 5064
rect 6380 5056 6388 5064
rect 6652 5056 6660 5064
rect 6668 5056 6676 5064
rect 6716 5056 6724 5064
rect 6860 5056 6868 5064
rect 6924 5056 6932 5064
rect 7036 5076 7044 5084
rect 7084 5076 7092 5084
rect 7164 5076 7172 5084
rect 7228 5076 7236 5084
rect 7004 5056 7012 5064
rect 7100 5056 7108 5064
rect 7132 5056 7140 5064
rect 7196 5056 7204 5064
rect 7324 5076 7332 5084
rect 7436 5076 7444 5084
rect 7276 5056 7284 5064
rect 7340 5056 7348 5064
rect 7388 5056 7396 5064
rect 7404 5056 7412 5064
rect 7516 5056 7524 5064
rect 4204 5036 4212 5044
rect 4828 5036 4836 5044
rect 4956 5036 4964 5044
rect 4972 5036 4980 5044
rect 5036 5036 5044 5044
rect 5436 5036 5444 5044
rect 5596 5036 5604 5044
rect 5692 5036 5700 5044
rect 5868 5036 5876 5044
rect 6012 5036 6020 5044
rect 6028 5036 6036 5044
rect 6188 5036 6196 5044
rect 6396 5036 6404 5044
rect 6428 5036 6436 5044
rect 6540 5036 6548 5044
rect 6636 5036 6644 5044
rect 6972 5036 6980 5044
rect 7244 5036 7252 5044
rect 7420 5036 7428 5044
rect 7532 5036 7540 5044
rect 2243 5006 2251 5014
rect 2253 5006 2261 5014
rect 2263 5006 2271 5014
rect 2273 5006 2281 5014
rect 2283 5006 2291 5014
rect 2293 5006 2301 5014
rect 5251 5006 5259 5014
rect 5261 5006 5269 5014
rect 5271 5006 5279 5014
rect 5281 5006 5289 5014
rect 5291 5006 5299 5014
rect 5301 5006 5309 5014
rect 188 4976 196 4984
rect 988 4976 996 4984
rect 1052 4976 1060 4984
rect 1404 4976 1412 4984
rect 2172 4976 2180 4984
rect 2476 4976 2484 4984
rect 2636 4976 2644 4984
rect 2892 4976 2900 4984
rect 3052 4976 3060 4984
rect 3628 4976 3636 4984
rect 4092 4976 4100 4984
rect 4556 4976 4564 4984
rect 5372 4976 5380 4984
rect 6124 4976 6132 4984
rect 6156 4976 6164 4984
rect 6620 4976 6628 4984
rect 6668 4976 6676 4984
rect 6844 4976 6852 4984
rect 6940 4976 6948 4984
rect 7244 4976 7252 4984
rect 7340 4976 7348 4984
rect 236 4956 244 4964
rect 220 4936 228 4944
rect 268 4956 276 4964
rect 1660 4956 1668 4964
rect 1724 4956 1732 4964
rect 1756 4956 1764 4964
rect 2460 4956 2468 4964
rect 2700 4956 2708 4964
rect 3004 4956 3012 4964
rect 3116 4956 3124 4964
rect 3516 4956 3524 4964
rect 3964 4956 3972 4964
rect 4828 4956 4836 4964
rect 5020 4956 5028 4964
rect 5036 4956 5044 4964
rect 5164 4956 5172 4964
rect 5564 4956 5572 4964
rect 5596 4956 5604 4964
rect 5612 4956 5620 4964
rect 6092 4956 6100 4964
rect 6108 4956 6116 4964
rect 6236 4956 6244 4964
rect 524 4936 532 4944
rect 76 4916 84 4924
rect 124 4916 132 4924
rect 204 4916 212 4924
rect 300 4916 308 4924
rect 316 4916 324 4924
rect 380 4916 388 4924
rect 412 4916 420 4924
rect 428 4916 436 4924
rect 476 4916 484 4924
rect 492 4916 500 4924
rect 572 4916 580 4924
rect 700 4916 708 4924
rect 716 4916 724 4924
rect 764 4916 772 4924
rect 860 4916 868 4924
rect 876 4916 884 4924
rect 924 4916 932 4924
rect 1004 4936 1012 4944
rect 1100 4936 1108 4944
rect 1164 4936 1172 4944
rect 1180 4936 1188 4944
rect 1212 4936 1220 4944
rect 1244 4936 1252 4944
rect 1292 4936 1300 4944
rect 1628 4936 1636 4944
rect 1724 4936 1732 4944
rect 2284 4936 2292 4944
rect 2620 4936 2628 4944
rect 2908 4936 2916 4944
rect 2940 4936 2948 4944
rect 3036 4936 3044 4944
rect 3596 4936 3604 4944
rect 3788 4936 3796 4944
rect 3948 4936 3956 4944
rect 4044 4936 4052 4944
rect 4076 4936 4084 4944
rect 4172 4936 4180 4944
rect 4396 4936 4404 4944
rect 4588 4936 4596 4944
rect 4860 4936 4868 4944
rect 4892 4936 4900 4944
rect 4988 4936 4996 4944
rect 5148 4936 5156 4944
rect 5196 4936 5204 4944
rect 5228 4936 5236 4944
rect 5324 4936 5332 4944
rect 5484 4936 5492 4944
rect 5500 4936 5508 4944
rect 5644 4936 5652 4944
rect 5724 4936 5732 4944
rect 5740 4936 5748 4944
rect 5836 4936 5844 4944
rect 5852 4936 5860 4944
rect 5948 4936 5956 4944
rect 6060 4936 6068 4944
rect 6076 4936 6084 4944
rect 1020 4916 1028 4924
rect 1132 4916 1140 4924
rect 1148 4916 1156 4924
rect 1068 4896 1076 4904
rect 1116 4896 1124 4904
rect 1292 4916 1300 4924
rect 1340 4916 1348 4924
rect 1484 4916 1492 4924
rect 1500 4916 1508 4924
rect 1532 4916 1540 4924
rect 1580 4916 1588 4924
rect 1596 4916 1604 4924
rect 1612 4916 1620 4924
rect 1660 4916 1668 4924
rect 1676 4916 1684 4924
rect 1820 4918 1828 4926
rect 1884 4916 1892 4924
rect 1964 4916 1972 4924
rect 1980 4916 1988 4924
rect 2044 4916 2052 4924
rect 2060 4916 2068 4924
rect 2076 4916 2084 4924
rect 2124 4916 2132 4924
rect 2364 4916 2372 4924
rect 2380 4916 2388 4924
rect 2444 4916 2452 4924
rect 2492 4916 2500 4924
rect 2524 4916 2532 4924
rect 2572 4916 2580 4924
rect 2588 4916 2596 4924
rect 2604 4916 2612 4924
rect 2668 4916 2676 4924
rect 2780 4916 2788 4924
rect 2828 4916 2836 4924
rect 2908 4916 2916 4924
rect 2972 4916 2980 4924
rect 3020 4916 3028 4924
rect 3084 4916 3092 4924
rect 3132 4916 3140 4924
rect 3148 4916 3156 4924
rect 3196 4916 3204 4924
rect 3228 4916 3236 4924
rect 3244 4916 3252 4924
rect 3292 4916 3300 4924
rect 3340 4916 3348 4924
rect 3388 4916 3396 4924
rect 3404 4916 3412 4924
rect 3420 4916 3428 4924
rect 3484 4916 3492 4924
rect 3500 4916 3508 4924
rect 3548 4916 3556 4924
rect 3580 4916 3588 4924
rect 3612 4916 3620 4924
rect 3740 4916 3748 4924
rect 3852 4916 3860 4924
rect 3932 4916 3940 4924
rect 4028 4916 4036 4924
rect 4060 4916 4068 4924
rect 4172 4916 4180 4924
rect 4236 4918 4244 4926
rect 4300 4916 4308 4924
rect 4428 4918 4436 4926
rect 4620 4918 4628 4926
rect 4796 4916 4804 4924
rect 4876 4916 4884 4924
rect 6188 4932 6196 4940
rect 6364 4936 6372 4944
rect 6428 4936 6436 4944
rect 7004 4956 7012 4964
rect 7116 4956 7124 4964
rect 7196 4956 7204 4964
rect 7484 4956 7492 4964
rect 6492 4936 6500 4944
rect 6636 4936 6644 4944
rect 6684 4936 6692 4944
rect 6892 4936 6900 4944
rect 7004 4936 7012 4944
rect 7020 4936 7028 4944
rect 7100 4936 7108 4944
rect 7148 4936 7156 4944
rect 7292 4936 7300 4944
rect 7308 4936 7316 4944
rect 7404 4936 7412 4944
rect 7500 4936 7508 4944
rect 5340 4916 5348 4924
rect 5516 4916 5524 4924
rect 5564 4916 5572 4924
rect 5596 4916 5604 4924
rect 5628 4916 5636 4924
rect 5660 4916 5668 4924
rect 5708 4916 5716 4924
rect 5772 4916 5780 4924
rect 6140 4916 6148 4924
rect 6204 4916 6212 4924
rect 6284 4916 6292 4924
rect 6316 4916 6324 4924
rect 6348 4916 6356 4924
rect 6364 4916 6372 4924
rect 6412 4916 6420 4924
rect 6460 4916 6468 4924
rect 6556 4916 6564 4924
rect 6652 4916 6660 4924
rect 6732 4916 6740 4924
rect 6908 4916 6916 4924
rect 6956 4916 6964 4924
rect 7068 4916 7076 4924
rect 7116 4916 7124 4924
rect 7148 4916 7156 4924
rect 7212 4916 7220 4924
rect 7452 4916 7460 4924
rect 7516 4916 7524 4924
rect 3996 4896 4004 4904
rect 4124 4896 4132 4904
rect 4764 4896 4772 4904
rect 5548 4896 5556 4904
rect 5740 4896 5748 4904
rect 5804 4896 5812 4904
rect 6604 4896 6612 4904
rect 6860 4896 6868 4904
rect 7068 4896 7076 4904
rect 7260 4896 7268 4904
rect 7548 4896 7556 4904
rect 748 4876 756 4884
rect 1948 4876 1956 4884
rect 2860 4876 2868 4884
rect 3916 4876 3924 4884
rect 6540 4876 6548 4884
rect 5884 4856 5892 4864
rect 364 4836 372 4844
rect 460 4836 468 4844
rect 684 4836 692 4844
rect 908 4836 916 4844
rect 1468 4836 1476 4844
rect 1564 4836 1572 4844
rect 1996 4836 2004 4844
rect 2108 4836 2116 4844
rect 2412 4836 2420 4844
rect 2556 4836 2564 4844
rect 3180 4836 3188 4844
rect 3276 4836 3284 4844
rect 3356 4836 3364 4844
rect 3452 4836 3460 4844
rect 4364 4836 4372 4844
rect 4748 4836 4756 4844
rect 4796 4836 4804 4844
rect 4828 4836 4836 4844
rect 4924 4836 4932 4844
rect 5084 4836 5092 4844
rect 5452 4836 5460 4844
rect 5676 4836 5684 4844
rect 5996 4836 6004 4844
rect 6316 4836 6324 4844
rect 6556 4836 6564 4844
rect 6844 4836 6852 4844
rect 6876 4836 6884 4844
rect 7132 4836 7140 4844
rect 7196 4836 7204 4844
rect 7276 4836 7284 4844
rect 7420 4836 7428 4844
rect 7468 4836 7476 4844
rect 7516 4836 7524 4844
rect 739 4806 747 4814
rect 749 4806 757 4814
rect 759 4806 767 4814
rect 769 4806 777 4814
rect 779 4806 787 4814
rect 789 4806 797 4814
rect 3747 4806 3755 4814
rect 3757 4806 3765 4814
rect 3767 4806 3775 4814
rect 3777 4806 3785 4814
rect 3787 4806 3795 4814
rect 3797 4806 3805 4814
rect 6755 4806 6763 4814
rect 6765 4806 6773 4814
rect 6775 4806 6783 4814
rect 6785 4806 6793 4814
rect 6795 4806 6803 4814
rect 6805 4806 6813 4814
rect 396 4776 404 4784
rect 812 4776 820 4784
rect 1196 4776 1204 4784
rect 1276 4776 1284 4784
rect 2092 4776 2100 4784
rect 2220 4776 2228 4784
rect 2828 4776 2836 4784
rect 3628 4776 3636 4784
rect 5052 4776 5060 4784
rect 5068 4776 5076 4784
rect 5308 4776 5316 4784
rect 6588 4776 6596 4784
rect 7564 4776 7572 4784
rect 492 4756 500 4764
rect 4092 4756 4100 4764
rect 4748 4756 4756 4764
rect 5996 4756 6004 4764
rect 1900 4736 1908 4744
rect 2684 4736 2692 4744
rect 3164 4736 3172 4744
rect 3820 4736 3828 4744
rect 4076 4736 4084 4744
rect 4348 4736 4356 4744
rect 5036 4736 5044 4744
rect 5772 4736 5780 4744
rect 524 4716 532 4724
rect 636 4716 644 4724
rect 76 4696 84 4704
rect 124 4696 132 4704
rect 252 4694 260 4702
rect 428 4696 436 4704
rect 460 4696 468 4704
rect 492 4696 500 4704
rect 572 4696 580 4704
rect 604 4696 612 4704
rect 668 4696 676 4704
rect 700 4696 708 4704
rect 812 4696 820 4704
rect 860 4716 868 4724
rect 1052 4716 1060 4724
rect 908 4696 916 4704
rect 924 4696 932 4704
rect 972 4696 980 4704
rect 1020 4696 1028 4704
rect 1084 4696 1092 4704
rect 1116 4696 1124 4704
rect 1148 4696 1156 4704
rect 1164 4696 1172 4704
rect 1212 4696 1220 4704
rect 1228 4696 1236 4704
rect 1308 4696 1316 4704
rect 1356 4716 1364 4724
rect 1452 4694 1460 4702
rect 1516 4696 1524 4704
rect 1644 4694 1652 4702
rect 1708 4696 1716 4704
rect 1804 4696 1812 4704
rect 1820 4696 1828 4704
rect 1980 4716 1988 4724
rect 1868 4696 1876 4704
rect 1900 4696 1908 4704
rect 1948 4696 1956 4704
rect 1964 4696 1972 4704
rect 2028 4696 2036 4704
rect 2060 4696 2068 4704
rect 2092 4696 2100 4704
rect 2156 4696 2164 4704
rect 2172 4696 2180 4704
rect 2188 4696 2196 4704
rect 2236 4696 2244 4704
rect 2396 4696 2404 4704
rect 2524 4696 2532 4704
rect 2620 4696 2628 4704
rect 3260 4716 3268 4724
rect 3388 4716 3396 4724
rect 3500 4716 3508 4724
rect 3516 4716 3524 4724
rect 3644 4716 3652 4724
rect 3836 4716 3844 4724
rect 4140 4716 4148 4724
rect 5420 4716 5428 4724
rect 5532 4716 5540 4724
rect 5740 4716 5748 4724
rect 2684 4696 2692 4704
rect 2892 4696 2900 4704
rect 2956 4696 2964 4704
rect 3052 4696 3060 4704
rect 3068 4696 3076 4704
rect 3164 4696 3172 4704
rect 3228 4696 3236 4704
rect 3292 4696 3300 4704
rect 3324 4696 3332 4704
rect 3372 4696 3380 4704
rect 3420 4696 3428 4704
rect 3436 4696 3444 4704
rect 3452 4696 3460 4704
rect 3548 4696 3556 4704
rect 3580 4696 3588 4704
rect 3676 4696 3684 4704
rect 3708 4696 3716 4704
rect 3868 4696 3876 4704
rect 3948 4694 3956 4702
rect 4124 4696 4132 4704
rect 4172 4696 4180 4704
rect 4252 4694 4260 4702
rect 4444 4694 4452 4702
rect 4588 4696 4596 4704
rect 4780 4696 4788 4704
rect 4812 4696 4820 4704
rect 4860 4696 4868 4704
rect 4972 4696 4980 4704
rect 5164 4696 5172 4704
rect 5196 4696 5204 4704
rect 5340 4696 5348 4704
rect 5532 4696 5540 4704
rect 5660 4696 5668 4704
rect 5756 4696 5764 4704
rect 5836 4696 5844 4704
rect 6028 4696 6036 4704
rect 6076 4696 6084 4704
rect 6396 4716 6404 4724
rect 6924 4716 6932 4724
rect 7052 4716 7060 4724
rect 7116 4716 7124 4724
rect 7132 4716 7140 4724
rect 7244 4716 7252 4724
rect 7356 4716 7364 4724
rect 6460 4696 6468 4704
rect 6492 4696 6500 4704
rect 6508 4696 6516 4704
rect 6556 4696 6564 4704
rect 6652 4696 6660 4704
rect 6668 4696 6676 4704
rect 6716 4696 6724 4704
rect 6956 4696 6964 4704
rect 7148 4696 7156 4704
rect 7212 4696 7220 4704
rect 7276 4696 7284 4704
rect 7404 4696 7412 4704
rect 7420 4696 7428 4704
rect 7516 4696 7524 4704
rect 268 4676 276 4684
rect 444 4676 452 4684
rect 572 4676 580 4684
rect 716 4676 724 4684
rect 732 4676 740 4684
rect 892 4676 900 4684
rect 1004 4676 1012 4684
rect 1132 4676 1140 4684
rect 1292 4676 1300 4684
rect 1356 4676 1364 4684
rect 1388 4676 1396 4684
rect 1788 4676 1796 4684
rect 1852 4676 1860 4684
rect 1916 4676 1924 4684
rect 1932 4676 1940 4684
rect 2044 4676 2052 4684
rect 2108 4676 2116 4684
rect 2348 4676 2356 4684
rect 2444 4676 2452 4684
rect 2572 4676 2580 4684
rect 2636 4676 2644 4684
rect 2700 4676 2708 4684
rect 2716 4676 2724 4684
rect 2940 4676 2948 4684
rect 2988 4676 2996 4684
rect 3212 4676 3220 4684
rect 3340 4676 3348 4684
rect 3468 4676 3476 4684
rect 3564 4676 3572 4684
rect 3596 4676 3604 4684
rect 3692 4676 3700 4684
rect 3724 4676 3732 4684
rect 3884 4676 3892 4684
rect 3980 4676 3988 4684
rect 4188 4676 4196 4684
rect 4220 4676 4228 4684
rect 4636 4676 4644 4684
rect 4732 4676 4740 4684
rect 4796 4676 4804 4684
rect 4908 4676 4916 4684
rect 4972 4676 4980 4684
rect 5100 4676 5108 4684
rect 5212 4676 5220 4684
rect 5388 4676 5396 4684
rect 5468 4676 5476 4684
rect 5548 4676 5556 4684
rect 1996 4656 2004 4664
rect 2124 4656 2132 4664
rect 2556 4656 2564 4664
rect 2860 4656 2868 4664
rect 3196 4656 3204 4664
rect 3324 4656 3332 4664
rect 4444 4656 4452 4664
rect 4908 4656 4916 4664
rect 5036 4656 5044 4664
rect 5116 4656 5124 4664
rect 5228 4656 5236 4664
rect 5244 4656 5252 4664
rect 5436 4656 5444 4664
rect 5484 4656 5492 4664
rect 5580 4656 5588 4664
rect 5628 4676 5636 4684
rect 5692 4676 5700 4684
rect 5804 4676 5812 4684
rect 5900 4676 5908 4684
rect 5660 4656 5668 4664
rect 5724 4656 5732 4664
rect 5980 4676 5988 4684
rect 6060 4676 6068 4684
rect 6108 4676 6116 4684
rect 6124 4676 6132 4684
rect 6220 4676 6228 4684
rect 6236 4676 6244 4684
rect 6284 4676 6292 4684
rect 6380 4676 6388 4684
rect 6444 4676 6452 4684
rect 6540 4676 6548 4684
rect 6620 4676 6628 4684
rect 6732 4676 6740 4684
rect 6764 4676 6772 4684
rect 6892 4676 6900 4684
rect 6956 4676 6964 4684
rect 6012 4656 6020 4664
rect 6460 4656 6468 4664
rect 6604 4656 6612 4664
rect 6700 4656 6708 4664
rect 6908 4656 6916 4664
rect 7020 4676 7028 4684
rect 7068 4676 7076 4684
rect 7196 4676 7204 4684
rect 7260 4676 7268 4684
rect 7324 4676 7332 4684
rect 7372 4676 7380 4684
rect 7436 4676 7444 4684
rect 7532 4676 7540 4684
rect 7116 4656 7124 4664
rect 7180 4656 7188 4664
rect 7404 4656 7412 4664
rect 7468 4656 7476 4664
rect 7484 4656 7492 4664
rect 7516 4656 7524 4664
rect 188 4636 196 4644
rect 380 4636 388 4644
rect 396 4636 404 4644
rect 700 4636 708 4644
rect 956 4636 964 4644
rect 1116 4636 1124 4644
rect 1580 4636 1588 4644
rect 1772 4636 1780 4644
rect 2012 4636 2020 4644
rect 2140 4636 2148 4644
rect 2508 4636 2516 4644
rect 2620 4636 2628 4644
rect 2924 4636 2932 4644
rect 3148 4636 3156 4644
rect 4140 4636 4148 4644
rect 4380 4636 4388 4644
rect 4572 4636 4580 4644
rect 4620 4636 4628 4644
rect 4668 4636 4676 4644
rect 4844 4636 4852 4644
rect 4956 4636 4964 4644
rect 5132 4636 5140 4644
rect 5420 4636 5428 4644
rect 5612 4636 5620 4644
rect 5772 4636 5780 4644
rect 5964 4636 5972 4644
rect 6188 4636 6196 4644
rect 6252 4636 6260 4644
rect 6396 4636 6404 4644
rect 6476 4636 6484 4644
rect 6748 4636 6756 4644
rect 6924 4636 6932 4644
rect 6988 4636 6996 4644
rect 7052 4636 7060 4644
rect 7084 4636 7092 4644
rect 7164 4636 7172 4644
rect 7244 4636 7252 4644
rect 7308 4636 7316 4644
rect 7452 4636 7460 4644
rect 2243 4606 2251 4614
rect 2253 4606 2261 4614
rect 2263 4606 2271 4614
rect 2273 4606 2281 4614
rect 2283 4606 2291 4614
rect 2293 4606 2301 4614
rect 5251 4606 5259 4614
rect 5261 4606 5269 4614
rect 5271 4606 5279 4614
rect 5281 4606 5289 4614
rect 5291 4606 5299 4614
rect 5301 4606 5309 4614
rect 76 4576 84 4584
rect 252 4576 260 4584
rect 556 4576 564 4584
rect 620 4576 628 4584
rect 828 4576 836 4584
rect 924 4576 932 4584
rect 1388 4576 1396 4584
rect 1580 4576 1588 4584
rect 1740 4576 1748 4584
rect 1980 4576 1988 4584
rect 2316 4576 2324 4584
rect 2860 4576 2868 4584
rect 3404 4576 3412 4584
rect 3612 4576 3620 4584
rect 3980 4576 3988 4584
rect 4044 4576 4052 4584
rect 4108 4576 4116 4584
rect 4172 4576 4180 4584
rect 4652 4576 4660 4584
rect 5196 4576 5204 4584
rect 5388 4576 5396 4584
rect 5500 4576 5508 4584
rect 5852 4576 5860 4584
rect 6492 4576 6500 4584
rect 7132 4576 7140 4584
rect 12 4556 20 4564
rect 92 4536 100 4544
rect 220 4536 228 4544
rect 236 4536 244 4544
rect 460 4556 468 4564
rect 492 4556 500 4564
rect 604 4556 612 4564
rect 908 4556 916 4564
rect 1644 4556 1652 4564
rect 1708 4556 1716 4564
rect 2044 4556 2052 4564
rect 2060 4556 2068 4564
rect 2124 4556 2132 4564
rect 2444 4556 2452 4564
rect 2668 4556 2676 4564
rect 2988 4556 2996 4564
rect 3196 4556 3204 4564
rect 3532 4556 3540 4564
rect 332 4536 340 4544
rect 396 4536 404 4544
rect 508 4536 516 4544
rect 652 4536 660 4544
rect 844 4536 852 4544
rect 860 4536 868 4544
rect 1116 4536 1124 4544
rect 1148 4536 1156 4544
rect 1212 4536 1220 4544
rect 1532 4536 1540 4544
rect 1564 4536 1572 4544
rect 1660 4536 1668 4544
rect 1724 4536 1732 4544
rect 1788 4536 1796 4544
rect 1948 4536 1956 4544
rect 1964 4536 1972 4544
rect 2028 4536 2036 4544
rect 2076 4536 2084 4544
rect 2252 4536 2260 4544
rect 2508 4536 2516 4544
rect 2540 4536 2548 4544
rect 2604 4536 2612 4544
rect 2668 4536 2676 4544
rect 2716 4536 2724 4544
rect 3052 4536 3060 4544
rect 3148 4536 3156 4544
rect 3212 4536 3220 4544
rect 3340 4536 3348 4544
rect 3356 4536 3364 4544
rect 3420 4536 3428 4544
rect 3436 4536 3444 4544
rect 3484 4536 3492 4544
rect 4060 4556 4068 4564
rect 4124 4556 4132 4564
rect 4188 4556 4196 4564
rect 4556 4556 4564 4564
rect 4780 4556 4788 4564
rect 4940 4556 4948 4564
rect 5036 4556 5044 4564
rect 3580 4536 3588 4544
rect 3772 4536 3780 4544
rect 3868 4536 3876 4544
rect 4028 4536 4036 4544
rect 4092 4536 4100 4544
rect 4156 4536 4164 4544
rect 4220 4536 4228 4544
rect 4316 4536 4324 4544
rect 4348 4536 4356 4544
rect 4444 4536 4452 4544
rect 4668 4536 4676 4544
rect 4764 4536 4772 4544
rect 4876 4536 4884 4544
rect 5020 4536 5028 4544
rect 5036 4536 5044 4544
rect 5116 4536 5124 4544
rect 5180 4536 5188 4544
rect 5228 4532 5236 4540
rect 5244 4536 5252 4544
rect 5372 4556 5380 4564
rect 5564 4556 5572 4564
rect 5644 4556 5652 4564
rect 5788 4556 5796 4564
rect 5804 4556 5812 4564
rect 5868 4556 5876 4564
rect 5948 4556 5956 4564
rect 5980 4556 5988 4564
rect 6028 4556 6036 4564
rect 6236 4556 6244 4564
rect 6300 4556 6308 4564
rect 6620 4556 6628 4564
rect 7212 4556 7220 4564
rect 7340 4556 7348 4564
rect 7372 4556 7380 4564
rect 5404 4536 5412 4544
rect 5484 4536 5492 4544
rect 5516 4536 5524 4544
rect 5676 4536 5684 4544
rect 5708 4536 5716 4544
rect 5772 4536 5780 4544
rect 5932 4536 5940 4544
rect 5996 4536 6004 4544
rect 6156 4536 6164 4544
rect 6268 4536 6276 4544
rect 6332 4536 6340 4544
rect 6364 4536 6372 4544
rect 6380 4536 6388 4544
rect 6412 4536 6420 4544
rect 6444 4536 6452 4544
rect 6540 4536 6548 4544
rect 6636 4536 6644 4544
rect 6684 4536 6692 4544
rect 6844 4536 6852 4544
rect 6876 4536 6884 4544
rect 6908 4536 6916 4544
rect 6972 4536 6980 4544
rect 7196 4536 7204 4544
rect 7260 4536 7268 4544
rect 7308 4536 7316 4544
rect 7356 4536 7364 4544
rect 7452 4536 7460 4544
rect 44 4516 52 4524
rect 108 4516 116 4524
rect 156 4516 164 4524
rect 172 4516 180 4524
rect 220 4516 228 4524
rect 284 4516 292 4524
rect 348 4516 356 4524
rect 412 4516 420 4524
rect 428 4516 436 4524
rect 492 4516 500 4524
rect 540 4516 548 4524
rect 588 4516 596 4524
rect 636 4516 644 4524
rect 668 4516 676 4524
rect 796 4516 804 4524
rect 828 4516 836 4524
rect 860 4516 868 4524
rect 940 4516 948 4524
rect 1068 4516 1076 4524
rect 1164 4516 1172 4524
rect 1276 4516 1284 4524
rect 1324 4516 1332 4524
rect 1340 4516 1348 4524
rect 1356 4516 1364 4524
rect 1420 4516 1428 4524
rect 1468 4516 1476 4524
rect 1484 4516 1492 4524
rect 1500 4516 1508 4524
rect 1548 4516 1556 4524
rect 1612 4516 1620 4524
rect 1676 4516 1684 4524
rect 1740 4516 1748 4524
rect 1772 4516 1780 4524
rect 1788 4516 1796 4524
rect 1820 4516 1828 4524
rect 1868 4516 1876 4524
rect 1932 4516 1940 4524
rect 1980 4516 1988 4524
rect 2012 4516 2020 4524
rect 2092 4516 2100 4524
rect 380 4496 388 4504
rect 444 4496 452 4504
rect 700 4496 708 4504
rect 1244 4496 1252 4504
rect 1708 4496 1716 4504
rect 1900 4496 1908 4504
rect 1932 4496 1940 4504
rect 2172 4496 2180 4504
rect 2204 4516 2212 4524
rect 2236 4516 2244 4524
rect 2428 4516 2436 4524
rect 2524 4516 2532 4524
rect 2620 4516 2628 4524
rect 2684 4516 2692 4524
rect 2700 4516 2708 4524
rect 2732 4516 2740 4524
rect 2764 4516 2772 4524
rect 2844 4516 2852 4524
rect 2940 4516 2948 4524
rect 3052 4516 3060 4524
rect 2572 4496 2580 4504
rect 2796 4496 2804 4504
rect 3068 4496 3076 4504
rect 3148 4516 3156 4524
rect 3228 4516 3236 4524
rect 3292 4516 3300 4524
rect 3324 4516 3332 4524
rect 3372 4516 3380 4524
rect 3404 4516 3412 4524
rect 3116 4496 3124 4504
rect 3180 4496 3188 4504
rect 3260 4496 3268 4504
rect 3468 4516 3476 4524
rect 3500 4516 3508 4524
rect 3564 4516 3572 4524
rect 3596 4516 3604 4524
rect 3724 4516 3732 4524
rect 4012 4516 4020 4524
rect 4076 4516 4084 4524
rect 4140 4516 4148 4524
rect 4204 4516 4212 4524
rect 4268 4516 4276 4524
rect 4300 4516 4308 4524
rect 4412 4516 4420 4524
rect 4524 4516 4532 4524
rect 4572 4516 4580 4524
rect 4620 4516 4628 4524
rect 4828 4516 4836 4524
rect 4876 4516 4884 4524
rect 4988 4516 4996 4524
rect 5004 4516 5012 4524
rect 5132 4516 5140 4524
rect 5164 4516 5172 4524
rect 5260 4516 5268 4524
rect 5356 4516 5364 4524
rect 5420 4516 5428 4524
rect 5436 4516 5444 4524
rect 5516 4516 5524 4524
rect 5612 4516 5620 4524
rect 5660 4516 5668 4524
rect 5900 4516 5908 4524
rect 5948 4516 5956 4524
rect 5980 4516 5988 4524
rect 6076 4516 6084 4524
rect 6156 4516 6164 4524
rect 6188 4516 6196 4524
rect 6284 4516 6292 4524
rect 6396 4516 6404 4524
rect 6524 4516 6532 4524
rect 6572 4516 6580 4524
rect 6700 4516 6708 4524
rect 6828 4516 6836 4524
rect 6924 4516 6932 4524
rect 6956 4516 6964 4524
rect 7020 4516 7028 4524
rect 7052 4516 7060 4524
rect 7100 4516 7108 4524
rect 7212 4516 7220 4524
rect 7308 4516 7316 4524
rect 7404 4516 7412 4524
rect 7484 4536 7492 4544
rect 4268 4496 4276 4504
rect 5100 4496 5108 4504
rect 5548 4496 5556 4504
rect 5884 4496 5892 4504
rect 6108 4496 6116 4504
rect 6172 4496 6180 4504
rect 6332 4496 6340 4504
rect 6428 4496 6436 4504
rect 6476 4496 6484 4504
rect 6492 4496 6500 4504
rect 6556 4496 6564 4504
rect 6668 4496 6676 4504
rect 6796 4496 6804 4504
rect 6828 4496 6836 4504
rect 6908 4496 6916 4504
rect 6924 4496 6932 4504
rect 7036 4496 7044 4504
rect 7148 4496 7156 4504
rect 7436 4498 7444 4506
rect 7532 4496 7540 4504
rect 1164 4476 1172 4484
rect 2348 4476 2356 4484
rect 2892 4476 2900 4484
rect 4508 4476 4516 4484
rect 4860 4476 4868 4484
rect 6012 4476 6020 4484
rect 6204 4476 6212 4484
rect 6588 4476 6596 4484
rect 6796 4476 6804 4484
rect 7068 4476 7076 4484
rect 6220 4456 6228 4464
rect 6572 4456 6580 4464
rect 348 4436 356 4444
rect 956 4436 964 4444
rect 1292 4436 1300 4444
rect 1452 4436 1460 4444
rect 1852 4436 1860 4444
rect 2764 4436 2772 4444
rect 3324 4436 3332 4444
rect 4604 4436 4612 4444
rect 4700 4436 4708 4444
rect 4956 4436 4964 4444
rect 5132 4436 5140 4444
rect 5564 4436 5572 4444
rect 5708 4436 5716 4444
rect 6028 4436 6036 4444
rect 6236 4436 6244 4444
rect 6348 4436 6356 4444
rect 6988 4436 6996 4444
rect 7052 4436 7060 4444
rect 7180 4436 7188 4444
rect 7292 4436 7300 4444
rect 7500 4436 7508 4444
rect 739 4406 747 4414
rect 749 4406 757 4414
rect 759 4406 767 4414
rect 769 4406 777 4414
rect 779 4406 787 4414
rect 789 4406 797 4414
rect 3747 4406 3755 4414
rect 3757 4406 3765 4414
rect 3767 4406 3775 4414
rect 3777 4406 3785 4414
rect 3787 4406 3795 4414
rect 3797 4406 3805 4414
rect 6755 4406 6763 4414
rect 6765 4406 6773 4414
rect 6775 4406 6783 4414
rect 6785 4406 6793 4414
rect 6795 4406 6803 4414
rect 6805 4406 6813 4414
rect 556 4376 564 4384
rect 844 4376 852 4384
rect 1020 4376 1028 4384
rect 1228 4376 1236 4384
rect 1740 4376 1748 4384
rect 1836 4376 1844 4384
rect 2268 4376 2276 4384
rect 2332 4376 2340 4384
rect 2348 4376 2356 4384
rect 2716 4376 2724 4384
rect 3132 4376 3140 4384
rect 3436 4376 3444 4384
rect 3852 4376 3860 4384
rect 3932 4376 3940 4384
rect 3980 4376 3988 4384
rect 4028 4376 4036 4384
rect 4236 4376 4244 4384
rect 4284 4376 4292 4384
rect 4972 4376 4980 4384
rect 5036 4376 5044 4384
rect 5468 4376 5476 4384
rect 5676 4376 5684 4384
rect 5948 4376 5956 4384
rect 5980 4376 5988 4384
rect 6444 4376 6452 4384
rect 6492 4376 6500 4384
rect 6588 4376 6596 4384
rect 6652 4376 6660 4384
rect 6972 4376 6980 4384
rect 7404 4376 7412 4384
rect 7468 4376 7476 4384
rect 460 4356 468 4364
rect 1644 4356 1652 4364
rect 5836 4356 5844 4364
rect 588 4336 596 4344
rect 956 4336 964 4344
rect 1180 4336 1188 4344
rect 1356 4336 1364 4344
rect 1516 4336 1524 4344
rect 3180 4336 3188 4344
rect 4812 4336 4820 4344
rect 4908 4336 4916 4344
rect 5548 4336 5556 4344
rect 5964 4336 5972 4344
rect 6572 4336 6580 4344
rect 1052 4316 1060 4324
rect 1212 4316 1220 4324
rect 76 4296 84 4304
rect 124 4296 132 4304
rect 204 4296 212 4304
rect 300 4296 308 4304
rect 332 4296 340 4304
rect 380 4296 388 4304
rect 396 4296 404 4304
rect 412 4296 420 4304
rect 428 4296 436 4304
rect 476 4296 484 4304
rect 524 4296 532 4304
rect 572 4296 580 4304
rect 588 4296 596 4304
rect 636 4296 644 4304
rect 652 4296 660 4304
rect 732 4296 740 4304
rect 812 4296 820 4304
rect 908 4296 916 4304
rect 956 4296 964 4304
rect 972 4296 980 4304
rect 1020 4296 1028 4304
rect 1100 4296 1108 4304
rect 1148 4296 1156 4304
rect 1180 4296 1188 4304
rect 1260 4296 1268 4304
rect 1292 4296 1300 4304
rect 1340 4296 1348 4304
rect 1356 4296 1364 4304
rect 1404 4296 1412 4304
rect 2396 4316 2404 4324
rect 2780 4316 2788 4324
rect 3644 4316 3652 4324
rect 3708 4316 3716 4324
rect 3996 4316 4004 4324
rect 4252 4316 4260 4324
rect 4780 4316 4788 4324
rect 4844 4316 4852 4324
rect 4860 4316 4868 4324
rect 5820 4316 5828 4324
rect 5852 4316 5860 4324
rect 6028 4316 6036 4324
rect 6060 4316 6068 4324
rect 6348 4316 6356 4324
rect 6540 4316 6548 4324
rect 6764 4316 6772 4324
rect 6844 4316 6852 4324
rect 7036 4316 7044 4324
rect 7228 4316 7236 4324
rect 1484 4296 1492 4304
rect 1580 4296 1588 4304
rect 1596 4296 1604 4304
rect 1612 4296 1620 4304
rect 1660 4296 1668 4304
rect 1692 4296 1700 4304
rect 1708 4296 1716 4304
rect 1756 4296 1764 4304
rect 1804 4296 1812 4304
rect 1852 4296 1860 4304
rect 1868 4296 1876 4304
rect 2012 4294 2020 4302
rect 2076 4296 2084 4304
rect 2172 4296 2180 4304
rect 2188 4296 2196 4304
rect 2300 4296 2308 4304
rect 2396 4296 2404 4304
rect 2428 4296 2436 4304
rect 2476 4296 2484 4304
rect 2508 4296 2516 4304
rect 2524 4296 2532 4304
rect 2556 4296 2564 4304
rect 2604 4296 2612 4304
rect 2652 4296 2660 4304
rect 2668 4296 2676 4304
rect 2684 4296 2692 4304
rect 2748 4296 2756 4304
rect 2828 4296 2836 4304
rect 2860 4296 2868 4304
rect 2876 4296 2884 4304
rect 2892 4296 2900 4304
rect 2940 4296 2948 4304
rect 2988 4296 2996 4304
rect 3004 4296 3012 4304
rect 3020 4296 3028 4304
rect 3036 4296 3044 4304
rect 3084 4296 3092 4304
rect 3116 4296 3124 4304
rect 3196 4296 3204 4304
rect 3308 4296 3316 4304
rect 3324 4296 3332 4304
rect 3404 4296 3412 4304
rect 3420 4296 3428 4304
rect 3468 4296 3476 4304
rect 3500 4296 3508 4304
rect 3516 4296 3524 4304
rect 3564 4296 3572 4304
rect 3612 4296 3620 4304
rect 3676 4296 3684 4304
rect 3724 4296 3732 4304
rect 3804 4296 3812 4304
rect 3820 4296 3828 4304
rect 3868 4296 3876 4304
rect 3900 4296 3908 4304
rect 3948 4296 3956 4304
rect 4028 4296 4036 4304
rect 4108 4294 4116 4302
rect 4172 4296 4180 4304
rect 4252 4296 4260 4304
rect 4284 4296 4292 4304
rect 4316 4296 4324 4304
rect 4364 4296 4372 4304
rect 4428 4294 4436 4302
rect 4588 4296 4596 4304
rect 4652 4296 4660 4304
rect 4748 4296 4756 4304
rect 4828 4296 4836 4304
rect 4860 4296 4868 4304
rect 4940 4296 4948 4304
rect 4988 4296 4996 4304
rect 5068 4296 5076 4304
rect 5100 4296 5108 4304
rect 5132 4296 5140 4304
rect 5148 4296 5156 4304
rect 5212 4296 5220 4304
rect 5244 4296 5252 4304
rect 5340 4296 5348 4304
rect 5388 4296 5396 4304
rect 5436 4296 5444 4304
rect 5724 4296 5732 4304
rect 5948 4296 5956 4304
rect 6076 4296 6084 4304
rect 6140 4296 6148 4304
rect 6220 4296 6228 4304
rect 6268 4296 6276 4304
rect 6524 4296 6532 4304
rect 6556 4296 6564 4304
rect 6620 4296 6628 4304
rect 6908 4296 6916 4304
rect 6924 4296 6932 4304
rect 6988 4296 6996 4304
rect 7052 4296 7060 4304
rect 7084 4296 7092 4304
rect 7180 4296 7188 4304
rect 7292 4296 7300 4304
rect 7340 4296 7348 4304
rect 7372 4296 7380 4304
rect 7404 4296 7412 4304
rect 7436 4296 7444 4304
rect 7564 4296 7572 4304
rect 220 4276 228 4284
rect 236 4276 244 4284
rect 508 4276 516 4284
rect 572 4276 580 4284
rect 780 4276 788 4284
rect 796 4276 804 4284
rect 860 4276 868 4284
rect 972 4276 980 4284
rect 1036 4276 1044 4284
rect 1100 4276 1108 4284
rect 1116 4276 1124 4284
rect 1164 4276 1172 4284
rect 1276 4276 1284 4284
rect 1340 4276 1348 4284
rect 1388 4276 1396 4284
rect 1452 4276 1460 4284
rect 1468 4276 1476 4284
rect 1532 4276 1540 4284
rect 2044 4276 2052 4284
rect 2092 4276 2100 4284
rect 268 4256 276 4264
rect 364 4256 372 4264
rect 620 4256 628 4264
rect 876 4256 884 4264
rect 924 4256 932 4264
rect 1052 4256 1060 4264
rect 1388 4256 1396 4264
rect 1548 4256 1556 4264
rect 2412 4276 2420 4284
rect 2444 4276 2452 4284
rect 2460 4276 2468 4284
rect 2492 4276 2500 4284
rect 2524 4276 2532 4284
rect 2572 4276 2580 4284
rect 2732 4276 2740 4284
rect 2796 4276 2804 4284
rect 2844 4276 2852 4284
rect 2924 4276 2932 4284
rect 3116 4276 3124 4284
rect 3580 4276 3588 4284
rect 3660 4276 3668 4284
rect 3724 4276 3732 4284
rect 4044 4276 4052 4284
rect 4300 4276 4308 4284
rect 4332 4276 4340 4284
rect 4444 4276 4452 4284
rect 4572 4276 4580 4284
rect 4636 4276 4644 4284
rect 4748 4276 4756 4284
rect 4780 4276 4788 4284
rect 5020 4276 5028 4284
rect 5084 4276 5092 4284
rect 5484 4276 5492 4284
rect 5820 4276 5828 4284
rect 5852 4276 5860 4284
rect 6028 4276 6036 4284
rect 6348 4276 6356 4284
rect 6364 4276 6372 4284
rect 6412 4276 6420 4284
rect 6444 4276 6452 4284
rect 6604 4276 6612 4284
rect 6716 4276 6724 4284
rect 6812 4276 6820 4284
rect 6892 4276 6900 4284
rect 6924 4276 6932 4284
rect 6972 4276 6980 4284
rect 6988 4276 6996 4284
rect 7036 4276 7044 4284
rect 7228 4276 7236 4284
rect 7260 4276 7268 4284
rect 7276 4276 7284 4284
rect 7452 4276 7460 4284
rect 7500 4276 7508 4284
rect 2140 4256 2148 4264
rect 2572 4256 2580 4264
rect 2796 4256 2804 4264
rect 2828 4256 2836 4264
rect 2956 4256 2964 4264
rect 3148 4256 3156 4264
rect 3548 4256 3556 4264
rect 3644 4256 3652 4264
rect 4364 4256 4372 4264
rect 4700 4256 4708 4264
rect 4908 4256 4916 4264
rect 5180 4256 5188 4264
rect 5244 4256 5252 4264
rect 5372 4256 5380 4264
rect 5596 4256 5604 4264
rect 5628 4256 5636 4264
rect 5644 4256 5652 4264
rect 5676 4256 5684 4264
rect 5740 4256 5748 4264
rect 5788 4256 5796 4264
rect 5868 4256 5876 4264
rect 5996 4256 6004 4264
rect 6172 4256 6180 4264
rect 6236 4256 6244 4264
rect 6284 4256 6292 4264
rect 6476 4256 6484 4264
rect 6508 4256 6516 4264
rect 6668 4256 6676 4264
rect 6716 4256 6724 4264
rect 6860 4256 6868 4264
rect 6972 4256 6980 4264
rect 7084 4256 7092 4264
rect 7116 4256 7124 4264
rect 7132 4256 7140 4264
rect 7164 4256 7172 4264
rect 7340 4256 7348 4264
rect 7468 4256 7476 4264
rect 188 4236 196 4244
rect 1292 4236 1300 4244
rect 1884 4236 1892 4244
rect 2108 4236 2116 4244
rect 3388 4236 3396 4244
rect 3980 4236 3988 4244
rect 4556 4236 4564 4244
rect 4620 4236 4628 4244
rect 4684 4236 4692 4244
rect 4780 4236 4788 4244
rect 4972 4236 4980 4244
rect 5036 4236 5044 4244
rect 5420 4236 5428 4244
rect 6108 4236 6116 4244
rect 6188 4236 6196 4244
rect 6252 4236 6260 4244
rect 6828 4236 6836 4244
rect 6876 4236 6884 4244
rect 7020 4236 7028 4244
rect 7228 4236 7236 4244
rect 2243 4206 2251 4214
rect 2253 4206 2261 4214
rect 2263 4206 2271 4214
rect 2273 4206 2281 4214
rect 2283 4206 2291 4214
rect 2293 4206 2301 4214
rect 5251 4206 5259 4214
rect 5261 4206 5269 4214
rect 5271 4206 5279 4214
rect 5281 4206 5289 4214
rect 5291 4206 5299 4214
rect 5301 4206 5309 4214
rect 188 4176 196 4184
rect 364 4176 372 4184
rect 1068 4176 1076 4184
rect 1596 4176 1604 4184
rect 1868 4176 1876 4184
rect 1980 4176 1988 4184
rect 2236 4176 2244 4184
rect 2428 4176 2436 4184
rect 2588 4176 2596 4184
rect 2812 4176 2820 4184
rect 2828 4176 2836 4184
rect 3308 4176 3316 4184
rect 3772 4176 3780 4184
rect 4060 4176 4068 4184
rect 4300 4176 4308 4184
rect 4380 4176 4388 4184
rect 4908 4176 4916 4184
rect 5148 4176 5156 4184
rect 5196 4176 5204 4184
rect 5260 4176 5268 4184
rect 5372 4176 5380 4184
rect 5804 4176 5812 4184
rect 5836 4176 5844 4184
rect 6092 4176 6100 4184
rect 6204 4176 6212 4184
rect 6540 4176 6548 4184
rect 6636 4176 6644 4184
rect 6716 4176 6724 4184
rect 6828 4176 6836 4184
rect 7404 4176 7412 4184
rect 7484 4176 7492 4184
rect 7516 4176 7524 4184
rect 220 4136 228 4144
rect 268 4156 276 4164
rect 348 4156 356 4164
rect 812 4156 820 4164
rect 1196 4156 1204 4164
rect 1612 4156 1620 4164
rect 1660 4156 1668 4164
rect 1900 4156 1908 4164
rect 2364 4156 2372 4164
rect 3372 4156 3380 4164
rect 4076 4156 4084 4164
rect 4140 4156 4148 4164
rect 4396 4156 4404 4164
rect 4476 4156 4484 4164
rect 4524 4156 4532 4164
rect 4604 4156 4612 4164
rect 460 4136 468 4144
rect 556 4136 564 4144
rect 652 4136 660 4144
rect 796 4136 804 4144
rect 876 4136 884 4144
rect 940 4136 948 4144
rect 956 4136 964 4144
rect 1004 4136 1012 4144
rect 1052 4136 1060 4144
rect 1260 4136 1268 4144
rect 1372 4136 1380 4144
rect 1468 4136 1476 4144
rect 1532 4136 1540 4144
rect 1676 4136 1684 4144
rect 1708 4136 1716 4144
rect 1740 4136 1748 4144
rect 1756 4136 1764 4144
rect 1804 4136 1812 4144
rect 1820 4136 1828 4144
rect 1884 4136 1892 4144
rect 1948 4136 1956 4144
rect 2028 4136 2036 4144
rect 2044 4136 2052 4144
rect 2156 4136 2164 4144
rect 2476 4136 2484 4144
rect 2572 4136 2580 4144
rect 2748 4136 2756 4144
rect 3020 4136 3028 4144
rect 3132 4136 3140 4144
rect 76 4116 84 4124
rect 124 4116 132 4124
rect 204 4116 212 4124
rect 236 4116 244 4124
rect 300 4116 308 4124
rect 316 4116 324 4124
rect 476 4116 484 4124
rect 572 4116 580 4124
rect 572 4096 580 4104
rect 668 4116 676 4124
rect 684 4116 692 4124
rect 732 4116 740 4124
rect 860 4116 868 4124
rect 892 4116 900 4124
rect 924 4116 932 4124
rect 988 4116 996 4124
rect 1036 4116 1044 4124
rect 1196 4118 1204 4126
rect 1276 4116 1284 4124
rect 1292 4116 1300 4124
rect 620 4096 628 4104
rect 844 4096 852 4104
rect 1004 4096 1012 4104
rect 1356 4116 1364 4124
rect 1388 4116 1396 4124
rect 1404 4116 1412 4124
rect 1452 4116 1460 4124
rect 1516 4116 1524 4124
rect 1564 4116 1572 4124
rect 1580 4116 1588 4124
rect 1628 4116 1636 4124
rect 1724 4116 1732 4124
rect 1324 4096 1332 4104
rect 1788 4116 1796 4124
rect 1836 4116 1844 4124
rect 1868 4116 1876 4124
rect 1932 4116 1940 4124
rect 2060 4116 2068 4124
rect 1900 4096 1908 4104
rect 2092 4096 2100 4104
rect 2124 4116 2132 4124
rect 2140 4116 2148 4124
rect 2348 4116 2356 4124
rect 2460 4116 2468 4124
rect 2508 4096 2516 4104
rect 2556 4116 2564 4124
rect 2700 4116 2708 4124
rect 2780 4116 2788 4124
rect 2908 4116 2916 4124
rect 2956 4118 2964 4126
rect 3292 4136 3300 4144
rect 3484 4136 3492 4144
rect 3548 4136 3556 4144
rect 3580 4136 3588 4144
rect 3612 4136 3620 4144
rect 3916 4136 3924 4144
rect 4012 4136 4020 4144
rect 4044 4136 4052 4144
rect 4124 4136 4132 4144
rect 4188 4136 4196 4144
rect 4284 4136 4292 4144
rect 4348 4136 4356 4144
rect 4412 4136 4420 4144
rect 4748 4156 4756 4164
rect 4972 4156 4980 4164
rect 5484 4156 5492 4164
rect 5692 4156 5700 4164
rect 5852 4156 5860 4164
rect 6252 4156 6260 4164
rect 6284 4156 6292 4164
rect 6380 4156 6388 4164
rect 6492 4156 6500 4164
rect 6988 4156 6996 4164
rect 7180 4156 7188 4164
rect 7340 4156 7348 4164
rect 7420 4156 7428 4164
rect 7500 4156 7508 4164
rect 4428 4132 4436 4140
rect 4828 4132 4836 4140
rect 4860 4136 4868 4144
rect 5212 4136 5220 4144
rect 5228 4132 5236 4140
rect 5484 4136 5492 4144
rect 5500 4136 5508 4144
rect 5532 4136 5540 4144
rect 5548 4136 5556 4144
rect 5612 4136 5620 4144
rect 5660 4136 5668 4144
rect 5756 4136 5764 4144
rect 5916 4136 5924 4144
rect 6012 4136 6020 4144
rect 6028 4136 6036 4144
rect 6124 4136 6132 4144
rect 6140 4136 6148 4144
rect 6188 4136 6196 4144
rect 6300 4136 6308 4144
rect 6332 4136 6340 4144
rect 6396 4136 6404 4144
rect 6556 4136 6564 4144
rect 3020 4116 3028 4124
rect 3036 4096 3044 4104
rect 3148 4116 3156 4124
rect 3084 4096 3092 4104
rect 3196 4096 3204 4104
rect 3244 4116 3252 4124
rect 3276 4116 3284 4124
rect 3340 4116 3348 4124
rect 3388 4116 3396 4124
rect 3404 4116 3412 4124
rect 3452 4116 3460 4124
rect 3500 4116 3508 4124
rect 3644 4118 3652 4126
rect 3852 4116 3860 4124
rect 3900 4116 3908 4124
rect 3996 4116 4004 4124
rect 4028 4116 4036 4124
rect 4092 4116 4100 4124
rect 4172 4116 4180 4124
rect 4236 4116 4244 4124
rect 4252 4116 4260 4124
rect 4332 4116 4340 4124
rect 4364 4116 4372 4124
rect 4508 4116 4516 4124
rect 4556 4116 4564 4124
rect 4620 4116 4628 4124
rect 4652 4116 4660 4124
rect 4700 4116 4708 4124
rect 4748 4116 4756 4124
rect 5004 4116 5012 4124
rect 5052 4116 5060 4124
rect 5100 4116 5108 4124
rect 5116 4116 5124 4124
rect 5164 4116 5172 4124
rect 5308 4116 5316 4124
rect 5388 4116 5396 4124
rect 5436 4116 5444 4124
rect 5628 4116 5636 4124
rect 5708 4116 5716 4124
rect 5740 4116 5748 4124
rect 5772 4116 5780 4124
rect 5820 4116 5828 4124
rect 5868 4116 5876 4124
rect 6172 4116 6180 4124
rect 6236 4116 6244 4124
rect 6284 4116 6292 4124
rect 6348 4116 6356 4124
rect 6412 4116 6420 4124
rect 6556 4116 6564 4124
rect 6668 4136 6676 4144
rect 6844 4136 6852 4144
rect 6940 4136 6948 4144
rect 7004 4136 7012 4144
rect 7164 4136 7172 4144
rect 7244 4136 7252 4144
rect 7308 4136 7316 4144
rect 7356 4136 7364 4144
rect 7452 4136 7460 4144
rect 6684 4116 6692 4124
rect 6732 4116 6740 4124
rect 6860 4116 6868 4124
rect 6892 4116 6900 4124
rect 7020 4116 7028 4124
rect 7212 4116 7220 4124
rect 7292 4116 7300 4124
rect 7372 4116 7380 4124
rect 7548 4116 7556 4124
rect 3548 4096 3556 4104
rect 3964 4096 3972 4104
rect 4140 4096 4148 4104
rect 4300 4096 4308 4104
rect 5580 4096 5588 4104
rect 5708 4096 5716 4104
rect 5740 4096 5748 4104
rect 6140 4096 6148 4104
rect 6492 4096 6500 4104
rect 6892 4096 6900 4104
rect 7052 4096 7060 4104
rect 7260 4096 7268 4104
rect 7452 4096 7460 4104
rect 7484 4096 7492 4104
rect 924 4076 932 4084
rect 2556 4076 2564 4084
rect 5068 4076 5076 4084
rect 7244 4076 7252 4084
rect 332 4036 340 4044
rect 1436 4036 1444 4044
rect 1980 4036 1988 4044
rect 3244 4036 3252 4044
rect 3436 4036 3444 4044
rect 3884 4036 3892 4044
rect 3948 4036 3956 4044
rect 4204 4036 4212 4044
rect 4460 4036 4468 4044
rect 4476 4036 4484 4044
rect 4604 4036 4612 4044
rect 4684 4036 4692 4044
rect 5020 4036 5028 4044
rect 5196 4036 5204 4044
rect 5420 4036 5428 4044
rect 5900 4036 5908 4044
rect 5964 4036 5972 4044
rect 6300 4036 6308 4044
rect 6908 4036 6916 4044
rect 7132 4036 7140 4044
rect 7292 4036 7300 4044
rect 739 4006 747 4014
rect 749 4006 757 4014
rect 759 4006 767 4014
rect 769 4006 777 4014
rect 779 4006 787 4014
rect 789 4006 797 4014
rect 3747 4006 3755 4014
rect 3757 4006 3765 4014
rect 3767 4006 3775 4014
rect 3777 4006 3785 4014
rect 3787 4006 3795 4014
rect 3797 4006 3805 4014
rect 6755 4006 6763 4014
rect 6765 4006 6773 4014
rect 6775 4006 6783 4014
rect 6785 4006 6793 4014
rect 6795 4006 6803 4014
rect 6805 4006 6813 4014
rect 492 3976 500 3984
rect 1068 3976 1076 3984
rect 1788 3976 1796 3984
rect 1964 3976 1972 3984
rect 3052 3976 3060 3984
rect 4076 3976 4084 3984
rect 5068 3976 5076 3984
rect 5164 3976 5172 3984
rect 5660 3976 5668 3984
rect 6860 3976 6868 3984
rect 7260 3976 7268 3984
rect 2668 3956 2676 3964
rect 204 3936 212 3944
rect 460 3936 468 3944
rect 764 3936 772 3944
rect 1356 3936 1364 3944
rect 1548 3936 1556 3944
rect 1580 3936 1588 3944
rect 1772 3936 1780 3944
rect 2396 3936 2404 3944
rect 2620 3936 2628 3944
rect 2972 3936 2980 3944
rect 3756 3936 3764 3944
rect 5116 3936 5124 3944
rect 5340 3936 5348 3944
rect 5804 3936 5812 3944
rect 7100 3936 7108 3944
rect 7244 3936 7252 3944
rect 236 3916 244 3924
rect 76 3896 84 3904
rect 124 3896 132 3904
rect 556 3916 564 3924
rect 860 3916 868 3924
rect 1516 3916 1524 3924
rect 2252 3916 2260 3924
rect 284 3896 292 3904
rect 364 3894 372 3902
rect 524 3896 532 3904
rect 540 3896 548 3904
rect 636 3896 644 3904
rect 908 3896 916 3904
rect 956 3896 964 3904
rect 972 3896 980 3904
rect 988 3896 996 3904
rect 1036 3896 1044 3904
rect 1100 3896 1108 3904
rect 1116 3896 1124 3904
rect 1292 3894 1300 3902
rect 1404 3896 1412 3904
rect 1420 3896 1428 3904
rect 1484 3896 1492 3904
rect 1548 3896 1556 3904
rect 1644 3894 1652 3902
rect 1820 3896 1828 3904
rect 1852 3896 1860 3904
rect 1900 3896 1908 3904
rect 1916 3896 1924 3904
rect 1948 3896 1956 3904
rect 1996 3896 2004 3904
rect 2012 3896 2020 3904
rect 2140 3896 2148 3904
rect 2364 3916 2372 3924
rect 2716 3916 2724 3924
rect 2364 3896 2372 3904
rect 2508 3896 2516 3904
rect 2588 3896 2596 3904
rect 2636 3896 2644 3904
rect 3036 3916 3044 3924
rect 3884 3916 3892 3924
rect 4204 3916 4212 3924
rect 4444 3916 4452 3924
rect 4828 3916 4836 3924
rect 4876 3916 4884 3924
rect 4924 3916 4932 3924
rect 5212 3916 5220 3924
rect 5436 3916 5444 3924
rect 5788 3916 5796 3924
rect 5836 3916 5844 3924
rect 5884 3916 5892 3924
rect 5948 3916 5956 3924
rect 5964 3916 5972 3924
rect 6988 3916 6996 3924
rect 7180 3916 7188 3924
rect 7276 3916 7284 3924
rect 7356 3916 7364 3924
rect 7388 3916 7396 3924
rect 7452 3916 7460 3924
rect 2748 3896 2756 3904
rect 2780 3896 2788 3904
rect 2844 3894 2852 3902
rect 2908 3896 2916 3904
rect 2988 3896 2996 3904
rect 3116 3896 3124 3904
rect 3180 3894 3188 3902
rect 3260 3896 3268 3904
rect 3308 3896 3316 3904
rect 3388 3896 3396 3904
rect 3420 3896 3428 3904
rect 3516 3896 3524 3904
rect 3564 3896 3572 3904
rect 3628 3894 3636 3902
rect 3820 3896 3828 3904
rect 3948 3894 3956 3902
rect 4124 3896 4132 3904
rect 4188 3896 4196 3904
rect 4236 3896 4244 3904
rect 4396 3896 4404 3904
rect 4476 3896 4484 3904
rect 4524 3896 4532 3904
rect 4668 3896 4676 3904
rect 4732 3896 4740 3904
rect 4988 3896 4996 3904
rect 5036 3896 5044 3904
rect 5084 3896 5092 3904
rect 5132 3896 5140 3904
rect 5532 3896 5540 3904
rect 5644 3896 5652 3904
rect 5692 3896 5700 3904
rect 5740 3896 5748 3904
rect 5820 3896 5828 3904
rect 204 3876 212 3884
rect 252 3876 260 3884
rect 300 3876 308 3884
rect 332 3876 340 3884
rect 508 3876 516 3884
rect 588 3876 596 3884
rect 764 3876 772 3884
rect 828 3876 836 3884
rect 1052 3876 1060 3884
rect 1260 3876 1268 3884
rect 1388 3876 1396 3884
rect 1468 3876 1476 3884
rect 1516 3876 1524 3884
rect 1532 3876 1540 3884
rect 1612 3876 1620 3884
rect 1836 3876 1844 3884
rect 2220 3876 2228 3884
rect 2380 3876 2388 3884
rect 2684 3876 2692 3884
rect 2780 3876 2788 3884
rect 2988 3876 2996 3884
rect 3212 3876 3220 3884
rect 3244 3876 3252 3884
rect 3308 3876 3316 3884
rect 3532 3876 3540 3884
rect 3644 3876 3652 3884
rect 3836 3876 3844 3884
rect 3868 3876 3876 3884
rect 3964 3876 3972 3884
rect 4092 3876 4100 3884
rect 4156 3876 4164 3884
rect 4268 3876 4276 3884
rect 4284 3876 4292 3884
rect 4348 3876 4356 3884
rect 4396 3876 4404 3884
rect 4412 3876 4420 3884
rect 4460 3876 4468 3884
rect 4540 3876 4548 3884
rect 4572 3876 4580 3884
rect 4636 3880 4644 3888
rect 4652 3876 4660 3884
rect 4700 3876 4708 3884
rect 4716 3876 4724 3884
rect 4780 3876 4788 3884
rect 4860 3876 4868 3884
rect 4908 3876 4916 3884
rect 4956 3876 4964 3884
rect 4972 3876 4980 3884
rect 5180 3876 5188 3884
rect 5228 3876 5236 3884
rect 5388 3876 5396 3884
rect 5404 3876 5412 3884
rect 5436 3876 5444 3884
rect 5484 3876 5492 3884
rect 5596 3876 5604 3884
rect 5628 3876 5636 3884
rect 5708 3876 5716 3884
rect 5916 3896 5924 3904
rect 5932 3876 5940 3884
rect 6124 3896 6132 3904
rect 6188 3896 6196 3904
rect 6252 3896 6260 3904
rect 6428 3896 6436 3904
rect 6476 3896 6484 3904
rect 6732 3896 6740 3904
rect 6748 3896 6756 3904
rect 6892 3896 6900 3904
rect 6940 3896 6948 3904
rect 7036 3896 7044 3904
rect 7100 3896 7108 3904
rect 7260 3896 7268 3904
rect 6012 3876 6020 3884
rect 6108 3876 6116 3884
rect 6380 3876 6388 3884
rect 6412 3876 6420 3884
rect 6508 3876 6516 3884
rect 6572 3876 6580 3884
rect 6620 3876 6628 3884
rect 6668 3880 6676 3888
rect 6684 3876 6692 3884
rect 6908 3876 6916 3884
rect 6956 3876 6964 3884
rect 7212 3876 7220 3884
rect 7308 3896 7316 3904
rect 7404 3896 7412 3904
rect 7516 3896 7524 3904
rect 7356 3876 7364 3884
rect 7500 3876 7508 3884
rect 7564 3876 7572 3884
rect 876 3856 884 3864
rect 924 3856 932 3864
rect 1148 3856 1156 3864
rect 1356 3856 1364 3864
rect 2156 3856 2164 3864
rect 2524 3856 2532 3864
rect 3036 3856 3044 3864
rect 3564 3856 3572 3864
rect 4140 3856 4148 3864
rect 4268 3856 4276 3864
rect 5500 3856 5508 3864
rect 5548 3856 5556 3864
rect 5724 3856 5732 3864
rect 5772 3856 5780 3864
rect 6124 3856 6132 3864
rect 6188 3856 6196 3864
rect 6204 3856 6212 3864
rect 6268 3856 6276 3864
rect 6316 3856 6324 3864
rect 6348 3856 6356 3864
rect 6380 3856 6388 3864
rect 6444 3856 6452 3864
rect 6492 3856 6500 3864
rect 6972 3856 6980 3864
rect 7004 3856 7012 3864
rect 7052 3856 7060 3864
rect 7164 3856 7172 3864
rect 7436 3856 7444 3864
rect 7500 3856 7508 3864
rect 844 3836 852 3844
rect 892 3836 900 3844
rect 940 3836 948 3844
rect 1132 3836 1140 3844
rect 1164 3836 1172 3844
rect 1452 3836 1460 3844
rect 2028 3836 2036 3844
rect 3260 3836 3268 3844
rect 3324 3836 3332 3844
rect 4364 3836 4372 3844
rect 4428 3836 4436 3844
rect 4508 3836 4516 3844
rect 4556 3836 4564 3844
rect 4764 3836 4772 3844
rect 4812 3836 4820 3844
rect 4828 3836 4836 3844
rect 4876 3836 4884 3844
rect 4924 3836 4932 3844
rect 5020 3836 5028 3844
rect 5164 3836 5172 3844
rect 5228 3836 5236 3844
rect 5420 3836 5428 3844
rect 5516 3836 5524 3844
rect 5628 3836 5636 3844
rect 5964 3836 5972 3844
rect 6396 3836 6404 3844
rect 6460 3836 6468 3844
rect 6588 3836 6596 3844
rect 6844 3836 6852 3844
rect 7180 3836 7188 3844
rect 7340 3836 7348 3844
rect 7372 3836 7380 3844
rect 2243 3806 2251 3814
rect 2253 3806 2261 3814
rect 2263 3806 2271 3814
rect 2273 3806 2281 3814
rect 2283 3806 2291 3814
rect 2293 3806 2301 3814
rect 5251 3806 5259 3814
rect 5261 3806 5269 3814
rect 5271 3806 5279 3814
rect 5281 3806 5289 3814
rect 5291 3806 5299 3814
rect 5301 3806 5309 3814
rect 188 3776 196 3784
rect 348 3776 356 3784
rect 716 3776 724 3784
rect 908 3776 916 3784
rect 1420 3776 1428 3784
rect 1500 3776 1508 3784
rect 1692 3776 1700 3784
rect 1820 3776 1828 3784
rect 1884 3776 1892 3784
rect 2124 3776 2132 3784
rect 2252 3776 2260 3784
rect 2636 3776 2644 3784
rect 3132 3776 3140 3784
rect 3356 3776 3364 3784
rect 3420 3776 3428 3784
rect 3612 3776 3620 3784
rect 4092 3776 4100 3784
rect 5836 3776 5844 3784
rect 6604 3776 6612 3784
rect 204 3756 212 3764
rect 364 3756 372 3764
rect 1996 3756 2004 3764
rect 2076 3756 2084 3764
rect 3212 3756 3220 3764
rect 3340 3756 3348 3764
rect 284 3736 292 3744
rect 332 3736 340 3744
rect 412 3736 420 3744
rect 428 3736 436 3744
rect 492 3736 500 3744
rect 524 3736 532 3744
rect 556 3736 564 3744
rect 796 3736 804 3744
rect 924 3736 932 3744
rect 940 3736 948 3744
rect 1004 3736 1012 3744
rect 1020 3736 1028 3744
rect 1052 3736 1060 3744
rect 1116 3736 1124 3744
rect 1132 3736 1140 3744
rect 1196 3736 1204 3744
rect 1228 3736 1236 3744
rect 1260 3736 1268 3744
rect 1484 3736 1492 3744
rect 1612 3736 1620 3744
rect 1628 3736 1636 3744
rect 1836 3736 1844 3744
rect 1932 3736 1940 3744
rect 1996 3736 2004 3744
rect 2140 3736 2148 3744
rect 2348 3736 2356 3744
rect 2396 3736 2404 3744
rect 2444 3736 2452 3744
rect 2476 3736 2484 3744
rect 2524 3736 2532 3744
rect 2876 3736 2884 3744
rect 2940 3736 2948 3744
rect 2972 3736 2980 3744
rect 3148 3736 3156 3744
rect 3212 3736 3220 3744
rect 3260 3736 3268 3744
rect 3324 3736 3332 3744
rect 3404 3736 3412 3744
rect 3452 3756 3460 3764
rect 3964 3756 3972 3764
rect 4124 3756 4132 3764
rect 4172 3756 4180 3764
rect 3500 3736 3508 3744
rect 3596 3736 3604 3744
rect 3852 3736 3860 3744
rect 3932 3736 3940 3744
rect 4364 3756 4372 3764
rect 4444 3756 4452 3764
rect 4636 3756 4644 3764
rect 4668 3756 4676 3764
rect 4684 3756 4692 3764
rect 4716 3756 4724 3764
rect 4956 3756 4964 3764
rect 5148 3756 5156 3764
rect 5404 3756 5412 3764
rect 5468 3756 5476 3764
rect 5564 3756 5572 3764
rect 5580 3756 5588 3764
rect 5660 3756 5668 3764
rect 5724 3756 5732 3764
rect 5740 3756 5748 3764
rect 5996 3756 6004 3764
rect 6028 3756 6036 3764
rect 6124 3756 6132 3764
rect 6252 3756 6260 3764
rect 6412 3756 6420 3764
rect 6876 3756 6884 3764
rect 7196 3756 7204 3764
rect 7260 3756 7268 3764
rect 4268 3732 4276 3740
rect 4284 3736 4292 3744
rect 4380 3736 4388 3744
rect 4444 3736 4452 3744
rect 4476 3736 4484 3744
rect 4556 3736 4564 3744
rect 4620 3736 4628 3744
rect 4732 3736 4740 3744
rect 4796 3736 4804 3744
rect 4844 3736 4852 3744
rect 4972 3736 4980 3744
rect 5036 3736 5044 3744
rect 5068 3736 5076 3744
rect 5100 3736 5108 3744
rect 5164 3736 5172 3744
rect 5260 3736 5268 3744
rect 5388 3736 5396 3744
rect 5644 3736 5652 3744
rect 5772 3736 5780 3744
rect 5868 3736 5876 3744
rect 5884 3736 5892 3744
rect 5980 3736 5988 3744
rect 6076 3736 6084 3744
rect 6156 3736 6164 3744
rect 6188 3736 6196 3744
rect 6300 3736 6308 3744
rect 6556 3736 6564 3744
rect 6636 3736 6644 3744
rect 6668 3736 6676 3744
rect 6748 3736 6756 3744
rect 6860 3736 6868 3744
rect 6988 3736 6996 3744
rect 76 3716 84 3724
rect 124 3716 132 3724
rect 236 3716 244 3724
rect 252 3716 260 3724
rect 300 3716 308 3724
rect 316 3716 324 3724
rect 380 3716 388 3724
rect 428 3716 436 3724
rect 588 3718 596 3726
rect 812 3716 820 3724
rect 876 3716 884 3724
rect 908 3716 916 3724
rect 956 3716 964 3724
rect 988 3716 996 3724
rect 1036 3716 1044 3724
rect 1084 3716 1092 3724
rect 1132 3716 1140 3724
rect 1292 3718 1300 3726
rect 492 3696 500 3704
rect 844 3696 852 3704
rect 1068 3696 1076 3704
rect 1468 3716 1476 3724
rect 1612 3716 1620 3724
rect 1724 3716 1732 3724
rect 1740 3716 1748 3724
rect 1788 3716 1796 3724
rect 1196 3696 1204 3704
rect 1436 3696 1444 3704
rect 1468 3696 1476 3704
rect 1868 3696 1876 3704
rect 1916 3716 1924 3724
rect 1948 3716 1956 3724
rect 2028 3716 2036 3724
rect 2044 3716 2052 3724
rect 2076 3716 2084 3724
rect 2092 3716 2100 3724
rect 2364 3716 2372 3724
rect 2508 3718 2516 3726
rect 2716 3716 2724 3724
rect 2732 3716 2740 3724
rect 2748 3716 2756 3724
rect 2812 3716 2820 3724
rect 2828 3716 2836 3724
rect 2908 3716 2916 3724
rect 2924 3716 2932 3724
rect 3004 3718 3012 3726
rect 7212 3736 7220 3744
rect 7276 3736 7284 3744
rect 7372 3736 7380 3744
rect 7420 3736 7428 3744
rect 7436 3736 7444 3744
rect 7564 3736 7572 3744
rect 3164 3716 3172 3724
rect 3244 3716 3252 3724
rect 3260 3716 3268 3724
rect 3308 3716 3316 3724
rect 3372 3716 3380 3724
rect 3388 3716 3396 3724
rect 3500 3716 3508 3724
rect 2412 3696 2420 3704
rect 2844 3696 2852 3704
rect 3196 3696 3204 3704
rect 3532 3696 3540 3704
rect 3580 3716 3588 3724
rect 3676 3716 3684 3724
rect 3724 3716 3732 3724
rect 3900 3716 3908 3724
rect 3980 3716 3988 3724
rect 4140 3716 4148 3724
rect 4172 3716 4180 3724
rect 4332 3716 4340 3724
rect 4492 3716 4500 3724
rect 4508 3716 4516 3724
rect 4844 3716 4852 3724
rect 4892 3716 4900 3724
rect 4940 3716 4948 3724
rect 5084 3716 5092 3724
rect 5132 3716 5140 3724
rect 5212 3716 5220 3724
rect 5452 3716 5460 3724
rect 5516 3716 5524 3724
rect 5612 3716 5620 3724
rect 5628 3716 5636 3724
rect 5692 3716 5700 3724
rect 6028 3716 6036 3724
rect 6060 3716 6068 3724
rect 6204 3716 6212 3724
rect 6220 3716 6228 3724
rect 3580 3696 3588 3704
rect 5132 3696 5140 3704
rect 6108 3696 6116 3704
rect 6156 3696 6164 3704
rect 6188 3696 6196 3704
rect 6332 3716 6340 3724
rect 6444 3716 6452 3724
rect 6476 3716 6484 3724
rect 6508 3716 6516 3724
rect 6572 3716 6580 3724
rect 6604 3716 6612 3724
rect 6684 3716 6692 3724
rect 6700 3716 6708 3724
rect 6732 3716 6740 3724
rect 6764 3716 6772 3724
rect 6924 3716 6932 3724
rect 6972 3716 6980 3724
rect 7004 3716 7012 3724
rect 7036 3716 7044 3724
rect 7164 3716 7172 3724
rect 7212 3716 7220 3724
rect 7452 3716 7460 3724
rect 7500 3716 7508 3724
rect 6268 3696 6276 3704
rect 6364 3696 6372 3704
rect 6492 3696 6500 3704
rect 6604 3696 6612 3704
rect 7388 3696 7396 3704
rect 1836 3676 1844 3684
rect 3100 3676 3108 3684
rect 3244 3676 3252 3684
rect 3644 3676 3652 3684
rect 4668 3676 4676 3684
rect 4860 3676 4868 3684
rect 6076 3676 6084 3684
rect 6524 3676 6532 3684
rect 956 3636 964 3644
rect 1500 3636 1508 3644
rect 1772 3636 1780 3644
rect 2012 3636 2020 3644
rect 2684 3636 2692 3644
rect 2796 3636 2804 3644
rect 3308 3636 3316 3644
rect 3868 3636 3876 3644
rect 4108 3636 4116 3644
rect 4300 3636 4308 3644
rect 4556 3636 4564 3644
rect 4700 3636 4708 3644
rect 4796 3636 4804 3644
rect 4908 3636 4916 3644
rect 5036 3636 5044 3644
rect 5228 3636 5236 3644
rect 5420 3636 5428 3644
rect 5612 3636 5620 3644
rect 5756 3636 5764 3644
rect 5948 3636 5956 3644
rect 6044 3636 6052 3644
rect 6396 3636 6404 3644
rect 6508 3636 6516 3644
rect 6668 3636 6676 3644
rect 6956 3636 6964 3644
rect 7116 3636 7124 3644
rect 7260 3636 7268 3644
rect 7308 3636 7316 3644
rect 7404 3636 7412 3644
rect 7484 3636 7492 3644
rect 739 3606 747 3614
rect 749 3606 757 3614
rect 759 3606 767 3614
rect 769 3606 777 3614
rect 779 3606 787 3614
rect 789 3606 797 3614
rect 3747 3606 3755 3614
rect 3757 3606 3765 3614
rect 3767 3606 3775 3614
rect 3777 3606 3785 3614
rect 3787 3606 3795 3614
rect 3797 3606 3805 3614
rect 6755 3606 6763 3614
rect 6765 3606 6773 3614
rect 6775 3606 6783 3614
rect 6785 3606 6793 3614
rect 6795 3606 6803 3614
rect 6805 3606 6813 3614
rect 124 3576 132 3584
rect 508 3576 516 3584
rect 604 3576 612 3584
rect 684 3576 692 3584
rect 940 3576 948 3584
rect 1436 3576 1444 3584
rect 1660 3576 1668 3584
rect 1820 3576 1828 3584
rect 2700 3576 2708 3584
rect 3148 3576 3156 3584
rect 3884 3576 3892 3584
rect 6476 3576 6484 3584
rect 7516 3576 7524 3584
rect 796 3556 804 3564
rect 6012 3556 6020 3564
rect 6316 3556 6324 3564
rect 332 3536 340 3544
rect 1116 3536 1124 3544
rect 1468 3536 1476 3544
rect 1628 3536 1636 3544
rect 2364 3536 2372 3544
rect 2668 3536 2676 3544
rect 3564 3536 3572 3544
rect 4444 3536 4452 3544
rect 6316 3536 6324 3544
rect 6332 3536 6340 3544
rect 6892 3536 6900 3544
rect 860 3516 868 3524
rect 988 3516 996 3524
rect 1052 3516 1060 3524
rect 1340 3516 1348 3524
rect 220 3496 228 3504
rect 348 3496 356 3504
rect 412 3496 420 3504
rect 444 3496 452 3504
rect 476 3496 484 3504
rect 524 3496 532 3504
rect 620 3496 628 3504
rect 636 3496 644 3504
rect 652 3496 660 3504
rect 700 3496 708 3504
rect 828 3496 836 3504
rect 860 3496 868 3504
rect 892 3496 900 3504
rect 908 3496 916 3504
rect 956 3496 964 3504
rect 1036 3496 1044 3504
rect 1084 3496 1092 3504
rect 1180 3496 1188 3504
rect 1724 3516 1732 3524
rect 1868 3516 1876 3524
rect 2092 3516 2100 3524
rect 1244 3494 1252 3502
rect 1388 3496 1396 3504
rect 1436 3496 1444 3504
rect 1548 3496 1556 3504
rect 1676 3496 1684 3504
rect 1692 3496 1700 3504
rect 1740 3496 1748 3504
rect 1836 3496 1844 3504
rect 1852 3496 1860 3504
rect 1900 3496 1908 3504
rect 1948 3496 1956 3504
rect 1980 3496 1988 3504
rect 2028 3496 2036 3504
rect 2076 3496 2084 3504
rect 2124 3496 2132 3504
rect 2156 3496 2164 3504
rect 2220 3496 2228 3504
rect 2332 3496 2340 3504
rect 2396 3496 2404 3504
rect 2444 3516 2452 3524
rect 2860 3516 2868 3524
rect 3100 3516 3108 3524
rect 3212 3516 3220 3524
rect 2540 3494 2548 3502
rect 2748 3496 2756 3504
rect 2844 3496 2852 3504
rect 2892 3496 2900 3504
rect 2956 3496 2964 3504
rect 2988 3496 2996 3504
rect 3020 3496 3028 3504
rect 3068 3496 3076 3504
rect 3116 3496 3124 3504
rect 3212 3496 3220 3504
rect 3244 3496 3252 3504
rect 3292 3496 3300 3504
rect 3340 3516 3348 3524
rect 3628 3516 3636 3524
rect 4236 3516 4244 3524
rect 4332 3516 4340 3524
rect 4380 3516 4388 3524
rect 4572 3516 4580 3524
rect 4860 3516 4868 3524
rect 4892 3516 4900 3524
rect 5436 3516 5444 3524
rect 5756 3516 5764 3524
rect 5948 3516 5956 3524
rect 6156 3516 6164 3524
rect 6204 3516 6212 3524
rect 3436 3494 3444 3502
rect 3580 3496 3588 3504
rect 3692 3494 3700 3502
rect 3900 3496 3908 3504
rect 3932 3496 3940 3504
rect 3964 3496 3972 3504
rect 4012 3496 4020 3504
rect 4060 3496 4068 3504
rect 4140 3496 4148 3504
rect 4204 3496 4212 3504
rect 4252 3496 4260 3504
rect 4316 3496 4324 3504
rect 4428 3496 4436 3504
rect 4492 3496 4500 3504
rect 4604 3496 4612 3504
rect 4684 3496 4692 3504
rect 4716 3496 4724 3504
rect 4780 3496 4788 3504
rect 4844 3496 4852 3504
rect 4940 3496 4948 3504
rect 5036 3496 5044 3504
rect 5068 3496 5076 3504
rect 5164 3496 5172 3504
rect 5196 3496 5204 3504
rect 5244 3496 5252 3504
rect 5404 3496 5412 3504
rect 5516 3496 5524 3504
rect 5548 3496 5556 3504
rect 5772 3496 5780 3504
rect 5980 3496 5988 3504
rect 6124 3496 6132 3504
rect 6300 3516 6308 3524
rect 6364 3516 6372 3524
rect 6316 3496 6324 3504
rect 6364 3496 6372 3504
rect 6396 3496 6404 3504
rect 6460 3496 6468 3504
rect 6524 3516 6532 3524
rect 6844 3516 6852 3524
rect 6860 3516 6868 3524
rect 6956 3516 6964 3524
rect 7068 3516 7076 3524
rect 7100 3516 7108 3524
rect 7308 3516 7316 3524
rect 7452 3516 7460 3524
rect 7484 3516 7492 3524
rect 6620 3496 6628 3504
rect 6652 3496 6660 3504
rect 6732 3496 6740 3504
rect 6940 3496 6948 3504
rect 7004 3496 7012 3504
rect 7020 3496 7028 3504
rect 7084 3496 7092 3504
rect 7132 3496 7140 3504
rect 7212 3496 7220 3504
rect 7228 3496 7236 3504
rect 7292 3496 7300 3504
rect 7356 3496 7364 3504
rect 7420 3496 7428 3504
rect 7436 3496 7444 3504
rect 12 3476 20 3484
rect 172 3476 180 3484
rect 364 3476 372 3484
rect 812 3476 820 3484
rect 876 3476 884 3484
rect 1036 3476 1044 3484
rect 1276 3476 1284 3484
rect 1308 3476 1316 3484
rect 1404 3476 1412 3484
rect 1420 3476 1428 3484
rect 1500 3476 1508 3484
rect 1644 3476 1652 3484
rect 1916 3476 1924 3484
rect 1932 3476 1940 3484
rect 1964 3476 1972 3484
rect 1996 3476 2004 3484
rect 2012 3476 2020 3484
rect 2044 3476 2052 3484
rect 2140 3476 2148 3484
rect 2172 3476 2180 3484
rect 2380 3476 2388 3484
rect 2444 3476 2452 3484
rect 2476 3476 2484 3484
rect 2508 3476 2516 3484
rect 2684 3476 2692 3484
rect 2732 3476 2740 3484
rect 2796 3476 2804 3484
rect 2860 3476 2868 3484
rect 2908 3476 2916 3484
rect 2956 3476 2964 3484
rect 2972 3476 2980 3484
rect 3004 3476 3012 3484
rect 3036 3476 3044 3484
rect 3052 3476 3060 3484
rect 3084 3476 3092 3484
rect 3164 3476 3172 3484
rect 3260 3476 3268 3484
rect 3276 3476 3284 3484
rect 3324 3476 3332 3484
rect 3372 3476 3380 3484
rect 3404 3476 3412 3484
rect 3580 3476 3588 3484
rect 3660 3476 3668 3484
rect 3756 3476 3764 3484
rect 3948 3476 3956 3484
rect 444 3456 452 3464
rect 988 3456 996 3464
rect 1356 3456 1364 3464
rect 2252 3456 2260 3464
rect 2748 3456 2756 3464
rect 2812 3456 2820 3464
rect 2924 3456 2932 3464
rect 3628 3456 3636 3464
rect 4044 3456 4052 3464
rect 4092 3456 4100 3464
rect 4268 3476 4276 3484
rect 4300 3476 4308 3484
rect 4364 3476 4372 3484
rect 4412 3476 4420 3484
rect 4444 3476 4452 3484
rect 4476 3476 4484 3484
rect 4524 3476 4532 3484
rect 4540 3476 4548 3484
rect 4588 3476 4596 3484
rect 4652 3476 4660 3484
rect 4668 3476 4676 3484
rect 4700 3476 4708 3484
rect 4796 3476 4804 3484
rect 4828 3476 4836 3484
rect 4892 3476 4900 3484
rect 5052 3476 5060 3484
rect 5116 3476 5124 3484
rect 5148 3476 5156 3484
rect 5196 3476 5204 3484
rect 5228 3476 5236 3484
rect 5500 3476 5508 3484
rect 5532 3476 5540 3484
rect 5612 3476 5620 3484
rect 5708 3476 5716 3484
rect 5724 3476 5732 3484
rect 5788 3476 5796 3484
rect 5932 3476 5940 3484
rect 5980 3476 5988 3484
rect 6028 3476 6036 3484
rect 6108 3476 6116 3484
rect 6156 3476 6164 3484
rect 6172 3476 6180 3484
rect 6252 3476 6260 3484
rect 6412 3476 6420 3484
rect 6556 3476 6564 3484
rect 6684 3476 6692 3484
rect 6716 3476 6724 3484
rect 6828 3476 6836 3484
rect 6844 3476 6852 3484
rect 6892 3476 6900 3484
rect 6956 3476 6964 3484
rect 7036 3476 7044 3484
rect 7068 3476 7076 3484
rect 7132 3476 7140 3484
rect 7164 3476 7172 3484
rect 380 3436 388 3444
rect 684 3436 692 3444
rect 1052 3436 1060 3444
rect 1868 3436 1876 3444
rect 2188 3436 2196 3444
rect 3212 3436 3220 3444
rect 3980 3436 3988 3444
rect 4124 3436 4132 3444
rect 4252 3456 4260 3464
rect 4284 3456 4292 3464
rect 4428 3456 4436 3464
rect 4508 3456 4516 3464
rect 4764 3456 4772 3464
rect 4828 3456 4836 3464
rect 4844 3456 4852 3464
rect 4988 3456 4996 3464
rect 5004 3456 5012 3464
rect 5036 3456 5044 3464
rect 5196 3456 5204 3464
rect 5228 3456 5236 3464
rect 5340 3456 5348 3464
rect 5356 3456 5364 3464
rect 5484 3456 5492 3464
rect 5596 3456 5604 3464
rect 5820 3456 5828 3464
rect 5996 3456 6004 3464
rect 6028 3456 6036 3464
rect 6076 3456 6084 3464
rect 6268 3456 6276 3464
rect 6428 3456 6436 3464
rect 6572 3456 6580 3464
rect 6652 3456 6660 3464
rect 6924 3456 6932 3464
rect 6940 3456 6948 3464
rect 7084 3456 7092 3464
rect 7244 3476 7252 3484
rect 7292 3476 7300 3484
rect 7372 3476 7380 3484
rect 7404 3476 7412 3484
rect 7436 3476 7444 3484
rect 7308 3456 7316 3464
rect 7372 3456 7380 3464
rect 7500 3456 7508 3464
rect 4236 3436 4244 3444
rect 4316 3436 4324 3444
rect 4332 3436 4340 3444
rect 4396 3436 4404 3444
rect 4492 3436 4500 3444
rect 4572 3436 4580 3444
rect 4604 3436 4612 3444
rect 4780 3436 4788 3444
rect 4860 3436 4868 3444
rect 4908 3436 4916 3444
rect 5468 3436 5476 3444
rect 5644 3436 5652 3444
rect 5756 3436 5764 3444
rect 5868 3436 5876 3444
rect 6220 3436 6228 3444
rect 6524 3436 6532 3444
rect 6588 3436 6596 3444
rect 6684 3436 6692 3444
rect 7004 3436 7012 3444
rect 7020 3436 7028 3444
rect 7100 3436 7108 3444
rect 7164 3436 7172 3444
rect 7260 3436 7268 3444
rect 7292 3436 7300 3444
rect 7388 3436 7396 3444
rect 4764 3416 4772 3424
rect 4988 3416 4996 3424
rect 5356 3416 5364 3424
rect 5596 3416 5604 3424
rect 2243 3406 2251 3414
rect 2253 3406 2261 3414
rect 2263 3406 2271 3414
rect 2273 3406 2281 3414
rect 2283 3406 2291 3414
rect 2293 3406 2301 3414
rect 5251 3406 5259 3414
rect 5261 3406 5269 3414
rect 5271 3406 5279 3414
rect 5281 3406 5289 3414
rect 5291 3406 5299 3414
rect 5301 3406 5309 3414
rect 4140 3396 4148 3404
rect 4364 3396 4372 3404
rect 4636 3396 4644 3404
rect 124 3376 132 3384
rect 220 3376 228 3384
rect 444 3376 452 3384
rect 460 3376 468 3384
rect 684 3376 692 3384
rect 748 3376 756 3384
rect 972 3376 980 3384
rect 1436 3376 1444 3384
rect 1708 3376 1716 3384
rect 1756 3376 1764 3384
rect 2060 3376 2068 3384
rect 2348 3376 2356 3384
rect 2684 3376 2692 3384
rect 2732 3376 2740 3384
rect 3916 3376 3924 3384
rect 3964 3376 3972 3384
rect 4508 3376 4516 3384
rect 4540 3376 4548 3384
rect 4956 3376 4964 3384
rect 5052 3376 5060 3384
rect 5084 3376 5092 3384
rect 5180 3376 5188 3384
rect 5212 3376 5220 3384
rect 5580 3376 5588 3384
rect 5612 3376 5620 3384
rect 6380 3376 6388 3384
rect 6540 3376 6548 3384
rect 6716 3376 6724 3384
rect 6988 3376 6996 3384
rect 7212 3376 7220 3384
rect 7292 3376 7300 3384
rect 7388 3376 7396 3384
rect 7452 3376 7460 3384
rect 188 3356 196 3364
rect 12 3336 20 3344
rect 316 3356 324 3364
rect 556 3356 564 3364
rect 1644 3356 1652 3364
rect 1948 3356 1956 3364
rect 2924 3356 2932 3364
rect 3132 3356 3140 3364
rect 3324 3356 3332 3364
rect 3484 3356 3492 3364
rect 4108 3356 4116 3364
rect 4140 3356 4148 3364
rect 4172 3356 4180 3364
rect 4236 3356 4244 3364
rect 4348 3356 4356 3364
rect 4364 3356 4372 3364
rect 4460 3356 4468 3364
rect 4492 3356 4500 3364
rect 4572 3356 4580 3364
rect 236 3336 244 3344
rect 284 3336 292 3344
rect 524 3336 532 3344
rect 956 3336 964 3344
rect 1020 3336 1028 3344
rect 1036 3336 1044 3344
rect 1068 3336 1076 3344
rect 1132 3336 1140 3344
rect 156 3316 164 3324
rect 252 3316 260 3324
rect 364 3316 372 3324
rect 492 3316 500 3324
rect 572 3316 580 3324
rect 700 3316 708 3324
rect 716 3316 724 3324
rect 764 3316 772 3324
rect 844 3316 852 3324
rect 876 3316 884 3324
rect 940 3316 948 3324
rect 972 3316 980 3324
rect 1036 3316 1044 3324
rect 1068 3316 1076 3324
rect 1116 3316 1124 3324
rect 1132 3316 1140 3324
rect 1196 3336 1204 3344
rect 1244 3336 1252 3344
rect 1276 3336 1284 3344
rect 1724 3336 1732 3344
rect 1916 3336 1924 3344
rect 2028 3336 2036 3344
rect 2220 3336 2228 3344
rect 2364 3336 2372 3344
rect 2492 3336 2500 3344
rect 2748 3336 2756 3344
rect 2828 3336 2836 3344
rect 3148 3336 3156 3344
rect 3212 3336 3220 3344
rect 3372 3336 3380 3344
rect 3500 3336 3508 3344
rect 3612 3336 3620 3344
rect 3644 3336 3652 3344
rect 3756 3336 3764 3344
rect 3948 3336 3956 3344
rect 4044 3336 4052 3344
rect 4060 3336 4068 3344
rect 4492 3336 4500 3344
rect 4556 3336 4564 3344
rect 4636 3356 4644 3364
rect 4780 3356 4788 3364
rect 4892 3356 4900 3364
rect 4940 3356 4948 3364
rect 5020 3356 5028 3364
rect 5148 3356 5156 3364
rect 5276 3356 5284 3364
rect 5388 3356 5396 3364
rect 5404 3356 5412 3364
rect 5564 3356 5572 3364
rect 4636 3336 4644 3344
rect 4732 3336 4740 3344
rect 4956 3336 4964 3344
rect 5004 3336 5012 3344
rect 5036 3336 5044 3344
rect 5084 3336 5092 3344
rect 5132 3336 5140 3344
rect 5164 3336 5172 3344
rect 5292 3336 5300 3344
rect 5372 3336 5380 3344
rect 5404 3336 5412 3344
rect 5580 3336 5588 3344
rect 5628 3336 5636 3344
rect 5708 3336 5716 3344
rect 5820 3356 5828 3364
rect 6492 3356 6500 3364
rect 6508 3356 6516 3364
rect 6652 3356 6660 3364
rect 6924 3356 6932 3364
rect 6940 3356 6948 3364
rect 7068 3356 7076 3364
rect 7116 3356 7124 3364
rect 7180 3356 7188 3364
rect 7468 3356 7476 3364
rect 7484 3356 7492 3364
rect 5788 3336 5796 3344
rect 5948 3332 5956 3340
rect 5964 3336 5972 3344
rect 6076 3336 6084 3344
rect 6156 3336 6164 3344
rect 6252 3336 6260 3344
rect 6268 3336 6276 3344
rect 1164 3316 1172 3324
rect 1308 3318 1316 3326
rect 908 3296 916 3304
rect 1052 3296 1060 3304
rect 1084 3296 1092 3304
rect 1452 3316 1460 3324
rect 1468 3316 1476 3324
rect 1532 3316 1540 3324
rect 1612 3316 1620 3324
rect 1628 3316 1636 3324
rect 1676 3316 1684 3324
rect 1740 3316 1748 3324
rect 1884 3318 1892 3326
rect 1980 3316 1988 3324
rect 2044 3316 2052 3324
rect 2188 3318 2196 3326
rect 2316 3316 2324 3324
rect 2508 3316 2516 3324
rect 2572 3316 2580 3324
rect 2620 3316 2628 3324
rect 2636 3316 2644 3324
rect 2652 3316 2660 3324
rect 2700 3316 2708 3324
rect 2764 3316 2772 3324
rect 2796 3316 2804 3324
rect 2860 3318 2868 3326
rect 2908 3316 2916 3324
rect 3004 3316 3012 3324
rect 3020 3316 3028 3324
rect 3068 3316 3076 3324
rect 3100 3316 3108 3324
rect 3196 3316 3204 3324
rect 3228 3316 3236 3324
rect 3244 3316 3252 3324
rect 3308 3316 3316 3324
rect 3356 3316 3364 3324
rect 3388 3316 3396 3324
rect 3420 3316 3428 3324
rect 3484 3316 3492 3324
rect 3516 3316 3524 3324
rect 3532 3316 3540 3324
rect 3596 3316 3604 3324
rect 3628 3316 3636 3324
rect 3788 3318 3796 3326
rect 3852 3316 3860 3324
rect 3932 3316 3940 3324
rect 4060 3316 4068 3324
rect 4076 3316 4084 3324
rect 4108 3316 4116 3324
rect 4204 3316 4212 3324
rect 4268 3316 4276 3324
rect 4316 3316 4324 3324
rect 4412 3316 4420 3324
rect 4508 3316 4516 3324
rect 4572 3316 4580 3324
rect 4588 3316 4596 3324
rect 4604 3316 4612 3324
rect 4684 3316 4692 3324
rect 4716 3316 4724 3324
rect 4732 3316 4740 3324
rect 4780 3316 4788 3324
rect 4812 3316 4820 3324
rect 4860 3316 4868 3324
rect 4908 3316 4916 3324
rect 4924 3316 4932 3324
rect 4956 3316 4964 3324
rect 5020 3316 5028 3324
rect 5084 3316 5092 3324
rect 5148 3316 5156 3324
rect 5244 3316 5252 3324
rect 5388 3316 5396 3324
rect 5452 3316 5460 3324
rect 5484 3316 5492 3324
rect 5532 3316 5540 3324
rect 5580 3316 5588 3324
rect 5644 3316 5652 3324
rect 5660 3316 5668 3324
rect 5692 3316 5700 3324
rect 5724 3316 5732 3324
rect 5740 3316 5748 3324
rect 5804 3316 5812 3324
rect 5852 3316 5860 3324
rect 6076 3316 6084 3324
rect 6124 3316 6132 3324
rect 6156 3316 6164 3324
rect 6476 3336 6484 3344
rect 6572 3336 6580 3344
rect 6700 3336 6708 3344
rect 6732 3336 6740 3344
rect 6908 3336 6916 3344
rect 6940 3336 6948 3344
rect 6988 3336 6996 3344
rect 7052 3336 7060 3344
rect 7132 3336 7140 3344
rect 7148 3336 7156 3344
rect 7212 3336 7220 3344
rect 7260 3336 7268 3344
rect 7340 3336 7348 3344
rect 7436 3336 7444 3344
rect 7468 3336 7476 3344
rect 7516 3336 7524 3344
rect 6412 3316 6420 3324
rect 6604 3316 6612 3324
rect 6748 3316 6756 3324
rect 6828 3316 6836 3324
rect 6924 3316 6932 3324
rect 6988 3316 6996 3324
rect 7068 3316 7076 3324
rect 7084 3316 7092 3324
rect 7212 3316 7220 3324
rect 7244 3316 7252 3324
rect 7276 3316 7284 3324
rect 7324 3316 7332 3324
rect 7388 3316 7396 3324
rect 7420 3316 7428 3324
rect 7532 3316 7540 3324
rect 1212 3296 1220 3304
rect 2796 3296 2804 3304
rect 3196 3296 3204 3304
rect 3420 3296 3428 3304
rect 3660 3296 3668 3304
rect 3996 3296 4004 3304
rect 4220 3296 4228 3304
rect 4252 3296 4260 3304
rect 4444 3296 4452 3304
rect 4796 3296 4804 3304
rect 5004 3296 5012 3304
rect 5068 3296 5076 3304
rect 5132 3296 5140 3304
rect 5196 3296 5204 3304
rect 5340 3296 5348 3304
rect 5468 3296 5476 3304
rect 5548 3296 5556 3304
rect 6140 3296 6148 3304
rect 6524 3296 6532 3304
rect 6540 3296 6548 3304
rect 6588 3296 6596 3304
rect 6876 3296 6884 3304
rect 7052 3296 7060 3304
rect 7164 3296 7172 3304
rect 7404 3296 7412 3304
rect 412 3276 420 3284
rect 1788 3276 1796 3284
rect 2604 3276 2612 3284
rect 3356 3276 3364 3284
rect 4172 3276 4180 3284
rect 4284 3276 4292 3284
rect 4828 3276 4836 3284
rect 4860 3276 4868 3284
rect 5500 3276 5508 3284
rect 6108 3276 6116 3284
rect 6300 3276 6308 3284
rect 6620 3276 6628 3284
rect 7372 3276 7380 3284
rect 4812 3256 4820 3264
rect 5788 3256 5796 3264
rect 7084 3256 7092 3264
rect 1484 3236 1492 3244
rect 1580 3236 1588 3244
rect 1996 3236 2004 3244
rect 2476 3236 2484 3244
rect 2540 3236 2548 3244
rect 2988 3236 2996 3244
rect 3036 3236 3044 3244
rect 3276 3236 3284 3244
rect 3548 3236 3556 3244
rect 4268 3236 4276 3244
rect 4332 3236 4340 3244
rect 4716 3236 4724 3244
rect 5484 3236 5492 3244
rect 5884 3236 5892 3244
rect 6124 3236 6132 3244
rect 6636 3236 6644 3244
rect 6764 3236 6772 3244
rect 7196 3236 7204 3244
rect 739 3206 747 3214
rect 749 3206 757 3214
rect 759 3206 767 3214
rect 769 3206 777 3214
rect 779 3206 787 3214
rect 789 3206 797 3214
rect 3747 3206 3755 3214
rect 3757 3206 3765 3214
rect 3767 3206 3775 3214
rect 3777 3206 3785 3214
rect 3787 3206 3795 3214
rect 3797 3206 3805 3214
rect 6755 3206 6763 3214
rect 6765 3206 6773 3214
rect 6775 3206 6783 3214
rect 6785 3206 6793 3214
rect 6795 3206 6803 3214
rect 6805 3206 6813 3214
rect 124 3176 132 3184
rect 892 3176 900 3184
rect 956 3176 964 3184
rect 1356 3176 1364 3184
rect 1628 3176 1636 3184
rect 2012 3176 2020 3184
rect 2108 3176 2116 3184
rect 2732 3176 2740 3184
rect 4060 3176 4068 3184
rect 4876 3176 4884 3184
rect 4988 3176 4996 3184
rect 6060 3176 6068 3184
rect 7500 3176 7508 3184
rect 2204 3156 2212 3164
rect 3420 3156 3428 3164
rect 4316 3156 4324 3164
rect 6364 3156 6372 3164
rect 7276 3156 7284 3164
rect 636 3136 644 3144
rect 1196 3136 1204 3144
rect 1596 3136 1604 3144
rect 3036 3136 3044 3144
rect 3068 3136 3076 3144
rect 3100 3136 3108 3144
rect 4268 3136 4276 3144
rect 4332 3136 4340 3144
rect 4524 3136 4532 3144
rect 6428 3136 6436 3144
rect 6972 3136 6980 3144
rect 572 3116 580 3124
rect 604 3116 612 3124
rect 668 3116 676 3124
rect 1244 3116 1252 3124
rect 44 3096 52 3104
rect 108 3096 116 3104
rect 156 3096 164 3104
rect 236 3096 244 3104
rect 284 3096 292 3104
rect 428 3096 436 3104
rect 572 3096 580 3104
rect 636 3096 644 3104
rect 684 3096 692 3104
rect 844 3096 852 3104
rect 860 3096 868 3104
rect 908 3096 916 3104
rect 1004 3096 1012 3104
rect 2572 3116 2580 3124
rect 2764 3116 2772 3124
rect 2828 3116 2836 3124
rect 1068 3094 1076 3102
rect 1292 3096 1300 3104
rect 1324 3096 1332 3104
rect 1468 3096 1476 3104
rect 1564 3096 1572 3104
rect 1660 3096 1668 3104
rect 1772 3096 1780 3104
rect 1900 3096 1908 3104
rect 1932 3096 1940 3104
rect 1996 3096 2004 3104
rect 2044 3096 2052 3104
rect 2060 3096 2068 3104
rect 2124 3096 2132 3104
rect 2140 3096 2148 3104
rect 2156 3096 2164 3104
rect 2252 3096 2260 3104
rect 2380 3094 2388 3102
rect 2444 3096 2452 3104
rect 2540 3096 2548 3104
rect 2588 3096 2596 3104
rect 2636 3096 2644 3104
rect 2668 3096 2676 3104
rect 2732 3096 2740 3104
rect 2796 3096 2804 3104
rect 2876 3096 2884 3104
rect 2956 3096 2964 3104
rect 3100 3096 3108 3104
rect 3148 3116 3156 3124
rect 3260 3116 3268 3124
rect 3324 3116 3332 3124
rect 3996 3116 4004 3124
rect 4300 3116 4308 3124
rect 4412 3116 4420 3124
rect 4588 3116 4596 3124
rect 4748 3116 4756 3124
rect 4780 3116 4788 3124
rect 4796 3116 4804 3124
rect 3180 3096 3188 3104
rect 3244 3096 3252 3104
rect 3276 3096 3284 3104
rect 3356 3096 3364 3104
rect 3388 3096 3396 3104
rect 3452 3096 3460 3104
rect 3468 3096 3476 3104
rect 3500 3096 3508 3104
rect 3548 3096 3556 3104
rect 3564 3096 3572 3104
rect 3580 3096 3588 3104
rect 3708 3096 3716 3104
rect 3836 3096 3844 3104
rect 3932 3096 3940 3104
rect 4044 3096 4052 3104
rect 4092 3096 4100 3104
rect 4188 3096 4196 3104
rect 4220 3096 4228 3104
rect 4252 3096 4260 3104
rect 4316 3096 4324 3104
rect 4364 3096 4372 3104
rect 4396 3096 4404 3104
rect 4444 3096 4452 3104
rect 4476 3096 4484 3104
rect 4540 3096 4548 3104
rect 4604 3096 4612 3104
rect 4652 3096 4660 3104
rect 4748 3096 4756 3104
rect 4876 3096 4884 3104
rect 4988 3096 4996 3104
rect 5036 3116 5044 3124
rect 5196 3116 5204 3124
rect 5212 3116 5220 3124
rect 5372 3116 5380 3124
rect 5500 3116 5508 3124
rect 5084 3096 5092 3104
rect 5148 3096 5156 3104
rect 5420 3096 5428 3104
rect 5500 3096 5508 3104
rect 5644 3116 5652 3124
rect 5548 3096 5556 3104
rect 5692 3096 5700 3104
rect 5772 3096 5780 3104
rect 5820 3116 5828 3124
rect 5868 3116 5876 3124
rect 5964 3116 5972 3124
rect 6220 3116 6228 3124
rect 6268 3116 6276 3124
rect 6396 3116 6404 3124
rect 6460 3116 6468 3124
rect 6908 3116 6916 3124
rect 7084 3116 7092 3124
rect 7388 3116 7396 3124
rect 7484 3116 7492 3124
rect 5900 3096 5908 3104
rect 6012 3096 6020 3104
rect 6092 3096 6100 3104
rect 6124 3096 6132 3104
rect 6316 3096 6324 3104
rect 6380 3096 6388 3104
rect 6428 3096 6436 3104
rect 6572 3096 6580 3104
rect 6636 3096 6644 3104
rect 6652 3096 6660 3104
rect 6732 3096 6740 3104
rect 6860 3096 6868 3104
rect 6956 3096 6964 3104
rect 7020 3096 7028 3104
rect 7052 3096 7060 3104
rect 7132 3096 7140 3104
rect 7180 3096 7188 3104
rect 7436 3096 7444 3104
rect 92 3076 100 3084
rect 412 3076 420 3084
rect 556 3076 564 3084
rect 620 3076 628 3084
rect 700 3076 708 3084
rect 12 3056 20 3064
rect 748 3056 756 3064
rect 940 3056 948 3064
rect 988 3076 996 3084
rect 1100 3076 1108 3084
rect 1212 3076 1220 3084
rect 1308 3076 1316 3084
rect 1388 3076 1396 3084
rect 1644 3076 1652 3084
rect 1756 3056 1764 3064
rect 1948 3076 1956 3084
rect 1980 3076 1988 3084
rect 1948 3056 1956 3064
rect 2188 3056 2196 3064
rect 2236 3076 2244 3084
rect 2396 3076 2404 3084
rect 2652 3076 2660 3084
rect 2716 3076 2724 3084
rect 2780 3076 2788 3084
rect 2908 3076 2916 3084
rect 3084 3076 3092 3084
rect 3196 3076 3204 3084
rect 3372 3076 3380 3084
rect 3484 3076 3492 3084
rect 3852 3076 3860 3084
rect 3932 3076 3940 3084
rect 3948 3076 3956 3084
rect 3980 3076 3988 3084
rect 4044 3076 4052 3084
rect 4204 3076 4212 3084
rect 4236 3076 4244 3084
rect 4364 3076 4372 3084
rect 4460 3076 4468 3084
rect 4492 3076 4500 3084
rect 4524 3076 4532 3084
rect 4556 3076 4564 3084
rect 4828 3076 4836 3084
rect 5068 3076 5076 3084
rect 5100 3076 5108 3084
rect 5132 3076 5140 3084
rect 5164 3076 5172 3084
rect 5244 3076 5252 3084
rect 5468 3076 5476 3084
rect 5516 3076 5524 3084
rect 5612 3076 5620 3084
rect 5660 3076 5668 3084
rect 5756 3076 5764 3084
rect 5788 3076 5796 3084
rect 5852 3076 5860 3084
rect 5996 3076 6004 3084
rect 6012 3076 6020 3084
rect 6076 3076 6084 3084
rect 6124 3076 6132 3084
rect 6252 3076 6260 3084
rect 6300 3076 6308 3084
rect 6316 3076 6324 3084
rect 6364 3076 6372 3084
rect 6444 3076 6452 3084
rect 6540 3076 6548 3084
rect 6556 3076 6564 3084
rect 6620 3076 6628 3084
rect 2844 3056 2852 3064
rect 2876 3056 2884 3064
rect 3308 3056 3316 3064
rect 3612 3056 3620 3064
rect 3628 3056 3636 3064
rect 3692 3056 3700 3064
rect 4108 3056 4116 3064
rect 4140 3056 4148 3064
rect 4284 3056 4292 3064
rect 4396 3056 4404 3064
rect 4540 3056 4548 3064
rect 4604 3056 4612 3064
rect 4636 3056 4644 3064
rect 4652 3056 4660 3064
rect 4684 3056 4692 3064
rect 4700 3056 4708 3064
rect 4924 3056 4932 3064
rect 4940 3056 4948 3064
rect 5132 3056 5140 3064
rect 5260 3056 5268 3064
rect 5356 3056 5364 3064
rect 5452 3056 5460 3064
rect 5580 3056 5588 3064
rect 5740 3056 5748 3064
rect 5948 3056 5956 3064
rect 6108 3056 6116 3064
rect 6556 3056 6564 3064
rect 6716 3076 6724 3084
rect 6796 3076 6804 3084
rect 6892 3076 6900 3084
rect 6940 3076 6948 3084
rect 6972 3076 6980 3084
rect 7020 3076 7028 3084
rect 7036 3076 7044 3084
rect 7100 3076 7108 3084
rect 7132 3076 7140 3084
rect 7164 3076 7172 3084
rect 7244 3076 7252 3084
rect 7340 3076 7348 3084
rect 7356 3076 7364 3084
rect 7516 3076 7524 3084
rect 6956 3056 6964 3064
rect 7164 3056 7172 3064
rect 7228 3056 7236 3064
rect 7404 3056 7412 3064
rect 7420 3056 7428 3064
rect 7468 3056 7476 3064
rect 76 3036 84 3044
rect 348 3036 356 3044
rect 540 3036 548 3044
rect 716 3036 724 3044
rect 892 3036 900 3044
rect 1260 3036 1268 3044
rect 1356 3036 1364 3044
rect 1548 3036 1556 3044
rect 1692 3036 1700 3044
rect 1884 3036 1892 3044
rect 1964 3036 1972 3044
rect 2508 3036 2516 3044
rect 2636 3036 2644 3044
rect 2828 3036 2836 3044
rect 3292 3036 3300 3044
rect 3324 3036 3332 3044
rect 3596 3036 3604 3044
rect 3740 3036 3748 3044
rect 4124 3036 4132 3044
rect 4476 3036 4484 3044
rect 4588 3036 4596 3044
rect 4828 3036 4836 3044
rect 5068 3036 5076 3044
rect 5148 3036 5156 3044
rect 5196 3036 5204 3044
rect 5372 3036 5380 3044
rect 5468 3036 5476 3044
rect 5484 3036 5492 3044
rect 5612 3036 5620 3044
rect 5852 3036 5860 3044
rect 5868 3036 5876 3044
rect 5964 3036 5972 3044
rect 6012 3036 6020 3044
rect 6124 3036 6132 3044
rect 6204 3036 6212 3044
rect 6268 3036 6276 3044
rect 6316 3036 6324 3044
rect 6460 3036 6468 3044
rect 6604 3036 6612 3044
rect 6684 3036 6692 3044
rect 6828 3036 6836 3044
rect 7020 3036 7028 3044
rect 7084 3036 7092 3044
rect 7212 3036 7220 3044
rect 7372 3036 7380 3044
rect 7500 3036 7508 3044
rect 4140 3016 4148 3024
rect 4700 3016 4708 3024
rect 4924 3016 4932 3024
rect 4940 3016 4948 3024
rect 5452 3016 5460 3024
rect 5580 3016 5588 3024
rect 5740 3016 5748 3024
rect 5948 3016 5956 3024
rect 2243 3006 2251 3014
rect 2253 3006 2261 3014
rect 2263 3006 2271 3014
rect 2273 3006 2281 3014
rect 2283 3006 2291 3014
rect 2293 3006 2301 3014
rect 5251 3006 5259 3014
rect 5261 3006 5269 3014
rect 5271 3006 5279 3014
rect 5281 3006 5289 3014
rect 5291 3006 5299 3014
rect 5301 3006 5309 3014
rect 4332 2996 4340 3004
rect 4364 2996 4372 3004
rect 4668 2996 4676 3004
rect 4892 2996 4900 3004
rect 5036 2996 5044 3004
rect 5468 2996 5476 3004
rect 12 2976 20 2984
rect 236 2976 244 2984
rect 748 2976 756 2984
rect 828 2976 836 2984
rect 1228 2976 1236 2984
rect 1292 2976 1300 2984
rect 1868 2976 1876 2984
rect 2092 2976 2100 2984
rect 2460 2976 2468 2984
rect 2588 2976 2596 2984
rect 2652 2976 2660 2984
rect 2972 2976 2980 2984
rect 3820 2976 3828 2984
rect 4252 2976 4260 2984
rect 4316 2976 4324 2984
rect 4444 2976 4452 2984
rect 4460 2976 4468 2984
rect 4492 2976 4500 2984
rect 4524 2976 4532 2984
rect 4540 2976 4548 2984
rect 4732 2976 4740 2984
rect 4748 2976 4756 2984
rect 4828 2976 4836 2984
rect 5196 2976 5204 2984
rect 5228 2976 5236 2984
rect 5356 2976 5364 2984
rect 5484 2976 5492 2984
rect 5500 2976 5508 2984
rect 300 2956 308 2964
rect 796 2956 804 2964
rect 1004 2956 1012 2964
rect 1036 2956 1044 2964
rect 1500 2956 1508 2964
rect 1740 2956 1748 2964
rect 124 2936 132 2944
rect 220 2936 228 2944
rect 300 2936 308 2944
rect 620 2936 628 2944
rect 668 2936 676 2944
rect 860 2936 868 2944
rect 924 2936 932 2944
rect 940 2936 948 2944
rect 972 2936 980 2944
rect 1068 2936 1076 2944
rect 1340 2936 1348 2944
rect 1420 2936 1428 2944
rect 1468 2936 1476 2944
rect 2156 2956 2164 2964
rect 2604 2956 2612 2964
rect 2668 2956 2676 2964
rect 2892 2956 2900 2964
rect 3324 2956 3332 2964
rect 3740 2956 3748 2964
rect 4332 2956 4340 2964
rect 4364 2956 4372 2964
rect 4476 2956 4484 2964
rect 4668 2956 4676 2964
rect 4876 2956 4884 2964
rect 4892 2956 4900 2964
rect 1788 2936 1796 2944
rect 2076 2936 2084 2944
rect 2572 2936 2580 2944
rect 2716 2936 2724 2944
rect 2844 2936 2852 2944
rect 2956 2936 2964 2944
rect 3228 2936 3236 2944
rect 3260 2936 3268 2944
rect 3276 2936 3284 2944
rect 3340 2936 3348 2944
rect 3548 2936 3556 2944
rect 3676 2936 3684 2944
rect 3708 2936 3716 2944
rect 3932 2936 3940 2944
rect 4204 2936 4212 2944
rect 4268 2936 4276 2944
rect 4332 2936 4340 2944
rect 4524 2936 4532 2944
rect 4540 2936 4548 2944
rect 4748 2936 4756 2944
rect 4780 2936 4788 2944
rect 4828 2936 4836 2944
rect 5036 2956 5044 2964
rect 5260 2956 5268 2964
rect 5036 2936 5044 2944
rect 5100 2936 5108 2944
rect 5212 2936 5220 2944
rect 5244 2936 5252 2944
rect 92 2916 100 2924
rect 204 2916 212 2924
rect 268 2916 276 2924
rect 364 2916 372 2924
rect 380 2916 388 2924
rect 428 2916 436 2924
rect 444 2916 452 2924
rect 476 2916 484 2924
rect 524 2916 532 2924
rect 540 2916 548 2924
rect 636 2916 644 2924
rect 844 2916 852 2924
rect 876 2916 884 2924
rect 924 2916 932 2924
rect 956 2916 964 2924
rect 1036 2916 1044 2924
rect 1116 2916 1124 2924
rect 1164 2916 1172 2924
rect 1244 2916 1252 2924
rect 1308 2916 1316 2924
rect 1324 2916 1332 2924
rect 1356 2916 1364 2924
rect 1404 2916 1412 2924
rect 1468 2916 1476 2924
rect 1500 2916 1508 2924
rect 1532 2916 1540 2924
rect 1580 2916 1588 2924
rect 1676 2916 1684 2924
rect 1692 2916 1700 2924
rect 1708 2916 1716 2924
rect 1772 2916 1780 2924
rect 1804 2916 1812 2924
rect 1820 2916 1828 2924
rect 1932 2916 1940 2924
rect 1948 2916 1956 2924
rect 2060 2916 2068 2924
rect 2124 2916 2132 2924
rect 2172 2916 2180 2924
rect 2348 2916 2356 2924
rect 2396 2916 2404 2924
rect 2476 2916 2484 2924
rect 2492 2916 2500 2924
rect 2540 2916 2548 2924
rect 2556 2916 2564 2924
rect 2620 2916 2628 2924
rect 2700 2916 2708 2924
rect 2732 2916 2740 2924
rect 2764 2916 2772 2924
rect 2844 2916 2852 2924
rect 2860 2916 2868 2924
rect 2924 2916 2932 2924
rect 2940 2916 2948 2924
rect 3036 2916 3044 2924
rect 3068 2916 3076 2924
rect 3164 2916 3172 2924
rect 3244 2916 3252 2924
rect 3292 2916 3300 2924
rect 3324 2916 3332 2924
rect 3356 2916 3364 2924
rect 3372 2916 3380 2924
rect 3420 2916 3428 2924
rect 3468 2916 3476 2924
rect 3516 2916 3524 2924
rect 3532 2916 3540 2924
rect 3564 2916 3572 2924
rect 3612 2916 3620 2924
rect 3660 2916 3668 2924
rect 3692 2916 3700 2924
rect 3804 2916 3812 2924
rect 3916 2916 3924 2924
rect 4060 2918 4068 2926
rect 4220 2916 4228 2924
rect 4252 2916 4260 2924
rect 4284 2916 4292 2924
rect 4412 2916 4420 2924
rect 4524 2916 4532 2924
rect 988 2896 996 2904
rect 1196 2896 1204 2904
rect 1388 2896 1396 2904
rect 2796 2896 2804 2904
rect 2908 2896 2916 2904
rect 3212 2896 3220 2904
rect 3596 2896 3604 2904
rect 3628 2896 3636 2904
rect 4444 2896 4452 2904
rect 4492 2896 4500 2904
rect 4572 2896 4580 2904
rect 2268 2876 2276 2884
rect 2700 2876 2708 2884
rect 4188 2876 4196 2884
rect 4604 2876 4612 2884
rect 4700 2916 4708 2924
rect 4844 2916 4852 2924
rect 4924 2916 4932 2924
rect 4972 2916 4980 2924
rect 5084 2916 5092 2924
rect 5148 2916 5156 2924
rect 5196 2916 5204 2924
rect 5260 2916 5268 2924
rect 5340 2916 5348 2924
rect 5452 2956 5460 2964
rect 5468 2956 5476 2964
rect 5660 2976 5668 2984
rect 5756 2976 5764 2984
rect 6284 2976 6292 2984
rect 6684 2976 6692 2984
rect 6732 2976 6740 2984
rect 6908 2976 6916 2984
rect 6924 2976 6932 2984
rect 7340 2976 7348 2984
rect 5692 2956 5700 2964
rect 5708 2956 5716 2964
rect 5772 2956 5780 2964
rect 5884 2956 5892 2964
rect 5916 2956 5924 2964
rect 5932 2956 5940 2964
rect 6028 2956 6036 2964
rect 6252 2956 6260 2964
rect 6300 2956 6308 2964
rect 6572 2956 6580 2964
rect 6604 2956 6612 2964
rect 6636 2956 6644 2964
rect 6668 2956 6676 2964
rect 6860 2956 6868 2964
rect 7020 2956 7028 2964
rect 7100 2956 7108 2964
rect 5388 2936 5396 2944
rect 5484 2936 5492 2944
rect 5532 2936 5540 2944
rect 5676 2936 5684 2944
rect 5708 2936 5716 2944
rect 5756 2936 5764 2944
rect 5980 2936 5988 2944
rect 6012 2936 6020 2944
rect 6156 2936 6164 2944
rect 6172 2936 6180 2944
rect 6284 2936 6292 2944
rect 6380 2936 6388 2944
rect 6460 2936 6468 2944
rect 6492 2936 6500 2944
rect 6524 2936 6532 2944
rect 6620 2936 6628 2944
rect 6684 2936 6692 2944
rect 6716 2936 6724 2944
rect 6844 2936 6852 2944
rect 7036 2936 7044 2944
rect 7068 2936 7076 2944
rect 7100 2936 7108 2944
rect 7148 2936 7156 2944
rect 7164 2936 7172 2944
rect 7212 2936 7220 2944
rect 7228 2936 7236 2944
rect 7324 2936 7332 2944
rect 5388 2916 5396 2924
rect 5404 2916 5412 2924
rect 5420 2916 5428 2924
rect 5548 2916 5556 2924
rect 5580 2916 5588 2924
rect 5692 2916 5700 2924
rect 5756 2916 5764 2924
rect 5804 2916 5812 2924
rect 5836 2916 5844 2924
rect 5948 2916 5956 2924
rect 5996 2916 6004 2924
rect 6060 2916 6068 2924
rect 6204 2916 6212 2924
rect 6300 2916 6308 2924
rect 6396 2916 6404 2924
rect 6508 2916 6516 2924
rect 6668 2916 6676 2924
rect 6732 2916 6740 2924
rect 6748 2916 6756 2924
rect 6876 2916 6884 2924
rect 6988 2916 6996 2924
rect 7052 2916 7060 2924
rect 7196 2916 7204 2924
rect 7388 2936 7396 2944
rect 7484 2936 7492 2944
rect 4636 2896 4644 2904
rect 4780 2896 4788 2904
rect 4796 2896 4804 2904
rect 4972 2896 4980 2904
rect 5004 2896 5012 2904
rect 5116 2896 5124 2904
rect 5132 2896 5140 2904
rect 5436 2896 5444 2904
rect 5516 2896 5524 2904
rect 5580 2896 5588 2904
rect 5644 2896 5652 2904
rect 4636 2876 4644 2884
rect 5164 2876 5172 2884
rect 5964 2896 5972 2904
rect 6028 2896 6036 2904
rect 6124 2896 6132 2904
rect 6652 2896 6660 2904
rect 7164 2896 7172 2904
rect 7532 2916 7540 2924
rect 5852 2876 5860 2884
rect 6492 2876 6500 2884
rect 6556 2876 6564 2884
rect 2764 2856 2772 2864
rect 3500 2856 3508 2864
rect 412 2836 420 2844
rect 508 2836 516 2844
rect 892 2836 900 2844
rect 1356 2836 1364 2844
rect 1564 2836 1572 2844
rect 1660 2836 1668 2844
rect 1852 2836 1860 2844
rect 2204 2836 2212 2844
rect 2860 2836 2868 2844
rect 3196 2836 3204 2844
rect 3404 2836 3412 2844
rect 4316 2836 4324 2844
rect 4588 2836 4596 2844
rect 4860 2836 4868 2844
rect 4940 2836 4948 2844
rect 5148 2836 5156 2844
rect 5836 2836 5844 2844
rect 5900 2836 5908 2844
rect 7500 2836 7508 2844
rect 739 2806 747 2814
rect 749 2806 757 2814
rect 759 2806 767 2814
rect 769 2806 777 2814
rect 779 2806 787 2814
rect 789 2806 797 2814
rect 3747 2806 3755 2814
rect 3757 2806 3765 2814
rect 3767 2806 3775 2814
rect 3777 2806 3785 2814
rect 3787 2806 3795 2814
rect 3797 2806 3805 2814
rect 6755 2806 6763 2814
rect 6765 2806 6773 2814
rect 6775 2806 6783 2814
rect 6785 2806 6793 2814
rect 6795 2806 6803 2814
rect 6805 2806 6813 2814
rect 460 2776 468 2784
rect 556 2776 564 2784
rect 924 2776 932 2784
rect 1532 2776 1540 2784
rect 1868 2776 1876 2784
rect 2124 2776 2132 2784
rect 2668 2776 2676 2784
rect 2716 2776 2724 2784
rect 3532 2776 3540 2784
rect 3996 2776 4004 2784
rect 4988 2776 4996 2784
rect 5180 2776 5188 2784
rect 5420 2776 5428 2784
rect 5564 2776 5572 2784
rect 6028 2776 6036 2784
rect 6236 2776 6244 2784
rect 6540 2776 6548 2784
rect 6700 2776 6708 2784
rect 4428 2756 4436 2764
rect 4620 2756 4628 2764
rect 5580 2756 5588 2764
rect 7292 2756 7300 2764
rect 1484 2736 1492 2744
rect 1916 2736 1924 2744
rect 2300 2736 2308 2744
rect 3148 2736 3156 2744
rect 4124 2736 4132 2744
rect 860 2716 868 2724
rect 1004 2716 1012 2724
rect 1244 2716 1252 2724
rect 1436 2716 1444 2724
rect 1788 2716 1796 2724
rect 2076 2716 2084 2724
rect 140 2694 148 2702
rect 236 2696 244 2704
rect 252 2696 260 2704
rect 300 2696 308 2704
rect 364 2696 372 2704
rect 428 2696 436 2704
rect 476 2696 484 2704
rect 508 2696 516 2704
rect 524 2696 532 2704
rect 572 2696 580 2704
rect 588 2696 596 2704
rect 652 2694 660 2702
rect 908 2696 916 2704
rect 940 2696 948 2704
rect 956 2696 964 2704
rect 1020 2696 1028 2704
rect 1036 2696 1044 2704
rect 1052 2696 1060 2704
rect 1084 2696 1092 2704
rect 1116 2696 1124 2704
rect 1148 2696 1156 2704
rect 1212 2696 1220 2704
rect 1292 2696 1300 2704
rect 1308 2696 1316 2704
rect 1356 2696 1364 2704
rect 1404 2696 1412 2704
rect 1484 2696 1492 2704
rect 1500 2696 1508 2704
rect 1548 2696 1556 2704
rect 1596 2696 1604 2704
rect 1628 2696 1636 2704
rect 1660 2696 1668 2704
rect 1692 2696 1700 2704
rect 1724 2696 1732 2704
rect 1756 2696 1764 2704
rect 1820 2696 1828 2704
rect 1884 2696 1892 2704
rect 1900 2696 1908 2704
rect 1964 2696 1972 2704
rect 2012 2696 2020 2704
rect 2044 2696 2052 2704
rect 2092 2696 2100 2704
rect 2140 2696 2148 2704
rect 2156 2696 2164 2704
rect 2204 2696 2212 2704
rect 2412 2696 2420 2704
rect 124 2676 132 2684
rect 316 2676 324 2684
rect 620 2676 628 2684
rect 892 2676 900 2684
rect 2540 2694 2548 2702
rect 2684 2696 2692 2704
rect 2748 2696 2756 2704
rect 3452 2716 3460 2724
rect 4060 2716 4068 2724
rect 4316 2716 4324 2724
rect 4636 2716 4644 2724
rect 4780 2716 4788 2724
rect 4860 2716 4868 2724
rect 5004 2736 5012 2744
rect 5164 2736 5172 2744
rect 5852 2736 5860 2744
rect 6588 2736 6596 2744
rect 6716 2736 6724 2744
rect 7100 2736 7108 2744
rect 5132 2716 5140 2724
rect 5228 2716 5236 2724
rect 2812 2696 2820 2704
rect 2860 2696 2868 2704
rect 2876 2696 2884 2704
rect 2924 2696 2932 2704
rect 2972 2696 2980 2704
rect 3020 2696 3028 2704
rect 3052 2696 3060 2704
rect 3068 2696 3076 2704
rect 3116 2696 3124 2704
rect 3132 2696 3140 2704
rect 3228 2696 3236 2704
rect 3276 2694 3284 2702
rect 3372 2696 3380 2704
rect 3436 2696 3444 2704
rect 3500 2696 3508 2704
rect 3516 2696 3524 2704
rect 3564 2696 3572 2704
rect 3580 2696 3588 2704
rect 3612 2696 3620 2704
rect 3660 2696 3668 2704
rect 3692 2696 3700 2704
rect 3868 2694 3876 2702
rect 4012 2696 4020 2704
rect 4092 2696 4100 2704
rect 4236 2696 4244 2704
rect 4348 2696 4356 2704
rect 4380 2696 4388 2704
rect 4492 2694 4500 2702
rect 4652 2696 4660 2704
rect 4668 2696 4676 2704
rect 4716 2696 4724 2704
rect 4764 2696 4772 2704
rect 4860 2696 4868 2704
rect 4924 2696 4932 2704
rect 4956 2696 4964 2704
rect 4988 2696 4996 2704
rect 5036 2696 5044 2704
rect 5116 2696 5124 2704
rect 5148 2696 5156 2704
rect 5436 2716 5444 2724
rect 5484 2716 5492 2724
rect 5756 2716 5764 2724
rect 5948 2716 5956 2724
rect 6044 2716 6052 2724
rect 6428 2716 6436 2724
rect 7164 2716 7172 2724
rect 7196 2716 7204 2724
rect 5356 2696 5364 2704
rect 5532 2696 5540 2704
rect 5788 2696 5796 2704
rect 5804 2696 5812 2704
rect 5852 2696 5860 2704
rect 5932 2696 5940 2704
rect 5948 2696 5956 2704
rect 5980 2696 5988 2704
rect 6124 2696 6132 2704
rect 6204 2696 6212 2704
rect 6236 2696 6244 2704
rect 6252 2696 6260 2704
rect 6316 2696 6324 2704
rect 6332 2696 6340 2704
rect 6348 2696 6356 2704
rect 6412 2696 6420 2704
rect 6524 2696 6532 2704
rect 6572 2696 6580 2704
rect 6636 2696 6644 2704
rect 6700 2696 6708 2704
rect 6844 2696 6852 2704
rect 7036 2696 7044 2704
rect 7068 2696 7076 2704
rect 7148 2696 7156 2704
rect 7212 2696 7220 2704
rect 7260 2696 7268 2704
rect 7308 2696 7316 2704
rect 7372 2696 7380 2704
rect 7420 2696 7428 2704
rect 956 2676 964 2684
rect 1068 2676 1076 2684
rect 1132 2676 1140 2684
rect 1180 2676 1188 2684
rect 1196 2676 1204 2684
rect 1260 2676 1268 2684
rect 1292 2676 1300 2684
rect 1372 2676 1380 2684
rect 1388 2676 1396 2684
rect 1500 2676 1508 2684
rect 1564 2676 1572 2684
rect 1580 2676 1588 2684
rect 1644 2676 1652 2684
rect 1708 2676 1716 2684
rect 1836 2676 1844 2684
rect 1948 2676 1956 2684
rect 2012 2676 2020 2684
rect 2028 2676 2036 2684
rect 2396 2676 2404 2684
rect 2732 2676 2740 2684
rect 2780 2676 2788 2684
rect 2796 2676 2804 2684
rect 2860 2676 2868 2684
rect 2876 2676 2884 2684
rect 2940 2676 2948 2684
rect 3052 2676 3060 2684
rect 3372 2676 3380 2684
rect 3420 2676 3428 2684
rect 3484 2676 3492 2684
rect 3676 2676 3684 2684
rect 3708 2676 3716 2684
rect 3836 2676 3844 2684
rect 4108 2676 4116 2684
rect 4364 2676 4372 2684
rect 4396 2676 4404 2684
rect 4508 2676 4516 2684
rect 4812 2676 4820 2684
rect 4860 2676 4868 2684
rect 4908 2676 4916 2684
rect 5036 2676 5044 2684
rect 5196 2676 5204 2684
rect 5276 2676 5284 2684
rect 5404 2676 5412 2684
rect 5452 2676 5460 2684
rect 5612 2676 5620 2684
rect 5724 2676 5732 2684
rect 5916 2676 5924 2684
rect 5996 2676 6004 2684
rect 6012 2676 6020 2684
rect 6060 2676 6068 2684
rect 6076 2680 6084 2688
rect 6460 2680 6468 2688
rect 6588 2676 6596 2684
rect 6876 2676 6884 2684
rect 6940 2676 6948 2684
rect 6972 2676 6980 2684
rect 7052 2676 7060 2684
rect 7116 2676 7124 2684
rect 7324 2676 7332 2684
rect 7404 2676 7412 2684
rect 7436 2676 7444 2684
rect 204 2656 212 2664
rect 396 2656 404 2664
rect 940 2656 948 2664
rect 1020 2656 1028 2664
rect 1260 2656 1268 2664
rect 1292 2656 1300 2664
rect 1452 2656 1460 2664
rect 1660 2656 1668 2664
rect 1852 2656 1860 2664
rect 1932 2656 1940 2664
rect 2988 2656 2996 2664
rect 3340 2656 3348 2664
rect 3756 2656 3764 2664
rect 4060 2656 4068 2664
rect 4252 2656 4260 2664
rect 4428 2656 4436 2664
rect 4716 2656 4724 2664
rect 4732 2656 4740 2664
rect 4828 2656 4836 2664
rect 4924 2656 4932 2664
rect 5068 2656 5076 2664
rect 5084 2656 5092 2664
rect 5372 2656 5380 2664
rect 5500 2656 5508 2664
rect 5548 2656 5556 2664
rect 5596 2656 5604 2664
rect 5772 2656 5780 2664
rect 5804 2656 5812 2664
rect 5884 2656 5892 2664
rect 6124 2656 6132 2664
rect 6204 2656 6212 2664
rect 6284 2656 6292 2664
rect 6380 2656 6388 2664
rect 6492 2656 6500 2664
rect 6652 2656 6660 2664
rect 6812 2656 6820 2664
rect 6860 2656 6868 2664
rect 7244 2656 7252 2664
rect 7340 2656 7348 2664
rect 7356 2656 7364 2664
rect 7452 2656 7460 2664
rect 7516 2656 7524 2664
rect 12 2636 20 2644
rect 220 2636 228 2644
rect 332 2636 340 2644
rect 780 2636 788 2644
rect 860 2636 868 2644
rect 1116 2636 1124 2644
rect 1356 2636 1364 2644
rect 1436 2636 1444 2644
rect 1628 2636 1636 2644
rect 1724 2636 1732 2644
rect 1964 2636 1972 2644
rect 2076 2636 2084 2644
rect 2188 2636 2196 2644
rect 2668 2636 2676 2644
rect 2812 2636 2820 2644
rect 2924 2636 2932 2644
rect 3452 2636 3460 2644
rect 3724 2636 3732 2644
rect 4316 2636 4324 2644
rect 4780 2636 4788 2644
rect 4812 2636 4820 2644
rect 5196 2636 5204 2644
rect 5404 2636 5412 2644
rect 5468 2636 5476 2644
rect 5516 2636 5524 2644
rect 5676 2636 5684 2644
rect 5740 2636 5748 2644
rect 6108 2636 6116 2644
rect 6156 2636 6164 2644
rect 6940 2636 6948 2644
rect 7468 2636 7476 2644
rect 4716 2616 4724 2624
rect 4828 2616 4836 2624
rect 5372 2616 5380 2624
rect 6124 2616 6132 2624
rect 2243 2606 2251 2614
rect 2253 2606 2261 2614
rect 2263 2606 2271 2614
rect 2273 2606 2281 2614
rect 2283 2606 2291 2614
rect 2293 2606 2301 2614
rect 5251 2606 5259 2614
rect 5261 2606 5269 2614
rect 5271 2606 5279 2614
rect 5281 2606 5289 2614
rect 5291 2606 5299 2614
rect 5301 2606 5309 2614
rect 4476 2596 4484 2604
rect 4492 2596 4500 2604
rect 5484 2596 5492 2604
rect 5500 2596 5508 2604
rect 5596 2596 5604 2604
rect 12 2576 20 2584
rect 220 2576 228 2584
rect 300 2576 308 2584
rect 556 2576 564 2584
rect 604 2576 612 2584
rect 924 2576 932 2584
rect 1356 2576 1364 2584
rect 1660 2576 1668 2584
rect 2220 2576 2228 2584
rect 2428 2576 2436 2584
rect 2988 2576 2996 2584
rect 3052 2576 3060 2584
rect 3404 2576 3412 2584
rect 3948 2576 3956 2584
rect 4028 2576 4036 2584
rect 4044 2576 4052 2584
rect 4380 2576 4388 2584
rect 4572 2576 4580 2584
rect 4620 2576 4628 2584
rect 4748 2576 4756 2584
rect 4908 2576 4916 2584
rect 5356 2576 5364 2584
rect 5580 2576 5588 2584
rect 5900 2576 5908 2584
rect 6396 2576 6404 2584
rect 6412 2576 6420 2584
rect 6588 2576 6596 2584
rect 6684 2576 6692 2584
rect 6716 2576 6724 2584
rect 6828 2576 6836 2584
rect 7244 2576 7252 2584
rect 204 2556 212 2564
rect 364 2556 372 2564
rect 716 2556 724 2564
rect 940 2556 948 2564
rect 1548 2556 1556 2564
rect 3340 2556 3348 2564
rect 3436 2556 3444 2564
rect 3452 2556 3460 2564
rect 3628 2556 3636 2564
rect 3660 2556 3668 2564
rect 3676 2556 3684 2564
rect 3980 2556 3988 2564
rect 4060 2556 4068 2564
rect 4252 2556 4260 2564
rect 4476 2556 4484 2564
rect 4492 2556 4500 2564
rect 4844 2556 4852 2564
rect 5052 2556 5060 2564
rect 5164 2556 5172 2564
rect 172 2536 180 2544
rect 236 2536 244 2544
rect 284 2536 292 2544
rect 588 2536 596 2544
rect 764 2536 772 2544
rect 988 2536 996 2544
rect 1020 2536 1028 2544
rect 1052 2536 1060 2544
rect 1116 2536 1124 2544
rect 1196 2536 1204 2544
rect 1372 2536 1380 2544
rect 1500 2536 1508 2544
rect 1772 2536 1780 2544
rect 1852 2536 1860 2544
rect 1916 2536 1924 2544
rect 2060 2536 2068 2544
rect 2124 2536 2132 2544
rect 2156 2536 2164 2544
rect 2172 2536 2180 2544
rect 2332 2536 2340 2544
rect 2444 2536 2452 2544
rect 2508 2536 2516 2544
rect 2700 2536 2708 2544
rect 2764 2536 2772 2544
rect 2796 2536 2804 2544
rect 2892 2536 2900 2544
rect 3004 2536 3012 2544
rect 3116 2536 3124 2544
rect 3148 2536 3156 2544
rect 140 2518 148 2526
rect 268 2516 276 2524
rect 332 2516 340 2524
rect 428 2518 436 2526
rect 492 2516 500 2524
rect 572 2516 580 2524
rect 636 2516 644 2524
rect 812 2516 820 2524
rect 972 2516 980 2524
rect 1068 2516 1076 2524
rect 1116 2516 1124 2524
rect 1132 2516 1140 2524
rect 1228 2518 1236 2526
rect 1388 2516 1396 2524
rect 1452 2516 1460 2524
rect 1484 2516 1492 2524
rect 1516 2516 1524 2524
rect 1532 2516 1540 2524
rect 1564 2516 1572 2524
rect 1580 2516 1588 2524
rect 1644 2516 1652 2524
rect 1788 2518 1796 2526
rect 1868 2516 1876 2524
rect 1996 2516 2004 2524
rect 2044 2516 2052 2524
rect 1100 2496 1108 2504
rect 1164 2496 1172 2504
rect 1420 2496 1428 2504
rect 1948 2496 1956 2504
rect 2092 2496 2100 2504
rect 2140 2516 2148 2524
rect 2348 2516 2356 2524
rect 2396 2516 2404 2524
rect 2444 2516 2452 2524
rect 2524 2516 2532 2524
rect 2572 2516 2580 2524
rect 2588 2516 2596 2524
rect 2620 2516 2628 2524
rect 2668 2516 2676 2524
rect 2684 2516 2692 2524
rect 2716 2516 2724 2524
rect 2860 2518 2868 2526
rect 2300 2496 2308 2504
rect 2492 2496 2500 2504
rect 3004 2516 3012 2524
rect 2764 2496 2772 2504
rect 3100 2516 3108 2524
rect 3260 2536 3268 2544
rect 3356 2536 3364 2544
rect 3500 2536 3508 2544
rect 3596 2536 3604 2544
rect 3788 2536 3796 2544
rect 4060 2536 4068 2544
rect 4092 2536 4100 2544
rect 4188 2536 4196 2544
rect 4412 2536 4420 2544
rect 4620 2536 4628 2544
rect 4684 2536 4692 2544
rect 4828 2536 4836 2544
rect 4876 2536 4884 2544
rect 4908 2536 4916 2544
rect 4988 2536 4996 2544
rect 5116 2536 5124 2544
rect 5484 2556 5492 2564
rect 5500 2556 5508 2564
rect 5596 2556 5604 2564
rect 5820 2556 5828 2564
rect 5948 2556 5956 2564
rect 6076 2556 6084 2564
rect 6220 2556 6228 2564
rect 6300 2556 6308 2564
rect 6476 2556 6484 2564
rect 6572 2556 6580 2564
rect 6652 2556 6660 2564
rect 6956 2556 6964 2564
rect 7052 2556 7060 2564
rect 7260 2556 7268 2564
rect 7340 2556 7348 2564
rect 5212 2536 5220 2544
rect 5340 2536 5348 2544
rect 5356 2536 5364 2544
rect 5836 2536 5844 2544
rect 5948 2536 5956 2544
rect 5980 2536 5988 2544
rect 6124 2536 6132 2544
rect 6428 2536 6436 2544
rect 6460 2536 6468 2544
rect 6492 2536 6500 2544
rect 6588 2536 6596 2544
rect 6620 2536 6628 2544
rect 6636 2536 6644 2544
rect 6668 2536 6676 2544
rect 6716 2536 6724 2544
rect 6780 2536 6788 2544
rect 7036 2536 7044 2544
rect 7100 2536 7108 2544
rect 7196 2536 7204 2544
rect 7308 2536 7316 2544
rect 7356 2536 7364 2544
rect 7452 2536 7460 2544
rect 3180 2516 3188 2524
rect 3068 2496 3076 2504
rect 3308 2516 3316 2524
rect 3372 2516 3380 2524
rect 3484 2516 3492 2524
rect 3548 2516 3556 2524
rect 3580 2516 3588 2524
rect 3596 2516 3604 2524
rect 3820 2518 3828 2526
rect 3996 2516 4004 2524
rect 4076 2516 4084 2524
rect 4124 2516 4132 2524
rect 4172 2516 4180 2524
rect 4252 2518 4260 2526
rect 4300 2516 4308 2524
rect 4428 2516 4436 2524
rect 4540 2516 4548 2524
rect 3228 2496 3236 2504
rect 3404 2496 3412 2504
rect 3548 2496 3556 2504
rect 3676 2496 3684 2504
rect 4140 2496 4148 2504
rect 4396 2496 4404 2504
rect 4636 2516 4644 2524
rect 4716 2516 4724 2524
rect 4812 2516 4820 2524
rect 4940 2516 4948 2524
rect 5084 2516 5092 2524
rect 5132 2516 5140 2524
rect 5196 2516 5204 2524
rect 5228 2516 5236 2524
rect 4588 2496 4596 2504
rect 4876 2496 4884 2504
rect 4908 2496 4916 2504
rect 5036 2496 5044 2504
rect 5116 2496 5124 2504
rect 5356 2496 5364 2504
rect 5388 2496 5396 2504
rect 5436 2516 5444 2524
rect 5548 2516 5556 2524
rect 5644 2516 5652 2524
rect 5676 2516 5684 2524
rect 5740 2516 5748 2524
rect 5788 2516 5796 2524
rect 6028 2516 6036 2524
rect 6156 2516 6164 2524
rect 6172 2516 6180 2524
rect 6252 2516 6260 2524
rect 6332 2516 6340 2524
rect 6364 2516 6372 2524
rect 6412 2516 6420 2524
rect 6476 2516 6484 2524
rect 6572 2516 6580 2524
rect 6652 2516 6660 2524
rect 6716 2516 6724 2524
rect 6748 2516 6756 2524
rect 6780 2516 6788 2524
rect 6924 2516 6932 2524
rect 6940 2516 6948 2524
rect 6972 2516 6980 2524
rect 7052 2516 7060 2524
rect 7084 2516 7092 2524
rect 7100 2516 7108 2524
rect 5596 2496 5604 2504
rect 6028 2496 6036 2504
rect 6284 2496 6292 2504
rect 6460 2496 6468 2504
rect 6524 2496 6532 2504
rect 6700 2496 6708 2504
rect 6988 2496 6996 2504
rect 7212 2516 7220 2524
rect 7484 2516 7492 2524
rect 7516 2516 7524 2524
rect 7164 2496 7172 2504
rect 7532 2496 7540 2504
rect 1132 2476 1140 2484
rect 1868 2476 1876 2484
rect 2012 2476 2020 2484
rect 3628 2476 3636 2484
rect 3916 2476 3924 2484
rect 5436 2476 5444 2484
rect 7084 2476 7092 2484
rect 7388 2476 7396 2484
rect 7116 2456 7124 2464
rect 1484 2436 1492 2444
rect 1596 2436 1604 2444
rect 1964 2436 1972 2444
rect 2380 2436 2388 2444
rect 2540 2436 2548 2444
rect 2636 2436 2644 2444
rect 3180 2436 3188 2444
rect 3276 2436 3284 2444
rect 3324 2436 3332 2444
rect 3420 2436 3428 2444
rect 3468 2436 3476 2444
rect 3964 2436 3972 2444
rect 5004 2436 5012 2444
rect 5644 2436 5652 2444
rect 6252 2436 6260 2444
rect 6540 2436 6548 2444
rect 7340 2436 7348 2444
rect 739 2406 747 2414
rect 749 2406 757 2414
rect 759 2406 767 2414
rect 769 2406 777 2414
rect 779 2406 787 2414
rect 789 2406 797 2414
rect 3747 2406 3755 2414
rect 3757 2406 3765 2414
rect 3767 2406 3775 2414
rect 3777 2406 3785 2414
rect 3787 2406 3795 2414
rect 3797 2406 3805 2414
rect 6755 2406 6763 2414
rect 6765 2406 6773 2414
rect 6775 2406 6783 2414
rect 6785 2406 6793 2414
rect 6795 2406 6803 2414
rect 6805 2406 6813 2414
rect 124 2376 132 2384
rect 364 2376 372 2384
rect 412 2376 420 2384
rect 1052 2376 1060 2384
rect 1452 2376 1460 2384
rect 1564 2376 1572 2384
rect 1708 2376 1716 2384
rect 1916 2376 1924 2384
rect 2028 2376 2036 2384
rect 2364 2376 2372 2384
rect 2508 2376 2516 2384
rect 3212 2376 3220 2384
rect 4156 2376 4164 2384
rect 4620 2376 4628 2384
rect 5196 2376 5204 2384
rect 5436 2376 5444 2384
rect 5580 2376 5588 2384
rect 6348 2376 6356 2384
rect 6620 2376 6628 2384
rect 6844 2376 6852 2384
rect 7052 2376 7060 2384
rect 7116 2376 7124 2384
rect 7532 2376 7540 2384
rect 3628 2356 3636 2364
rect 6572 2356 6580 2364
rect 268 2336 276 2344
rect 1292 2336 1300 2344
rect 1372 2336 1380 2344
rect 1964 2336 1972 2344
rect 2124 2336 2132 2344
rect 3180 2336 3188 2344
rect 4076 2336 4084 2344
rect 4092 2336 4100 2344
rect 5004 2336 5012 2344
rect 5404 2336 5412 2344
rect 5452 2336 5460 2344
rect 5708 2336 5716 2344
rect 5980 2336 5988 2344
rect 6796 2336 6804 2344
rect 6828 2336 6836 2344
rect 7132 2336 7140 2344
rect 860 2316 868 2324
rect 1324 2316 1332 2324
rect 156 2296 164 2304
rect 204 2296 212 2304
rect 300 2296 308 2304
rect 332 2296 340 2304
rect 508 2296 516 2304
rect 636 2296 644 2304
rect 828 2296 836 2304
rect 860 2296 868 2304
rect 924 2294 932 2302
rect 988 2296 996 2304
rect 1100 2296 1108 2304
rect 1180 2296 1188 2304
rect 1324 2296 1332 2304
rect 1404 2296 1412 2304
rect 1484 2296 1492 2304
rect 1772 2316 1780 2324
rect 2428 2316 2436 2324
rect 1564 2296 1572 2304
rect 1676 2296 1684 2304
rect 1708 2296 1716 2304
rect 1740 2296 1748 2304
rect 1788 2296 1796 2304
rect 1836 2296 1844 2304
rect 1868 2296 1876 2304
rect 1884 2296 1892 2304
rect 1932 2296 1940 2304
rect 1996 2296 2004 2304
rect 2092 2296 2100 2304
rect 2156 2296 2164 2304
rect 2172 2296 2180 2304
rect 2204 2296 2212 2304
rect 2252 2296 2260 2304
rect 2268 2296 2276 2304
rect 3452 2316 3460 2324
rect 3468 2316 3476 2324
rect 3644 2316 3652 2324
rect 3836 2316 3844 2324
rect 4172 2316 4180 2324
rect 2476 2296 2484 2304
rect 2620 2296 2628 2304
rect 2908 2296 2916 2304
rect 2972 2294 2980 2302
rect 3116 2296 3124 2304
rect 3228 2296 3236 2304
rect 3292 2296 3300 2304
rect 3388 2296 3396 2304
rect 3404 2296 3412 2304
rect 3500 2296 3508 2304
rect 3532 2296 3540 2304
rect 3596 2296 3604 2304
rect 3676 2296 3684 2304
rect 3692 2296 3700 2304
rect 3756 2296 3764 2304
rect 12 2276 20 2284
rect 188 2276 196 2284
rect 236 2280 244 2288
rect 252 2276 260 2284
rect 316 2276 324 2284
rect 620 2276 628 2284
rect 812 2276 820 2284
rect 1196 2276 1204 2284
rect 1228 2276 1236 2284
rect 1308 2276 1316 2284
rect 1436 2276 1444 2284
rect 1468 2276 1476 2284
rect 1484 2276 1492 2284
rect 1548 2276 1556 2284
rect 1612 2276 1620 2284
rect 1724 2276 1732 2284
rect 1820 2276 1828 2284
rect 1852 2276 1860 2284
rect 2012 2276 2020 2284
rect 2380 2276 2388 2284
rect 2396 2276 2404 2284
rect 2460 2276 2468 2284
rect 2492 2276 2500 2284
rect 2668 2276 2676 2284
rect 2700 2276 2708 2284
rect 2828 2276 2836 2284
rect 3244 2276 3252 2284
rect 3292 2276 3300 2284
rect 3324 2276 3332 2284
rect 3356 2276 3364 2284
rect 3420 2276 3428 2284
rect 3516 2276 3524 2284
rect 3548 2276 3556 2284
rect 3708 2276 3716 2284
rect 3724 2276 3732 2284
rect 188 2256 196 2264
rect 428 2256 436 2264
rect 540 2256 548 2264
rect 1628 2256 1636 2264
rect 1660 2256 1668 2264
rect 3276 2256 3284 2264
rect 3580 2256 3588 2264
rect 3884 2296 3892 2304
rect 3948 2294 3956 2302
rect 4124 2296 4132 2304
rect 4236 2296 4244 2304
rect 4284 2316 4292 2324
rect 4524 2316 4532 2324
rect 4940 2316 4948 2324
rect 5004 2316 5012 2324
rect 5164 2316 5172 2324
rect 5276 2316 5284 2324
rect 5420 2316 5428 2324
rect 5500 2316 5508 2324
rect 5676 2316 5684 2324
rect 5932 2316 5940 2324
rect 6092 2316 6100 2324
rect 6444 2316 6452 2324
rect 6460 2316 6468 2324
rect 6668 2316 6676 2324
rect 6860 2316 6868 2324
rect 6972 2316 6980 2324
rect 7164 2316 7172 2324
rect 7212 2316 7220 2324
rect 7276 2316 7284 2324
rect 4476 2296 4484 2304
rect 4572 2296 4580 2304
rect 3884 2276 3892 2284
rect 3916 2276 3924 2284
rect 4140 2276 4148 2284
rect 4316 2276 4324 2284
rect 4332 2276 4340 2284
rect 4348 2280 4356 2288
rect 4188 2256 4196 2264
rect 4492 2276 4500 2284
rect 4524 2276 4532 2284
rect 4444 2256 4452 2264
rect 4524 2256 4532 2264
rect 4652 2276 4660 2284
rect 4684 2296 4692 2304
rect 4780 2296 4788 2304
rect 4572 2256 4580 2264
rect 4604 2256 4612 2264
rect 4620 2256 4628 2264
rect 4716 2256 4724 2264
rect 4748 2276 4756 2284
rect 4764 2276 4772 2284
rect 4796 2276 4804 2284
rect 4892 2276 4900 2284
rect 4988 2296 4996 2304
rect 5020 2296 5028 2304
rect 5116 2296 5124 2304
rect 5244 2296 5252 2304
rect 5324 2296 5332 2304
rect 5436 2296 5444 2304
rect 5516 2296 5524 2304
rect 5532 2296 5540 2304
rect 5596 2296 5604 2304
rect 5756 2296 5764 2304
rect 5820 2296 5828 2304
rect 5900 2296 5908 2304
rect 5948 2296 5956 2304
rect 6012 2296 6020 2304
rect 6108 2296 6116 2304
rect 6172 2296 6180 2304
rect 6188 2296 6196 2304
rect 6476 2296 6484 2304
rect 6540 2296 6548 2304
rect 6588 2296 6596 2304
rect 6668 2296 6676 2304
rect 6844 2296 6852 2304
rect 6924 2296 6932 2304
rect 7100 2296 7108 2304
rect 7132 2296 7140 2304
rect 7180 2296 7188 2304
rect 7196 2296 7204 2304
rect 7244 2296 7252 2304
rect 4972 2276 4980 2284
rect 5036 2276 5044 2284
rect 5084 2276 5092 2284
rect 5228 2276 5236 2284
rect 5372 2276 5380 2284
rect 5548 2276 5556 2284
rect 5676 2276 5684 2284
rect 5708 2276 5716 2284
rect 5852 2276 5860 2284
rect 5916 2276 5924 2284
rect 6060 2276 6068 2284
rect 6156 2276 6164 2284
rect 6252 2276 6260 2284
rect 6316 2276 6324 2284
rect 6348 2276 6356 2284
rect 6444 2276 6452 2284
rect 6476 2276 6484 2284
rect 6636 2276 6644 2284
rect 6700 2276 6708 2284
rect 6908 2276 6916 2284
rect 6940 2276 6948 2284
rect 7036 2276 7044 2284
rect 7084 2276 7092 2284
rect 7260 2276 7268 2284
rect 7324 2276 7332 2284
rect 7436 2296 7444 2304
rect 7484 2296 7492 2304
rect 7516 2296 7524 2304
rect 7484 2276 7492 2284
rect 5068 2256 5076 2264
rect 5084 2256 5092 2264
rect 5212 2256 5220 2264
rect 5356 2256 5364 2264
rect 5484 2256 5492 2264
rect 5660 2256 5668 2264
rect 5772 2256 5780 2264
rect 5820 2256 5828 2264
rect 5900 2256 5908 2264
rect 5964 2256 5972 2264
rect 5996 2256 6004 2264
rect 6236 2256 6244 2264
rect 6428 2256 6436 2264
rect 6684 2256 6692 2264
rect 6876 2256 6884 2264
rect 7052 2256 7060 2264
rect 7196 2256 7204 2264
rect 7484 2256 7492 2264
rect 7548 2256 7556 2264
rect 476 2236 484 2244
rect 524 2236 532 2244
rect 732 2236 740 2244
rect 1068 2236 1076 2244
rect 1532 2236 1540 2244
rect 2028 2236 2036 2244
rect 2220 2236 2228 2244
rect 2844 2236 2852 2244
rect 3260 2236 3268 2244
rect 3564 2236 3572 2244
rect 3644 2236 3652 2244
rect 4140 2236 4148 2244
rect 4268 2236 4276 2244
rect 4316 2236 4324 2244
rect 4412 2236 4420 2244
rect 4940 2236 4948 2244
rect 5292 2236 5300 2244
rect 5324 2236 5332 2244
rect 5676 2236 5684 2244
rect 5724 2236 5732 2244
rect 6156 2236 6164 2244
rect 6524 2236 6532 2244
rect 6892 2236 6900 2244
rect 4188 2216 4196 2224
rect 5084 2216 5092 2224
rect 2243 2206 2251 2214
rect 2253 2206 2261 2214
rect 2263 2206 2271 2214
rect 2273 2206 2281 2214
rect 2283 2206 2291 2214
rect 2293 2206 2301 2214
rect 5251 2206 5259 2214
rect 5261 2206 5269 2214
rect 5271 2206 5279 2214
rect 5281 2206 5289 2214
rect 5291 2206 5299 2214
rect 5301 2206 5309 2214
rect 5516 2196 5524 2204
rect 5836 2196 5844 2204
rect 220 2176 228 2184
rect 460 2176 468 2184
rect 556 2176 564 2184
rect 636 2176 644 2184
rect 844 2176 852 2184
rect 1388 2176 1396 2184
rect 1724 2176 1732 2184
rect 2492 2176 2500 2184
rect 2620 2176 2628 2184
rect 2972 2176 2980 2184
rect 3340 2176 3348 2184
rect 4044 2176 4052 2184
rect 4060 2176 4068 2184
rect 12 2156 20 2164
rect 44 2156 52 2164
rect 156 2156 164 2164
rect 204 2156 212 2164
rect 300 2156 308 2164
rect 1100 2156 1108 2164
rect 2556 2156 2564 2164
rect 2748 2156 2756 2164
rect 2892 2156 2900 2164
rect 2908 2156 2916 2164
rect 2988 2156 2996 2164
rect 3148 2156 3156 2164
rect 3404 2156 3412 2164
rect 3612 2156 3620 2164
rect 3916 2156 3924 2164
rect 4076 2156 4084 2164
rect 4524 2156 4532 2164
rect 4684 2176 4692 2184
rect 4892 2176 4900 2184
rect 5052 2176 5060 2184
rect 5196 2176 5204 2184
rect 5596 2176 5604 2184
rect 5644 2176 5652 2184
rect 5660 2176 5668 2184
rect 5692 2176 5700 2184
rect 5708 2176 5716 2184
rect 5868 2176 5876 2184
rect 5948 2176 5956 2184
rect 6236 2176 6244 2184
rect 6332 2176 6340 2184
rect 6396 2176 6404 2184
rect 6508 2176 6516 2184
rect 6716 2176 6724 2184
rect 6892 2176 6900 2184
rect 6988 2176 6996 2184
rect 7084 2176 7092 2184
rect 7164 2176 7172 2184
rect 7356 2176 7364 2184
rect 7388 2176 7396 2184
rect 7468 2176 7476 2184
rect 4620 2156 4628 2164
rect 4700 2156 4708 2164
rect 4732 2156 4740 2164
rect 4748 2156 4756 2164
rect 4956 2156 4964 2164
rect 4988 2156 4996 2164
rect 5148 2156 5156 2164
rect 5212 2156 5220 2164
rect 5516 2156 5524 2164
rect 5836 2156 5844 2164
rect 6284 2156 6292 2164
rect 6412 2156 6420 2164
rect 6428 2156 6436 2164
rect 6588 2156 6596 2164
rect 6700 2156 6708 2164
rect 6956 2156 6964 2164
rect 6972 2156 6980 2164
rect 7068 2156 7076 2164
rect 7100 2156 7108 2164
rect 44 2136 52 2144
rect 268 2136 276 2144
rect 284 2136 292 2144
rect 332 2136 340 2144
rect 396 2136 404 2144
rect 476 2136 484 2144
rect 572 2136 580 2144
rect 588 2136 596 2144
rect 684 2136 692 2144
rect 956 2136 964 2144
rect 1180 2136 1188 2144
rect 1228 2136 1236 2144
rect 1708 2136 1716 2144
rect 1772 2136 1780 2144
rect 1884 2136 1892 2144
rect 1996 2136 2004 2144
rect 2108 2136 2116 2144
rect 2332 2136 2340 2144
rect 2508 2136 2516 2144
rect 2604 2136 2612 2144
rect 2700 2136 2708 2144
rect 2764 2136 2772 2144
rect 2876 2136 2884 2144
rect 76 2116 84 2124
rect 92 2116 100 2124
rect 124 2116 132 2124
rect 172 2116 180 2124
rect 188 2116 196 2124
rect 252 2116 260 2124
rect 348 2116 356 2124
rect 380 2116 388 2124
rect 540 2116 548 2124
rect 604 2116 612 2124
rect 316 2096 324 2104
rect 444 2096 452 2104
rect 524 2096 532 2104
rect 540 2096 548 2104
rect 684 2116 692 2124
rect 812 2116 820 2124
rect 860 2116 868 2124
rect 876 2116 884 2124
rect 924 2116 932 2124
rect 972 2116 980 2124
rect 988 2116 996 2124
rect 1004 2116 1012 2124
rect 1068 2116 1076 2124
rect 1132 2116 1140 2124
rect 1164 2116 1172 2124
rect 1196 2116 1204 2124
rect 1260 2118 1268 2126
rect 1420 2116 1428 2124
rect 1436 2116 1444 2124
rect 1532 2116 1540 2124
rect 1596 2118 1604 2126
rect 1692 2116 1700 2124
rect 1756 2116 1764 2124
rect 1820 2116 1828 2124
rect 1836 2116 1844 2124
rect 1900 2116 1908 2124
rect 652 2096 660 2104
rect 1036 2096 1044 2104
rect 1452 2096 1460 2104
rect 1692 2096 1700 2104
rect 1724 2096 1732 2104
rect 1980 2116 1988 2124
rect 2124 2116 2132 2124
rect 2300 2116 2308 2124
rect 2380 2116 2388 2124
rect 1980 2096 1988 2104
rect 2540 2096 2548 2104
rect 2588 2116 2596 2124
rect 2652 2116 2660 2124
rect 2668 2116 2676 2124
rect 2716 2116 2724 2124
rect 2780 2116 2788 2124
rect 2860 2116 2868 2124
rect 2956 2136 2964 2144
rect 2988 2136 2996 2144
rect 3068 2136 3076 2144
rect 3180 2136 3188 2144
rect 3372 2136 3380 2144
rect 3436 2136 3444 2144
rect 3676 2136 3684 2144
rect 3692 2136 3700 2144
rect 3852 2136 3860 2144
rect 4108 2136 4116 2144
rect 4300 2136 4308 2144
rect 2940 2116 2948 2124
rect 3036 2116 3044 2124
rect 3052 2116 3060 2124
rect 3116 2116 3124 2124
rect 3212 2118 3220 2126
rect 3356 2116 3364 2124
rect 3468 2118 3476 2126
rect 3644 2116 3652 2124
rect 3660 2116 3668 2124
rect 3836 2116 3844 2124
rect 3932 2116 3940 2124
rect 4140 2118 4148 2126
rect 4332 2118 4340 2126
rect 4508 2116 4516 2124
rect 4572 2136 4580 2144
rect 4668 2136 4676 2144
rect 4780 2136 4788 2144
rect 4844 2136 4852 2144
rect 4908 2136 4916 2144
rect 5004 2136 5012 2144
rect 5132 2136 5140 2144
rect 5180 2136 5188 2144
rect 5292 2136 5300 2144
rect 5388 2136 5396 2144
rect 5404 2136 5412 2144
rect 5452 2136 5460 2144
rect 5644 2136 5652 2144
rect 5692 2136 5700 2144
rect 5708 2136 5716 2144
rect 5884 2136 5892 2144
rect 5900 2136 5908 2144
rect 5996 2136 6004 2144
rect 6012 2136 6020 2144
rect 6028 2132 6036 2140
rect 6220 2136 6228 2144
rect 6268 2136 6276 2144
rect 6380 2136 6388 2144
rect 6460 2136 6468 2144
rect 6572 2136 6580 2144
rect 6652 2136 6660 2144
rect 6764 2136 6772 2144
rect 6780 2136 6788 2144
rect 6860 2136 6868 2144
rect 7148 2136 7156 2144
rect 7196 2156 7204 2164
rect 7244 2156 7252 2164
rect 7308 2156 7316 2164
rect 7372 2156 7380 2164
rect 7340 2136 7348 2144
rect 7420 2136 7428 2144
rect 7436 2136 7444 2144
rect 7532 2136 7540 2144
rect 4620 2116 4628 2124
rect 4652 2116 4660 2124
rect 4780 2116 4788 2124
rect 4828 2116 4836 2124
rect 4860 2116 4868 2124
rect 4956 2116 4964 2124
rect 5212 2116 5220 2124
rect 5564 2116 5572 2124
rect 3100 2096 3108 2104
rect 3612 2096 3620 2104
rect 3772 2096 3780 2104
rect 3788 2096 3796 2104
rect 4700 2096 4708 2104
rect 5100 2096 5108 2104
rect 5148 2096 5156 2104
rect 5436 2096 5444 2104
rect 5500 2096 5508 2104
rect 5612 2096 5620 2104
rect 5660 2096 5668 2104
rect 5740 2096 5748 2104
rect 5788 2116 5796 2124
rect 6076 2116 6084 2124
rect 5852 2096 5860 2104
rect 6332 2116 6340 2124
rect 6476 2116 6484 2124
rect 6572 2116 6580 2124
rect 6668 2116 6676 2124
rect 6748 2116 6756 2124
rect 6924 2116 6932 2124
rect 7004 2116 7012 2124
rect 7020 2116 7028 2124
rect 7132 2116 7140 2124
rect 7228 2116 7236 2124
rect 6428 2096 6436 2104
rect 6524 2096 6532 2104
rect 6556 2096 6564 2104
rect 6620 2096 6628 2104
rect 6684 2096 6692 2104
rect 6716 2096 6724 2104
rect 6876 2096 6884 2104
rect 6940 2096 6948 2104
rect 7116 2096 7124 2104
rect 7388 2096 7396 2104
rect 76 2076 84 2084
rect 108 2076 116 2084
rect 732 2076 740 2084
rect 908 2076 916 2084
rect 1660 2076 1668 2084
rect 1932 2076 1940 2084
rect 2012 2076 2020 2084
rect 2812 2076 2820 2084
rect 3308 2076 3316 2084
rect 4012 2076 4020 2084
rect 4460 2076 4468 2084
rect 4476 2076 4484 2084
rect 6108 2076 6116 2084
rect 6652 2076 6660 2084
rect 412 2036 420 2044
rect 844 2036 852 2044
rect 1468 2036 1476 2044
rect 1788 2036 1796 2044
rect 1868 2036 1876 2044
rect 2204 2036 2212 2044
rect 2860 2036 2868 2044
rect 3404 2036 3412 2044
rect 3596 2036 3604 2044
rect 4268 2036 4276 2044
rect 4556 2036 4564 2044
rect 4972 2036 4980 2044
rect 5468 2036 5476 2044
rect 5788 2036 5796 2044
rect 6060 2036 6068 2044
rect 739 2006 747 2014
rect 749 2006 757 2014
rect 759 2006 767 2014
rect 769 2006 777 2014
rect 779 2006 787 2014
rect 789 2006 797 2014
rect 3747 2006 3755 2014
rect 3757 2006 3765 2014
rect 3767 2006 3775 2014
rect 3777 2006 3785 2014
rect 3787 2006 3795 2014
rect 3797 2006 3805 2014
rect 6755 2006 6763 2014
rect 6765 2006 6773 2014
rect 6775 2006 6783 2014
rect 6785 2006 6793 2014
rect 6795 2006 6803 2014
rect 6805 2006 6813 2014
rect 556 1976 564 1984
rect 1516 1976 1524 1984
rect 1548 1976 1556 1984
rect 2892 1976 2900 1984
rect 2940 1976 2948 1984
rect 2988 1976 2996 1984
rect 3036 1976 3044 1984
rect 3068 1976 3076 1984
rect 3276 1976 3284 1984
rect 3580 1976 3588 1984
rect 4156 1976 4164 1984
rect 4236 1976 4244 1984
rect 4364 1976 4372 1984
rect 4428 1976 4436 1984
rect 4524 1976 4532 1984
rect 4572 1976 4580 1984
rect 4700 1976 4708 1984
rect 5148 1976 5156 1984
rect 5900 1976 5908 1984
rect 5964 1976 5972 1984
rect 6316 1976 6324 1984
rect 6428 1976 6436 1984
rect 6716 1976 6724 1984
rect 6988 1976 6996 1984
rect 7468 1976 7476 1984
rect 492 1956 500 1964
rect 652 1956 660 1964
rect 12 1936 20 1944
rect 4108 1936 4116 1944
rect 4140 1936 4148 1944
rect 4636 1936 4644 1944
rect 4716 1936 4724 1944
rect 4748 1936 4756 1944
rect 140 1894 148 1902
rect 220 1896 228 1904
rect 236 1896 244 1904
rect 268 1916 276 1924
rect 1052 1916 1060 1924
rect 1260 1916 1268 1924
rect 1292 1916 1300 1924
rect 1324 1916 1332 1924
rect 1916 1916 1924 1924
rect 396 1896 404 1904
rect 508 1896 516 1904
rect 524 1896 532 1904
rect 572 1896 580 1904
rect 668 1896 676 1904
rect 684 1896 692 1904
rect 828 1896 836 1904
rect 972 1896 980 1904
rect 988 1896 996 1904
rect 1132 1896 1140 1904
rect 1340 1896 1348 1904
rect 1388 1896 1396 1904
rect 1420 1896 1428 1904
rect 1452 1896 1460 1904
rect 1468 1896 1476 1904
rect 1532 1896 1540 1904
rect 1580 1896 1588 1904
rect 1596 1896 1604 1904
rect 1660 1896 1668 1904
rect 1692 1896 1700 1904
rect 1820 1896 1828 1904
rect 1900 1896 1908 1904
rect 1964 1916 1972 1924
rect 2796 1916 2804 1924
rect 2060 1894 2068 1902
rect 2204 1896 2212 1904
rect 2220 1896 2228 1904
rect 2268 1896 2276 1904
rect 2428 1896 2436 1904
rect 2460 1896 2468 1904
rect 2492 1896 2500 1904
rect 2556 1896 2564 1904
rect 3324 1916 3332 1924
rect 3356 1916 3364 1924
rect 3420 1916 3428 1924
rect 3484 1916 3492 1924
rect 3548 1916 3556 1924
rect 3612 1916 3620 1924
rect 3644 1916 3652 1924
rect 3676 1916 3684 1924
rect 3740 1916 3748 1924
rect 4412 1916 4420 1924
rect 4460 1916 4468 1924
rect 4492 1916 4500 1924
rect 4636 1916 4644 1924
rect 4668 1916 4676 1924
rect 4684 1916 4692 1924
rect 4876 1916 4884 1924
rect 5020 1916 5028 1924
rect 5372 1916 5380 1924
rect 5436 1916 5444 1924
rect 5532 1916 5540 1924
rect 5612 1916 5620 1924
rect 6364 1916 6372 1924
rect 6700 1916 6708 1924
rect 6828 1916 6836 1924
rect 6940 1916 6948 1924
rect 7052 1916 7060 1924
rect 2620 1894 2628 1902
rect 2844 1896 2852 1904
rect 3164 1896 3172 1904
rect 3292 1896 3300 1904
rect 3388 1896 3396 1904
rect 3452 1896 3460 1904
rect 3516 1896 3524 1904
rect 3580 1896 3588 1904
rect 3644 1896 3652 1904
rect 3708 1896 3716 1904
rect 4028 1896 4036 1904
rect 4188 1896 4196 1904
rect 4204 1896 4212 1904
rect 4284 1896 4292 1904
rect 4364 1896 4372 1904
rect 4540 1896 4548 1904
rect 4700 1896 4708 1904
rect 4748 1896 4756 1904
rect 4796 1896 4804 1904
rect 4860 1896 4868 1904
rect 4908 1896 4916 1904
rect 5052 1896 5060 1904
rect 5340 1896 5348 1904
rect 5468 1896 5476 1904
rect 5692 1896 5700 1904
rect 5740 1896 5748 1904
rect 5804 1896 5812 1904
rect 5836 1896 5844 1904
rect 5852 1896 5860 1904
rect 5932 1896 5940 1904
rect 5964 1896 5972 1904
rect 5996 1896 6004 1904
rect 6060 1896 6068 1904
rect 6092 1896 6100 1904
rect 6108 1896 6116 1904
rect 6172 1896 6180 1904
rect 6220 1896 6228 1904
rect 6252 1896 6260 1904
rect 6300 1896 6308 1904
rect 6348 1896 6356 1904
rect 6364 1896 6372 1904
rect 6396 1896 6404 1904
rect 6460 1896 6468 1904
rect 6508 1896 6516 1904
rect 6540 1896 6548 1904
rect 6652 1896 6660 1904
rect 6812 1896 6820 1904
rect 6876 1896 6884 1904
rect 6908 1896 6916 1904
rect 6924 1896 6932 1904
rect 6956 1896 6964 1904
rect 7004 1896 7012 1904
rect 7068 1896 7076 1904
rect 7196 1896 7204 1904
rect 7260 1896 7268 1904
rect 7308 1896 7316 1904
rect 7388 1896 7396 1904
rect 7452 1896 7460 1904
rect 7516 1896 7524 1904
rect 172 1876 180 1884
rect 204 1876 212 1884
rect 300 1876 308 1884
rect 332 1876 340 1884
rect 780 1876 788 1884
rect 956 1876 964 1884
rect 1020 1876 1028 1884
rect 1084 1876 1092 1884
rect 1308 1876 1316 1884
rect 1356 1876 1364 1884
rect 1372 1876 1380 1884
rect 1436 1876 1444 1884
rect 460 1856 468 1864
rect 1484 1856 1492 1864
rect 1628 1856 1636 1864
rect 1676 1876 1684 1884
rect 1804 1876 1812 1884
rect 1900 1876 1908 1884
rect 1996 1876 2004 1884
rect 2348 1876 2356 1884
rect 2540 1876 2548 1884
rect 2764 1876 2772 1884
rect 2860 1876 2868 1884
rect 2876 1876 2884 1884
rect 2956 1876 2964 1884
rect 2972 1876 2980 1884
rect 3052 1876 3060 1884
rect 3180 1876 3188 1884
rect 3260 1876 3268 1884
rect 3308 1876 3316 1884
rect 3372 1876 3380 1884
rect 3404 1876 3412 1884
rect 3436 1876 3444 1884
rect 3500 1876 3508 1884
rect 3532 1876 3540 1884
rect 3564 1876 3572 1884
rect 3628 1876 3636 1884
rect 3692 1876 3700 1884
rect 3820 1876 3828 1884
rect 3948 1876 3956 1884
rect 4012 1876 4020 1884
rect 4444 1876 4452 1884
rect 4492 1876 4500 1884
rect 4556 1876 4564 1884
rect 4588 1876 4596 1884
rect 2060 1856 2068 1864
rect 2460 1856 2468 1864
rect 2524 1856 2532 1864
rect 2620 1856 2628 1864
rect 4300 1856 4308 1864
rect 4332 1856 4340 1864
rect 4364 1856 4372 1864
rect 4508 1856 4516 1864
rect 4636 1876 4644 1884
rect 4812 1876 4820 1884
rect 4844 1876 4852 1884
rect 4892 1876 4900 1884
rect 5116 1876 5124 1884
rect 5212 1876 5220 1884
rect 5516 1876 5524 1884
rect 5564 1876 5572 1884
rect 5580 1876 5588 1884
rect 5660 1876 5668 1884
rect 5676 1876 5684 1884
rect 5756 1876 5764 1884
rect 5868 1876 5876 1884
rect 5916 1876 5924 1884
rect 4780 1856 4788 1864
rect 4796 1856 4804 1864
rect 4956 1856 4964 1864
rect 4972 1856 4980 1864
rect 5084 1856 5092 1864
rect 5228 1856 5236 1864
rect 5516 1856 5524 1864
rect 5772 1856 5780 1864
rect 5900 1856 5908 1864
rect 6044 1876 6052 1884
rect 6124 1876 6132 1884
rect 6156 1876 6164 1884
rect 6220 1876 6228 1884
rect 6236 1876 6244 1884
rect 6348 1876 6356 1884
rect 6412 1876 6420 1884
rect 6492 1876 6500 1884
rect 6524 1876 6532 1884
rect 6604 1876 6612 1884
rect 6732 1876 6740 1884
rect 6748 1876 6756 1884
rect 6876 1876 6884 1884
rect 6892 1876 6900 1884
rect 7004 1876 7012 1884
rect 7052 1876 7060 1884
rect 7084 1876 7092 1884
rect 7212 1876 7220 1884
rect 7244 1876 7252 1884
rect 7404 1876 7412 1884
rect 6108 1856 6116 1864
rect 6188 1856 6196 1864
rect 6300 1856 6308 1864
rect 6476 1856 6484 1864
rect 6588 1856 6596 1864
rect 6684 1856 6692 1864
rect 6812 1856 6820 1864
rect 7244 1856 7252 1864
rect 7340 1856 7348 1864
rect 7500 1876 7508 1884
rect 7452 1856 7460 1864
rect 7484 1856 7492 1864
rect 940 1836 948 1844
rect 1244 1836 1252 1844
rect 1388 1836 1396 1844
rect 1548 1836 1556 1844
rect 1708 1836 1716 1844
rect 2188 1836 2196 1844
rect 2236 1836 2244 1844
rect 2748 1836 2756 1844
rect 2812 1836 2820 1844
rect 3484 1836 3492 1844
rect 3740 1836 3748 1844
rect 4156 1836 4164 1844
rect 4252 1836 4260 1844
rect 4316 1836 4324 1844
rect 4524 1836 4532 1844
rect 4572 1836 4580 1844
rect 4652 1836 4660 1844
rect 4812 1836 4820 1844
rect 4860 1836 4868 1844
rect 4988 1836 4996 1844
rect 5404 1836 5412 1844
rect 5564 1836 5572 1844
rect 5580 1836 5588 1844
rect 5596 1836 5604 1844
rect 5628 1836 5636 1844
rect 5660 1836 5668 1844
rect 5724 1836 5732 1844
rect 6124 1836 6132 1844
rect 6172 1836 6180 1844
rect 6572 1836 6580 1844
rect 6636 1836 6644 1844
rect 6876 1836 6884 1844
rect 7004 1836 7012 1844
rect 7116 1836 7124 1844
rect 7228 1836 7236 1844
rect 7356 1836 7364 1844
rect 7468 1836 7476 1844
rect 7548 1836 7556 1844
rect 4956 1816 4964 1824
rect 5084 1816 5092 1824
rect 5228 1816 5236 1824
rect 5516 1816 5524 1824
rect 2243 1806 2251 1814
rect 2253 1806 2261 1814
rect 2263 1806 2271 1814
rect 2273 1806 2281 1814
rect 2283 1806 2291 1814
rect 2293 1806 2301 1814
rect 5251 1806 5259 1814
rect 5261 1806 5269 1814
rect 5271 1806 5279 1814
rect 5281 1806 5289 1814
rect 5291 1806 5299 1814
rect 5301 1806 5309 1814
rect 4940 1796 4948 1804
rect 5340 1796 5348 1804
rect 5852 1796 5860 1804
rect 12 1776 20 1784
rect 396 1776 404 1784
rect 588 1776 596 1784
rect 1516 1776 1524 1784
rect 1644 1776 1652 1784
rect 2412 1776 2420 1784
rect 2460 1776 2468 1784
rect 2668 1776 2676 1784
rect 2796 1776 2804 1784
rect 2892 1776 2900 1784
rect 2956 1776 2964 1784
rect 3180 1776 3188 1784
rect 3228 1776 3236 1784
rect 3324 1776 3332 1784
rect 3692 1776 3700 1784
rect 3740 1776 3748 1784
rect 3900 1776 3908 1784
rect 4044 1776 4052 1784
rect 4140 1776 4148 1784
rect 4300 1776 4308 1784
rect 4412 1776 4420 1784
rect 4540 1776 4548 1784
rect 4604 1776 4612 1784
rect 4700 1776 4708 1784
rect 4732 1776 4740 1784
rect 4764 1776 4772 1784
rect 4796 1776 4804 1784
rect 4812 1776 4820 1784
rect 5148 1776 5156 1784
rect 5628 1776 5636 1784
rect 5644 1776 5652 1784
rect 5916 1776 5924 1784
rect 5964 1776 5972 1784
rect 6188 1776 6196 1784
rect 6268 1776 6276 1784
rect 6284 1776 6292 1784
rect 6460 1776 6468 1784
rect 6556 1776 6564 1784
rect 6876 1776 6884 1784
rect 6988 1776 6996 1784
rect 7020 1776 7028 1784
rect 7116 1776 7124 1784
rect 7532 1776 7540 1784
rect 300 1756 308 1764
rect 460 1756 468 1764
rect 1228 1756 1236 1764
rect 1276 1756 1284 1764
rect 1356 1756 1364 1764
rect 1388 1756 1396 1764
rect 1580 1756 1588 1764
rect 1836 1756 1844 1764
rect 1932 1756 1940 1764
rect 2028 1756 2036 1764
rect 3340 1756 3348 1764
rect 3596 1756 3604 1764
rect 3644 1756 3652 1764
rect 4060 1756 4068 1764
rect 4092 1756 4100 1764
rect 4172 1756 4180 1764
rect 4284 1756 4292 1764
rect 4428 1756 4436 1764
rect 172 1736 180 1744
rect 220 1736 228 1744
rect 236 1736 244 1744
rect 380 1736 388 1744
rect 476 1736 484 1744
rect 572 1736 580 1744
rect 748 1736 756 1744
rect 844 1736 852 1744
rect 972 1736 980 1744
rect 988 1736 996 1744
rect 1116 1736 1124 1744
rect 1260 1736 1268 1744
rect 1420 1736 1428 1744
rect 1484 1736 1492 1744
rect 1500 1736 1508 1744
rect 1564 1736 1572 1744
rect 1628 1736 1636 1744
rect 1692 1736 1700 1744
rect 1852 1736 1860 1744
rect 1916 1736 1924 1744
rect 1980 1736 1988 1744
rect 2044 1736 2052 1744
rect 2172 1736 2180 1744
rect 2316 1736 2324 1744
rect 2444 1736 2452 1744
rect 2620 1736 2628 1744
rect 2652 1736 2660 1744
rect 2764 1736 2772 1744
rect 2908 1736 2916 1744
rect 140 1718 148 1726
rect 204 1716 212 1724
rect 268 1716 276 1724
rect 316 1716 324 1724
rect 364 1716 372 1724
rect 428 1716 436 1724
rect 508 1696 516 1704
rect 540 1716 548 1724
rect 556 1716 564 1724
rect 700 1716 708 1724
rect 812 1716 820 1724
rect 908 1716 916 1724
rect 956 1716 964 1724
rect 1004 1716 1012 1724
rect 1068 1716 1076 1724
rect 1100 1716 1108 1724
rect 1132 1716 1140 1724
rect 1148 1716 1156 1724
rect 1196 1716 1204 1724
rect 1228 1716 1236 1724
rect 1324 1716 1332 1724
rect 1404 1716 1412 1724
rect 1436 1716 1444 1724
rect 1468 1716 1476 1724
rect 1516 1716 1524 1724
rect 1548 1716 1556 1724
rect 1612 1716 1620 1724
rect 1708 1716 1716 1724
rect 1724 1716 1732 1724
rect 1772 1716 1780 1724
rect 1788 1716 1796 1724
rect 1804 1716 1812 1724
rect 1900 1716 1908 1724
rect 1964 1716 1972 1724
rect 1996 1716 2004 1724
rect 2044 1716 2052 1724
rect 2060 1716 2068 1724
rect 2108 1716 2116 1724
rect 2156 1716 2164 1724
rect 2188 1716 2196 1724
rect 2204 1716 2212 1724
rect 2252 1716 2260 1724
rect 2380 1716 2388 1724
rect 2588 1718 2596 1726
rect 2732 1716 2740 1724
rect 2844 1716 2852 1724
rect 2908 1716 2916 1724
rect 3196 1736 3204 1744
rect 3244 1736 3252 1744
rect 3260 1736 3268 1744
rect 3564 1736 3572 1744
rect 3724 1736 3732 1744
rect 3884 1736 3892 1744
rect 3948 1736 3956 1744
rect 4188 1736 4196 1744
rect 4396 1736 4404 1744
rect 4540 1756 4548 1764
rect 4940 1756 4948 1764
rect 4956 1756 4964 1764
rect 5084 1756 5092 1764
rect 5340 1756 5348 1764
rect 5356 1756 5364 1764
rect 5404 1756 5412 1764
rect 5580 1756 5588 1764
rect 5692 1756 5700 1764
rect 5852 1756 5860 1764
rect 6108 1756 6116 1764
rect 6124 1756 6132 1764
rect 6140 1756 6148 1764
rect 6204 1756 6212 1764
rect 6348 1756 6356 1764
rect 6428 1756 6436 1764
rect 6732 1756 6740 1764
rect 6812 1756 6820 1764
rect 6828 1756 6836 1764
rect 6940 1756 6948 1764
rect 6956 1756 6964 1764
rect 7100 1756 7108 1764
rect 7372 1756 7380 1764
rect 7388 1756 7396 1764
rect 7452 1756 7460 1764
rect 7516 1756 7524 1764
rect 7548 1756 7556 1764
rect 4476 1736 4484 1744
rect 4492 1736 4500 1744
rect 4572 1736 4580 1744
rect 4700 1736 4708 1744
rect 4748 1736 4756 1744
rect 4764 1736 4772 1744
rect 4812 1736 4820 1744
rect 4876 1736 4884 1744
rect 5004 1736 5012 1744
rect 5148 1736 5156 1744
rect 5420 1736 5428 1744
rect 5628 1736 5636 1744
rect 5644 1736 5652 1744
rect 5692 1736 5700 1744
rect 5756 1736 5764 1744
rect 5804 1736 5812 1744
rect 5964 1736 5972 1744
rect 6012 1736 6020 1744
rect 6060 1736 6068 1744
rect 6140 1736 6148 1744
rect 6172 1736 6180 1744
rect 6220 1736 6228 1744
rect 6252 1736 6260 1744
rect 6332 1736 6340 1744
rect 6348 1736 6356 1744
rect 6412 1736 6420 1744
rect 6444 1736 6452 1744
rect 6508 1736 6516 1744
rect 6556 1736 6564 1744
rect 6588 1736 6596 1744
rect 6620 1736 6628 1744
rect 6684 1736 6692 1744
rect 6828 1736 6836 1744
rect 6860 1736 6868 1744
rect 6876 1736 6884 1744
rect 6940 1736 6948 1744
rect 6972 1736 6980 1744
rect 7020 1736 7028 1744
rect 7068 1736 7076 1744
rect 7132 1736 7140 1744
rect 7260 1736 7268 1744
rect 7420 1736 7428 1744
rect 3004 1716 3012 1724
rect 3068 1716 3076 1724
rect 3116 1716 3124 1724
rect 3276 1716 3284 1724
rect 3292 1716 3300 1724
rect 3404 1718 3412 1726
rect 3468 1716 3476 1724
rect 3548 1716 3556 1724
rect 3612 1716 3620 1724
rect 3660 1716 3668 1724
rect 3708 1716 3716 1724
rect 3868 1716 3876 1724
rect 3932 1716 3940 1724
rect 4028 1716 4036 1724
rect 4236 1716 4244 1724
rect 4284 1716 4292 1724
rect 4316 1716 4324 1724
rect 4396 1716 4404 1724
rect 892 1696 900 1704
rect 924 1696 932 1704
rect 1036 1696 1044 1704
rect 1340 1696 1348 1704
rect 1580 1696 1588 1704
rect 1644 1696 1652 1704
rect 1932 1696 1940 1704
rect 2092 1696 2100 1704
rect 2156 1696 2164 1704
rect 2396 1696 2404 1704
rect 2412 1696 2420 1704
rect 2748 1696 2756 1704
rect 2860 1696 2868 1704
rect 2876 1696 2884 1704
rect 3020 1696 3028 1704
rect 3084 1696 3092 1704
rect 3212 1696 3220 1704
rect 3308 1696 3316 1704
rect 3820 1696 3828 1704
rect 3900 1696 3908 1704
rect 4588 1716 4596 1724
rect 4668 1696 4676 1704
rect 4716 1696 4724 1704
rect 4796 1696 4804 1704
rect 4844 1696 4852 1704
rect 4892 1716 4900 1724
rect 5004 1716 5012 1724
rect 5020 1716 5028 1724
rect 5052 1716 5060 1724
rect 5228 1716 5236 1724
rect 5372 1716 5380 1724
rect 5436 1716 5444 1724
rect 5500 1716 5508 1724
rect 5548 1716 5556 1724
rect 5564 1716 5572 1724
rect 5820 1716 5828 1724
rect 5884 1716 5892 1724
rect 5020 1696 5028 1704
rect 5116 1696 5124 1704
rect 5164 1696 5172 1704
rect 5196 1696 5204 1704
rect 5436 1696 5444 1704
rect 5468 1696 5476 1704
rect 5484 1696 5492 1704
rect 5596 1696 5604 1704
rect 5676 1696 5684 1704
rect 6092 1716 6100 1724
rect 6124 1716 6132 1724
rect 6188 1716 6196 1724
rect 6204 1716 6212 1724
rect 6268 1716 6276 1724
rect 6284 1716 6292 1724
rect 6348 1716 6356 1724
rect 6364 1716 6372 1724
rect 6428 1716 6436 1724
rect 6492 1716 6500 1724
rect 6556 1716 6564 1724
rect 6572 1716 6580 1724
rect 6636 1716 6644 1724
rect 6812 1716 6820 1724
rect 6876 1716 6884 1724
rect 6892 1716 6900 1724
rect 6956 1716 6964 1724
rect 7004 1716 7012 1724
rect 7084 1716 7092 1724
rect 7164 1716 7172 1724
rect 7292 1716 7300 1724
rect 7340 1716 7348 1724
rect 7484 1716 7492 1724
rect 5932 1696 5940 1704
rect 5980 1696 5988 1704
rect 6028 1696 6036 1704
rect 6476 1696 6484 1704
rect 6508 1696 6516 1704
rect 6652 1696 6660 1704
rect 7004 1696 7012 1704
rect 7276 1696 7284 1704
rect 1084 1676 1092 1684
rect 1868 1676 1876 1684
rect 2364 1676 2372 1684
rect 2716 1676 2724 1684
rect 2828 1676 2836 1684
rect 2988 1676 2996 1684
rect 3052 1676 3060 1684
rect 3132 1676 3140 1684
rect 3500 1676 3508 1684
rect 5132 1676 5140 1684
rect 5244 1676 5252 1684
rect 5388 1676 5396 1684
rect 5516 1676 5524 1684
rect 6412 1676 6420 1684
rect 6620 1676 6628 1684
rect 7068 1676 7076 1684
rect 7196 1676 7204 1684
rect 7308 1676 7316 1684
rect 7340 1676 7348 1684
rect 1468 1656 1476 1664
rect 2380 1656 2388 1664
rect 3068 1656 3076 1664
rect 4988 1656 4996 1664
rect 6700 1656 6708 1664
rect 7292 1656 7300 1664
rect 7388 1656 7396 1664
rect 1180 1636 1188 1644
rect 1756 1636 1764 1644
rect 3532 1636 3540 1644
rect 3596 1636 3604 1644
rect 4220 1636 4228 1644
rect 4684 1636 4692 1644
rect 5180 1636 5188 1644
rect 5228 1636 5236 1644
rect 5500 1636 5508 1644
rect 5612 1636 5620 1644
rect 5660 1636 5668 1644
rect 5772 1636 5780 1644
rect 5996 1636 6004 1644
rect 6220 1636 6228 1644
rect 6332 1636 6340 1644
rect 7532 1636 7540 1644
rect 739 1606 747 1614
rect 749 1606 757 1614
rect 759 1606 767 1614
rect 769 1606 777 1614
rect 779 1606 787 1614
rect 789 1606 797 1614
rect 3747 1606 3755 1614
rect 3757 1606 3765 1614
rect 3767 1606 3775 1614
rect 3777 1606 3785 1614
rect 3787 1606 3795 1614
rect 3797 1606 3805 1614
rect 6755 1606 6763 1614
rect 6765 1606 6773 1614
rect 6775 1606 6783 1614
rect 6785 1606 6793 1614
rect 6795 1606 6803 1614
rect 6805 1606 6813 1614
rect 1052 1576 1060 1584
rect 1148 1576 1156 1584
rect 1308 1576 1316 1584
rect 1836 1576 1844 1584
rect 1868 1576 1876 1584
rect 1916 1576 1924 1584
rect 2076 1576 2084 1584
rect 2108 1576 2116 1584
rect 2140 1576 2148 1584
rect 2300 1576 2308 1584
rect 2476 1576 2484 1584
rect 2572 1576 2580 1584
rect 2684 1576 2692 1584
rect 2732 1576 2740 1584
rect 2908 1576 2916 1584
rect 3148 1576 3156 1584
rect 3660 1576 3668 1584
rect 3724 1576 3732 1584
rect 3852 1576 3860 1584
rect 4108 1576 4116 1584
rect 4156 1576 4164 1584
rect 4284 1576 4292 1584
rect 4732 1576 4740 1584
rect 4924 1576 4932 1584
rect 6188 1576 6196 1584
rect 7388 1576 7396 1584
rect 7484 1576 7492 1584
rect 2524 1556 2532 1564
rect 3036 1556 3044 1564
rect 412 1536 420 1544
rect 1004 1536 1012 1544
rect 1996 1536 2004 1544
rect 2060 1536 2068 1544
rect 2156 1536 2164 1544
rect 2172 1536 2180 1544
rect 220 1516 228 1524
rect 44 1496 52 1504
rect 140 1496 148 1504
rect 300 1496 308 1504
rect 332 1496 340 1504
rect 428 1496 436 1504
rect 492 1496 500 1504
rect 540 1496 548 1504
rect 604 1496 612 1504
rect 652 1496 660 1504
rect 716 1496 724 1504
rect 908 1496 916 1504
rect 1020 1496 1028 1504
rect 1036 1496 1044 1504
rect 1084 1496 1092 1504
rect 1116 1496 1124 1504
rect 1132 1496 1140 1504
rect 1180 1496 1188 1504
rect 1244 1496 1252 1504
rect 1260 1496 1268 1504
rect 1276 1496 1284 1504
rect 1340 1496 1348 1504
rect 1356 1496 1364 1504
rect 1372 1496 1380 1504
rect 1436 1496 1444 1504
rect 1548 1516 1556 1524
rect 2028 1516 2036 1524
rect 2092 1516 2100 1524
rect 2188 1516 2196 1524
rect 2236 1536 2244 1544
rect 2380 1536 2388 1544
rect 2428 1536 2436 1544
rect 2444 1536 2452 1544
rect 2508 1536 2516 1544
rect 2668 1536 2676 1544
rect 2956 1536 2964 1544
rect 3020 1536 3028 1544
rect 3276 1536 3284 1544
rect 4124 1536 4132 1544
rect 4508 1536 4516 1544
rect 4748 1536 4756 1544
rect 5372 1536 5380 1544
rect 5404 1536 5412 1544
rect 6236 1536 6244 1544
rect 6908 1536 6916 1544
rect 7212 1536 7220 1544
rect 2428 1516 2436 1524
rect 2540 1516 2548 1524
rect 2556 1516 2564 1524
rect 2620 1516 2628 1524
rect 2700 1516 2708 1524
rect 2764 1516 2772 1524
rect 2876 1516 2884 1524
rect 2924 1516 2932 1524
rect 2988 1516 2996 1524
rect 3052 1516 3060 1524
rect 3084 1516 3092 1524
rect 3116 1516 3124 1524
rect 3132 1516 3140 1524
rect 3244 1516 3252 1524
rect 3676 1516 3684 1524
rect 3804 1516 3812 1524
rect 3980 1514 3988 1522
rect 4108 1516 4116 1524
rect 4364 1516 4372 1524
rect 4620 1516 4628 1524
rect 4700 1516 4708 1524
rect 4972 1516 4980 1524
rect 5116 1516 5124 1524
rect 5260 1516 5268 1524
rect 5420 1516 5428 1524
rect 5500 1516 5508 1524
rect 5564 1516 5572 1524
rect 5660 1516 5668 1524
rect 5692 1516 5700 1524
rect 6140 1516 6148 1524
rect 6316 1516 6324 1524
rect 6332 1516 6340 1524
rect 6396 1516 6404 1524
rect 6460 1516 6468 1524
rect 6700 1516 6708 1524
rect 6732 1516 6740 1524
rect 7132 1516 7140 1524
rect 7468 1516 7476 1524
rect 1516 1496 1524 1504
rect 1660 1496 1668 1504
rect 1756 1496 1764 1504
rect 1804 1496 1812 1504
rect 2044 1496 2052 1504
rect 2172 1496 2180 1504
rect 2220 1496 2228 1504
rect 2380 1496 2388 1504
rect 2444 1496 2452 1504
rect 2524 1496 2532 1504
rect 2684 1496 2692 1504
rect 2844 1496 2852 1504
rect 2860 1496 2868 1504
rect 2956 1496 2964 1504
rect 3036 1496 3044 1504
rect 3084 1496 3092 1504
rect 3212 1496 3220 1504
rect 3356 1496 3364 1504
rect 3468 1496 3476 1504
rect 3500 1496 3508 1504
rect 3596 1496 3604 1504
rect 3724 1496 3732 1504
rect 3868 1496 3876 1504
rect 4028 1496 4036 1504
rect 4108 1496 4116 1504
rect 4172 1496 4180 1504
rect 4188 1496 4196 1504
rect 4252 1496 4260 1504
rect 4300 1496 4308 1504
rect 4396 1496 4404 1504
rect 4476 1496 4484 1504
rect 4508 1496 4516 1504
rect 4572 1496 4580 1504
rect 4620 1496 4628 1504
rect 4652 1496 4660 1504
rect 4732 1496 4740 1504
rect 4796 1496 4804 1504
rect 4876 1496 4884 1504
rect 4924 1496 4932 1504
rect 5036 1496 5044 1504
rect 5116 1496 5124 1504
rect 5148 1496 5156 1504
rect 5228 1496 5236 1504
rect 5372 1496 5380 1504
rect 5420 1496 5428 1504
rect 5500 1496 5508 1504
rect 5532 1496 5540 1504
rect 5596 1496 5604 1504
rect 5708 1496 5716 1504
rect 5836 1496 5844 1504
rect 5916 1496 5924 1504
rect 5948 1496 5956 1504
rect 6092 1496 6100 1504
rect 6124 1496 6132 1504
rect 6236 1496 6244 1504
rect 6332 1496 6340 1504
rect 6380 1496 6388 1504
rect 6444 1496 6452 1504
rect 6508 1496 6516 1504
rect 6572 1496 6580 1504
rect 6652 1496 6660 1504
rect 6716 1496 6724 1504
rect 6860 1496 6868 1504
rect 6924 1496 6932 1504
rect 6940 1496 6948 1504
rect 6972 1496 6980 1504
rect 7004 1496 7012 1504
rect 108 1476 116 1484
rect 124 1476 132 1484
rect 188 1476 196 1484
rect 444 1476 452 1484
rect 524 1476 532 1484
rect 668 1476 676 1484
rect 700 1476 708 1484
rect 892 1476 900 1484
rect 1196 1476 1204 1484
rect 1420 1476 1428 1484
rect 1452 1476 1460 1484
rect 1500 1476 1508 1484
rect 1676 1476 1684 1484
rect 1884 1476 1892 1484
rect 1932 1476 1940 1484
rect 2124 1476 2132 1484
rect 2588 1476 2596 1484
rect 2636 1476 2644 1484
rect 2748 1476 2756 1484
rect 2764 1476 2772 1484
rect 2828 1476 2836 1484
rect 2892 1476 2900 1484
rect 2940 1476 2948 1484
rect 3068 1476 3076 1484
rect 3164 1476 3172 1484
rect 3244 1476 3252 1484
rect 3324 1476 3332 1484
rect 3644 1476 3652 1484
rect 3868 1476 3876 1484
rect 3884 1476 3892 1484
rect 3948 1476 3956 1484
rect 4044 1476 4052 1484
rect 4300 1476 4308 1484
rect 4412 1476 4420 1484
rect 4780 1476 4788 1484
rect 5164 1476 5172 1484
rect 5548 1476 5556 1484
rect 5740 1476 5748 1484
rect 5820 1476 5828 1484
rect 5948 1476 5956 1484
rect 6012 1476 6020 1484
rect 6060 1476 6068 1484
rect 6108 1476 6116 1484
rect 6172 1476 6180 1484
rect 6284 1476 6292 1484
rect 6300 1476 6308 1484
rect 6364 1476 6372 1484
rect 6396 1476 6404 1484
rect 6444 1476 6452 1484
rect 6492 1476 6500 1484
rect 6524 1476 6532 1484
rect 6572 1476 6580 1484
rect 6636 1476 6644 1484
rect 6668 1476 6676 1484
rect 6732 1476 6740 1484
rect 6780 1476 6788 1484
rect 6860 1476 6868 1484
rect 6908 1476 6916 1484
rect 12 1456 20 1464
rect 284 1456 292 1464
rect 524 1456 532 1464
rect 572 1456 580 1464
rect 636 1456 644 1464
rect 748 1456 756 1464
rect 1212 1456 1220 1464
rect 1484 1456 1492 1464
rect 1788 1456 1796 1464
rect 1948 1456 1956 1464
rect 2012 1456 2020 1464
rect 2332 1456 2340 1464
rect 3180 1456 3188 1464
rect 3276 1456 3284 1464
rect 3340 1456 3348 1464
rect 3692 1456 3700 1464
rect 3740 1456 3748 1464
rect 3964 1456 3972 1464
rect 4012 1456 4020 1464
rect 4140 1456 4148 1464
rect 4220 1456 4228 1464
rect 4428 1456 4436 1464
rect 4540 1456 4548 1464
rect 4844 1456 4852 1464
rect 4972 1456 4980 1464
rect 5068 1456 5076 1464
rect 5084 1456 5092 1464
rect 5180 1456 5188 1464
rect 5628 1456 5636 1464
rect 5740 1456 5748 1464
rect 5772 1456 5780 1464
rect 5788 1456 5796 1464
rect 5980 1456 5988 1464
rect 5996 1456 6004 1464
rect 6236 1456 6244 1464
rect 6268 1456 6276 1464
rect 6380 1456 6388 1464
rect 6508 1456 6516 1464
rect 6524 1456 6532 1464
rect 6636 1456 6644 1464
rect 6652 1456 6660 1464
rect 6988 1476 6996 1484
rect 7020 1476 7028 1484
rect 7116 1476 7124 1484
rect 7180 1496 7188 1504
rect 7292 1496 7300 1504
rect 7516 1496 7524 1504
rect 7180 1476 7188 1484
rect 7292 1476 7300 1484
rect 7356 1476 7364 1484
rect 7468 1476 7476 1484
rect 7500 1476 7508 1484
rect 7564 1476 7572 1484
rect 7340 1456 7348 1464
rect 76 1436 84 1444
rect 172 1436 180 1444
rect 460 1436 468 1444
rect 1548 1436 1556 1444
rect 1564 1436 1572 1444
rect 1772 1436 1780 1444
rect 1836 1436 1844 1444
rect 3292 1436 3300 1444
rect 3388 1436 3396 1444
rect 3580 1436 3588 1444
rect 3628 1436 3636 1444
rect 4332 1436 4340 1444
rect 4828 1436 4836 1444
rect 4988 1436 4996 1444
rect 5116 1436 5124 1444
rect 5388 1436 5396 1444
rect 5564 1436 5572 1444
rect 5964 1436 5972 1444
rect 6444 1436 6452 1444
rect 6460 1436 6468 1444
rect 6572 1436 6580 1444
rect 6684 1436 6692 1444
rect 6780 1436 6788 1444
rect 6860 1436 6868 1444
rect 7052 1436 7060 1444
rect 7132 1436 7140 1444
rect 7324 1436 7332 1444
rect 4428 1416 4436 1424
rect 4972 1416 4980 1424
rect 5068 1416 5076 1424
rect 5180 1416 5188 1424
rect 5628 1416 5636 1424
rect 5740 1416 5748 1424
rect 2243 1406 2251 1414
rect 2253 1406 2261 1414
rect 2263 1406 2271 1414
rect 2273 1406 2281 1414
rect 2283 1406 2291 1414
rect 2293 1406 2301 1414
rect 5251 1406 5259 1414
rect 5261 1406 5269 1414
rect 5271 1406 5279 1414
rect 5281 1406 5289 1414
rect 5291 1406 5299 1414
rect 5301 1406 5309 1414
rect 5084 1396 5092 1404
rect 5212 1396 5220 1404
rect 5580 1396 5588 1404
rect 5676 1396 5684 1404
rect 5804 1396 5812 1404
rect 12 1376 20 1384
rect 380 1376 388 1384
rect 572 1376 580 1384
rect 1020 1376 1028 1384
rect 1068 1376 1076 1384
rect 1452 1376 1460 1384
rect 1724 1376 1732 1384
rect 1948 1376 1956 1384
rect 2140 1376 2148 1384
rect 2380 1376 2388 1384
rect 2652 1376 2660 1384
rect 2700 1376 2708 1384
rect 2764 1376 2772 1384
rect 2844 1376 2852 1384
rect 2908 1376 2916 1384
rect 2956 1376 2964 1384
rect 3052 1376 3060 1384
rect 3164 1376 3172 1384
rect 3196 1376 3204 1384
rect 3260 1376 3268 1384
rect 3884 1376 3892 1384
rect 4172 1376 4180 1384
rect 4268 1376 4276 1384
rect 4284 1376 4292 1384
rect 4540 1376 4548 1384
rect 4684 1376 4692 1384
rect 4764 1376 4772 1384
rect 4972 1376 4980 1384
rect 5180 1376 5188 1384
rect 5500 1376 5508 1384
rect 5708 1376 5716 1384
rect 5836 1376 5844 1384
rect 5932 1376 5940 1384
rect 6076 1376 6084 1384
rect 6220 1376 6228 1384
rect 6428 1376 6436 1384
rect 6732 1376 6740 1384
rect 6956 1376 6964 1384
rect 7052 1376 7060 1384
rect 7116 1376 7124 1384
rect 892 1356 900 1364
rect 1132 1356 1140 1364
rect 1228 1356 1236 1364
rect 1740 1356 1748 1364
rect 2540 1356 2548 1364
rect 3564 1356 3572 1364
rect 3596 1356 3604 1364
rect 3628 1356 3636 1364
rect 4092 1356 4100 1364
rect 4188 1356 4196 1364
rect 4316 1356 4324 1364
rect 4444 1356 4452 1364
rect 4700 1356 4708 1364
rect 4860 1356 4868 1364
rect 124 1336 132 1344
rect 220 1336 228 1344
rect 284 1336 292 1344
rect 412 1336 420 1344
rect 476 1336 484 1344
rect 908 1336 916 1344
rect 1052 1336 1060 1344
rect 1148 1336 1156 1344
rect 1212 1336 1220 1344
rect 1276 1336 1284 1344
rect 1340 1336 1348 1344
rect 1404 1336 1412 1344
rect 1468 1336 1476 1344
rect 1532 1336 1540 1344
rect 1612 1336 1620 1344
rect 1644 1336 1652 1344
rect 1756 1336 1764 1344
rect 1820 1336 1828 1344
rect 1964 1336 1972 1344
rect 1980 1336 1988 1344
rect 2284 1336 2292 1344
rect 2364 1336 2372 1344
rect 2620 1336 2628 1344
rect 2684 1336 2692 1344
rect 2732 1336 2740 1344
rect 2876 1336 2884 1344
rect 2924 1336 2932 1344
rect 3132 1336 3140 1344
rect 3244 1336 3252 1344
rect 3276 1336 3284 1344
rect 3292 1336 3300 1344
rect 3356 1336 3364 1344
rect 3420 1336 3428 1344
rect 3484 1336 3492 1344
rect 3644 1336 3652 1344
rect 3916 1336 3924 1344
rect 4124 1336 4132 1344
rect 4156 1336 4164 1344
rect 4364 1336 4372 1344
rect 4428 1336 4436 1344
rect 4460 1336 4468 1344
rect 4524 1336 4532 1344
rect 4556 1336 4564 1344
rect 4588 1336 4596 1344
rect 4844 1336 4852 1344
rect 4908 1356 4916 1364
rect 4956 1356 4964 1364
rect 5084 1356 5092 1364
rect 5196 1356 5204 1364
rect 5212 1356 5220 1364
rect 5484 1356 5492 1364
rect 5580 1356 5588 1364
rect 5676 1356 5684 1364
rect 5692 1356 5700 1364
rect 5804 1356 5812 1364
rect 6012 1356 6020 1364
rect 6124 1356 6132 1364
rect 6284 1356 6292 1364
rect 6524 1356 6532 1364
rect 5100 1336 5108 1344
rect 5372 1336 5380 1344
rect 5452 1336 5460 1344
rect 5900 1336 5908 1344
rect 5932 1336 5940 1344
rect 5996 1336 6004 1344
rect 6028 1336 6036 1344
rect 6204 1336 6212 1344
rect 6332 1336 6340 1344
rect 6412 1336 6420 1344
rect 6444 1336 6452 1344
rect 6508 1336 6516 1344
rect 6652 1356 6660 1364
rect 6684 1356 6692 1364
rect 6876 1356 6884 1364
rect 6972 1356 6980 1364
rect 7068 1356 7076 1364
rect 7244 1356 7252 1364
rect 7324 1356 7332 1364
rect 7340 1356 7348 1364
rect 6556 1336 6564 1344
rect 6604 1336 6612 1344
rect 6908 1336 6916 1344
rect 92 1316 100 1324
rect 252 1318 260 1326
rect 460 1316 468 1324
rect 604 1316 612 1324
rect 652 1316 660 1324
rect 668 1316 676 1324
rect 684 1316 692 1324
rect 748 1316 756 1324
rect 812 1316 820 1324
rect 892 1318 900 1326
rect 1036 1316 1044 1324
rect 1100 1316 1108 1324
rect 1164 1316 1172 1324
rect 1260 1316 1268 1324
rect 1276 1316 1284 1324
rect 1324 1316 1332 1324
rect 1388 1316 1396 1324
rect 1420 1316 1428 1324
rect 1484 1316 1492 1324
rect 1516 1316 1524 1324
rect 1548 1316 1556 1324
rect 1564 1316 1572 1324
rect 1612 1316 1620 1324
rect 1660 1316 1668 1324
rect 1708 1316 1716 1324
rect 1772 1316 1780 1324
rect 1804 1316 1812 1324
rect 1836 1316 1844 1324
rect 1852 1316 1860 1324
rect 1900 1316 1908 1324
rect 2156 1316 2164 1324
rect 2220 1316 2228 1324
rect 2332 1316 2340 1324
rect 2444 1316 2452 1324
rect 2508 1316 2516 1324
rect 2812 1316 2820 1324
rect 3020 1316 3028 1324
rect 3308 1316 3316 1324
rect 3372 1316 3380 1324
rect 3436 1316 3444 1324
rect 3468 1316 3476 1324
rect 3532 1316 3540 1324
rect 3580 1316 3588 1324
rect 3772 1316 3780 1324
rect 3836 1316 3844 1324
rect 3948 1318 3956 1326
rect 4012 1316 4020 1324
rect 4220 1316 4228 1324
rect 4332 1316 4340 1324
rect 4428 1316 4436 1324
rect 4572 1316 4580 1324
rect 4604 1316 4612 1324
rect 4636 1316 4644 1324
rect 4652 1316 4660 1324
rect 4732 1316 4740 1324
rect 4828 1316 4836 1324
rect 4860 1316 4868 1324
rect 4940 1316 4948 1324
rect 5036 1316 5044 1324
rect 5116 1316 5124 1324
rect 5164 1316 5172 1324
rect 5324 1316 5332 1324
rect 5356 1316 5364 1324
rect 5404 1316 5412 1324
rect 5452 1316 5460 1324
rect 5532 1316 5540 1324
rect 5580 1316 5588 1324
rect 5628 1316 5636 1324
rect 5772 1316 5780 1324
rect 5868 1316 5876 1324
rect 5884 1316 5892 1324
rect 6044 1316 6052 1324
rect 6092 1316 6100 1324
rect 6124 1316 6132 1324
rect 6156 1316 6164 1324
rect 6188 1316 6196 1324
rect 6220 1316 6228 1324
rect 6252 1316 6260 1324
rect 6316 1316 6324 1324
rect 6348 1316 6356 1324
rect 6652 1316 6660 1324
rect 7004 1316 7012 1324
rect 7036 1336 7044 1344
rect 7084 1336 7092 1344
rect 7132 1336 7140 1344
rect 7164 1336 7172 1344
rect 7228 1336 7236 1344
rect 7404 1336 7412 1344
rect 7436 1356 7444 1364
rect 7484 1356 7492 1364
rect 7148 1316 7156 1324
rect 7180 1316 7188 1324
rect 7292 1316 7300 1324
rect 7308 1316 7316 1324
rect 7340 1316 7348 1324
rect 7388 1316 7396 1324
rect 7452 1316 7460 1324
rect 7500 1316 7508 1324
rect 716 1296 724 1304
rect 1452 1296 1460 1304
rect 1516 1296 1524 1304
rect 1660 1296 1668 1304
rect 1692 1296 1700 1304
rect 2172 1296 2180 1304
rect 2188 1296 2196 1304
rect 2348 1296 2356 1304
rect 2460 1296 2468 1304
rect 2524 1296 2532 1304
rect 2540 1296 2548 1304
rect 2828 1296 2836 1304
rect 2844 1296 2852 1304
rect 3036 1296 3044 1304
rect 3052 1296 3060 1304
rect 3244 1296 3252 1304
rect 3340 1296 3348 1304
rect 3404 1296 3412 1304
rect 3436 1296 3444 1304
rect 3468 1296 3476 1304
rect 3500 1296 3508 1304
rect 3532 1296 3540 1304
rect 3596 1296 3604 1304
rect 4124 1296 4132 1304
rect 4156 1296 4164 1304
rect 4332 1296 4340 1304
rect 4380 1296 4388 1304
rect 5004 1296 5012 1304
rect 5148 1296 5156 1304
rect 5324 1296 5332 1304
rect 5388 1296 5396 1304
rect 5500 1296 5508 1304
rect 5580 1296 5588 1304
rect 5740 1296 5748 1304
rect 6588 1296 6596 1304
rect 6636 1296 6644 1304
rect 6668 1296 6676 1304
rect 6956 1296 6964 1304
rect 7116 1296 7124 1304
rect 7180 1296 7188 1304
rect 7196 1296 7204 1304
rect 636 1276 644 1284
rect 1356 1276 1364 1284
rect 2140 1276 2148 1284
rect 2316 1276 2324 1284
rect 2428 1276 2436 1284
rect 2492 1276 2500 1284
rect 2588 1276 2596 1284
rect 2668 1276 2676 1284
rect 2732 1276 2740 1284
rect 2764 1276 2772 1284
rect 2796 1276 2804 1284
rect 2876 1276 2884 1284
rect 2972 1276 2980 1284
rect 3004 1276 3012 1284
rect 3100 1276 3108 1284
rect 3180 1276 3188 1284
rect 3196 1276 3204 1284
rect 3372 1276 3380 1284
rect 5420 1276 5428 1284
rect 7228 1276 7236 1284
rect 7564 1276 7572 1284
rect 1324 1256 1332 1264
rect 1804 1256 1812 1264
rect 2508 1256 2516 1264
rect 2812 1256 2820 1264
rect 3020 1256 3028 1264
rect 3308 1256 3316 1264
rect 4412 1256 4420 1264
rect 1196 1236 1204 1244
rect 1884 1236 1892 1244
rect 2092 1236 2100 1244
rect 2332 1236 2340 1244
rect 3884 1236 3892 1244
rect 4076 1236 4084 1244
rect 5436 1236 5444 1244
rect 5836 1236 5844 1244
rect 6892 1236 6900 1244
rect 7468 1236 7476 1244
rect 739 1206 747 1214
rect 749 1206 757 1214
rect 759 1206 767 1214
rect 769 1206 777 1214
rect 779 1206 787 1214
rect 789 1206 797 1214
rect 3747 1206 3755 1214
rect 3757 1206 3765 1214
rect 3767 1206 3775 1214
rect 3777 1206 3785 1214
rect 3787 1206 3795 1214
rect 3797 1206 3805 1214
rect 6755 1206 6763 1214
rect 6765 1206 6773 1214
rect 6775 1206 6783 1214
rect 6785 1206 6793 1214
rect 6795 1206 6803 1214
rect 6805 1206 6813 1214
rect 124 1176 132 1184
rect 364 1176 372 1184
rect 380 1176 388 1184
rect 652 1176 660 1184
rect 1180 1176 1188 1184
rect 1468 1176 1476 1184
rect 1916 1176 1924 1184
rect 2028 1176 2036 1184
rect 2156 1176 2164 1184
rect 2268 1176 2276 1184
rect 2396 1176 2404 1184
rect 2460 1176 2468 1184
rect 2524 1176 2532 1184
rect 2572 1176 2580 1184
rect 2668 1176 2676 1184
rect 2716 1176 2724 1184
rect 2732 1176 2740 1184
rect 2876 1176 2884 1184
rect 2924 1176 2932 1184
rect 3116 1176 3124 1184
rect 3196 1176 3204 1184
rect 4988 1176 4996 1184
rect 5052 1176 5060 1184
rect 5340 1176 5348 1184
rect 5660 1176 5668 1184
rect 6428 1176 6436 1184
rect 6796 1176 6804 1184
rect 7052 1176 7060 1184
rect 780 1136 788 1144
rect 972 1136 980 1144
rect 1724 1136 1732 1144
rect 2012 1136 2020 1144
rect 2076 1136 2084 1144
rect 2124 1136 2132 1144
rect 2140 1136 2148 1144
rect 2204 1136 2212 1144
rect 2364 1136 2372 1144
rect 2444 1136 2452 1144
rect 2508 1136 2516 1144
rect 4252 1136 4260 1144
rect 4812 1136 4820 1144
rect 5196 1136 5204 1144
rect 5500 1136 5508 1144
rect 6252 1136 6260 1144
rect 6316 1136 6324 1144
rect 6332 1136 6340 1144
rect 6588 1136 6596 1144
rect 7004 1136 7012 1144
rect 636 1116 644 1124
rect 1148 1116 1156 1124
rect 1212 1116 1220 1124
rect 1980 1116 1988 1124
rect 2044 1116 2052 1124
rect 2108 1116 2116 1124
rect 2172 1116 2180 1124
rect 2332 1116 2340 1124
rect 2348 1116 2356 1124
rect 2412 1116 2420 1124
rect 2476 1116 2484 1124
rect 2620 1116 2628 1124
rect 2828 1116 2836 1124
rect 3036 1116 3044 1124
rect 3276 1116 3284 1124
rect 3308 1116 3316 1124
rect 3500 1116 3508 1124
rect 3516 1116 3524 1124
rect 3692 1116 3700 1124
rect 3868 1116 3876 1124
rect 3932 1116 3940 1124
rect 3980 1116 3988 1124
rect 3996 1116 4004 1124
rect 4108 1116 4116 1124
rect 4204 1116 4212 1124
rect 4300 1116 4308 1124
rect 4380 1116 4388 1124
rect 5036 1116 5044 1124
rect 5468 1116 5476 1124
rect 5788 1116 5796 1124
rect 5868 1116 5876 1124
rect 6044 1116 6052 1124
rect 6348 1116 6356 1124
rect 6476 1116 6484 1124
rect 6620 1116 6628 1124
rect 6908 1116 6916 1124
rect 6972 1116 6980 1124
rect 7084 1116 7092 1124
rect 220 1096 228 1104
rect 284 1094 292 1102
rect 492 1096 500 1104
rect 684 1096 692 1104
rect 860 1096 868 1104
rect 908 1096 916 1104
rect 988 1096 996 1104
rect 1052 1096 1060 1104
rect 1116 1096 1124 1104
rect 1164 1096 1172 1104
rect 1180 1096 1188 1104
rect 1276 1094 1284 1102
rect 1340 1096 1348 1104
rect 1420 1096 1428 1104
rect 1436 1096 1444 1104
rect 1500 1096 1508 1104
rect 1548 1096 1556 1104
rect 1612 1096 1620 1104
rect 1628 1096 1636 1104
rect 1644 1096 1652 1104
rect 1708 1096 1716 1104
rect 1836 1096 1844 1104
rect 1964 1096 1972 1104
rect 1996 1096 2004 1104
rect 2060 1096 2068 1104
rect 2124 1096 2132 1104
rect 2188 1096 2196 1104
rect 2236 1096 2244 1104
rect 2364 1096 2372 1104
rect 2428 1096 2436 1104
rect 2492 1096 2500 1104
rect 2540 1096 2548 1104
rect 2636 1096 2644 1104
rect 2684 1096 2692 1104
rect 2764 1096 2772 1104
rect 3004 1096 3012 1104
rect 3020 1096 3028 1104
rect 3196 1096 3204 1104
rect 3356 1096 3364 1104
rect 3420 1096 3428 1104
rect 3612 1096 3620 1104
rect 3724 1096 3732 1104
rect 3772 1096 3780 1104
rect 3820 1096 3828 1104
rect 3900 1096 3908 1104
rect 4044 1096 4052 1104
rect 4140 1096 4148 1104
rect 4220 1096 4228 1104
rect 4316 1096 4324 1104
rect 4380 1096 4388 1104
rect 4428 1096 4436 1104
rect 4492 1094 4500 1102
rect 4684 1094 4692 1102
rect 4860 1096 4868 1104
rect 4876 1096 4884 1104
rect 5132 1096 5140 1104
rect 5244 1096 5252 1104
rect 5452 1096 5460 1104
rect 12 1076 20 1084
rect 476 1076 484 1084
rect 604 1076 612 1084
rect 636 1076 644 1084
rect 1004 1076 1012 1084
rect 348 1056 356 1064
rect 396 1056 404 1064
rect 700 1056 708 1064
rect 844 1056 852 1064
rect 1020 1056 1028 1064
rect 1100 1076 1108 1084
rect 1164 1076 1172 1084
rect 1244 1076 1252 1084
rect 1596 1076 1604 1084
rect 1692 1076 1700 1084
rect 1852 1076 1860 1084
rect 2300 1076 2308 1084
rect 2604 1076 2612 1084
rect 2780 1076 2788 1084
rect 2828 1076 2836 1084
rect 2844 1080 2852 1088
rect 3084 1080 3092 1088
rect 3164 1076 3172 1084
rect 3276 1076 3284 1084
rect 3308 1076 3316 1084
rect 3388 1076 3396 1084
rect 3404 1076 3412 1084
rect 3468 1076 3476 1084
rect 3548 1076 3556 1084
rect 3596 1076 3604 1084
rect 3660 1076 3668 1084
rect 3708 1076 3716 1084
rect 3820 1076 3828 1084
rect 3884 1076 3892 1084
rect 3948 1076 3956 1084
rect 3980 1076 3988 1084
rect 4028 1076 4036 1084
rect 4060 1076 4068 1084
rect 4092 1076 4100 1084
rect 4156 1076 4164 1084
rect 4172 1076 4180 1084
rect 4268 1076 4276 1084
rect 4332 1076 4340 1084
rect 4428 1076 4436 1084
rect 4508 1076 4516 1084
rect 4652 1076 4660 1084
rect 4748 1076 4756 1084
rect 4828 1076 4836 1084
rect 4924 1076 4932 1084
rect 5020 1076 5028 1084
rect 5068 1076 5076 1084
rect 5084 1076 5092 1084
rect 5292 1076 5300 1084
rect 5420 1076 5428 1084
rect 5468 1076 5476 1084
rect 5612 1096 5620 1104
rect 5884 1096 5892 1104
rect 6156 1096 6164 1104
rect 6204 1096 6212 1104
rect 6220 1096 6228 1104
rect 6268 1096 6276 1104
rect 6460 1096 6468 1104
rect 6508 1096 6516 1104
rect 6572 1096 6580 1104
rect 6636 1096 6644 1104
rect 6684 1096 6692 1104
rect 6748 1096 6756 1104
rect 6844 1096 6852 1104
rect 6892 1096 6900 1104
rect 6988 1096 6996 1104
rect 7100 1096 7108 1104
rect 7116 1096 7124 1104
rect 7148 1096 7156 1104
rect 7196 1096 7204 1104
rect 7244 1096 7252 1104
rect 7292 1096 7300 1104
rect 7484 1096 7492 1104
rect 7548 1096 7556 1104
rect 5516 1076 5524 1084
rect 5612 1076 5620 1084
rect 5772 1076 5780 1084
rect 5836 1076 5844 1084
rect 5932 1076 5940 1084
rect 6012 1076 6020 1084
rect 6108 1076 6116 1084
rect 6124 1076 6132 1084
rect 6364 1076 6372 1084
rect 6460 1076 6468 1084
rect 6620 1076 6628 1084
rect 6700 1076 6708 1084
rect 6940 1076 6948 1084
rect 7132 1076 7140 1084
rect 7180 1076 7188 1084
rect 1516 1056 1524 1064
rect 1932 1056 1940 1064
rect 1964 1056 1972 1064
rect 2796 1056 2804 1064
rect 2892 1056 2900 1064
rect 3052 1056 3060 1064
rect 3132 1056 3140 1064
rect 3164 1056 3172 1064
rect 3196 1056 3204 1064
rect 3244 1056 3252 1064
rect 3372 1056 3380 1064
rect 5420 1056 5428 1064
rect 6540 1056 6548 1064
rect 6668 1056 6676 1064
rect 6732 1056 6740 1064
rect 6812 1056 6820 1064
rect 6844 1056 6852 1064
rect 6956 1056 6964 1064
rect 7068 1056 7076 1064
rect 7228 1056 7236 1064
rect 7276 1056 7284 1064
rect 7292 1056 7300 1064
rect 7372 1076 7380 1084
rect 7468 1076 7476 1084
rect 7516 1056 7524 1064
rect 156 1036 164 1044
rect 588 1036 596 1044
rect 620 1036 628 1044
rect 1404 1036 1412 1044
rect 1580 1036 1588 1044
rect 2876 1036 2884 1044
rect 2972 1036 2980 1044
rect 3116 1036 3124 1044
rect 3228 1036 3236 1044
rect 3308 1036 3316 1044
rect 3452 1036 3460 1044
rect 3532 1036 3540 1044
rect 3580 1036 3588 1044
rect 3676 1036 3684 1044
rect 3756 1036 3764 1044
rect 3932 1036 3940 1044
rect 3980 1036 3988 1044
rect 4204 1036 4212 1044
rect 4300 1036 4308 1044
rect 4620 1036 4628 1044
rect 5708 1036 5716 1044
rect 5804 1036 5812 1044
rect 5852 1036 5860 1044
rect 5964 1036 5972 1044
rect 6172 1036 6180 1044
rect 7340 1036 7348 1044
rect 7404 1036 7412 1044
rect 2243 1006 2251 1014
rect 2253 1006 2261 1014
rect 2263 1006 2271 1014
rect 2273 1006 2281 1014
rect 2283 1006 2291 1014
rect 2293 1006 2301 1014
rect 5251 1006 5259 1014
rect 5261 1006 5269 1014
rect 5271 1006 5279 1014
rect 5281 1006 5289 1014
rect 5291 1006 5299 1014
rect 5301 1006 5309 1014
rect 444 976 452 984
rect 492 976 500 984
rect 940 976 948 984
rect 956 976 964 984
rect 1276 976 1284 984
rect 1708 976 1716 984
rect 1948 976 1956 984
rect 2060 976 2068 984
rect 2140 976 2148 984
rect 2172 976 2180 984
rect 2412 976 2420 984
rect 2444 976 2452 984
rect 2620 976 2628 984
rect 2684 976 2692 984
rect 2732 976 2740 984
rect 2892 976 2900 984
rect 3372 976 3380 984
rect 3868 976 3876 984
rect 4028 976 4036 984
rect 5596 976 5604 984
rect 5628 976 5636 984
rect 5740 976 5748 984
rect 5868 976 5876 984
rect 5916 976 5924 984
rect 5948 976 5956 984
rect 6188 976 6196 984
rect 6268 976 6276 984
rect 6428 976 6436 984
rect 6508 976 6516 984
rect 6572 976 6580 984
rect 6700 976 6708 984
rect 6716 976 6724 984
rect 6876 976 6884 984
rect 6956 976 6964 984
rect 7276 976 7284 984
rect 7308 976 7316 984
rect 7372 976 7380 984
rect 7516 976 7524 984
rect 252 956 260 964
rect 396 956 404 964
rect 412 956 420 964
rect 476 956 484 964
rect 700 956 708 964
rect 1196 956 1204 964
rect 1260 956 1268 964
rect 2076 956 2084 964
rect 2364 956 2372 964
rect 2540 956 2548 964
rect 12 936 20 944
rect 156 936 164 944
rect 220 936 228 944
rect 252 936 260 944
rect 300 936 308 944
rect 316 936 324 944
rect 380 936 388 944
rect 428 936 436 944
rect 508 936 516 944
rect 588 936 596 944
rect 636 936 644 944
rect 652 936 660 944
rect 844 936 852 944
rect 1116 936 1124 944
rect 1148 936 1156 944
rect 1180 936 1188 944
rect 1228 936 1236 944
rect 1292 936 1300 944
rect 1356 936 1364 944
rect 1372 936 1380 944
rect 1404 936 1412 944
rect 1420 936 1428 944
rect 1484 936 1492 944
rect 1516 936 1524 944
rect 1548 936 1556 944
rect 1756 936 1764 944
rect 1852 936 1860 944
rect 1964 936 1972 944
rect 2156 936 2164 944
rect 2220 936 2228 944
rect 2252 936 2260 944
rect 2380 936 2388 944
rect 2460 936 2468 944
rect 2636 956 2644 964
rect 2700 956 2708 964
rect 2748 956 2756 964
rect 2812 956 2820 964
rect 2908 956 2916 964
rect 2940 956 2948 964
rect 3068 956 3076 964
rect 3084 956 3092 964
rect 3116 956 3124 964
rect 3196 956 3204 964
rect 3228 956 3236 964
rect 3324 956 3332 964
rect 3356 956 3364 964
rect 3388 956 3396 964
rect 3596 956 3604 964
rect 4220 956 4228 964
rect 4364 956 4372 964
rect 4396 956 4404 964
rect 4412 956 4420 964
rect 4508 956 4516 964
rect 4780 956 4788 964
rect 4860 956 4868 964
rect 4924 956 4932 964
rect 5116 956 5124 964
rect 5244 956 5252 964
rect 5500 956 5508 964
rect 5676 956 5684 964
rect 5852 956 5860 964
rect 6140 956 6148 964
rect 6556 956 6564 964
rect 6652 956 6660 964
rect 6940 956 6948 964
rect 6972 956 6980 964
rect 7004 956 7012 964
rect 7100 956 7108 964
rect 7292 956 7300 964
rect 7420 956 7428 964
rect 7484 956 7492 964
rect 2572 936 2580 944
rect 2812 936 2820 944
rect 2844 936 2852 944
rect 2972 936 2980 944
rect 3004 936 3012 944
rect 3084 936 3092 944
rect 3148 936 3156 944
rect 3164 936 3172 944
rect 3260 936 3268 944
rect 3420 936 3428 944
rect 3484 936 3492 944
rect 3644 936 3652 944
rect 3692 936 3700 944
rect 3708 936 3716 944
rect 3740 936 3748 944
rect 3916 936 3924 944
rect 4108 936 4116 944
rect 4156 936 4164 944
rect 4252 936 4260 944
rect 4316 936 4324 944
rect 4364 936 4372 944
rect 4428 936 4436 944
rect 4652 936 4660 944
rect 4700 936 4708 944
rect 4716 936 4724 944
rect 4780 936 4788 944
rect 4828 936 4836 944
rect 5084 936 5092 944
rect 5148 936 5156 944
rect 5436 936 5444 944
rect 5580 936 5588 944
rect 5756 936 5764 944
rect 5788 936 5796 944
rect 5820 936 5828 944
rect 5900 936 5908 944
rect 6012 936 6020 944
rect 6108 936 6116 944
rect 6156 936 6164 944
rect 6252 936 6260 944
rect 6300 932 6308 940
rect 6316 936 6324 944
rect 6364 936 6372 944
rect 6380 936 6388 944
rect 6396 932 6404 940
rect 6444 936 6452 944
rect 6540 936 6548 944
rect 6668 936 6676 944
rect 748 916 756 924
rect 812 918 820 926
rect 1084 918 1092 926
rect 1180 916 1188 924
rect 1244 916 1252 924
rect 1308 916 1316 924
rect 1324 916 1332 924
rect 1436 916 1444 924
rect 1580 918 1588 926
rect 1820 918 1828 926
rect 188 896 196 904
rect 268 896 276 904
rect 348 896 356 904
rect 460 896 468 904
rect 540 896 548 904
rect 572 896 580 904
rect 1180 896 1188 904
rect 1324 896 1332 904
rect 1372 896 1380 904
rect 1996 916 2004 924
rect 2028 916 2036 924
rect 2076 916 2084 924
rect 2124 916 2132 924
rect 2316 916 2324 924
rect 2332 916 2340 924
rect 2348 916 2356 924
rect 2508 916 2516 924
rect 2524 916 2532 924
rect 2588 916 2596 924
rect 2716 916 2724 924
rect 2764 916 2772 924
rect 2860 916 2868 924
rect 3020 916 3028 924
rect 3148 916 3156 924
rect 3228 916 3236 924
rect 3260 916 3268 924
rect 3276 916 3284 924
rect 3292 916 3300 924
rect 3484 916 3492 924
rect 3548 916 3556 924
rect 3564 916 3572 924
rect 3628 916 3636 924
rect 3660 916 3668 924
rect 3820 916 3828 924
rect 3836 916 3844 924
rect 1484 896 1492 904
rect 1724 896 1732 904
rect 2012 896 2020 904
rect 2412 896 2420 904
rect 2940 896 2948 904
rect 3020 896 3028 904
rect 3180 896 3188 904
rect 3308 896 3316 904
rect 3516 896 3524 904
rect 3532 896 3540 904
rect 3692 896 3700 904
rect 3772 896 3780 904
rect 3948 916 3956 924
rect 3964 916 3972 924
rect 3996 916 4004 924
rect 4060 916 4068 924
rect 4076 916 4084 924
rect 4140 916 4148 924
rect 4188 916 4196 924
rect 4284 916 4292 924
rect 4316 916 4324 924
rect 4380 916 4388 924
rect 4444 916 4452 924
rect 4508 918 4516 926
rect 4572 916 4580 924
rect 4652 916 4660 924
rect 4716 916 4724 924
rect 4732 916 4740 924
rect 4796 916 4804 924
rect 4812 916 4820 924
rect 4860 916 4868 924
rect 4940 916 4948 924
rect 5068 916 5076 924
rect 5116 916 5124 924
rect 5180 918 5188 926
rect 5436 918 5444 926
rect 5708 916 5716 924
rect 5772 916 5780 924
rect 5836 916 5844 924
rect 5884 916 5892 924
rect 6028 916 6036 924
rect 6044 916 6052 924
rect 6108 916 6116 924
rect 6332 916 6340 924
rect 6588 916 6596 924
rect 6604 916 6612 924
rect 6828 936 6836 944
rect 6908 932 6916 940
rect 6924 936 6932 944
rect 7068 936 7076 944
rect 7132 936 7140 944
rect 7180 936 7188 944
rect 7356 936 7364 944
rect 7404 936 7412 944
rect 7532 936 7540 944
rect 6988 916 6996 924
rect 7036 916 7044 924
rect 7132 916 7140 924
rect 7196 916 7204 924
rect 7212 916 7220 924
rect 7260 916 7268 924
rect 7340 916 7348 924
rect 7548 916 7556 924
rect 3884 896 3892 904
rect 3980 896 3988 904
rect 4140 896 4148 904
rect 4204 896 4212 904
rect 4300 896 4308 904
rect 5612 896 5620 904
rect 5628 896 5636 904
rect 5724 896 5732 904
rect 5932 896 5940 904
rect 5948 896 5956 904
rect 6060 896 6068 904
rect 6076 896 6084 904
rect 6860 896 6868 904
rect 7052 896 7060 904
rect 7372 896 7380 904
rect 2044 876 2052 884
rect 2172 876 2180 884
rect 2220 876 2228 884
rect 2428 876 2436 884
rect 3356 876 3364 884
rect 4700 876 4708 884
rect 2828 856 2836 864
rect 7036 856 7044 864
rect 124 836 132 844
rect 252 836 260 844
rect 1740 836 1748 844
rect 2108 836 2116 844
rect 3100 836 3108 844
rect 4636 836 4644 844
rect 5052 836 5060 844
rect 5324 836 5332 844
rect 5564 836 5572 844
rect 5788 836 5796 844
rect 739 806 747 814
rect 749 806 757 814
rect 759 806 767 814
rect 769 806 777 814
rect 779 806 787 814
rect 789 806 797 814
rect 3747 806 3755 814
rect 3757 806 3765 814
rect 3767 806 3775 814
rect 3777 806 3785 814
rect 3787 806 3795 814
rect 3797 806 3805 814
rect 6755 806 6763 814
rect 6765 806 6773 814
rect 6775 806 6783 814
rect 6785 806 6793 814
rect 6795 806 6803 814
rect 6805 806 6813 814
rect 12 776 20 784
rect 524 776 532 784
rect 556 776 564 784
rect 604 776 612 784
rect 1196 776 1204 784
rect 1228 776 1236 784
rect 1260 776 1268 784
rect 1500 776 1508 784
rect 1644 776 1652 784
rect 1660 776 1668 784
rect 1980 776 1988 784
rect 2012 776 2020 784
rect 2076 776 2084 784
rect 2140 776 2148 784
rect 2236 776 2244 784
rect 2364 776 2372 784
rect 2428 776 2436 784
rect 2460 776 2468 784
rect 2476 776 2484 784
rect 2604 776 2612 784
rect 2636 776 2644 784
rect 2668 776 2676 784
rect 3372 776 3380 784
rect 3612 776 3620 784
rect 4668 776 4676 784
rect 4780 776 4788 784
rect 4908 776 4916 784
rect 5084 776 5092 784
rect 5580 776 5588 784
rect 5692 776 5700 784
rect 5884 776 5892 784
rect 5932 776 5940 784
rect 6508 776 6516 784
rect 7132 776 7140 784
rect 7180 776 7188 784
rect 7500 776 7508 784
rect 4364 756 4372 764
rect 4604 756 4612 764
rect 1052 736 1060 744
rect 1100 736 1108 744
rect 1308 736 1316 744
rect 2060 736 2068 744
rect 2124 736 2132 744
rect 2204 736 2212 744
rect 2348 736 2356 744
rect 2492 736 2500 744
rect 3164 736 3172 744
rect 3388 736 3396 744
rect 3948 736 3956 744
rect 4572 736 4580 744
rect 4668 736 4676 744
rect 4860 736 4868 744
rect 4924 736 4932 744
rect 4940 736 4948 744
rect 4988 736 4996 744
rect 5052 736 5060 744
rect 5068 736 5076 744
rect 5308 736 5316 744
rect 6876 736 6884 744
rect 6908 736 6916 744
rect 268 716 276 724
rect 412 716 420 724
rect 428 716 436 724
rect 684 716 692 724
rect 828 716 836 724
rect 1116 716 1124 724
rect 1580 716 1588 724
rect 2028 716 2036 724
rect 2092 716 2100 724
rect 2268 716 2276 724
rect 2524 716 2532 724
rect 2988 716 2996 724
rect 3020 716 3028 724
rect 3084 716 3092 724
rect 3196 716 3204 724
rect 3228 716 3236 724
rect 3292 716 3300 724
rect 3356 716 3364 724
rect 3468 716 3476 724
rect 3628 716 3636 724
rect 3676 716 3684 724
rect 3820 716 3828 724
rect 3884 716 3892 724
rect 3996 716 4004 724
rect 4380 716 4388 724
rect 4652 716 4660 724
rect 4796 716 4804 724
rect 4892 716 4900 724
rect 4956 716 4964 724
rect 5020 716 5028 724
rect 5036 716 5044 724
rect 5196 716 5204 724
rect 5388 716 5396 724
rect 5404 716 5412 724
rect 5452 716 5460 724
rect 5500 716 5508 724
rect 5900 716 5908 724
rect 5964 716 5972 724
rect 6044 716 6052 724
rect 6348 716 6356 724
rect 6412 716 6420 724
rect 6940 716 6948 724
rect 7212 716 7220 724
rect 7388 716 7396 724
rect 140 694 148 702
rect 204 696 212 704
rect 364 696 372 704
rect 412 696 420 704
rect 588 696 596 704
rect 652 696 660 704
rect 924 694 932 702
rect 988 696 996 704
rect 1068 696 1076 704
rect 1164 696 1172 704
rect 1276 696 1284 704
rect 1388 696 1396 704
rect 1724 696 1732 704
rect 1740 696 1748 704
rect 1852 694 1860 702
rect 1916 696 1924 704
rect 2044 696 2052 704
rect 2108 696 2116 704
rect 2204 696 2212 704
rect 2332 696 2340 704
rect 2396 696 2404 704
rect 2508 696 2516 704
rect 2572 696 2580 704
rect 2604 696 2612 704
rect 2748 696 2756 704
rect 2876 696 2884 704
rect 2908 696 2916 704
rect 2940 696 2948 704
rect 3004 696 3012 704
rect 3020 696 3028 704
rect 3052 696 3060 704
rect 3180 696 3188 704
rect 3212 696 3220 704
rect 3276 696 3284 704
rect 3324 696 3332 704
rect 3372 696 3380 704
rect 3436 696 3444 704
rect 3484 696 3492 704
rect 3516 696 3524 704
rect 3548 696 3556 704
rect 3580 696 3588 704
rect 3852 696 3860 704
rect 3916 696 3924 704
rect 4092 694 4100 702
rect 4236 696 4244 704
rect 4268 696 4276 704
rect 4300 696 4308 704
rect 4316 696 4324 704
rect 4492 696 4500 704
rect 4636 696 4644 704
rect 4684 696 4692 704
rect 4828 696 4836 704
rect 124 676 132 684
rect 220 676 228 684
rect 300 676 308 684
rect 348 676 356 684
rect 380 676 388 684
rect 396 676 404 684
rect 460 676 468 684
rect 476 676 484 684
rect 652 676 660 684
rect 716 676 724 684
rect 860 676 868 684
rect 1148 676 1156 684
rect 1340 676 1348 684
rect 1516 676 1524 684
rect 1580 676 1588 684
rect 1612 676 1620 684
rect 1692 676 1700 684
rect 1788 676 1796 684
rect 2380 676 2388 684
rect 2700 676 2708 684
rect 2940 676 2948 684
rect 2956 676 2964 684
rect 2988 676 2996 684
rect 3068 676 3076 684
rect 3116 676 3124 684
rect 3228 676 3236 684
rect 3260 676 3268 684
rect 3340 676 3348 684
rect 3420 676 3428 684
rect 3468 676 3476 684
rect 3500 676 3508 684
rect 3532 676 3540 684
rect 3564 676 3572 684
rect 3676 676 3684 684
rect 3708 676 3716 684
rect 3868 676 3876 684
rect 3932 676 3940 684
rect 4028 676 4036 684
rect 4108 676 4116 684
rect 4252 676 4260 684
rect 4284 676 4292 684
rect 4332 676 4340 684
rect 4412 676 4420 684
rect 4444 676 4452 684
rect 4540 676 4548 684
rect 4716 676 4724 684
rect 4828 676 4836 684
rect 4860 696 4868 704
rect 4940 696 4948 704
rect 5004 696 5012 704
rect 5052 696 5060 704
rect 5116 696 5124 704
rect 5340 696 5348 704
rect 5804 696 5812 704
rect 5100 676 5108 684
rect 5228 676 5236 684
rect 5356 676 5364 684
rect 5436 676 5444 684
rect 5484 676 5492 684
rect 5532 676 5540 684
rect 5548 676 5556 684
rect 5644 676 5652 684
rect 5660 676 5668 684
rect 5756 676 5764 684
rect 5932 696 5940 704
rect 5980 696 5988 704
rect 6012 696 6020 704
rect 6076 696 6084 704
rect 6140 696 6148 704
rect 6188 696 6196 704
rect 6236 696 6244 704
rect 6316 696 6324 704
rect 6364 696 6372 704
rect 6412 696 6420 704
rect 6444 696 6452 704
rect 6476 696 6484 704
rect 6556 696 6564 704
rect 6572 696 6580 704
rect 6636 696 6644 704
rect 6716 696 6724 704
rect 6748 696 6756 704
rect 6924 696 6932 704
rect 6956 696 6964 704
rect 7100 696 7108 704
rect 7148 696 7156 704
rect 7228 696 7236 704
rect 7308 696 7316 704
rect 7340 696 7348 704
rect 7388 696 7396 704
rect 5868 676 5876 684
rect 5996 676 6004 684
rect 6028 676 6036 684
rect 6092 676 6100 684
rect 6172 676 6180 684
rect 6348 676 6356 684
rect 6460 676 6468 684
rect 6620 676 6628 684
rect 6700 676 6708 684
rect 6732 676 6740 684
rect 7020 676 7028 684
rect 7052 676 7060 684
rect 7164 676 7172 684
rect 7276 676 7284 684
rect 7420 676 7428 684
rect 7532 676 7540 684
rect 252 656 260 664
rect 316 656 324 664
rect 764 656 772 664
rect 1212 656 1220 664
rect 1244 656 1252 664
rect 1516 656 1524 664
rect 1628 656 1636 664
rect 1660 656 1668 664
rect 1996 656 2004 664
rect 2156 656 2164 664
rect 2444 656 2452 664
rect 2556 656 2564 664
rect 2572 656 2580 664
rect 2620 656 2628 664
rect 2652 656 2660 664
rect 3084 656 3092 664
rect 3724 656 3732 664
rect 4364 656 4372 664
rect 4764 656 4772 664
rect 5164 656 5172 664
rect 5772 656 5780 664
rect 5804 656 5812 664
rect 5852 656 5860 664
rect 6028 656 6036 664
rect 6124 656 6132 664
rect 6220 656 6228 664
rect 6284 656 6292 664
rect 6396 656 6404 664
rect 6620 656 6628 664
rect 6652 656 6660 664
rect 6828 656 6836 664
rect 6924 656 6932 664
rect 6988 656 6996 664
rect 7052 656 7060 664
rect 7116 656 7124 664
rect 236 636 244 644
rect 268 636 276 644
rect 332 636 340 644
rect 732 636 740 644
rect 844 636 852 644
rect 1116 636 1124 644
rect 1196 636 1204 644
rect 2860 636 2868 644
rect 3292 636 3300 644
rect 3644 636 3652 644
rect 3692 636 3700 644
rect 3804 636 3812 644
rect 3820 636 3828 644
rect 3884 636 3892 644
rect 4012 636 4020 644
rect 4220 636 4228 644
rect 4380 636 4388 644
rect 4732 636 4740 644
rect 4796 636 4804 644
rect 5148 636 5156 644
rect 5180 636 5188 644
rect 5196 636 5204 644
rect 5372 636 5380 644
rect 5420 636 5428 644
rect 5468 636 5476 644
rect 5516 636 5524 644
rect 5724 636 5732 644
rect 6268 636 6276 644
rect 6412 636 6420 644
rect 6524 636 6532 644
rect 7068 636 7076 644
rect 2243 606 2251 614
rect 2253 606 2261 614
rect 2263 606 2271 614
rect 2273 606 2281 614
rect 2283 606 2291 614
rect 2293 606 2301 614
rect 5251 606 5259 614
rect 5261 606 5269 614
rect 5271 606 5279 614
rect 5281 606 5289 614
rect 5291 606 5299 614
rect 5301 606 5309 614
rect 188 576 196 584
rect 380 576 388 584
rect 396 576 404 584
rect 716 576 724 584
rect 876 576 884 584
rect 1148 576 1156 584
rect 1388 576 1396 584
rect 1580 576 1588 584
rect 1676 576 1684 584
rect 1820 576 1828 584
rect 1852 576 1860 584
rect 1916 576 1924 584
rect 2060 576 2068 584
rect 2172 576 2180 584
rect 2316 576 2324 584
rect 2460 576 2468 584
rect 3068 576 3076 584
rect 3164 576 3172 584
rect 3420 576 3428 584
rect 3612 576 3620 584
rect 3900 576 3908 584
rect 5036 576 5044 584
rect 5164 576 5172 584
rect 5740 576 5748 584
rect 5788 576 5796 584
rect 5900 576 5908 584
rect 5996 576 6004 584
rect 6124 576 6132 584
rect 6508 576 6516 584
rect 6572 576 6580 584
rect 6844 576 6852 584
rect 6956 576 6964 584
rect 7036 576 7044 584
rect 7084 576 7092 584
rect 7436 576 7444 584
rect 892 556 900 564
rect 956 556 964 564
rect 1404 556 1412 564
rect 1532 556 1540 564
rect 1644 556 1652 564
rect 1660 556 1668 564
rect 1836 556 1844 564
rect 2076 556 2084 564
rect 2188 556 2196 564
rect 2204 556 2212 564
rect 2460 556 2468 564
rect 2556 556 2564 564
rect 3036 556 3044 564
rect 3052 556 3060 564
rect 3180 556 3188 564
rect 3260 556 3268 564
rect 3292 556 3300 564
rect 3308 556 3316 564
rect 3548 556 3556 564
rect 3612 556 3620 564
rect 3932 556 3940 564
rect 4076 556 4084 564
rect 4204 556 4212 564
rect 4396 556 4404 564
rect 4476 556 4484 564
rect 4540 556 4548 564
rect 4732 556 4740 564
rect 4812 556 4820 564
rect 5020 556 5028 564
rect 5116 556 5124 564
rect 5132 556 5140 564
rect 5212 556 5220 564
rect 5452 556 5460 564
rect 5564 556 5572 564
rect 5980 556 5988 564
rect 6044 556 6052 564
rect 6140 556 6148 564
rect 6156 556 6164 564
rect 6316 556 6324 564
rect 6460 556 6468 564
rect 6620 556 6628 564
rect 6652 556 6660 564
rect 6988 556 6996 564
rect 7052 556 7060 564
rect 7068 556 7076 564
rect 7180 556 7188 564
rect 7292 556 7300 564
rect 7356 556 7364 564
rect 7484 556 7492 564
rect 7500 556 7508 564
rect 220 536 228 544
rect 684 536 692 544
rect 812 536 820 544
rect 828 536 836 544
rect 860 536 868 544
rect 924 536 932 544
rect 988 536 996 544
rect 1196 536 1204 544
rect 1292 536 1300 544
rect 1436 536 1444 544
rect 1500 536 1508 544
rect 1516 536 1524 544
rect 1564 536 1572 544
rect 1612 536 1620 544
rect 1692 536 1700 544
rect 1772 536 1780 544
rect 1868 536 1876 544
rect 1932 536 1940 544
rect 1980 536 1988 544
rect 2172 536 2180 544
rect 2300 536 2308 544
rect 2364 536 2372 544
rect 2460 536 2468 544
rect 2700 536 2708 544
rect 2764 536 2772 544
rect 2828 536 2836 544
rect 3116 536 3124 544
rect 76 516 84 524
rect 124 516 132 524
rect 284 516 292 524
rect 460 516 468 524
rect 508 516 516 524
rect 620 516 628 524
rect 668 516 676 524
rect 844 516 852 524
rect 908 516 916 524
rect 1020 518 1028 526
rect 1164 516 1172 524
rect 1276 516 1284 524
rect 1404 516 1412 524
rect 1788 516 1796 524
rect 1884 516 1892 524
rect 1996 516 2004 524
rect 2012 516 2020 524
rect 2044 516 2052 524
rect 2156 516 2164 524
rect 2364 516 2372 524
rect 2476 516 2484 524
rect 2556 518 2564 526
rect 2716 516 2724 524
rect 2732 516 2740 524
rect 2876 516 2884 524
rect 2924 516 2932 524
rect 3148 516 3156 524
rect 3164 516 3172 524
rect 3356 516 3364 524
rect 3500 536 3508 544
rect 3724 536 3732 544
rect 3756 536 3764 544
rect 3868 536 3876 544
rect 3900 536 3908 544
rect 3964 536 3972 544
rect 4044 536 4052 544
rect 4236 536 4244 544
rect 4348 536 4356 544
rect 4396 536 4404 544
rect 4412 536 4420 544
rect 4684 536 4692 544
rect 4732 536 4740 544
rect 4748 536 4756 544
rect 4908 536 4916 544
rect 5084 536 5092 544
rect 5308 536 5316 544
rect 5356 536 5364 544
rect 5420 536 5428 544
rect 5548 536 5556 544
rect 5644 536 5652 544
rect 5852 536 5860 544
rect 5868 536 5876 544
rect 5980 536 5988 544
rect 6108 536 6116 544
rect 6188 536 6196 544
rect 6252 536 6260 544
rect 6380 536 6388 544
rect 6412 536 6420 544
rect 6524 536 6532 544
rect 6540 536 6548 544
rect 6668 536 6676 544
rect 6700 536 6708 544
rect 6780 536 6788 544
rect 6876 536 6884 544
rect 6892 536 6900 544
rect 6940 536 6948 544
rect 7100 536 7108 544
rect 7164 536 7172 544
rect 7212 536 7220 544
rect 732 496 740 504
rect 796 496 804 504
rect 956 496 964 504
rect 1468 496 1476 504
rect 1548 496 1556 504
rect 1596 496 1604 504
rect 1644 496 1652 504
rect 1724 496 1732 504
rect 1964 496 1972 504
rect 2028 496 2036 504
rect 2316 496 2324 504
rect 2796 496 2804 504
rect 3036 496 3044 504
rect 3068 496 3076 504
rect 3372 496 3380 504
rect 3468 516 3476 524
rect 3484 516 3492 524
rect 3628 516 3636 524
rect 3708 516 3716 524
rect 3820 516 3828 524
rect 3852 516 3860 524
rect 3932 516 3940 524
rect 3996 516 4004 524
rect 4028 516 4036 524
rect 4108 516 4116 524
rect 4204 518 4212 526
rect 4348 516 4356 524
rect 4412 516 4420 524
rect 4428 516 4436 524
rect 4540 518 4548 526
rect 4684 516 4692 524
rect 4748 516 4756 524
rect 4764 516 4772 524
rect 4876 518 4884 526
rect 5068 516 5076 524
rect 5164 516 5172 524
rect 5388 516 5396 524
rect 5404 516 5412 524
rect 5500 516 5508 524
rect 5516 516 5524 524
rect 5532 516 5540 524
rect 5612 516 5620 524
rect 5628 516 5636 524
rect 5660 516 5668 524
rect 5708 516 5716 524
rect 6060 516 6068 524
rect 6108 516 6116 524
rect 6172 516 6180 524
rect 6204 516 6212 524
rect 6220 516 6228 524
rect 6236 516 6244 524
rect 6300 516 6308 524
rect 6364 516 6372 524
rect 6412 516 6420 524
rect 6428 516 6436 524
rect 6476 516 6484 524
rect 6556 516 6564 524
rect 6636 516 6644 524
rect 6924 516 6932 524
rect 7228 516 7236 524
rect 7324 516 7332 524
rect 7372 516 7380 524
rect 3436 496 3444 504
rect 3532 496 3540 504
rect 3548 496 3556 504
rect 4012 496 4020 504
rect 4076 496 4084 504
rect 4092 496 4100 504
rect 4476 496 4484 504
rect 4812 496 4820 504
rect 5100 496 5108 504
rect 5148 496 5156 504
rect 5356 496 5364 504
rect 5372 496 5380 504
rect 5500 496 5508 504
rect 5580 496 5588 504
rect 5596 496 5604 504
rect 7228 496 7236 504
rect 7292 496 7300 504
rect 3340 476 3348 484
rect 4124 476 4132 484
rect 5132 476 5140 484
rect 5468 476 5476 484
rect 7292 476 7300 484
rect 588 436 596 444
rect 636 436 644 444
rect 2684 436 2692 444
rect 2988 436 2996 444
rect 3276 436 3284 444
rect 3356 436 3364 444
rect 3756 436 3764 444
rect 4108 436 4116 444
rect 4332 436 4340 444
rect 4668 436 4676 444
rect 5004 436 5012 444
rect 5692 436 5700 444
rect 6268 436 6276 444
rect 6444 436 6452 444
rect 7404 436 7412 444
rect 7532 436 7540 444
rect 739 406 747 414
rect 749 406 757 414
rect 759 406 767 414
rect 769 406 777 414
rect 779 406 787 414
rect 789 406 797 414
rect 3747 406 3755 414
rect 3757 406 3765 414
rect 3767 406 3775 414
rect 3777 406 3785 414
rect 3787 406 3795 414
rect 3797 406 3805 414
rect 6755 406 6763 414
rect 6765 406 6773 414
rect 6775 406 6783 414
rect 6785 406 6793 414
rect 6795 406 6803 414
rect 6805 406 6813 414
rect 444 376 452 384
rect 524 376 532 384
rect 716 376 724 384
rect 1324 376 1332 384
rect 1356 376 1364 384
rect 1388 376 1396 384
rect 1420 376 1428 384
rect 1468 376 1476 384
rect 1500 376 1508 384
rect 1532 376 1540 384
rect 1836 376 1844 384
rect 2156 376 2164 384
rect 2380 376 2388 384
rect 2476 376 2484 384
rect 2556 376 2564 384
rect 3708 376 3716 384
rect 3884 376 3892 384
rect 4172 376 4180 384
rect 4268 376 4276 384
rect 4492 376 4500 384
rect 4780 376 4788 384
rect 5612 376 5620 384
rect 5804 376 5812 384
rect 6140 376 6148 384
rect 6236 376 6244 384
rect 6332 376 6340 384
rect 6572 376 6580 384
rect 6668 376 6676 384
rect 7004 376 7012 384
rect 7452 376 7460 384
rect 188 356 196 364
rect 3116 356 3124 364
rect 5132 356 5140 364
rect 1084 336 1092 344
rect 1292 336 1300 344
rect 2700 336 2708 344
rect 3068 336 3076 344
rect 3132 336 3140 344
rect 3900 336 3908 344
rect 4188 336 4196 344
rect 4508 336 4516 344
rect 4556 336 4564 344
rect 4636 336 4644 344
rect 4700 336 4708 344
rect 5260 336 5268 344
rect 5420 336 5428 344
rect 6556 336 6564 344
rect 7020 336 7028 344
rect 7164 336 7172 344
rect 620 316 628 324
rect 668 316 676 324
rect 1004 316 1012 324
rect 1100 316 1108 324
rect 1612 316 1620 324
rect 2076 316 2084 324
rect 60 294 68 302
rect 124 296 132 304
rect 252 294 260 302
rect 764 296 772 304
rect 876 296 884 304
rect 1004 296 1012 304
rect 1052 296 1060 304
rect 1196 294 1204 302
rect 1436 296 1444 304
rect 1564 296 1572 304
rect 1708 294 1716 302
rect 1772 296 1780 304
rect 1932 294 1940 302
rect 2108 296 2116 304
rect 220 276 228 284
rect 300 276 308 284
rect 540 276 548 284
rect 588 276 596 284
rect 652 276 660 284
rect 700 276 708 284
rect 860 276 868 284
rect 876 276 884 284
rect 924 276 932 284
rect 956 276 964 284
rect 1036 276 1044 284
rect 1132 276 1140 284
rect 1580 276 1588 284
rect 1644 276 1652 284
rect 1804 276 1812 284
rect 1852 276 1860 284
rect 1948 276 1956 284
rect 2092 276 2100 284
rect 2156 296 2164 304
rect 2300 316 2308 324
rect 2428 316 2436 324
rect 2508 316 2516 324
rect 3036 316 3044 324
rect 3116 316 3124 324
rect 3196 316 3204 324
rect 3212 316 3220 324
rect 2236 296 2244 304
rect 2364 296 2372 304
rect 2556 296 2564 304
rect 2604 296 2612 304
rect 2636 296 2644 304
rect 2700 296 2708 304
rect 2780 296 2788 304
rect 2892 296 2900 304
rect 2956 296 2964 304
rect 2972 296 2980 304
rect 3052 296 3060 304
rect 3116 296 3124 304
rect 3276 296 3284 304
rect 3324 316 3332 324
rect 3628 316 3636 324
rect 3692 316 3700 324
rect 3868 316 3876 324
rect 3932 316 3940 324
rect 3996 316 4004 324
rect 4092 316 4100 324
rect 4156 316 4164 324
rect 4428 314 4436 322
rect 4476 316 4484 324
rect 4588 316 4596 324
rect 4604 316 4612 324
rect 4732 316 4740 324
rect 5020 316 5028 324
rect 5228 316 5236 324
rect 5340 316 5348 324
rect 5692 316 5700 324
rect 5916 316 5924 324
rect 6028 316 6036 324
rect 6092 316 6100 324
rect 6172 316 6180 324
rect 6284 316 6292 324
rect 6476 316 6484 324
rect 6524 316 6532 324
rect 6716 316 6724 324
rect 6940 316 6948 324
rect 6988 316 6996 324
rect 7196 316 7204 324
rect 7292 316 7300 324
rect 7388 316 7396 324
rect 7484 316 7492 324
rect 3356 296 3364 304
rect 3436 296 3444 304
rect 3500 296 3508 304
rect 3548 296 3556 304
rect 3660 296 3668 304
rect 3836 296 3844 304
rect 3884 296 3892 304
rect 3964 296 3972 304
rect 4076 296 4084 304
rect 4092 296 4100 304
rect 4124 296 4132 304
rect 4172 296 4180 304
rect 4268 296 4276 304
rect 4396 296 4404 304
rect 4492 296 4500 304
rect 4540 296 4548 304
rect 4572 296 4580 304
rect 4636 296 4644 304
rect 4700 296 4708 304
rect 4748 296 4756 304
rect 4828 296 4836 304
rect 4892 296 4900 304
rect 5052 296 5060 304
rect 5084 296 5092 304
rect 5148 296 5156 304
rect 5212 296 5220 304
rect 5244 296 5252 304
rect 5388 296 5396 304
rect 5500 296 5508 304
rect 5644 296 5652 304
rect 5724 296 5732 304
rect 5756 296 5764 304
rect 5836 296 5844 304
rect 5964 296 5972 304
rect 5980 296 5988 304
rect 6060 296 6068 304
rect 6540 296 6548 304
rect 6588 296 6596 304
rect 6636 296 6644 304
rect 6876 296 6884 304
rect 7004 296 7012 304
rect 2140 276 2148 284
rect 2364 276 2372 284
rect 2444 276 2452 284
rect 2460 276 2468 284
rect 2620 276 2628 284
rect 2652 276 2660 284
rect 2812 276 2820 284
rect 2860 276 2868 284
rect 2908 276 2916 284
rect 2956 276 2964 284
rect 2988 276 2996 284
rect 3068 276 3076 284
rect 3164 276 3172 284
rect 3260 276 3268 284
rect 3292 276 3300 284
rect 3356 276 3364 284
rect 3388 276 3396 284
rect 3452 276 3460 284
rect 3468 276 3476 284
rect 3484 276 3492 284
rect 3580 276 3588 284
rect 3612 276 3620 284
rect 3644 276 3652 284
rect 3852 276 3860 284
rect 3932 276 3940 284
rect 3980 276 3988 284
rect 4140 276 4148 284
rect 4252 276 4260 284
rect 4380 276 4388 284
rect 4812 276 4820 284
rect 4908 276 4916 284
rect 4924 276 4932 284
rect 5036 276 5044 284
rect 5068 276 5076 284
rect 5084 276 5092 284
rect 5132 276 5140 284
rect 5196 276 5204 284
rect 5244 276 5252 284
rect 5292 276 5300 284
rect 5404 276 5412 284
rect 5484 276 5492 284
rect 5548 276 5556 284
rect 5596 276 5604 284
rect 5676 276 5684 284
rect 5740 276 5748 284
rect 5788 276 5796 284
rect 5884 276 5892 284
rect 5916 276 5924 284
rect 5964 276 5972 284
rect 6076 276 6084 284
rect 6124 276 6132 284
rect 6204 276 6212 284
rect 6252 276 6260 284
rect 6284 276 6292 284
rect 6396 276 6404 284
rect 6412 276 6420 284
rect 6508 276 6516 284
rect 6828 276 6836 284
rect 6844 276 6852 284
rect 6860 276 6868 284
rect 6876 276 6884 284
rect 6972 276 6980 284
rect 7052 276 7060 284
rect 7148 276 7156 284
rect 7212 296 7220 304
rect 7308 296 7316 304
rect 7372 296 7380 304
rect 7468 296 7476 304
rect 7420 276 7428 284
rect 7516 276 7524 284
rect 556 256 564 264
rect 684 256 692 264
rect 812 256 820 264
rect 892 256 900 264
rect 1196 256 1204 264
rect 1340 256 1348 264
rect 1372 256 1380 264
rect 1404 256 1412 264
rect 1484 256 1492 264
rect 1516 256 1524 264
rect 1548 256 1556 264
rect 1868 256 1876 264
rect 2204 256 2212 264
rect 2396 256 2404 264
rect 2524 256 2532 264
rect 2684 256 2692 264
rect 2732 256 2740 264
rect 2764 256 2772 264
rect 2828 256 2836 264
rect 2876 256 2884 264
rect 2940 256 2948 264
rect 3020 256 3028 264
rect 3180 256 3188 264
rect 3420 256 3428 264
rect 3532 256 3540 264
rect 3548 256 3556 264
rect 3724 256 3732 264
rect 4220 256 4228 264
rect 4332 256 4340 264
rect 4380 256 4388 264
rect 4668 256 4676 264
rect 4700 256 4708 264
rect 4796 256 4804 264
rect 4908 256 4916 264
rect 5164 256 5172 264
rect 5436 256 5444 264
rect 5468 256 5476 264
rect 5660 256 5668 264
rect 5820 256 5828 264
rect 5932 256 5940 264
rect 6012 256 6020 264
rect 6156 256 6164 264
rect 6220 256 6228 264
rect 6684 256 6692 264
rect 6716 256 6724 264
rect 6924 256 6932 264
rect 7340 256 7348 264
rect 7436 256 7444 264
rect 7532 256 7540 264
rect 380 236 388 244
rect 572 236 580 244
rect 844 236 852 244
rect 1116 236 1124 244
rect 1468 236 1476 244
rect 2060 236 2068 244
rect 2316 236 2324 244
rect 2572 236 2580 244
rect 2668 236 2676 244
rect 3004 236 3012 244
rect 3212 236 3220 244
rect 3404 236 3412 244
rect 3692 236 3700 244
rect 3740 236 3748 244
rect 3996 236 4004 244
rect 4044 236 4052 244
rect 4924 236 4932 244
rect 5180 236 5188 244
rect 5484 236 5492 244
rect 5692 236 5700 244
rect 5916 236 5924 244
rect 6108 236 6116 244
rect 6172 236 6180 244
rect 6284 236 6292 244
rect 6620 236 6628 244
rect 6940 236 6948 244
rect 7244 236 7252 244
rect 2243 206 2251 214
rect 2253 206 2261 214
rect 2263 206 2271 214
rect 2273 206 2281 214
rect 2283 206 2291 214
rect 2293 206 2301 214
rect 5251 206 5259 214
rect 5261 206 5269 214
rect 5271 206 5279 214
rect 5281 206 5289 214
rect 5291 206 5299 214
rect 5301 206 5309 214
rect 44 176 52 184
rect 140 176 148 184
rect 460 176 468 184
rect 652 176 660 184
rect 668 176 676 184
rect 956 176 964 184
rect 972 176 980 184
rect 1020 176 1028 184
rect 1148 176 1156 184
rect 1260 176 1268 184
rect 1884 176 1892 184
rect 2076 176 2084 184
rect 2412 176 2420 184
rect 2588 176 2596 184
rect 2748 176 2756 184
rect 2828 176 2836 184
rect 2876 176 2884 184
rect 3084 176 3092 184
rect 3116 176 3124 184
rect 3356 176 3364 184
rect 3548 176 3556 184
rect 3836 176 3844 184
rect 60 156 68 164
rect 124 156 132 164
rect 1164 156 1172 164
rect 1196 156 1204 164
rect 1468 156 1476 164
rect 1500 156 1508 164
rect 1516 156 1524 164
rect 1532 156 1540 164
rect 1660 156 1668 164
rect 1948 156 1956 164
rect 2108 156 2116 164
rect 2140 156 2148 164
rect 2156 156 2164 164
rect 2396 156 2404 164
rect 2428 156 2436 164
rect 2620 156 2628 164
rect 2700 156 2708 164
rect 2732 156 2740 164
rect 2796 156 2804 164
rect 2844 156 2852 164
rect 2860 156 2868 164
rect 3100 156 3108 164
rect 3132 156 3140 164
rect 3420 156 3428 164
rect 4284 176 4292 184
rect 4604 176 4612 184
rect 4668 176 4676 184
rect 5324 176 5332 184
rect 5644 176 5652 184
rect 6540 176 6548 184
rect 6748 176 6756 184
rect 6940 176 6948 184
rect 7260 176 7268 184
rect 7388 176 7396 184
rect 7500 176 7508 184
rect 4380 156 4388 164
rect 4444 156 4452 164
rect 4620 156 4628 164
rect 28 136 36 144
rect 108 136 116 144
rect 156 136 164 144
rect 220 136 228 144
rect 236 136 244 144
rect 268 136 276 144
rect 300 136 308 144
rect 492 136 500 144
rect 796 136 804 144
rect 1004 136 1012 144
rect 1052 136 1060 144
rect 1100 136 1108 144
rect 1132 136 1140 144
rect 1180 136 1188 144
rect 1228 136 1236 144
rect 1436 136 1444 144
rect 1644 136 1652 144
rect 1772 136 1780 144
rect 2172 136 2180 144
rect 2284 136 2292 144
rect 2460 136 2468 144
rect 2492 136 2500 144
rect 2556 136 2564 144
rect 2636 136 2644 144
rect 2716 136 2724 144
rect 2924 136 2932 144
rect 3164 136 3172 144
rect 3676 136 3684 144
rect 3948 136 3956 144
rect 3996 136 4004 144
rect 4188 136 4196 144
rect 4300 136 4308 144
rect 4348 136 4356 144
rect 4364 136 4372 144
rect 4412 136 4420 144
rect 4780 156 4788 164
rect 4988 156 4996 164
rect 5132 156 5140 164
rect 5196 156 5204 164
rect 5852 156 5860 164
rect 5948 156 5956 164
rect 6028 156 6036 164
rect 6236 156 6244 164
rect 6636 156 6644 164
rect 6780 156 6788 164
rect 6956 156 6964 164
rect 6972 156 6980 164
rect 7148 156 7156 164
rect 7212 156 7220 164
rect 4668 136 4676 144
rect 4732 136 4740 144
rect 4876 136 4884 144
rect 4940 136 4948 144
rect 4988 136 4996 144
rect 5052 136 5060 144
rect 5100 136 5108 144
rect 5484 136 5492 144
rect 5884 136 5892 144
rect 5932 136 5940 144
rect 6156 136 6164 144
rect 6220 136 6228 144
rect 6268 136 6276 144
rect 6316 136 6324 144
rect 6476 136 6484 144
rect 6572 136 6580 144
rect 6668 136 6676 144
rect 6684 136 6692 144
rect 6700 136 6708 144
rect 6844 136 6852 144
rect 6924 136 6932 144
rect 7036 136 7044 144
rect 7052 136 7060 144
rect 7100 136 7108 144
rect 7228 136 7236 144
rect 7276 136 7284 144
rect 7308 136 7316 144
rect 7356 136 7364 144
rect 7484 136 7492 144
rect 7516 136 7524 144
rect 12 116 20 124
rect 76 116 84 124
rect 348 116 356 124
rect 572 116 580 124
rect 764 116 772 124
rect 876 116 884 124
rect 1068 116 1076 124
rect 1116 116 1124 124
rect 1388 116 1396 124
rect 1468 116 1476 124
rect 1628 116 1636 124
rect 1692 116 1700 124
rect 1756 118 1764 126
rect 1964 116 1972 124
rect 2204 116 2212 124
rect 2236 116 2244 124
rect 2300 116 2308 124
rect 2540 116 2548 124
rect 2652 116 2660 124
rect 2684 116 2692 124
rect 2892 116 2900 124
rect 3004 116 3012 124
rect 3276 116 3284 124
rect 3324 116 3332 124
rect 3420 118 3428 126
rect 3596 116 3604 124
rect 3612 116 3620 124
rect 3740 116 3748 124
rect 4012 116 4020 124
rect 4060 116 4068 124
rect 4172 116 4180 124
rect 4300 116 4308 124
rect 4364 116 4372 124
rect 4428 116 4436 124
rect 4508 116 4516 124
rect 4588 116 4596 124
rect 4684 116 4692 124
rect 4844 116 4852 124
rect 4860 116 4868 124
rect 4876 116 4884 124
rect 4940 116 4948 124
rect 5004 116 5012 124
rect 5052 116 5060 124
rect 5084 116 5092 124
rect 5196 118 5204 126
rect 5420 116 5428 124
rect 5516 118 5524 126
rect 5660 116 5668 124
rect 5708 116 5716 124
rect 5756 116 5764 124
rect 5804 116 5812 124
rect 5980 116 5988 124
rect 6044 116 6052 124
rect 6140 116 6148 124
rect 6188 116 6196 124
rect 6204 116 6212 124
rect 6332 116 6340 124
rect 6380 116 6388 124
rect 6428 116 6436 124
rect 6588 116 6596 124
rect 6716 116 6724 124
rect 6780 116 6788 124
rect 6860 116 6868 124
rect 7004 116 7012 124
rect 7100 116 7108 124
rect 7116 116 7124 124
rect 7196 116 7204 124
rect 7468 116 7476 124
rect 7532 116 7540 124
rect 76 96 84 104
rect 188 96 196 104
rect 236 96 244 104
rect 972 96 980 104
rect 1020 96 1028 104
rect 1212 96 1220 104
rect 1260 96 1268 104
rect 1596 96 1604 104
rect 2140 96 2148 104
rect 2220 96 2228 104
rect 2332 96 2340 104
rect 3212 96 3220 104
rect 3996 96 4004 104
rect 4524 96 4532 104
rect 4540 96 4548 104
rect 4812 96 4820 104
rect 4828 96 4836 104
rect 5068 96 5076 104
rect 5132 96 5140 104
rect 5404 96 5412 104
rect 5932 96 5940 104
rect 5964 96 5972 104
rect 6108 96 6116 104
rect 6172 96 6180 104
rect 6316 96 6324 104
rect 6668 96 6676 104
rect 6700 96 6708 104
rect 6892 96 6900 104
rect 7276 96 7284 104
rect 7308 96 7316 104
rect 1276 76 1284 84
rect 1692 76 1700 84
rect 2092 76 2100 84
rect 2252 76 2260 84
rect 4348 76 4356 84
rect 4460 76 4468 84
rect 4492 76 4500 84
rect 4572 76 4580 84
rect 5036 76 5044 84
rect 5436 76 5444 84
rect 7116 76 7124 84
rect 4476 56 4484 64
rect 5420 56 5428 64
rect 1548 36 1556 44
rect 2508 36 2516 44
rect 3260 36 3268 44
rect 3308 36 3316 44
rect 3564 36 3572 44
rect 3644 36 3652 44
rect 4044 36 4052 44
rect 4092 36 4100 44
rect 4924 36 4932 44
rect 5692 36 5700 44
rect 5740 36 5748 44
rect 5788 36 5796 44
rect 5836 36 5844 44
rect 6012 36 6020 44
rect 6060 36 6068 44
rect 6364 36 6372 44
rect 6412 36 6420 44
rect 6460 36 6468 44
rect 6620 36 6628 44
rect 7164 36 7172 44
rect 739 6 747 14
rect 749 6 757 14
rect 759 6 767 14
rect 769 6 777 14
rect 779 6 787 14
rect 789 6 797 14
rect 3747 6 3755 14
rect 3757 6 3765 14
rect 3767 6 3775 14
rect 3777 6 3785 14
rect 3787 6 3795 14
rect 3797 6 3805 14
rect 6755 6 6763 14
rect 6765 6 6773 14
rect 6775 6 6783 14
rect 6785 6 6793 14
rect 6795 6 6803 14
rect 6805 6 6813 14
<< metal2 >>
rect 3885 5224 3891 5263
rect 4221 5257 4243 5263
rect 4461 5257 4483 5263
rect 4509 5257 4531 5263
rect 4669 5257 4691 5263
rect 762 5214 774 5216
rect 3770 5214 3782 5216
rect 747 5206 749 5214
rect 757 5206 759 5214
rect 767 5206 769 5214
rect 777 5206 779 5214
rect 787 5206 789 5214
rect 3755 5206 3757 5214
rect 3765 5206 3767 5214
rect 3775 5206 3777 5214
rect 3785 5206 3787 5214
rect 3795 5206 3797 5214
rect 762 5204 774 5206
rect 3770 5204 3782 5206
rect 381 5104 387 5116
rect 477 5102 483 5116
rect 77 5044 83 5096
rect 125 5084 131 5096
rect 77 4924 83 4956
rect 125 4924 131 5076
rect 189 5024 195 5036
rect 189 4944 195 4976
rect 205 4924 211 5096
rect 221 5064 227 5076
rect 269 5064 275 5096
rect 317 5064 323 5096
rect 397 5064 403 5076
rect 301 5024 307 5056
rect 349 5044 355 5056
rect 301 5003 307 5016
rect 301 4997 323 5003
rect 269 4944 275 4956
rect 221 4924 227 4936
rect 317 4924 323 4997
rect 381 4924 387 4936
rect 77 4584 83 4696
rect 93 4524 99 4536
rect 109 4524 115 4756
rect 125 4704 131 4916
rect 205 4764 211 4916
rect 125 4684 131 4696
rect 125 4304 131 4676
rect 189 4644 195 4656
rect 157 4524 163 4576
rect 189 4564 195 4636
rect 221 4544 227 4916
rect 301 4864 307 4916
rect 253 4584 259 4694
rect 237 4524 243 4536
rect 77 4284 83 4296
rect 125 4124 131 4296
rect 77 3904 83 3916
rect 125 3904 131 4116
rect 125 3884 131 3896
rect 125 3724 131 3876
rect 125 3584 131 3716
rect 173 3524 179 4516
rect 221 4423 227 4516
rect 205 4417 227 4423
rect 205 4304 211 4417
rect 301 4304 307 4536
rect 349 4524 355 4736
rect 365 4704 371 4836
rect 397 4784 403 5056
rect 413 4984 419 5096
rect 685 5084 691 5096
rect 525 4944 531 5076
rect 749 5044 755 5094
rect 477 4924 483 4936
rect 413 4744 419 4916
rect 461 4724 467 4836
rect 493 4824 499 4916
rect 573 4904 579 4916
rect 429 4644 435 4696
rect 381 4544 387 4636
rect 493 4564 499 4696
rect 525 4684 531 4716
rect 557 4704 563 4816
rect 605 4804 611 5036
rect 621 4944 627 5036
rect 717 4924 723 4936
rect 573 4704 579 4736
rect 637 4704 643 4716
rect 461 4544 467 4556
rect 509 4524 515 4536
rect 349 4464 355 4516
rect 308 4297 323 4303
rect 189 4244 195 4256
rect 189 4164 195 4176
rect 205 4124 211 4296
rect 221 4284 227 4296
rect 317 4124 323 4297
rect 333 4224 339 4296
rect 349 4244 355 4436
rect 397 4344 403 4456
rect 397 4304 403 4336
rect 413 4304 419 4516
rect 429 4324 435 4516
rect 445 4464 451 4496
rect 365 4264 371 4276
rect 381 4264 387 4296
rect 413 4264 419 4296
rect 333 4164 339 4216
rect 349 4164 355 4176
rect 365 4164 371 4176
rect 212 4117 227 4123
rect 205 3944 211 4076
rect 205 3884 211 3936
rect 221 3864 227 4117
rect 333 3924 339 4036
rect 237 3904 243 3916
rect 253 3884 259 3916
rect 301 3803 307 3876
rect 365 3823 371 3894
rect 349 3817 371 3823
rect 301 3797 316 3803
rect 196 3777 211 3783
rect 205 3764 211 3777
rect 237 3724 243 3736
rect 301 3724 307 3736
rect 317 3724 323 3796
rect 349 3784 355 3817
rect 365 3764 371 3776
rect 413 3744 419 3896
rect 429 3763 435 4256
rect 477 4224 483 4296
rect 493 4204 499 4516
rect 525 4504 531 4676
rect 557 4584 563 4696
rect 573 4664 579 4676
rect 621 4584 627 4676
rect 557 4564 563 4576
rect 605 4544 611 4556
rect 653 4544 659 4836
rect 701 4824 707 4916
rect 669 4684 675 4696
rect 509 4284 515 4496
rect 525 4284 531 4296
rect 541 4224 547 4516
rect 589 4323 595 4336
rect 573 4317 595 4323
rect 573 4304 579 4317
rect 573 4244 579 4276
rect 589 4204 595 4296
rect 461 3944 467 4136
rect 477 4104 483 4116
rect 493 3984 499 4176
rect 605 4164 611 4536
rect 669 4524 675 4556
rect 685 4344 691 4796
rect 701 4784 707 4816
rect 762 4814 774 4816
rect 747 4806 749 4814
rect 757 4806 759 4814
rect 767 4806 769 4814
rect 777 4806 779 4814
rect 787 4806 789 4814
rect 762 4804 774 4806
rect 813 4784 819 4896
rect 701 4704 707 4716
rect 813 4704 819 4716
rect 717 4684 723 4696
rect 733 4684 739 4696
rect 829 4683 835 4876
rect 845 4704 851 5096
rect 893 5064 899 5076
rect 973 5064 979 5096
rect 877 4924 883 4936
rect 861 4824 867 4916
rect 893 4903 899 5056
rect 925 4924 931 4996
rect 941 4944 947 5056
rect 989 4984 995 5116
rect 1101 5102 1107 5116
rect 2733 5104 2739 5116
rect 2893 5104 2899 5116
rect 3421 5104 3427 5116
rect 3581 5104 3587 5116
rect 1005 4944 1011 4956
rect 877 4897 899 4903
rect 861 4744 867 4816
rect 813 4677 835 4683
rect 717 4623 723 4676
rect 701 4617 723 4623
rect 701 4504 707 4617
rect 733 4583 739 4676
rect 717 4577 739 4583
rect 701 4484 707 4496
rect 637 4304 643 4336
rect 621 4224 627 4256
rect 653 4184 659 4296
rect 653 4144 659 4156
rect 557 4044 563 4136
rect 669 4124 675 4256
rect 685 4124 691 4176
rect 621 4104 627 4116
rect 541 3904 547 3916
rect 509 3864 515 3876
rect 557 3844 563 3916
rect 621 3904 627 4096
rect 669 4064 675 4116
rect 637 3904 643 3916
rect 429 3757 451 3763
rect 13 3444 19 3476
rect 13 3344 19 3436
rect 125 3384 131 3476
rect 221 3384 227 3496
rect 237 3344 243 3696
rect 301 3644 307 3716
rect 333 3704 339 3736
rect 413 3723 419 3736
rect 413 3717 428 3723
rect 381 3644 387 3716
rect 429 3704 435 3716
rect 333 3524 339 3536
rect 317 3364 323 3476
rect 333 3364 339 3516
rect 349 3504 355 3636
rect 13 3083 19 3336
rect 237 3324 243 3336
rect 125 3184 131 3316
rect 253 3104 259 3316
rect 285 3104 291 3336
rect 349 3104 355 3496
rect 365 3484 371 3496
rect 381 3464 387 3636
rect 445 3504 451 3757
rect 525 3744 531 3776
rect 493 3724 499 3736
rect 381 3323 387 3436
rect 445 3384 451 3456
rect 461 3384 467 3496
rect 461 3364 467 3376
rect 372 3317 387 3323
rect 413 3284 419 3336
rect 493 3324 499 3676
rect 509 3584 515 3696
rect 525 3464 531 3496
rect 557 3484 563 3736
rect 605 3584 611 3716
rect 685 3584 691 4096
rect 717 4044 723 4577
rect 797 4524 803 4536
rect 813 4523 819 4677
rect 829 4584 835 4656
rect 813 4517 828 4523
rect 845 4503 851 4536
rect 829 4497 851 4503
rect 829 4484 835 4497
rect 762 4414 774 4416
rect 747 4406 749 4414
rect 757 4406 759 4414
rect 767 4406 769 4414
rect 777 4406 779 4414
rect 787 4406 789 4414
rect 762 4404 774 4406
rect 733 4304 739 4336
rect 813 4304 819 4356
rect 733 4124 739 4296
rect 781 4284 787 4296
rect 765 4104 771 4276
rect 797 4264 803 4276
rect 829 4264 835 4476
rect 845 4384 851 4416
rect 861 4344 867 4516
rect 861 4284 867 4316
rect 877 4284 883 4897
rect 893 4704 899 4836
rect 909 4744 915 4836
rect 1005 4804 1011 4936
rect 1021 4924 1027 5096
rect 1037 5084 1043 5096
rect 1469 5064 1475 5096
rect 1517 5084 1523 5096
rect 1517 5064 1523 5076
rect 1053 4984 1059 5016
rect 1101 4944 1107 5036
rect 1229 5004 1235 5036
rect 1165 4944 1171 4976
rect 1117 4904 1123 4936
rect 1149 4904 1155 4916
rect 1021 4704 1027 4816
rect 893 4684 899 4696
rect 909 4684 915 4696
rect 925 4664 931 4696
rect 973 4664 979 4696
rect 1005 4684 1011 4696
rect 925 4584 931 4636
rect 957 4624 963 4636
rect 989 4564 995 4596
rect 909 4364 915 4556
rect 1021 4524 1027 4696
rect 1053 4664 1059 4716
rect 909 4304 915 4336
rect 941 4303 947 4516
rect 1053 4504 1059 4656
rect 1069 4623 1075 4896
rect 1197 4784 1203 4816
rect 1117 4704 1123 4736
rect 1213 4704 1219 4756
rect 1085 4644 1091 4696
rect 1133 4664 1139 4676
rect 1165 4644 1171 4696
rect 1069 4617 1091 4623
rect 1021 4384 1027 4396
rect 957 4323 963 4336
rect 1053 4324 1059 4496
rect 1069 4484 1075 4516
rect 957 4317 979 4323
rect 973 4304 979 4317
rect 941 4297 956 4303
rect 797 4184 803 4256
rect 797 4144 803 4156
rect 813 4144 819 4156
rect 813 4084 819 4136
rect 762 4014 774 4016
rect 747 4006 749 4014
rect 757 4006 759 4014
rect 767 4006 769 4014
rect 777 4006 779 4014
rect 787 4006 789 4014
rect 762 4004 774 4006
rect 765 3884 771 3936
rect 829 3884 835 4216
rect 861 4124 867 4236
rect 877 4224 883 4256
rect 909 4244 915 4296
rect 877 4144 883 4176
rect 877 4124 883 4136
rect 893 4124 899 4156
rect 925 4144 931 4256
rect 957 4204 963 4296
rect 1053 4283 1059 4316
rect 1044 4277 1059 4283
rect 973 4264 979 4276
rect 1069 4264 1075 4356
rect 1053 4144 1059 4216
rect 1069 4184 1075 4256
rect 1085 4163 1091 4617
rect 1149 4544 1155 4596
rect 1229 4564 1235 4696
rect 1245 4544 1251 4936
rect 1277 4784 1283 5016
rect 1293 4944 1299 5056
rect 1437 5044 1443 5056
rect 1405 4944 1411 4976
rect 1341 4904 1347 4916
rect 1309 4704 1315 4716
rect 1149 4524 1155 4536
rect 1213 4523 1219 4536
rect 1197 4517 1219 4523
rect 1117 4303 1123 4516
rect 1197 4444 1203 4517
rect 1245 4504 1251 4516
rect 1277 4504 1283 4516
rect 1108 4297 1123 4303
rect 1117 4284 1123 4297
rect 1101 4224 1107 4276
rect 1069 4157 1091 4163
rect 957 4124 963 4136
rect 861 3984 867 4116
rect 925 4104 931 4116
rect 989 4104 995 4116
rect 1005 4104 1011 4116
rect 1037 4064 1043 4116
rect 861 3824 867 3916
rect 957 3904 963 3976
rect 1053 3924 1059 4136
rect 1069 3984 1075 4157
rect 1149 3964 1155 4296
rect 1181 4064 1187 4296
rect 1197 4284 1203 4436
rect 1213 4423 1219 4496
rect 1213 4417 1235 4423
rect 1229 4384 1235 4417
rect 1245 4363 1251 4496
rect 1293 4464 1299 4676
rect 1309 4524 1315 4696
rect 1325 4524 1331 4596
rect 1341 4524 1347 4776
rect 1357 4684 1363 4696
rect 1357 4524 1363 4576
rect 1229 4357 1251 4363
rect 1213 4284 1219 4316
rect 1197 4164 1203 4176
rect 1117 3904 1123 3936
rect 989 3883 995 3896
rect 1037 3884 1043 3896
rect 973 3877 995 3883
rect 877 3784 883 3856
rect 797 3744 803 3756
rect 893 3723 899 3836
rect 909 3784 915 3876
rect 925 3784 931 3856
rect 941 3764 947 3836
rect 884 3717 899 3723
rect 762 3614 774 3616
rect 747 3606 749 3614
rect 757 3606 759 3614
rect 767 3606 769 3614
rect 777 3606 779 3614
rect 787 3606 789 3614
rect 762 3604 774 3606
rect 813 3544 819 3716
rect 845 3684 851 3696
rect 925 3684 931 3736
rect 637 3504 643 3536
rect 557 3364 563 3476
rect 653 3424 659 3496
rect 477 3317 492 3323
rect 93 3084 99 3096
rect 13 3077 35 3083
rect 13 2984 19 3056
rect 13 2644 19 2656
rect 13 2584 19 2596
rect 29 2283 35 3077
rect 77 2923 83 3036
rect 93 2944 99 3076
rect 77 2917 92 2923
rect 109 2864 115 3096
rect 237 2984 243 3096
rect 413 3084 419 3276
rect 429 3104 435 3116
rect 477 3044 483 3317
rect 605 3124 611 3136
rect 557 3084 563 3096
rect 349 2964 355 3036
rect 125 2684 131 2936
rect 221 2924 227 2936
rect 205 2864 211 2916
rect 237 2704 243 2916
rect 253 2704 259 2956
rect 125 2384 131 2676
rect 141 2584 147 2694
rect 221 2603 227 2636
rect 205 2597 227 2603
rect 205 2564 211 2597
rect 237 2444 243 2536
rect 253 2384 259 2696
rect 285 2544 291 2936
rect 301 2924 307 2936
rect 349 2924 355 2956
rect 365 2924 371 3036
rect 429 2944 435 2976
rect 429 2924 435 2936
rect 525 2924 531 2936
rect 301 2884 307 2916
rect 301 2704 307 2856
rect 365 2724 371 2916
rect 445 2904 451 2916
rect 413 2764 419 2836
rect 301 2663 307 2696
rect 317 2684 323 2696
rect 301 2657 323 2663
rect 285 2524 291 2536
rect 253 2304 259 2376
rect 269 2364 275 2516
rect 269 2304 275 2336
rect 301 2304 307 2556
rect 317 2464 323 2657
rect 333 2543 339 2636
rect 365 2624 371 2696
rect 429 2664 435 2696
rect 365 2564 371 2596
rect 397 2584 403 2656
rect 445 2644 451 2896
rect 541 2864 547 2916
rect 461 2784 467 2836
rect 333 2537 355 2543
rect 349 2524 355 2537
rect 461 2504 467 2736
rect 509 2724 515 2836
rect 541 2704 547 2856
rect 573 2744 579 3096
rect 621 3084 627 3116
rect 637 3084 643 3096
rect 621 2964 627 3076
rect 477 2664 483 2696
rect 509 2683 515 2696
rect 509 2677 531 2683
rect 477 2564 483 2656
rect 525 2644 531 2677
rect 573 2664 579 2696
rect 621 2684 627 2936
rect 653 2723 659 3416
rect 685 3403 691 3436
rect 669 3397 691 3403
rect 669 3144 675 3397
rect 749 3384 755 3496
rect 813 3464 819 3476
rect 765 3324 771 3376
rect 701 3284 707 3316
rect 717 3304 723 3316
rect 669 3044 675 3116
rect 685 3104 691 3236
rect 701 3084 707 3136
rect 717 3104 723 3296
rect 762 3214 774 3216
rect 747 3206 749 3214
rect 757 3206 759 3214
rect 767 3206 769 3214
rect 777 3206 779 3214
rect 787 3206 789 3214
rect 762 3204 774 3206
rect 749 3064 755 3096
rect 669 2944 675 2976
rect 717 2924 723 3036
rect 749 2984 755 3056
rect 797 3004 803 3036
rect 797 2964 803 2996
rect 829 2984 835 3496
rect 845 3324 851 3536
rect 877 3484 883 3616
rect 893 3504 899 3516
rect 925 3504 931 3676
rect 941 3624 947 3736
rect 957 3704 963 3716
rect 957 3504 963 3636
rect 861 3104 867 3396
rect 925 3344 931 3496
rect 973 3384 979 3877
rect 989 3724 995 3756
rect 1005 3744 1011 3756
rect 1053 3744 1059 3756
rect 1101 3723 1107 3896
rect 1149 3864 1155 3916
rect 1117 3763 1123 3856
rect 1149 3843 1155 3856
rect 1149 3837 1164 3843
rect 1117 3757 1139 3763
rect 1133 3744 1139 3757
rect 1092 3717 1107 3723
rect 1117 3723 1123 3736
rect 1181 3724 1187 4056
rect 1229 3804 1235 4357
rect 1261 4304 1267 4316
rect 1293 4304 1299 4436
rect 1325 4283 1331 4336
rect 1357 4323 1363 4336
rect 1341 4317 1363 4323
rect 1341 4304 1347 4317
rect 1373 4304 1379 4676
rect 1389 4644 1395 4676
rect 1325 4277 1340 4283
rect 1293 4144 1299 4236
rect 1261 4044 1267 4136
rect 1261 3924 1267 4036
rect 1277 4004 1283 4116
rect 1325 4104 1331 4256
rect 1357 4244 1363 4296
rect 1373 4163 1379 4296
rect 1389 4284 1395 4436
rect 1405 4304 1411 4536
rect 1421 4524 1427 5036
rect 1533 4964 1539 5096
rect 1661 5084 1667 5096
rect 1533 4924 1539 4936
rect 1469 4684 1475 4836
rect 1421 4504 1427 4516
rect 1373 4157 1395 4163
rect 1373 4024 1379 4136
rect 1389 4124 1395 4157
rect 1405 4124 1411 4136
rect 1437 4064 1443 4576
rect 1469 4524 1475 4596
rect 1501 4544 1507 4916
rect 1517 4724 1523 4896
rect 1517 4704 1523 4716
rect 1549 4604 1555 5036
rect 1581 4924 1587 5036
rect 1709 5004 1715 5076
rect 1773 5044 1779 5056
rect 1613 4924 1619 4976
rect 1565 4744 1571 4836
rect 1597 4784 1603 4916
rect 1565 4623 1571 4696
rect 1565 4617 1587 4623
rect 1581 4584 1587 4617
rect 1485 4524 1491 4536
rect 1533 4524 1539 4536
rect 1549 4524 1555 4556
rect 1565 4544 1571 4576
rect 1613 4564 1619 4916
rect 1629 4864 1635 4936
rect 1677 4804 1683 4916
rect 1709 4724 1715 4996
rect 1789 4984 1795 5096
rect 1805 5084 1811 5096
rect 1837 5064 1843 5076
rect 1885 5004 1891 5076
rect 1757 4904 1763 4956
rect 1885 4924 1891 4996
rect 2045 4984 2051 5096
rect 2061 5064 2067 5076
rect 2109 4924 2115 5056
rect 2141 5044 2147 5096
rect 2141 5024 2147 5036
rect 2157 4924 2163 5036
rect 2173 4984 2179 5076
rect 2349 5064 2355 5076
rect 2266 5014 2278 5016
rect 2251 5006 2253 5014
rect 2261 5006 2263 5014
rect 2271 5006 2273 5014
rect 2281 5006 2283 5014
rect 2291 5006 2293 5014
rect 2266 5004 2278 5006
rect 1949 4884 1955 4896
rect 1965 4884 1971 4916
rect 1981 4904 1987 4916
rect 1709 4704 1715 4716
rect 1805 4704 1811 4776
rect 1645 4564 1651 4616
rect 1661 4544 1667 4656
rect 1773 4644 1779 4676
rect 1789 4664 1795 4676
rect 1773 4624 1779 4636
rect 1773 4543 1779 4556
rect 1773 4537 1788 4543
rect 1677 4524 1683 4536
rect 1453 4344 1459 4436
rect 1469 4284 1475 4496
rect 1549 4464 1555 4516
rect 1485 4304 1491 4336
rect 1469 4144 1475 4276
rect 1469 4124 1475 4136
rect 1453 4084 1459 4116
rect 1293 3902 1299 3936
rect 1229 3744 1235 3776
rect 1261 3744 1267 3876
rect 1197 3724 1203 3736
rect 1117 3717 1132 3723
rect 989 3524 995 3616
rect 1037 3504 1043 3716
rect 1069 3624 1075 3696
rect 1101 3664 1107 3717
rect 1133 3704 1139 3716
rect 1204 3697 1219 3703
rect 1053 3504 1059 3516
rect 1085 3504 1091 3536
rect 1117 3504 1123 3536
rect 1037 3464 1043 3476
rect 1053 3404 1059 3436
rect 941 3324 947 3376
rect 1021 3344 1027 3396
rect 1037 3344 1043 3376
rect 1053 3337 1068 3343
rect 1053 3324 1059 3337
rect 877 3304 883 3316
rect 973 3304 979 3316
rect 893 3184 899 3276
rect 845 3064 851 3096
rect 861 2964 867 3096
rect 909 3064 915 3096
rect 941 3064 947 3116
rect 989 3064 995 3076
rect 1005 3064 1011 3096
rect 762 2814 774 2816
rect 747 2806 749 2814
rect 757 2806 759 2814
rect 767 2806 769 2814
rect 777 2806 779 2814
rect 787 2806 789 2814
rect 762 2804 774 2806
rect 653 2717 675 2723
rect 493 2524 499 2536
rect 365 2384 371 2396
rect 413 2384 419 2436
rect 20 2277 35 2283
rect 13 1784 19 1796
rect 13 1384 19 1456
rect 13 1364 19 1376
rect 29 1083 35 2277
rect 196 2257 211 2263
rect 205 2164 211 2257
rect 221 2184 227 2296
rect 260 2277 275 2283
rect 93 2124 99 2136
rect 173 2124 179 2136
rect 77 2084 83 2096
rect 205 2024 211 2156
rect 269 2144 275 2277
rect 301 2164 307 2296
rect 333 2284 339 2296
rect 317 2164 323 2276
rect 461 2184 467 2496
rect 493 2324 499 2516
rect 509 2304 515 2416
rect 525 2283 531 2636
rect 589 2544 595 2616
rect 605 2584 611 2636
rect 637 2524 643 2616
rect 573 2364 579 2516
rect 509 2277 531 2283
rect 477 2164 483 2236
rect 269 2124 275 2136
rect 317 2104 323 2156
rect 333 2124 339 2136
rect 381 2124 387 2136
rect 349 2104 355 2116
rect 397 2104 403 2136
rect 445 2104 451 2156
rect 477 2084 483 2136
rect 413 1984 419 2036
rect 221 1904 227 1916
rect 301 1884 307 1936
rect 509 1904 515 2277
rect 525 2124 531 2236
rect 557 2204 563 2236
rect 557 2184 563 2196
rect 573 2144 579 2256
rect 605 2143 611 2356
rect 621 2284 627 2316
rect 596 2137 611 2143
rect 525 2104 531 2116
rect 541 2084 547 2096
rect 557 1984 563 2096
rect 573 2084 579 2136
rect 605 2084 611 2116
rect 525 1904 531 1956
rect 173 1744 179 1876
rect 205 1864 211 1876
rect 141 1726 147 1736
rect 205 1724 211 1856
rect 301 1764 307 1796
rect 221 1724 227 1736
rect 317 1724 323 1836
rect 109 1504 115 1716
rect 221 1524 227 1696
rect 221 1504 227 1516
rect 333 1504 339 1876
rect 365 1724 371 1836
rect 397 1784 403 1896
rect 525 1864 531 1896
rect 461 1764 467 1856
rect 477 1744 483 1756
rect 381 1724 387 1736
rect 557 1724 563 1916
rect 573 1804 579 1896
rect 621 1884 627 2276
rect 637 2184 643 2296
rect 653 2124 659 2656
rect 669 2144 675 2717
rect 717 2564 723 2636
rect 781 2604 787 2636
rect 813 2524 819 2536
rect 762 2414 774 2416
rect 747 2406 749 2414
rect 757 2406 759 2414
rect 767 2406 769 2414
rect 777 2406 779 2414
rect 787 2406 789 2414
rect 762 2404 774 2406
rect 813 2284 819 2356
rect 829 2324 835 2956
rect 852 2917 867 2923
rect 733 2224 739 2236
rect 685 2144 691 2216
rect 845 2184 851 2796
rect 861 2764 867 2917
rect 877 2844 883 2916
rect 893 2864 899 3036
rect 925 2944 931 2956
rect 973 2944 979 2956
rect 909 2704 915 2916
rect 925 2784 931 2916
rect 941 2704 947 2936
rect 989 2923 995 3056
rect 1005 2964 1011 2996
rect 1037 2964 1043 3316
rect 1060 3297 1084 3303
rect 1069 3102 1075 3176
rect 1101 3084 1107 3476
rect 1117 3464 1123 3496
rect 1181 3484 1187 3496
rect 1140 3337 1155 3343
rect 1117 2983 1123 3136
rect 1133 3064 1139 3316
rect 1149 3284 1155 3337
rect 1197 3304 1203 3336
rect 1213 3324 1219 3697
rect 1261 3643 1267 3736
rect 1261 3637 1283 3643
rect 1245 3464 1251 3494
rect 1277 3484 1283 3637
rect 1325 3503 1331 3896
rect 1389 3884 1395 4056
rect 1421 3904 1427 3956
rect 1485 3904 1491 3996
rect 1357 3844 1363 3856
rect 1341 3564 1347 3796
rect 1389 3644 1395 3876
rect 1405 3744 1411 3896
rect 1469 3864 1475 3876
rect 1437 3584 1443 3696
rect 1341 3524 1347 3556
rect 1453 3544 1459 3836
rect 1485 3763 1491 3896
rect 1501 3784 1507 4256
rect 1517 4124 1523 4316
rect 1613 4304 1619 4336
rect 1661 4304 1667 4396
rect 1581 4284 1587 4296
rect 1533 4144 1539 4236
rect 1565 4124 1571 4236
rect 1597 4224 1603 4296
rect 1629 4204 1635 4276
rect 1677 4204 1683 4516
rect 1725 4503 1731 4536
rect 1821 4524 1827 4576
rect 1716 4497 1731 4503
rect 1741 4384 1747 4396
rect 1757 4304 1763 4376
rect 1693 4224 1699 4296
rect 1581 4124 1587 4136
rect 1517 3984 1523 4116
rect 1517 3924 1523 3936
rect 1533 3884 1539 4016
rect 1613 3944 1619 4156
rect 1629 4124 1635 4196
rect 1709 4144 1715 4296
rect 1789 4224 1795 4516
rect 1805 4304 1811 4416
rect 1837 4384 1843 4716
rect 1869 4704 1875 4736
rect 1949 4704 1955 4776
rect 1853 4664 1859 4676
rect 1901 4624 1907 4696
rect 1917 4684 1923 4696
rect 1940 4677 1955 4683
rect 1869 4524 1875 4576
rect 1853 4283 1859 4296
rect 1853 4277 1875 4283
rect 1741 4124 1747 4136
rect 1789 4124 1795 4196
rect 1869 4184 1875 4277
rect 1885 4224 1891 4236
rect 1821 4144 1827 4156
rect 1629 3984 1635 4116
rect 1725 4084 1731 4116
rect 1645 3884 1651 3894
rect 1469 3757 1491 3763
rect 1469 3724 1475 3757
rect 1501 3624 1507 3636
rect 1469 3544 1475 3616
rect 1453 3504 1459 3536
rect 1325 3497 1347 3503
rect 1309 3484 1315 3496
rect 1245 3344 1251 3376
rect 1277 3344 1283 3476
rect 1213 3304 1219 3316
rect 1309 3304 1315 3318
rect 1149 3244 1155 3276
rect 1197 3144 1203 3216
rect 1197 3124 1203 3136
rect 1101 2977 1123 2983
rect 1213 2983 1219 3076
rect 1213 2977 1228 2983
rect 1069 2944 1075 2976
rect 973 2917 995 2923
rect 957 2904 963 2916
rect 957 2704 963 2856
rect 973 2804 979 2917
rect 1053 2764 1059 2796
rect 909 2664 915 2696
rect 1005 2684 1011 2716
rect 1021 2704 1027 2716
rect 1053 2704 1059 2756
rect 1069 2684 1075 2716
rect 941 2664 947 2676
rect 941 2644 947 2656
rect 861 2324 867 2636
rect 957 2604 963 2676
rect 1021 2644 1027 2656
rect 1028 2637 1043 2643
rect 932 2577 947 2583
rect 941 2564 947 2577
rect 941 2444 947 2556
rect 973 2524 979 2616
rect 1021 2544 1027 2616
rect 1037 2383 1043 2637
rect 1053 2544 1059 2576
rect 1101 2543 1107 2977
rect 1229 2944 1235 2976
rect 1261 2924 1267 3036
rect 1117 2704 1123 2776
rect 1165 2664 1171 2916
rect 1197 2684 1203 2896
rect 1213 2704 1219 2856
rect 1245 2844 1251 2916
rect 1277 2724 1283 3196
rect 1293 3104 1299 3116
rect 1325 3104 1331 3196
rect 1341 3083 1347 3497
rect 1389 3404 1395 3496
rect 1357 3184 1363 3336
rect 1405 3284 1411 3476
rect 1421 3144 1427 3476
rect 1533 3464 1539 3876
rect 1613 3744 1619 3876
rect 1693 3824 1699 3856
rect 1693 3784 1699 3816
rect 1613 3704 1619 3716
rect 1629 3544 1635 3736
rect 1741 3724 1747 4096
rect 1805 3744 1811 4136
rect 1837 4124 1843 4176
rect 1892 4137 1907 4143
rect 1837 3884 1843 4076
rect 1853 4004 1859 4076
rect 1869 4004 1875 4116
rect 1901 4104 1907 4137
rect 1917 4103 1923 4656
rect 1949 4544 1955 4677
rect 1965 4563 1971 4676
rect 1981 4664 1987 4716
rect 1997 4684 2003 4836
rect 2061 4784 2067 4916
rect 2077 4904 2083 4916
rect 2109 4703 2115 4836
rect 2221 4784 2227 4856
rect 2189 4704 2195 4736
rect 2237 4704 2243 4776
rect 2100 4697 2115 4703
rect 2029 4684 2035 4696
rect 2045 4684 2051 4696
rect 1965 4557 1987 4563
rect 1933 4524 1939 4536
rect 1965 4524 1971 4536
rect 1981 4524 1987 4557
rect 1997 4544 2003 4656
rect 2013 4624 2019 4636
rect 2061 4624 2067 4696
rect 2157 4684 2163 4696
rect 2285 4684 2291 4936
rect 2349 4684 2355 5056
rect 2413 5044 2419 5096
rect 2493 5084 2499 5096
rect 2573 5084 2579 5094
rect 2445 5024 2451 5056
rect 2381 4924 2387 4956
rect 2445 4924 2451 5016
rect 2477 4984 2483 5036
rect 2493 5004 2499 5076
rect 2541 5064 2547 5076
rect 2493 4924 2499 4936
rect 2573 4924 2579 4956
rect 2605 4924 2611 5096
rect 2637 4984 2643 5076
rect 2717 5044 2723 5056
rect 2701 5024 2707 5036
rect 2717 5003 2723 5016
rect 2701 4997 2723 5003
rect 2701 4964 2707 4997
rect 2765 4964 2771 5076
rect 2781 4984 2787 5036
rect 2621 4924 2627 4936
rect 2589 4884 2595 4916
rect 2109 4664 2115 4676
rect 2045 4544 2051 4556
rect 2029 4504 2035 4536
rect 2077 4524 2083 4536
rect 2093 4424 2099 4516
rect 2109 4504 2115 4656
rect 2125 4584 2131 4656
rect 2141 4624 2147 4636
rect 2125 4564 2131 4576
rect 2157 4564 2163 4676
rect 1981 4184 1987 4236
rect 1908 4097 1923 4103
rect 1821 3784 1827 3876
rect 1853 3784 1859 3896
rect 1917 3883 1923 3896
rect 1933 3884 1939 4116
rect 1965 3984 1971 3996
rect 1901 3877 1923 3883
rect 1885 3784 1891 3816
rect 1725 3684 1731 3716
rect 1549 3484 1555 3496
rect 1325 3077 1347 3083
rect 1309 3064 1315 3076
rect 1309 3024 1315 3056
rect 1293 2984 1299 2996
rect 1325 2924 1331 3077
rect 1389 3044 1395 3076
rect 1357 2944 1363 3036
rect 1389 2984 1395 3036
rect 1309 2844 1315 2916
rect 1245 2684 1251 2716
rect 1293 2704 1299 2796
rect 1268 2677 1292 2683
rect 1309 2663 1315 2696
rect 1300 2657 1315 2663
rect 1117 2604 1123 2636
rect 1101 2537 1116 2543
rect 1069 2504 1075 2516
rect 1117 2504 1123 2516
rect 1165 2504 1171 2616
rect 1197 2544 1203 2656
rect 1261 2624 1267 2656
rect 1261 2584 1267 2616
rect 1037 2377 1052 2383
rect 989 2304 995 2336
rect 1069 2324 1075 2496
rect 1101 2484 1107 2496
rect 1101 2304 1107 2376
rect 1197 2344 1203 2536
rect 1229 2504 1235 2518
rect 1325 2503 1331 2916
rect 1389 2904 1395 2936
rect 1405 2924 1411 3016
rect 1405 2904 1411 2916
rect 1357 2824 1363 2836
rect 1341 2764 1347 2816
rect 1341 2544 1347 2736
rect 1357 2704 1363 2776
rect 1396 2677 1411 2683
rect 1357 2624 1363 2636
rect 1373 2544 1379 2556
rect 1389 2524 1395 2656
rect 1405 2564 1411 2677
rect 1421 2604 1427 2816
rect 1437 2744 1443 3316
rect 1453 2864 1459 3316
rect 1469 3224 1475 3316
rect 1469 2944 1475 3096
rect 1469 2884 1475 2916
rect 1437 2684 1443 2716
rect 1437 2624 1443 2636
rect 1453 2584 1459 2656
rect 1325 2497 1347 2503
rect 1181 2304 1187 2316
rect 1197 2284 1203 2336
rect 1309 2284 1315 2356
rect 1341 2284 1347 2497
rect 1389 2324 1395 2516
rect 1421 2404 1427 2496
rect 1453 2384 1459 2496
rect 1469 2384 1475 2836
rect 1485 2784 1491 3236
rect 1517 2944 1523 3356
rect 1533 3324 1539 3376
rect 1565 3244 1571 3376
rect 1629 3324 1635 3496
rect 1645 3364 1651 3476
rect 1565 3104 1571 3236
rect 1549 2964 1555 3036
rect 1581 2983 1587 3236
rect 1613 3224 1619 3316
rect 1629 3184 1635 3256
rect 1661 3164 1667 3556
rect 1677 3504 1683 3556
rect 1725 3544 1731 3676
rect 1773 3604 1779 3636
rect 1741 3504 1747 3576
rect 1709 3384 1715 3476
rect 1757 3384 1763 3496
rect 1757 3364 1763 3376
rect 1677 3324 1683 3356
rect 1725 3344 1731 3356
rect 1741 3264 1747 3316
rect 1789 3304 1795 3716
rect 1885 3703 1891 3716
rect 1876 3697 1891 3703
rect 1837 3523 1843 3676
rect 1837 3517 1859 3523
rect 1853 3504 1859 3517
rect 1869 3484 1875 3516
rect 1853 3477 1868 3483
rect 1853 3344 1859 3477
rect 1885 3404 1891 3697
rect 1901 3564 1907 3877
rect 1949 3784 1955 3896
rect 1981 3764 1987 4036
rect 1997 3904 2003 4216
rect 2013 4204 2019 4294
rect 2077 4264 2083 4296
rect 2093 4284 2099 4296
rect 2109 4204 2115 4236
rect 2125 4184 2131 4536
rect 2173 4484 2179 4496
rect 2141 4224 2147 4256
rect 2029 4124 2035 4136
rect 2045 4004 2051 4136
rect 2061 3924 2067 4116
rect 2093 4104 2099 4176
rect 2157 4144 2163 4456
rect 2141 4084 2147 4116
rect 2141 3984 2147 4076
rect 2013 3884 2019 3896
rect 1933 3704 1939 3736
rect 1949 3724 1955 3756
rect 2029 3744 2035 3836
rect 2125 3784 2131 3836
rect 2141 3824 2147 3896
rect 2157 3884 2163 4136
rect 2173 4044 2179 4296
rect 2189 4244 2195 4296
rect 2221 4164 2227 4676
rect 2266 4614 2278 4616
rect 2251 4606 2253 4614
rect 2261 4606 2263 4614
rect 2271 4606 2273 4614
rect 2281 4606 2283 4614
rect 2291 4606 2293 4614
rect 2266 4604 2278 4606
rect 2397 4604 2403 4696
rect 2237 4484 2243 4516
rect 2253 4464 2259 4536
rect 2269 4384 2275 4556
rect 2413 4544 2419 4836
rect 2557 4804 2563 4836
rect 2445 4564 2451 4676
rect 2509 4644 2515 4656
rect 2509 4544 2515 4616
rect 2525 4564 2531 4696
rect 2573 4684 2579 4736
rect 2589 4664 2595 4876
rect 2605 4764 2611 4916
rect 2541 4544 2547 4596
rect 2557 4564 2563 4656
rect 2605 4624 2611 4756
rect 2621 4704 2627 4796
rect 2621 4604 2627 4636
rect 2637 4624 2643 4676
rect 2605 4544 2611 4556
rect 2509 4524 2515 4536
rect 2525 4504 2531 4516
rect 2333 4424 2339 4456
rect 2333 4384 2339 4416
rect 2349 4403 2355 4476
rect 2349 4397 2371 4403
rect 2308 4297 2323 4303
rect 2266 4214 2278 4216
rect 2251 4206 2253 4214
rect 2261 4206 2263 4214
rect 2271 4206 2273 4214
rect 2281 4206 2283 4214
rect 2291 4206 2293 4214
rect 2266 4204 2278 4206
rect 2157 3784 2163 3856
rect 2189 3744 2195 4156
rect 2221 3884 2227 3936
rect 2221 3764 2227 3876
rect 2253 3864 2259 3916
rect 2266 3814 2278 3816
rect 2251 3806 2253 3814
rect 2261 3806 2263 3814
rect 2271 3806 2273 3814
rect 2281 3806 2283 3814
rect 2291 3806 2293 3814
rect 2266 3804 2278 3806
rect 2253 3744 2259 3776
rect 1997 3724 2003 3736
rect 1901 3504 1907 3556
rect 1949 3504 1955 3516
rect 1981 3504 1987 3536
rect 1997 3523 2003 3596
rect 2013 3544 2019 3636
rect 2029 3604 2035 3716
rect 2045 3584 2051 3716
rect 1997 3517 2012 3523
rect 2013 3484 2019 3516
rect 2029 3504 2035 3576
rect 2077 3504 2083 3716
rect 2093 3564 2099 3716
rect 2141 3684 2147 3736
rect 2093 3544 2099 3556
rect 2157 3504 2163 3516
rect 2173 3504 2179 3636
rect 1917 3424 1923 3476
rect 1965 3364 1971 3476
rect 1997 3444 2003 3476
rect 1597 3124 1603 3136
rect 1661 3104 1667 3156
rect 1645 3064 1651 3076
rect 1565 2977 1587 2983
rect 1501 2864 1507 2916
rect 1565 2863 1571 2977
rect 1581 2924 1587 2956
rect 1677 2924 1683 2956
rect 1693 2943 1699 3036
rect 1725 3004 1731 3236
rect 1757 3044 1763 3056
rect 1741 2964 1747 2996
rect 1773 2984 1779 3096
rect 1789 2964 1795 3276
rect 1693 2937 1708 2943
rect 1709 2924 1715 2936
rect 1821 2924 1827 3196
rect 1693 2903 1699 2916
rect 1805 2904 1811 2916
rect 1853 2904 1859 3296
rect 1885 3224 1891 3318
rect 1869 3023 1875 3176
rect 1869 3017 1891 3023
rect 1869 2984 1875 2996
rect 1549 2857 1571 2863
rect 1677 2897 1699 2903
rect 1485 2723 1491 2736
rect 1485 2717 1507 2723
rect 1501 2704 1507 2717
rect 1549 2704 1555 2857
rect 1661 2824 1667 2836
rect 1485 2644 1491 2696
rect 1565 2684 1571 2716
rect 1629 2704 1635 2756
rect 1501 2604 1507 2676
rect 1581 2643 1587 2676
rect 1677 2664 1683 2897
rect 1693 2704 1699 2796
rect 1709 2684 1715 2736
rect 1725 2704 1731 2836
rect 1757 2704 1763 2776
rect 1789 2724 1795 2736
rect 1533 2637 1587 2643
rect 1485 2524 1491 2536
rect 1517 2524 1523 2636
rect 1533 2624 1539 2637
rect 1549 2564 1555 2616
rect 1581 2524 1587 2556
rect 1565 2484 1571 2516
rect 1485 2424 1491 2436
rect 1485 2304 1491 2316
rect 1405 2284 1411 2296
rect 813 2124 819 2136
rect 861 2124 867 2276
rect 1069 2144 1075 2236
rect 1101 2164 1107 2176
rect 1229 2144 1235 2276
rect 653 2084 659 2096
rect 733 2044 739 2076
rect 762 2014 774 2016
rect 747 2006 749 2014
rect 757 2006 759 2014
rect 767 2006 769 2014
rect 777 2006 779 2014
rect 787 2006 789 2014
rect 762 2004 774 2006
rect 669 1864 675 1896
rect 589 1784 595 1796
rect 573 1744 579 1776
rect 589 1764 595 1776
rect 436 1717 451 1723
rect 445 1504 451 1717
rect 557 1704 563 1716
rect 109 1484 115 1496
rect 77 1323 83 1436
rect 125 1424 131 1476
rect 77 1317 92 1323
rect 125 1184 131 1336
rect 173 1324 179 1436
rect 189 1384 195 1476
rect 301 1464 307 1496
rect 285 1344 291 1456
rect 381 1384 387 1436
rect 429 1424 435 1496
rect 445 1484 451 1496
rect 221 1104 227 1336
rect 461 1324 467 1436
rect 365 1184 371 1236
rect 20 1077 35 1083
rect 13 944 19 1076
rect 237 957 252 963
rect 125 684 131 836
rect 157 784 163 936
rect 189 884 195 896
rect 237 824 243 957
rect 269 924 275 996
rect 285 964 291 1094
rect 317 944 323 1036
rect 349 924 355 1056
rect 397 1004 403 1056
rect 461 1024 467 1156
rect 477 1084 483 1336
rect 509 1324 515 1636
rect 605 1504 611 1516
rect 525 1484 531 1496
rect 637 1464 643 1536
rect 653 1504 659 1776
rect 685 1744 691 1896
rect 845 1824 851 2036
rect 845 1744 851 1756
rect 685 1463 691 1736
rect 749 1684 755 1736
rect 762 1614 774 1616
rect 747 1606 749 1614
rect 757 1606 759 1614
rect 767 1606 769 1614
rect 777 1606 779 1614
rect 787 1606 789 1614
rect 762 1604 774 1606
rect 813 1504 819 1716
rect 861 1644 867 2116
rect 877 2064 883 2116
rect 957 2064 963 2136
rect 1133 2124 1139 2136
rect 973 2104 979 2116
rect 893 1704 899 1716
rect 909 1704 915 1716
rect 925 1704 931 2056
rect 973 1924 979 2036
rect 1005 2004 1011 2116
rect 1037 2064 1043 2096
rect 973 1904 979 1916
rect 941 1844 947 1856
rect 957 1844 963 1876
rect 1021 1864 1027 1876
rect 973 1744 979 1816
rect 989 1764 995 1856
rect 1037 1824 1043 2056
rect 1133 1904 1139 1916
rect 989 1744 995 1756
rect 973 1724 979 1736
rect 1005 1724 1011 1736
rect 1069 1724 1075 1736
rect 717 1484 723 1496
rect 669 1457 691 1463
rect 525 1404 531 1456
rect 605 1324 611 1336
rect 653 1324 659 1356
rect 669 1324 675 1457
rect 701 1344 707 1476
rect 749 1404 755 1456
rect 685 1324 691 1336
rect 749 1324 755 1356
rect 813 1324 819 1496
rect 893 1484 899 1676
rect 957 1664 963 1716
rect 1005 1564 1011 1716
rect 1085 1703 1091 1876
rect 1117 1744 1123 1876
rect 1181 1864 1187 2136
rect 1197 2083 1203 2116
rect 1197 2077 1219 2083
rect 1213 1844 1219 2077
rect 1261 1904 1267 1916
rect 1069 1697 1091 1703
rect 1069 1684 1075 1697
rect 1101 1664 1107 1716
rect 1117 1704 1123 1736
rect 1197 1724 1203 1816
rect 1005 1524 1011 1536
rect 1021 1504 1027 1636
rect 1053 1584 1059 1656
rect 893 1364 899 1476
rect 909 1384 915 1496
rect 1069 1444 1075 1616
rect 1133 1584 1139 1716
rect 1149 1684 1155 1716
rect 1149 1584 1155 1656
rect 1181 1604 1187 1636
rect 1213 1624 1219 1836
rect 1277 1764 1283 1956
rect 1325 1924 1331 2036
rect 1373 2024 1379 2256
rect 1405 2204 1411 2276
rect 1389 1904 1395 1916
rect 1229 1684 1235 1716
rect 1117 1524 1123 1556
rect 1117 1504 1123 1516
rect 1245 1504 1251 1676
rect 1309 1603 1315 1876
rect 1357 1844 1363 1876
rect 1389 1824 1395 1836
rect 1357 1764 1363 1796
rect 1405 1743 1411 2156
rect 1421 2124 1427 2256
rect 1437 2164 1443 2276
rect 1469 2184 1475 2276
rect 1485 2244 1491 2276
rect 1485 2224 1491 2236
rect 1437 1884 1443 2116
rect 1501 2104 1507 2476
rect 1549 2284 1555 2396
rect 1565 2304 1571 2336
rect 1533 2204 1539 2236
rect 1533 2124 1539 2136
rect 1453 2044 1459 2096
rect 1549 2064 1555 2276
rect 1469 1964 1475 2036
rect 1517 1984 1523 1996
rect 1549 1984 1555 2056
rect 1453 1904 1459 1916
rect 1421 1744 1427 1796
rect 1453 1744 1459 1896
rect 1485 1864 1491 1936
rect 1565 1924 1571 2216
rect 1597 2203 1603 2436
rect 1629 2404 1635 2636
rect 1661 2624 1667 2656
rect 1645 2524 1651 2536
rect 1613 2204 1619 2276
rect 1629 2264 1635 2316
rect 1661 2264 1667 2316
rect 1677 2304 1683 2636
rect 1725 2544 1731 2636
rect 1741 2324 1747 2676
rect 1773 2544 1779 2696
rect 1805 2663 1811 2896
rect 1885 2864 1891 3017
rect 1901 2944 1907 3096
rect 1933 3063 1939 3096
rect 1949 3084 1955 3096
rect 1981 3084 1987 3316
rect 1997 3224 2003 3236
rect 2013 3184 2019 3456
rect 2045 3343 2051 3476
rect 2141 3444 2147 3476
rect 2061 3384 2067 3416
rect 2045 3337 2067 3343
rect 2029 3324 2035 3336
rect 2045 3264 2051 3316
rect 2061 3224 2067 3337
rect 2157 3324 2163 3496
rect 2173 3484 2179 3496
rect 2189 3484 2195 3736
rect 2045 3104 2051 3136
rect 1933 3057 1948 3063
rect 1933 2924 1939 3016
rect 1965 2924 1971 3036
rect 1981 2944 1987 3076
rect 1997 2944 2003 3096
rect 2061 3044 2067 3096
rect 2061 3024 2067 3036
rect 2077 2963 2083 3136
rect 2173 3124 2179 3476
rect 2253 3444 2259 3456
rect 2189 3326 2195 3436
rect 2266 3414 2278 3416
rect 2251 3406 2253 3414
rect 2261 3406 2263 3414
rect 2271 3406 2273 3414
rect 2281 3406 2283 3414
rect 2291 3406 2293 3414
rect 2266 3404 2278 3406
rect 2317 3324 2323 4297
rect 2365 4284 2371 4397
rect 2397 4344 2403 4496
rect 2509 4444 2515 4476
rect 2397 4324 2403 4336
rect 2365 4164 2371 4276
rect 2397 4124 2403 4296
rect 2461 4284 2467 4336
rect 2525 4304 2531 4416
rect 2477 4284 2483 4296
rect 2429 4184 2435 4256
rect 2445 4184 2451 4276
rect 2461 4264 2467 4276
rect 2493 4224 2499 4276
rect 2525 4264 2531 4276
rect 2477 4144 2483 4176
rect 2541 4164 2547 4516
rect 2621 4424 2627 4516
rect 2573 4204 2579 4256
rect 2589 4184 2595 4256
rect 2573 4144 2579 4156
rect 2333 3824 2339 3976
rect 2397 3964 2403 4116
rect 2461 4104 2467 4116
rect 2557 4104 2563 4116
rect 2365 3864 2371 3896
rect 2381 3764 2387 3876
rect 2349 3744 2355 3756
rect 2333 3464 2339 3496
rect 2077 2957 2099 2963
rect 2061 2924 2067 2936
rect 1821 2684 1827 2696
rect 1837 2684 1843 2836
rect 1853 2684 1859 2836
rect 1885 2704 1891 2796
rect 1901 2684 1907 2696
rect 1933 2684 1939 2916
rect 1949 2684 1955 2716
rect 1965 2704 1971 2816
rect 1805 2657 1827 2663
rect 1821 2544 1827 2657
rect 1837 2604 1843 2676
rect 1853 2584 1859 2656
rect 1901 2644 1907 2676
rect 1933 2643 1939 2656
rect 1917 2637 1939 2643
rect 1917 2584 1923 2637
rect 1917 2544 1923 2576
rect 1965 2564 1971 2636
rect 1789 2484 1795 2518
rect 1821 2443 1827 2536
rect 1805 2437 1827 2443
rect 1773 2343 1779 2376
rect 1773 2337 1795 2343
rect 1741 2304 1747 2316
rect 1773 2304 1779 2316
rect 1789 2304 1795 2337
rect 1709 2284 1715 2296
rect 1581 2197 1603 2203
rect 1581 2024 1587 2197
rect 1597 2126 1603 2176
rect 1629 2004 1635 2196
rect 1693 2144 1699 2276
rect 1709 2224 1715 2276
rect 1725 2244 1731 2276
rect 1741 2264 1747 2296
rect 1709 2144 1715 2156
rect 1693 2124 1699 2136
rect 1709 2083 1715 2136
rect 1741 2124 1747 2236
rect 1757 2124 1763 2296
rect 1709 2077 1724 2083
rect 1581 1904 1587 1996
rect 1661 1964 1667 2076
rect 1661 1917 1715 1923
rect 1661 1904 1667 1917
rect 1517 1784 1523 1856
rect 1389 1737 1411 1743
rect 1325 1724 1331 1736
rect 1309 1597 1331 1603
rect 1261 1504 1267 1516
rect 1277 1504 1283 1516
rect 1085 1484 1091 1496
rect 893 1326 899 1336
rect 509 1163 515 1316
rect 669 1283 675 1316
rect 653 1277 675 1283
rect 653 1184 659 1277
rect 762 1214 774 1216
rect 747 1206 749 1214
rect 757 1206 759 1214
rect 767 1206 769 1214
rect 777 1206 779 1214
rect 787 1206 789 1214
rect 762 1204 774 1206
rect 509 1157 531 1163
rect 381 944 387 976
rect 269 904 275 916
rect 349 884 355 896
rect 253 704 259 836
rect 269 724 275 876
rect 77 524 83 596
rect 125 544 131 676
rect 205 644 211 696
rect 301 644 307 676
rect 317 664 323 816
rect 381 684 387 916
rect 413 824 419 956
rect 429 924 435 936
rect 461 904 467 1016
rect 493 984 499 1096
rect 477 924 483 956
rect 509 944 515 956
rect 413 724 419 796
rect 365 677 380 683
rect 237 604 243 636
rect 125 524 131 536
rect 61 223 67 294
rect 45 217 67 223
rect 45 184 51 217
rect 61 164 67 176
rect 109 144 115 356
rect 125 304 131 516
rect 141 184 147 216
rect 125 164 131 176
rect 189 104 195 316
rect 221 284 227 536
rect 285 524 291 596
rect 301 584 307 636
rect 333 604 339 636
rect 365 484 371 677
rect 381 584 387 596
rect 429 504 435 716
rect 461 684 467 856
rect 525 784 531 1157
rect 589 1044 595 1056
rect 589 944 595 1036
rect 605 944 611 1076
rect 621 964 627 1036
rect 637 944 643 1076
rect 701 1064 707 1116
rect 813 1024 819 1316
rect 909 1104 915 1336
rect 973 1104 979 1136
rect 989 1104 995 1416
rect 1021 1384 1027 1396
rect 1037 1324 1043 1436
rect 1085 1124 1091 1436
rect 1133 1364 1139 1496
rect 1149 1404 1155 1496
rect 1181 1484 1187 1496
rect 1101 1324 1107 1336
rect 1101 1124 1107 1316
rect 1149 1124 1155 1336
rect 1165 1284 1171 1316
rect 1197 1284 1203 1476
rect 1220 1457 1235 1463
rect 1229 1364 1235 1457
rect 1261 1384 1267 1496
rect 1181 1184 1187 1256
rect 1213 1184 1219 1336
rect 1245 1304 1251 1356
rect 1284 1337 1299 1343
rect 1261 1304 1267 1316
rect 1277 1284 1283 1316
rect 1293 1264 1299 1337
rect 1309 1224 1315 1536
rect 1325 1424 1331 1597
rect 1357 1504 1363 1636
rect 1373 1504 1379 1516
rect 1325 1324 1331 1356
rect 1341 1344 1347 1396
rect 1357 1304 1363 1336
rect 1389 1324 1395 1737
rect 1469 1724 1475 1756
rect 1485 1744 1491 1756
rect 1421 1717 1436 1723
rect 1405 1684 1411 1716
rect 1405 1344 1411 1656
rect 1421 1484 1427 1717
rect 1501 1484 1507 1616
rect 1517 1584 1523 1716
rect 1533 1684 1539 1896
rect 1597 1884 1603 1896
rect 1549 1804 1555 1836
rect 1565 1744 1571 1796
rect 1629 1764 1635 1856
rect 1645 1784 1651 1796
rect 1629 1744 1635 1756
rect 1549 1704 1555 1716
rect 1613 1704 1619 1716
rect 1645 1704 1651 1736
rect 1533 1403 1539 1556
rect 1549 1464 1555 1516
rect 1565 1444 1571 1476
rect 1581 1404 1587 1696
rect 1597 1423 1603 1456
rect 1597 1417 1619 1423
rect 1533 1397 1555 1403
rect 1357 1284 1363 1296
rect 861 1084 867 1096
rect 653 944 659 956
rect 548 897 572 903
rect 541 884 547 896
rect 557 784 563 897
rect 605 784 611 916
rect 660 697 675 703
rect 461 604 467 676
rect 477 644 483 676
rect 461 524 467 536
rect 509 524 515 636
rect 589 524 595 696
rect 653 584 659 676
rect 669 664 675 697
rect 669 524 675 656
rect 701 564 707 956
rect 845 944 851 1056
rect 762 814 774 816
rect 747 806 749 814
rect 757 806 759 814
rect 767 806 769 814
rect 777 806 779 814
rect 787 806 789 814
rect 762 804 774 806
rect 861 744 867 1016
rect 909 1004 915 1096
rect 1005 1084 1011 1116
rect 1053 1104 1059 1116
rect 1165 1104 1171 1176
rect 1341 1104 1347 1216
rect 989 1063 995 1076
rect 989 1057 1020 1063
rect 1181 1063 1187 1096
rect 1165 1057 1187 1063
rect 1117 944 1123 996
rect 861 684 867 736
rect 1053 724 1059 736
rect 1101 723 1107 736
rect 1117 724 1123 776
rect 1165 744 1171 1057
rect 1197 784 1203 956
rect 1213 904 1219 1016
rect 1245 1004 1251 1076
rect 1277 984 1283 1094
rect 1357 944 1363 996
rect 1389 984 1395 1316
rect 1405 1284 1411 1336
rect 1421 1324 1427 1376
rect 1421 1104 1427 1316
rect 1469 1303 1475 1336
rect 1517 1324 1523 1356
rect 1533 1344 1539 1376
rect 1549 1324 1555 1397
rect 1581 1384 1587 1396
rect 1597 1363 1603 1396
rect 1572 1357 1603 1363
rect 1613 1344 1619 1417
rect 1460 1297 1475 1303
rect 1437 1084 1443 1096
rect 1405 944 1411 1036
rect 1453 1004 1459 1296
rect 1485 1283 1491 1316
rect 1565 1304 1571 1316
rect 1469 1277 1491 1283
rect 1469 1184 1475 1277
rect 1613 1244 1619 1316
rect 1501 1043 1507 1096
rect 1517 1084 1523 1116
rect 1517 1064 1523 1076
rect 1501 1037 1523 1043
rect 1517 1004 1523 1037
rect 1421 944 1427 956
rect 1517 944 1523 996
rect 1533 983 1539 1216
rect 1629 1123 1635 1416
rect 1645 1363 1651 1636
rect 1661 1444 1667 1496
rect 1677 1484 1683 1816
rect 1693 1784 1699 1896
rect 1709 1884 1715 1917
rect 1709 1763 1715 1836
rect 1700 1757 1715 1763
rect 1693 1744 1699 1756
rect 1709 1724 1715 1736
rect 1725 1664 1731 1716
rect 1741 1584 1747 2096
rect 1773 2004 1779 2136
rect 1805 2104 1811 2437
rect 1853 2323 1859 2516
rect 1869 2504 1875 2516
rect 1981 2503 1987 2896
rect 1997 2524 2003 2856
rect 2061 2844 2067 2916
rect 2077 2884 2083 2936
rect 2013 2704 2019 2736
rect 2029 2684 2035 2836
rect 2013 2624 2019 2676
rect 2045 2664 2051 2696
rect 2029 2657 2044 2663
rect 1981 2497 2003 2503
rect 1917 2384 1923 2476
rect 1853 2317 1875 2323
rect 1869 2304 1875 2317
rect 1837 2224 1843 2296
rect 1853 2284 1859 2296
rect 1885 2284 1891 2296
rect 1837 2124 1843 2196
rect 1821 2044 1827 2116
rect 1853 2064 1859 2276
rect 1933 2244 1939 2296
rect 1885 2104 1891 2136
rect 1901 2124 1907 2136
rect 1789 1743 1795 2036
rect 1821 1884 1827 1896
rect 1805 1824 1811 1876
rect 1837 1764 1843 1976
rect 1869 1924 1875 2036
rect 1869 1904 1875 1916
rect 1933 1884 1939 2076
rect 1901 1784 1907 1876
rect 1917 1763 1923 1796
rect 1901 1757 1923 1763
rect 1853 1744 1859 1756
rect 1789 1737 1811 1743
rect 1805 1724 1811 1737
rect 1901 1724 1907 1757
rect 1924 1737 1939 1743
rect 1773 1664 1779 1716
rect 1805 1684 1811 1716
rect 1933 1704 1939 1737
rect 1805 1523 1811 1676
rect 1821 1657 1836 1663
rect 1821 1604 1827 1657
rect 1933 1604 1939 1696
rect 1837 1584 1843 1596
rect 1949 1584 1955 2416
rect 1965 2404 1971 2436
rect 1965 2324 1971 2336
rect 1965 2264 1971 2316
rect 1997 2304 2003 2497
rect 2013 2484 2019 2496
rect 2029 2423 2035 2657
rect 2045 2524 2051 2636
rect 2061 2604 2067 2736
rect 2093 2704 2099 2957
rect 2109 2863 2115 3116
rect 2173 3103 2179 3116
rect 2164 3097 2179 3103
rect 2125 2964 2131 3096
rect 2141 3044 2147 3096
rect 2157 2964 2163 3016
rect 2125 2944 2131 2956
rect 2173 2924 2179 3056
rect 2125 2884 2131 2916
rect 2173 2864 2179 2916
rect 2221 2864 2227 3276
rect 2317 3204 2323 3316
rect 2333 3143 2339 3456
rect 2349 3444 2355 3596
rect 2381 3524 2387 3756
rect 2397 3704 2403 3736
rect 2413 3704 2419 3716
rect 2429 3684 2435 4076
rect 2461 3904 2467 4096
rect 2509 4084 2515 4096
rect 2573 4063 2579 4136
rect 2557 4057 2579 4063
rect 2509 3904 2515 3916
rect 2557 3864 2563 4057
rect 2605 3944 2611 4296
rect 2637 4284 2643 4616
rect 2653 4424 2659 4796
rect 2669 4584 2675 4916
rect 2701 4804 2707 4956
rect 2765 4944 2771 4956
rect 2781 4924 2787 4936
rect 2829 4784 2835 4916
rect 2861 4884 2867 5096
rect 2973 5024 2979 5036
rect 3053 4984 3059 5096
rect 3085 5084 3091 5096
rect 3357 5084 3363 5096
rect 3453 5084 3459 5096
rect 3661 5084 3667 5096
rect 3005 4964 3011 4976
rect 3037 4944 3043 4956
rect 2893 4937 2908 4943
rect 2893 4924 2899 4937
rect 2893 4704 2899 4916
rect 2909 4804 2915 4916
rect 3021 4804 3027 4916
rect 2957 4704 2963 4756
rect 3069 4704 3075 5076
rect 3149 4984 3155 5036
rect 3117 4964 3123 4976
rect 3085 4924 3091 4956
rect 3149 4924 3155 4976
rect 3197 4924 3203 4936
rect 3245 4924 3251 5036
rect 3293 4924 3299 4936
rect 3341 4924 3347 4976
rect 3357 4964 3363 5076
rect 3389 4924 3395 5056
rect 3469 5044 3475 5056
rect 3476 5037 3491 5043
rect 3421 4924 3427 4976
rect 3485 4924 3491 5037
rect 3517 4944 3523 4956
rect 3549 4924 3555 4996
rect 3597 4944 3603 4996
rect 3629 4944 3635 4976
rect 3133 4884 3139 4916
rect 3229 4903 3235 4916
rect 3229 4897 3251 4903
rect 2685 4664 2691 4696
rect 2701 4664 2707 4676
rect 2685 4543 2691 4656
rect 2717 4564 2723 4676
rect 2861 4584 2867 4656
rect 2893 4644 2899 4696
rect 3053 4683 3059 4696
rect 3165 4684 3171 4696
rect 3053 4677 3075 4683
rect 2941 4644 2947 4676
rect 2676 4537 2691 4543
rect 2653 4304 2659 4416
rect 2669 4304 2675 4536
rect 2701 4464 2707 4516
rect 2717 4504 2723 4536
rect 2733 4524 2739 4536
rect 2925 4523 2931 4636
rect 2989 4564 2995 4676
rect 2925 4517 2940 4523
rect 2717 4384 2723 4496
rect 2765 4344 2771 4436
rect 2781 4324 2787 4496
rect 2829 4364 2835 4456
rect 2685 4304 2691 4316
rect 2829 4304 2835 4356
rect 2845 4304 2851 4516
rect 3053 4504 3059 4516
rect 3069 4504 3075 4677
rect 3149 4644 3155 4656
rect 3149 4544 3155 4636
rect 3181 4523 3187 4836
rect 3229 4704 3235 4876
rect 3197 4564 3203 4656
rect 3213 4584 3219 4676
rect 3213 4544 3219 4576
rect 3181 4517 3203 4523
rect 2893 4323 2899 4476
rect 2925 4464 2931 4496
rect 2893 4317 2915 4323
rect 2669 3964 2675 4276
rect 2621 3924 2627 3936
rect 2445 3744 2451 3776
rect 2525 3744 2531 3856
rect 2589 3843 2595 3896
rect 2573 3837 2595 3843
rect 2509 3704 2515 3718
rect 2429 3544 2435 3676
rect 2573 3664 2579 3837
rect 2621 3724 2627 3916
rect 2621 3604 2627 3716
rect 2445 3524 2451 3536
rect 2381 3484 2387 3516
rect 2349 3384 2355 3436
rect 2349 3324 2355 3356
rect 2365 3344 2371 3476
rect 2381 3424 2387 3476
rect 2397 3384 2403 3496
rect 2445 3484 2451 3496
rect 2477 3484 2483 3536
rect 2509 3443 2515 3476
rect 2493 3437 2515 3443
rect 2365 3204 2371 3336
rect 2381 3304 2387 3356
rect 2493 3344 2499 3437
rect 2509 3324 2515 3376
rect 2637 3343 2643 3456
rect 2621 3337 2643 3343
rect 2621 3324 2627 3337
rect 2653 3324 2659 3896
rect 2669 3883 2675 3936
rect 2685 3904 2691 4296
rect 2733 4264 2739 4276
rect 2813 4264 2819 4296
rect 2861 4263 2867 4296
rect 2893 4284 2899 4296
rect 2836 4257 2867 4263
rect 2797 4204 2803 4256
rect 2813 4184 2819 4256
rect 2829 4184 2835 4196
rect 2909 4144 2915 4317
rect 2925 4284 2931 4456
rect 2989 4304 2995 4416
rect 2909 4124 2915 4136
rect 2701 4084 2707 4116
rect 2781 4083 2787 4116
rect 2765 4077 2787 4083
rect 2669 3877 2684 3883
rect 2685 3524 2691 3636
rect 2701 3584 2707 3876
rect 2717 3724 2723 3796
rect 2749 3724 2755 3776
rect 2749 3504 2755 3516
rect 2733 3484 2739 3496
rect 2765 3484 2771 4077
rect 2781 3904 2787 3916
rect 2781 3864 2787 3876
rect 2813 3823 2819 3976
rect 2909 3904 2915 4116
rect 2941 3944 2947 4296
rect 2957 4264 2963 4276
rect 3005 4264 3011 4296
rect 3021 4184 3027 4296
rect 3037 4284 3043 4296
rect 3053 4244 3059 4496
rect 3085 4304 3091 4336
rect 3117 4304 3123 4436
rect 3133 4384 3139 4436
rect 3149 4364 3155 4516
rect 3197 4424 3203 4517
rect 3245 4523 3251 4897
rect 3405 4884 3411 4916
rect 3261 4624 3267 4716
rect 3236 4517 3251 4523
rect 3197 4304 3203 4356
rect 3229 4324 3235 4516
rect 3261 4464 3267 4496
rect 3117 4224 3123 4276
rect 3021 4144 3027 4156
rect 2957 4104 2963 4118
rect 2989 3904 2995 3976
rect 2813 3817 2835 3823
rect 2669 3477 2684 3483
rect 2669 3363 2675 3477
rect 2685 3384 2691 3396
rect 2669 3357 2691 3363
rect 2333 3137 2355 3143
rect 2237 3084 2243 3116
rect 2266 3014 2278 3016
rect 2251 3006 2253 3014
rect 2261 3006 2263 3014
rect 2271 3006 2273 3014
rect 2281 3006 2283 3014
rect 2291 3006 2293 3014
rect 2266 3004 2278 3006
rect 2349 2943 2355 3137
rect 2381 3102 2387 3156
rect 2477 3124 2483 3236
rect 2445 3104 2451 3116
rect 2509 3083 2515 3316
rect 2541 3144 2547 3236
rect 2573 3124 2579 3136
rect 2509 3077 2531 3083
rect 2333 2937 2355 2943
rect 2109 2857 2131 2863
rect 2125 2784 2131 2857
rect 2157 2704 2163 2756
rect 2077 2624 2083 2636
rect 2061 2544 2067 2596
rect 2013 2417 2035 2423
rect 2013 2324 2019 2417
rect 2013 2284 2019 2316
rect 1981 2124 1987 2196
rect 1997 2124 2003 2136
rect 2013 2103 2019 2116
rect 1988 2097 2019 2103
rect 2029 2044 2035 2236
rect 1965 1904 1971 1916
rect 1965 1724 1971 1876
rect 1997 1864 2003 1876
rect 2029 1764 2035 1976
rect 2061 1902 2067 1916
rect 2061 1824 2067 1856
rect 1981 1744 1987 1756
rect 2045 1744 2051 1756
rect 2061 1724 2067 1736
rect 2077 1723 2083 2256
rect 2093 2244 2099 2296
rect 2109 2144 2115 2676
rect 2125 2544 2131 2676
rect 2141 2544 2147 2696
rect 2173 2584 2179 2836
rect 2205 2804 2211 2836
rect 2173 2544 2179 2576
rect 2141 2504 2147 2516
rect 2157 2464 2163 2536
rect 2189 2404 2195 2636
rect 2205 2564 2211 2696
rect 2221 2584 2227 2696
rect 2266 2614 2278 2616
rect 2251 2606 2253 2614
rect 2261 2606 2263 2614
rect 2271 2606 2273 2614
rect 2281 2606 2283 2614
rect 2291 2606 2293 2614
rect 2266 2604 2278 2606
rect 2333 2583 2339 2937
rect 2333 2577 2355 2583
rect 2333 2544 2339 2556
rect 2349 2524 2355 2577
rect 2173 2304 2179 2316
rect 2189 2204 2195 2336
rect 2205 2244 2211 2296
rect 2269 2264 2275 2296
rect 2221 2224 2227 2236
rect 2266 2214 2278 2216
rect 2251 2206 2253 2214
rect 2261 2206 2263 2214
rect 2271 2206 2273 2214
rect 2281 2206 2283 2214
rect 2291 2206 2293 2214
rect 2266 2204 2278 2206
rect 2317 2183 2323 2496
rect 2365 2384 2371 2856
rect 2381 2523 2387 2976
rect 2397 2924 2403 3076
rect 2509 3044 2515 3056
rect 2461 2944 2467 2976
rect 2493 2924 2499 2936
rect 2397 2684 2403 2916
rect 2413 2684 2419 2696
rect 2429 2664 2435 2916
rect 2525 2784 2531 3077
rect 2541 3044 2547 3096
rect 2589 2984 2595 3096
rect 2541 2924 2547 2956
rect 2573 2924 2579 2936
rect 2621 2924 2627 3296
rect 2637 3264 2643 3316
rect 2653 3204 2659 3316
rect 2637 3104 2643 3176
rect 2653 3144 2659 3176
rect 2653 3084 2659 3136
rect 2669 3104 2675 3116
rect 2637 3024 2643 3036
rect 2557 2884 2563 2916
rect 2621 2904 2627 2916
rect 2429 2584 2435 2656
rect 2509 2544 2515 2676
rect 2452 2537 2467 2543
rect 2381 2517 2396 2523
rect 2381 2504 2387 2517
rect 2381 2324 2387 2436
rect 2397 2284 2403 2376
rect 2381 2263 2387 2276
rect 2445 2264 2451 2516
rect 2461 2384 2467 2537
rect 2573 2524 2579 2596
rect 2589 2524 2595 2836
rect 2477 2304 2483 2316
rect 2493 2284 2499 2456
rect 2525 2424 2531 2516
rect 2621 2444 2627 2516
rect 2637 2504 2643 2996
rect 2653 2984 2659 3036
rect 2669 3004 2675 3096
rect 2653 2624 2659 2936
rect 2669 2784 2675 2956
rect 2685 2944 2691 3357
rect 2701 3324 2707 3476
rect 2733 3404 2739 3476
rect 2781 3463 2787 3816
rect 2813 3724 2819 3796
rect 2829 3724 2835 3817
rect 2845 3704 2851 3836
rect 3021 3824 3027 4116
rect 3085 4104 3091 4196
rect 3133 4004 3139 4136
rect 3149 4104 3155 4116
rect 3197 4104 3203 4256
rect 3197 3984 3203 4096
rect 3037 3924 3043 3956
rect 3245 3944 3251 4036
rect 3181 3902 3187 3936
rect 3245 3884 3251 3916
rect 3261 3904 3267 4416
rect 3277 4184 3283 4836
rect 3293 4704 3299 4736
rect 3309 4523 3315 4836
rect 3357 4724 3363 4836
rect 3325 4704 3331 4716
rect 3341 4624 3347 4676
rect 3373 4664 3379 4696
rect 3405 4624 3411 4876
rect 3517 4724 3523 4776
rect 3453 4704 3459 4716
rect 3309 4517 3324 4523
rect 3293 4504 3299 4516
rect 3341 4464 3347 4536
rect 3373 4444 3379 4516
rect 3389 4504 3395 4616
rect 3421 4603 3427 4696
rect 3549 4684 3555 4696
rect 3565 4684 3571 4836
rect 3613 4804 3619 4916
rect 3629 4784 3635 4876
rect 3581 4704 3587 4736
rect 3645 4724 3651 4776
rect 3661 4664 3667 5076
rect 3677 5004 3683 5076
rect 3725 5004 3731 5096
rect 3757 4984 3763 5056
rect 3789 4944 3795 4956
rect 3725 4824 3731 4936
rect 3853 4924 3859 5216
rect 4221 5184 4227 5257
rect 4461 5184 4467 5257
rect 4509 5184 4515 5257
rect 4685 5184 4691 5257
rect 4765 5224 4771 5263
rect 5325 5257 5347 5263
rect 7469 5257 7491 5263
rect 5325 5184 5331 5257
rect 6778 5214 6790 5216
rect 6763 5206 6765 5214
rect 6773 5206 6775 5214
rect 6783 5206 6785 5214
rect 6793 5206 6795 5214
rect 6803 5206 6805 5214
rect 6778 5204 6790 5206
rect 7469 5184 7475 5257
rect 5533 5144 5539 5156
rect 4637 5104 4643 5136
rect 4957 5124 4963 5136
rect 5437 5124 5443 5136
rect 5133 5117 5148 5123
rect 4781 5104 4787 5116
rect 3901 4964 3907 5076
rect 4093 4984 4099 5056
rect 4141 4944 4147 5096
rect 4253 5084 4259 5096
rect 4173 4944 4179 4976
rect 3949 4924 3955 4936
rect 3770 4814 3782 4816
rect 3755 4806 3757 4814
rect 3765 4806 3767 4814
rect 3775 4806 3777 4814
rect 3785 4806 3787 4814
rect 3795 4806 3797 4814
rect 3770 4804 3782 4806
rect 3837 4784 3843 4896
rect 3677 4684 3683 4696
rect 3693 4684 3699 4736
rect 3709 4704 3715 4756
rect 3837 4724 3843 4776
rect 3853 4703 3859 4916
rect 3917 4884 3923 4896
rect 3933 4864 3939 4916
rect 4045 4903 4051 4936
rect 4061 4924 4067 4936
rect 4077 4924 4083 4936
rect 4045 4897 4067 4903
rect 3997 4864 4003 4896
rect 3837 4697 3859 4703
rect 3725 4684 3731 4696
rect 3405 4597 3427 4603
rect 3405 4584 3411 4597
rect 3421 4504 3427 4536
rect 3325 4424 3331 4436
rect 3437 4384 3443 4516
rect 3405 4304 3411 4356
rect 3309 4184 3315 4296
rect 3277 4124 3283 4156
rect 3325 4144 3331 4296
rect 3421 4284 3427 4296
rect 3389 4244 3395 4276
rect 3373 4237 3388 4243
rect 3373 4164 3379 4237
rect 3293 4124 3299 4136
rect 2877 3744 2883 3776
rect 2941 3744 2947 3756
rect 3149 3744 3155 3876
rect 3261 3824 3267 3836
rect 3213 3764 3219 3776
rect 2797 3544 2803 3636
rect 2861 3504 2867 3516
rect 2765 3457 2787 3463
rect 2749 3344 2755 3416
rect 2701 2984 2707 3316
rect 2733 3184 2739 3296
rect 2749 3144 2755 3336
rect 2765 3324 2771 3457
rect 2845 3444 2851 3496
rect 2765 3204 2771 3316
rect 2781 3104 2787 3156
rect 2717 3084 2723 3096
rect 2733 3084 2739 3096
rect 2781 3084 2787 3096
rect 2797 3084 2803 3096
rect 2829 3063 2835 3116
rect 2829 3057 2844 3063
rect 2797 2964 2803 3056
rect 2701 2924 2707 2936
rect 2717 2904 2723 2936
rect 2717 2784 2723 2896
rect 2765 2884 2771 2916
rect 2829 2904 2835 3036
rect 2845 2984 2851 3056
rect 2845 2944 2851 2956
rect 2861 2944 2867 3296
rect 2877 3104 2883 3576
rect 2893 3504 2899 3716
rect 2925 3704 2931 3716
rect 2893 3384 2899 3496
rect 2909 3484 2915 3556
rect 2941 3464 2947 3736
rect 3229 3717 3244 3723
rect 3197 3704 3203 3716
rect 2957 3504 2963 3576
rect 2989 3504 2995 3536
rect 2973 3484 2979 3496
rect 3021 3484 3027 3496
rect 3053 3484 3059 3556
rect 3101 3544 3107 3676
rect 3149 3584 3155 3696
rect 3101 3504 3107 3516
rect 2925 3364 2931 3456
rect 2909 3084 2915 3316
rect 2941 3104 2947 3196
rect 2973 3184 2979 3476
rect 3005 3343 3011 3476
rect 3069 3463 3075 3496
rect 3053 3457 3075 3463
rect 3005 3337 3027 3343
rect 3021 3324 3027 3337
rect 2957 3104 2963 3136
rect 2989 3124 2995 3236
rect 2861 2924 2867 2936
rect 2717 2724 2723 2776
rect 2669 2603 2675 2636
rect 2653 2597 2675 2603
rect 2653 2564 2659 2597
rect 2685 2563 2691 2636
rect 2669 2557 2691 2563
rect 2669 2524 2675 2557
rect 2685 2524 2691 2536
rect 2701 2504 2707 2536
rect 2381 2257 2403 2263
rect 2301 2177 2323 2183
rect 2301 2124 2307 2177
rect 2381 2124 2387 2156
rect 2068 1717 2083 1723
rect 1965 1704 1971 1716
rect 1789 1517 1811 1523
rect 1789 1504 1795 1517
rect 1645 1357 1667 1363
rect 1645 1284 1651 1336
rect 1661 1324 1667 1357
rect 1677 1224 1683 1476
rect 1725 1384 1731 1396
rect 1757 1384 1763 1456
rect 1693 1304 1699 1376
rect 1709 1324 1715 1356
rect 1773 1324 1779 1436
rect 1789 1364 1795 1456
rect 1805 1344 1811 1496
rect 1885 1484 1891 1496
rect 1837 1343 1843 1436
rect 1828 1337 1843 1343
rect 1613 1117 1635 1123
rect 1613 1104 1619 1117
rect 1645 1104 1651 1116
rect 1597 1084 1603 1096
rect 1581 984 1587 1036
rect 1533 977 1555 983
rect 1549 944 1555 977
rect 1613 964 1619 1096
rect 1492 937 1507 943
rect 1309 924 1315 936
rect 1229 784 1235 876
rect 1261 784 1267 816
rect 1325 784 1331 896
rect 1469 884 1475 936
rect 1485 904 1491 916
rect 1501 883 1507 937
rect 1581 884 1587 918
rect 1501 877 1532 883
rect 1101 717 1116 723
rect 1277 704 1283 716
rect 717 584 723 676
rect 445 384 451 416
rect 525 384 531 516
rect 685 504 691 536
rect 733 504 739 616
rect 765 564 771 656
rect 893 643 899 696
rect 877 637 899 643
rect 589 444 595 496
rect 221 144 227 236
rect 253 224 259 294
rect 269 144 275 276
rect 301 144 307 276
rect 461 184 467 376
rect 589 324 595 436
rect 637 304 643 436
rect 557 264 563 296
rect 653 284 659 456
rect 685 284 691 496
rect 829 484 835 536
rect 845 524 851 636
rect 877 584 883 637
rect 909 524 915 596
rect 717 384 723 476
rect 762 414 774 416
rect 747 406 749 414
rect 757 406 759 414
rect 767 406 769 414
rect 777 406 779 414
rect 787 406 789 414
rect 762 404 774 406
rect 589 264 595 276
rect 557 184 563 256
rect 573 124 579 236
rect 653 184 659 276
rect 669 184 675 276
rect 237 63 243 96
rect 237 57 252 63
rect 253 -23 259 56
rect 717 24 723 316
rect 765 124 771 296
rect 813 264 819 296
rect 765 104 771 116
rect 829 24 835 476
rect 861 244 867 276
rect 845 124 851 236
rect 877 124 883 276
rect 941 44 947 616
rect 989 544 995 696
rect 957 284 963 316
rect 957 184 963 276
rect 973 184 979 236
rect 989 224 995 536
rect 1069 524 1075 696
rect 1149 644 1155 676
rect 1165 664 1171 696
rect 1389 684 1395 696
rect 1117 604 1123 636
rect 1149 584 1155 636
rect 1165 524 1171 656
rect 1197 564 1203 636
rect 1213 584 1219 656
rect 1245 624 1251 656
rect 1293 544 1299 676
rect 1021 504 1027 518
rect 1005 324 1011 336
rect 1037 284 1043 376
rect 1053 304 1059 516
rect 1085 323 1091 336
rect 1085 317 1100 323
rect 1133 284 1139 416
rect 1197 404 1203 536
rect 989 144 995 216
rect 1021 184 1027 276
rect 1165 264 1171 396
rect 1293 344 1299 536
rect 1325 384 1331 416
rect 1357 384 1363 596
rect 1405 564 1411 656
rect 1405 544 1411 556
rect 1437 544 1443 556
rect 1485 523 1491 876
rect 1501 784 1507 836
rect 1501 544 1507 576
rect 1485 517 1507 523
rect 1389 384 1395 456
rect 1421 384 1427 516
rect 1476 497 1491 503
rect 1469 384 1475 396
rect 1485 344 1491 497
rect 1501 384 1507 517
rect 1517 404 1523 536
rect 1549 504 1555 796
rect 1581 584 1587 676
rect 1597 584 1603 876
rect 1613 684 1619 836
rect 1629 764 1635 1096
rect 1693 1084 1699 1276
rect 1725 1124 1731 1136
rect 1645 784 1651 1076
rect 1709 1004 1715 1096
rect 1709 984 1715 996
rect 1757 944 1763 1296
rect 1805 1284 1811 1316
rect 1821 1304 1827 1336
rect 1853 1264 1859 1316
rect 1901 1244 1907 1316
rect 1837 964 1843 1096
rect 1853 1084 1859 1216
rect 1853 944 1859 1076
rect 1741 723 1747 836
rect 1821 784 1827 918
rect 1725 717 1747 723
rect 1725 704 1731 717
rect 1629 504 1635 656
rect 1661 564 1667 656
rect 1677 584 1683 616
rect 1693 544 1699 556
rect 1709 544 1715 656
rect 1789 643 1795 676
rect 1789 637 1811 643
rect 1773 544 1779 556
rect 1645 504 1651 536
rect 1533 384 1539 476
rect 1117 124 1123 236
rect 1149 184 1155 236
rect 1165 164 1171 256
rect 1197 224 1203 256
rect 1133 144 1139 156
rect 1069 104 1075 116
rect 1213 104 1219 196
rect 1261 184 1267 276
rect 1277 104 1283 216
rect 685 -23 691 16
rect 762 14 774 16
rect 747 6 749 14
rect 757 6 759 14
rect 767 6 769 14
rect 777 6 779 14
rect 787 6 789 14
rect 762 4 774 6
rect 845 -17 851 36
rect 973 23 979 96
rect 1021 83 1027 96
rect 1021 77 1036 83
rect 973 17 988 23
rect 829 -23 851 -17
rect 861 -23 867 16
rect 989 -23 995 16
rect 1037 -23 1043 76
rect 1165 -23 1171 36
rect 1213 -23 1219 96
rect 1261 44 1267 96
rect 1277 84 1283 96
rect 1341 44 1347 256
rect 1373 84 1379 256
rect 1389 124 1395 156
rect 1261 -23 1267 36
rect 1405 24 1411 256
rect 1437 224 1443 296
rect 1549 283 1555 496
rect 1597 404 1603 496
rect 1613 324 1619 336
rect 1549 277 1571 283
rect 1469 184 1475 236
rect 1485 204 1491 256
rect 1517 244 1523 256
rect 1517 164 1523 176
rect 1501 104 1507 156
rect 1549 -17 1555 36
rect 1565 24 1571 277
rect 1597 104 1603 156
rect 1629 124 1635 196
rect 1645 144 1651 236
rect 1549 -23 1571 -17
rect 1597 -23 1603 16
rect 1645 -23 1651 36
rect 1677 -23 1683 536
rect 1709 364 1715 516
rect 1725 344 1731 496
rect 1805 324 1811 637
rect 1821 624 1827 696
rect 1853 584 1859 616
rect 1869 564 1875 936
rect 1885 604 1891 1236
rect 1917 1184 1923 1476
rect 1933 1404 1939 1476
rect 1965 1443 1971 1616
rect 1981 1544 1987 1576
rect 1997 1564 2003 1716
rect 2093 1704 2099 1736
rect 2157 1724 2163 1816
rect 2173 1744 2179 2056
rect 2205 1904 2211 2036
rect 2301 1924 2307 2116
rect 2205 1884 2211 1896
rect 2221 1884 2227 1896
rect 2269 1864 2275 1896
rect 2189 1844 2195 1856
rect 2221 1837 2236 1843
rect 2189 1744 2195 1816
rect 2221 1804 2227 1837
rect 2266 1814 2278 1816
rect 2251 1806 2253 1814
rect 2261 1806 2263 1814
rect 2271 1806 2273 1814
rect 2281 1806 2283 1814
rect 2291 1806 2293 1814
rect 2266 1804 2278 1806
rect 2205 1704 2211 1716
rect 2013 1504 2019 1596
rect 2077 1584 2083 1676
rect 2109 1584 2115 1696
rect 2029 1524 2035 1576
rect 1949 1437 1971 1443
rect 1949 1384 1955 1437
rect 1965 1344 1971 1356
rect 1933 804 1939 1056
rect 1949 984 1955 1336
rect 1981 1084 1987 1116
rect 1997 1104 2003 1336
rect 2013 1324 2019 1456
rect 2029 1303 2035 1436
rect 2045 1344 2051 1496
rect 2013 1297 2035 1303
rect 2013 1163 2019 1297
rect 2029 1184 2035 1276
rect 2013 1157 2035 1163
rect 2029 1103 2035 1157
rect 2045 1124 2051 1256
rect 2061 1123 2067 1376
rect 2077 1203 2083 1556
rect 2093 1524 2099 1576
rect 2125 1384 2131 1476
rect 2157 1444 2163 1536
rect 2173 1524 2179 1536
rect 2173 1464 2179 1496
rect 2173 1423 2179 1436
rect 2157 1417 2179 1423
rect 2157 1324 2163 1417
rect 2189 1403 2195 1516
rect 2173 1397 2195 1403
rect 2173 1304 2179 1397
rect 2189 1304 2195 1376
rect 2125 1277 2140 1283
rect 2093 1224 2099 1236
rect 2077 1197 2099 1203
rect 2061 1117 2083 1123
rect 2029 1097 2051 1103
rect 1997 1084 2003 1096
rect 1965 1024 1971 1056
rect 2045 963 2051 1097
rect 2061 1084 2067 1096
rect 2061 984 2067 1016
rect 2077 1004 2083 1117
rect 2093 1024 2099 1197
rect 2109 1124 2115 1196
rect 2125 1144 2131 1277
rect 2157 1184 2163 1296
rect 2173 1204 2179 1236
rect 2189 1184 2195 1236
rect 2205 1144 2211 1536
rect 2221 1523 2227 1696
rect 2253 1624 2259 1716
rect 2269 1604 2275 1656
rect 2301 1584 2307 1656
rect 2221 1517 2243 1523
rect 2237 1464 2243 1517
rect 2253 1464 2259 1576
rect 2285 1484 2291 1576
rect 2301 1444 2307 1476
rect 2317 1444 2323 1736
rect 2333 1644 2339 1816
rect 2349 1744 2355 1876
rect 2381 1724 2387 1956
rect 2397 1724 2403 2257
rect 2452 2257 2467 2263
rect 2461 1904 2467 2257
rect 2541 2244 2547 2436
rect 2637 2364 2643 2436
rect 2733 2384 2739 2676
rect 2749 2664 2755 2696
rect 2781 2684 2787 2696
rect 2797 2684 2803 2896
rect 2845 2784 2851 2916
rect 2813 2684 2819 2696
rect 2797 2544 2803 2556
rect 2765 2504 2771 2516
rect 2493 2184 2499 2236
rect 2500 2177 2515 2183
rect 2509 2144 2515 2177
rect 2589 2124 2595 2156
rect 2605 2144 2611 2356
rect 2621 2284 2627 2296
rect 2621 2184 2627 2256
rect 2541 2104 2547 2116
rect 2525 2024 2531 2076
rect 2605 2064 2611 2136
rect 2653 2124 2659 2216
rect 2669 2124 2675 2136
rect 2717 2124 2723 2196
rect 2765 2163 2771 2496
rect 2756 2157 2771 2163
rect 2541 1904 2547 2016
rect 2429 1884 2435 1896
rect 2541 1884 2547 1896
rect 2461 1864 2467 1876
rect 2413 1784 2419 1836
rect 2557 1804 2563 1896
rect 2589 1864 2595 1896
rect 2557 1784 2563 1796
rect 2461 1764 2467 1776
rect 2381 1664 2387 1676
rect 2397 1524 2403 1696
rect 2413 1684 2419 1696
rect 2413 1523 2419 1576
rect 2429 1544 2435 1696
rect 2477 1584 2483 1676
rect 2557 1584 2563 1776
rect 2589 1726 2595 1836
rect 2669 1784 2675 2096
rect 2797 1924 2803 2316
rect 2829 2284 2835 2776
rect 2861 2704 2867 2836
rect 2877 2704 2883 3056
rect 2893 2964 2899 2976
rect 2941 2964 2947 3096
rect 2941 2924 2947 2956
rect 2845 2683 2851 2696
rect 2845 2677 2860 2683
rect 2877 2664 2883 2676
rect 2893 2544 2899 2756
rect 2925 2664 2931 2696
rect 2941 2684 2947 2796
rect 2957 2704 2963 2936
rect 3005 2844 3011 3316
rect 3037 3204 3043 3236
rect 3053 3184 3059 3457
rect 3069 3224 3075 3316
rect 3037 2924 3043 3136
rect 3053 3044 3059 3176
rect 3069 3124 3075 3136
rect 3085 3084 3091 3456
rect 3101 3324 3107 3436
rect 3117 3364 3123 3496
rect 3181 3424 3187 3636
rect 3197 3524 3203 3696
rect 3092 3077 3107 3083
rect 3037 2764 3043 2916
rect 3021 2704 3027 2736
rect 3053 2704 3059 3036
rect 2925 2604 2931 2636
rect 2861 2526 2867 2536
rect 2957 2504 2963 2696
rect 2973 2644 2979 2696
rect 2973 2564 2979 2636
rect 3053 2584 3059 2656
rect 3069 2644 3075 2696
rect 2989 2564 2995 2576
rect 3005 2544 3011 2576
rect 3005 2504 3011 2516
rect 2829 2224 2835 2276
rect 2845 2244 2851 2296
rect 2813 1984 2819 2076
rect 2829 1944 2835 2216
rect 2845 2204 2851 2236
rect 2861 2124 2867 2336
rect 2909 2284 2915 2296
rect 2893 2164 2899 2196
rect 2877 2023 2883 2136
rect 2861 2017 2883 2023
rect 2797 1904 2803 1916
rect 2861 1884 2867 2017
rect 2893 1984 2899 2136
rect 2573 1584 2579 1716
rect 2509 1544 2515 1556
rect 2525 1544 2531 1556
rect 2557 1524 2563 1536
rect 2413 1517 2428 1523
rect 2266 1414 2278 1416
rect 2251 1406 2253 1414
rect 2261 1406 2263 1414
rect 2271 1406 2273 1414
rect 2281 1406 2283 1414
rect 2291 1406 2293 1414
rect 2266 1404 2278 1406
rect 2221 1324 2227 1396
rect 2333 1344 2339 1456
rect 2381 1384 2387 1456
rect 2141 1117 2172 1123
rect 2141 1104 2147 1117
rect 2125 1084 2131 1096
rect 2045 957 2067 963
rect 1997 924 2003 956
rect 1917 684 1923 696
rect 1917 584 1923 616
rect 1821 557 1836 563
rect 1821 524 1827 557
rect 1869 544 1875 556
rect 1933 544 1939 556
rect 1837 384 1843 536
rect 1885 464 1891 516
rect 1885 424 1891 456
rect 1933 444 1939 536
rect 1773 144 1779 296
rect 1853 124 1859 276
rect 1869 264 1875 316
rect 1949 304 1955 676
rect 1965 504 1971 896
rect 1997 783 2003 916
rect 2013 904 2019 916
rect 2061 903 2067 957
rect 2125 963 2131 1016
rect 2141 984 2147 1016
rect 2084 957 2099 963
rect 2125 957 2147 963
rect 2061 897 2083 903
rect 2052 877 2067 883
rect 2013 784 2019 796
rect 1988 777 2003 783
rect 2061 744 2067 877
rect 2077 784 2083 897
rect 2093 824 2099 957
rect 2029 724 2035 736
rect 2013 624 2019 656
rect 2077 583 2083 756
rect 2109 704 2115 836
rect 2125 763 2131 916
rect 2141 784 2147 957
rect 2157 944 2163 1096
rect 2189 1084 2195 1096
rect 2173 984 2179 996
rect 2189 924 2195 1076
rect 2125 757 2147 763
rect 2141 624 2147 757
rect 2068 577 2083 583
rect 1997 524 2003 556
rect 2077 524 2083 556
rect 2157 543 2163 656
rect 2173 603 2179 876
rect 2205 744 2211 1136
rect 2221 983 2227 1256
rect 2285 1063 2291 1336
rect 2301 1164 2307 1316
rect 2317 1284 2323 1296
rect 2333 1124 2339 1236
rect 2349 1124 2355 1196
rect 2397 1184 2403 1416
rect 2445 1324 2451 1396
rect 2477 1283 2483 1336
rect 2509 1324 2515 1476
rect 2541 1383 2547 1516
rect 2589 1384 2595 1476
rect 2637 1464 2643 1476
rect 2653 1384 2659 1736
rect 2685 1584 2691 1616
rect 2701 1604 2707 1776
rect 2733 1724 2739 1856
rect 2749 1844 2755 1876
rect 2765 1764 2771 1876
rect 2797 1784 2803 1876
rect 2861 1804 2867 1876
rect 2893 1784 2899 1876
rect 2765 1724 2771 1736
rect 2525 1377 2547 1383
rect 2525 1304 2531 1377
rect 2557 1324 2563 1356
rect 2669 1344 2675 1536
rect 2685 1504 2691 1536
rect 2701 1464 2707 1516
rect 2685 1344 2691 1456
rect 2717 1424 2723 1676
rect 2733 1604 2739 1696
rect 2749 1524 2755 1696
rect 2765 1584 2771 1616
rect 2781 1523 2787 1776
rect 2893 1737 2908 1743
rect 2877 1683 2883 1696
rect 2861 1677 2883 1683
rect 2829 1664 2835 1676
rect 2772 1517 2787 1523
rect 2749 1384 2755 1476
rect 2765 1384 2771 1416
rect 2621 1324 2627 1336
rect 2541 1284 2547 1296
rect 2461 1277 2483 1283
rect 2429 1244 2435 1276
rect 2461 1184 2467 1277
rect 2509 1264 2515 1276
rect 2413 1104 2419 1116
rect 2365 1084 2371 1096
rect 2429 1084 2435 1096
rect 2493 1084 2499 1096
rect 2308 1077 2355 1083
rect 2349 1063 2355 1077
rect 2509 1063 2515 1076
rect 2285 1057 2323 1063
rect 2349 1057 2515 1063
rect 2266 1014 2278 1016
rect 2251 1006 2253 1014
rect 2261 1006 2263 1014
rect 2271 1006 2273 1014
rect 2281 1006 2283 1014
rect 2291 1006 2293 1014
rect 2266 1004 2278 1006
rect 2221 977 2243 983
rect 2221 944 2227 956
rect 2221 664 2227 876
rect 2237 784 2243 977
rect 2253 944 2259 956
rect 2317 924 2323 1057
rect 2269 724 2275 796
rect 2333 784 2339 916
rect 2365 904 2371 956
rect 2381 944 2387 956
rect 2372 897 2387 903
rect 2381 684 2387 897
rect 2397 784 2403 996
rect 2413 984 2419 1016
rect 2445 984 2451 1016
rect 2541 984 2547 1096
rect 2557 1004 2563 1296
rect 2573 1184 2579 1196
rect 2589 1024 2595 1276
rect 2621 1204 2627 1316
rect 2653 1277 2668 1283
rect 2653 1224 2659 1277
rect 2685 1263 2691 1336
rect 2733 1324 2739 1336
rect 2797 1304 2803 1616
rect 2861 1584 2867 1677
rect 2877 1524 2883 1576
rect 2893 1563 2899 1737
rect 2909 1584 2915 1716
rect 2925 1584 2931 2336
rect 3005 2324 3011 2496
rect 2973 2184 2979 2294
rect 3085 2164 3091 2996
rect 3101 2524 3107 3077
rect 3117 3004 3123 3356
rect 3133 3344 3139 3356
rect 3149 3344 3155 3356
rect 3197 3343 3203 3516
rect 3213 3484 3219 3496
rect 3229 3444 3235 3717
rect 3261 3703 3267 3716
rect 3245 3697 3267 3703
rect 3245 3684 3251 3697
rect 3213 3364 3219 3436
rect 3245 3384 3251 3496
rect 3277 3484 3283 4116
rect 3293 4044 3299 4116
rect 3293 3704 3299 4036
rect 3325 3884 3331 4136
rect 3405 4124 3411 4196
rect 3453 4124 3459 4596
rect 3469 4524 3475 4616
rect 3469 4364 3475 4516
rect 3485 4444 3491 4536
rect 3501 4524 3507 4636
rect 3533 4564 3539 4576
rect 3581 4544 3587 4636
rect 3597 4524 3603 4656
rect 3677 4544 3683 4676
rect 3773 4544 3779 4676
rect 3501 4304 3507 4316
rect 3469 4284 3475 4296
rect 3517 4264 3523 4296
rect 3565 4284 3571 4296
rect 3581 4284 3587 4436
rect 3485 4164 3491 4236
rect 3485 4144 3491 4156
rect 3549 4124 3555 4136
rect 3389 4044 3395 4116
rect 3501 4104 3507 4116
rect 3565 4104 3571 4276
rect 3581 4184 3587 4276
rect 3597 4244 3603 4516
rect 3645 4324 3651 4456
rect 3770 4414 3782 4416
rect 3755 4406 3757 4414
rect 3765 4406 3767 4414
rect 3775 4406 3777 4414
rect 3785 4406 3787 4414
rect 3795 4406 3797 4414
rect 3770 4404 3782 4406
rect 3652 4317 3667 4323
rect 3613 4304 3619 4316
rect 3661 4284 3667 4317
rect 3725 4304 3731 4336
rect 3821 4304 3827 4316
rect 3677 4284 3683 4296
rect 3725 4264 3731 4276
rect 3581 4144 3587 4176
rect 3837 4124 3843 4697
rect 3949 4702 3955 4716
rect 3885 4664 3891 4676
rect 3981 4584 3987 4676
rect 4045 4584 4051 4876
rect 4061 4644 4067 4897
rect 3869 4544 3875 4556
rect 3853 4384 3859 4456
rect 3869 4304 3875 4436
rect 3933 4384 3939 4516
rect 3981 4384 3987 4536
rect 4013 4384 4019 4516
rect 4061 4504 4067 4556
rect 4093 4544 4099 4696
rect 4109 4584 4115 4896
rect 4125 4864 4131 4896
rect 4132 4857 4147 4863
rect 4125 4704 4131 4756
rect 4141 4724 4147 4857
rect 4157 4683 4163 4716
rect 4173 4704 4179 4916
rect 4189 4684 4195 4776
rect 4205 4764 4211 5036
rect 4237 4926 4243 4956
rect 4253 4784 4259 5076
rect 4317 5064 4323 5094
rect 4349 4944 4355 5076
rect 4493 4984 4499 5096
rect 4301 4924 4307 4936
rect 4349 4744 4355 4936
rect 4429 4904 4435 4918
rect 4365 4804 4371 4836
rect 4253 4702 4259 4716
rect 4157 4677 4179 4683
rect 4141 4563 4147 4636
rect 4173 4584 4179 4677
rect 4132 4557 4147 4563
rect 4093 4524 4099 4536
rect 4029 4384 4035 4496
rect 4077 4464 4083 4516
rect 4141 4484 4147 4516
rect 3901 4204 3907 4296
rect 3949 4204 3955 4296
rect 3437 3904 3443 4036
rect 3309 3864 3315 3876
rect 3325 3804 3331 3836
rect 3357 3784 3363 3896
rect 3389 3884 3395 3896
rect 3421 3784 3427 3896
rect 3341 3764 3347 3776
rect 3453 3764 3459 3836
rect 3501 3744 3507 3776
rect 3485 3737 3500 3743
rect 3309 3724 3315 3736
rect 3325 3724 3331 3736
rect 3405 3724 3411 3736
rect 3293 3504 3299 3596
rect 3261 3464 3267 3476
rect 3197 3337 3212 3343
rect 3133 3124 3139 3336
rect 3204 3317 3219 3323
rect 3213 3164 3219 3317
rect 3229 3264 3235 3316
rect 3245 3304 3251 3316
rect 3261 3163 3267 3436
rect 3309 3324 3315 3636
rect 3341 3524 3347 3596
rect 3373 3584 3379 3716
rect 3389 3644 3395 3716
rect 3325 3484 3331 3516
rect 3325 3344 3331 3356
rect 3357 3324 3363 3576
rect 3405 3484 3411 3536
rect 3437 3502 3443 3516
rect 3405 3464 3411 3476
rect 3373 3424 3379 3456
rect 3485 3424 3491 3737
rect 3549 3724 3555 4096
rect 3885 4044 3891 4096
rect 3901 4044 3907 4116
rect 3965 4104 3971 4176
rect 3981 4123 3987 4236
rect 3997 4184 4003 4316
rect 4045 4284 4051 4396
rect 4205 4364 4211 4516
rect 4237 4384 4243 4456
rect 4269 4323 4275 4496
rect 4285 4384 4291 4556
rect 4317 4544 4323 4556
rect 4349 4544 4355 4736
rect 4301 4524 4307 4536
rect 4260 4317 4275 4323
rect 4173 4304 4179 4316
rect 4045 4164 4051 4276
rect 4109 4244 4115 4294
rect 4061 4184 4067 4236
rect 3997 4124 4003 4136
rect 3981 4117 3996 4123
rect 3770 4014 3782 4016
rect 3755 4006 3757 4014
rect 3765 4006 3767 4014
rect 3775 4006 3777 4014
rect 3785 4006 3787 4014
rect 3795 4006 3797 4014
rect 3770 4004 3782 4006
rect 3885 3924 3891 4036
rect 3949 3902 3955 4036
rect 4013 3964 4019 4136
rect 4093 4124 4099 4196
rect 4125 4124 4131 4136
rect 4253 4124 4259 4296
rect 4029 4064 4035 4116
rect 4077 3984 4083 4076
rect 4093 3903 4099 4116
rect 4237 4084 4243 4116
rect 4269 4104 4275 4317
rect 4301 4304 4307 4516
rect 4381 4484 4387 4636
rect 4301 4264 4307 4276
rect 4301 4184 4307 4236
rect 4317 4224 4323 4296
rect 4333 4284 4339 4296
rect 4333 4124 4339 4276
rect 4365 4244 4371 4256
rect 4397 4164 4403 4556
rect 4445 4544 4451 4656
rect 4541 4564 4547 5096
rect 4589 5044 4595 5096
rect 4605 5084 4611 5096
rect 4653 5064 4659 5096
rect 4797 5084 4803 5116
rect 4765 5064 4771 5076
rect 4829 5064 4835 5116
rect 4877 5104 4883 5116
rect 4925 5064 4931 5076
rect 4557 4984 4563 5036
rect 4797 4924 4803 4936
rect 4621 4884 4627 4918
rect 4589 4704 4595 4796
rect 4749 4784 4755 4836
rect 4733 4684 4739 4696
rect 4573 4543 4579 4636
rect 4557 4537 4579 4543
rect 4445 4324 4451 4536
rect 4525 4483 4531 4516
rect 4516 4477 4531 4483
rect 4445 4284 4451 4316
rect 4525 4283 4531 4477
rect 4557 4444 4563 4537
rect 4589 4304 4595 4636
rect 4637 4544 4643 4676
rect 4653 4584 4659 4616
rect 4669 4584 4675 4636
rect 4765 4584 4771 4896
rect 4797 4724 4803 4836
rect 4813 4704 4819 5056
rect 4829 4964 4835 5036
rect 4957 5004 4963 5036
rect 4973 4984 4979 5036
rect 4861 4944 4867 4956
rect 4893 4944 4899 4976
rect 4989 4944 4995 4996
rect 5005 4984 5011 5096
rect 5069 5064 5075 5076
rect 5133 5064 5139 5117
rect 5229 5084 5235 5096
rect 5341 5084 5347 5096
rect 5373 5083 5379 5116
rect 5517 5104 5523 5116
rect 5469 5084 5475 5096
rect 5373 5077 5388 5083
rect 5389 5064 5395 5076
rect 5037 4964 5043 5036
rect 5274 5014 5286 5016
rect 5259 5006 5261 5014
rect 5269 5006 5271 5014
rect 5279 5006 5281 5014
rect 5289 5006 5291 5014
rect 5299 5006 5301 5014
rect 5274 5004 5286 5006
rect 4877 4904 4883 4916
rect 4797 4624 4803 4676
rect 4797 4584 4803 4616
rect 4669 4544 4675 4576
rect 4781 4564 4787 4576
rect 4765 4544 4771 4556
rect 4813 4524 4819 4696
rect 4829 4564 4835 4836
rect 4845 4604 4851 4636
rect 4861 4583 4867 4696
rect 4909 4644 4915 4656
rect 4845 4577 4867 4583
rect 4829 4524 4835 4556
rect 4621 4464 4627 4516
rect 4845 4484 4851 4577
rect 4884 4537 4899 4543
rect 4605 4304 4611 4436
rect 4701 4424 4707 4436
rect 4749 4304 4755 4476
rect 4813 4344 4819 4356
rect 4861 4343 4867 4476
rect 4845 4337 4867 4343
rect 4781 4304 4787 4316
rect 4829 4304 4835 4336
rect 4845 4324 4851 4337
rect 4877 4323 4883 4516
rect 4868 4317 4883 4323
rect 4893 4304 4899 4537
rect 4925 4384 4931 4836
rect 4973 4764 4979 4796
rect 5053 4784 5059 4916
rect 5149 4904 5155 4936
rect 5069 4784 5075 4876
rect 4973 4704 4979 4756
rect 4957 4624 4963 4636
rect 4941 4504 4947 4556
rect 4941 4304 4947 4436
rect 4957 4404 4963 4436
rect 4525 4277 4547 4283
rect 4349 4144 4355 4156
rect 4125 3944 4131 3976
rect 4205 3964 4211 4036
rect 4125 3904 4131 3936
rect 3821 3884 3827 3896
rect 4077 3897 4099 3903
rect 3501 3664 3507 3716
rect 3533 3704 3539 3716
rect 3533 3684 3539 3696
rect 3565 3544 3571 3796
rect 3597 3744 3603 3756
rect 3645 3684 3651 3876
rect 3677 3643 3683 3716
rect 3725 3704 3731 3716
rect 3661 3637 3683 3643
rect 3373 3344 3379 3416
rect 3364 3317 3379 3323
rect 3357 3284 3363 3296
rect 3277 3224 3283 3236
rect 3261 3157 3283 3163
rect 3181 3084 3187 3096
rect 3197 3084 3203 3156
rect 3245 3104 3251 3116
rect 3261 3064 3267 3116
rect 3277 3104 3283 3157
rect 3165 2924 3171 2996
rect 3229 2944 3235 2956
rect 3213 2904 3219 2936
rect 3245 2924 3251 3036
rect 3277 2944 3283 2956
rect 3261 2924 3267 2936
rect 3293 2924 3299 3036
rect 3325 3024 3331 3036
rect 3341 2963 3347 3256
rect 3373 3204 3379 3317
rect 3405 3317 3420 3323
rect 3389 3184 3395 3316
rect 3405 3304 3411 3317
rect 3341 2957 3363 2963
rect 3357 2924 3363 2957
rect 3373 2924 3379 2956
rect 3117 2704 3123 2736
rect 3133 2704 3139 2776
rect 3229 2764 3235 2816
rect 3245 2784 3251 2916
rect 3229 2704 3235 2756
rect 3261 2684 3267 2916
rect 3277 2684 3283 2694
rect 3117 2544 3123 2676
rect 3261 2544 3267 2596
rect 3229 2504 3235 2516
rect 3229 2464 3235 2496
rect 3181 2384 3187 2436
rect 3117 2304 3123 2376
rect 2941 2064 2947 2116
rect 2941 1984 2947 2056
rect 2957 2024 2963 2136
rect 3037 2124 3043 2156
rect 3181 2144 3187 2336
rect 3229 2304 3235 2396
rect 3261 2384 3267 2536
rect 3277 2444 3283 2536
rect 3309 2524 3315 2896
rect 3325 2884 3331 2916
rect 3341 2664 3347 2736
rect 3357 2643 3363 2736
rect 3373 2724 3379 2836
rect 3373 2704 3379 2716
rect 3341 2637 3363 2643
rect 3341 2564 3347 2637
rect 3357 2564 3363 2616
rect 3389 2604 3395 3096
rect 3421 2864 3427 2916
rect 3405 2784 3411 2836
rect 3437 2744 3443 3156
rect 3469 3104 3475 3376
rect 3485 3344 3491 3356
rect 3501 3344 3507 3496
rect 3565 3484 3571 3536
rect 3581 3504 3587 3616
rect 3453 3084 3459 3096
rect 3469 3044 3475 3096
rect 3485 3084 3491 3316
rect 3501 3304 3507 3336
rect 3533 3324 3539 3336
rect 3581 3324 3587 3476
rect 3613 3404 3619 3496
rect 3661 3484 3667 3637
rect 3693 3502 3699 3516
rect 3661 3464 3667 3476
rect 3629 3443 3635 3456
rect 3629 3437 3651 3443
rect 3597 3324 3603 3356
rect 3613 3344 3619 3396
rect 3645 3344 3651 3437
rect 3501 3144 3507 3296
rect 3476 3037 3491 3043
rect 3469 2924 3475 2996
rect 3485 2743 3491 3037
rect 3517 3003 3523 3316
rect 3549 3124 3555 3236
rect 3565 3104 3571 3176
rect 3581 3104 3587 3196
rect 3517 2997 3539 3003
rect 3517 2924 3523 2936
rect 3533 2924 3539 2997
rect 3549 2924 3555 2936
rect 3565 2924 3571 3096
rect 3629 3064 3635 3096
rect 3597 2943 3603 3036
rect 3597 2937 3619 2943
rect 3613 2924 3619 2937
rect 3533 2784 3539 2876
rect 3549 2804 3555 2916
rect 3565 2903 3571 2916
rect 3597 2904 3603 2916
rect 3629 2904 3635 2936
rect 3565 2897 3587 2903
rect 3565 2783 3571 2876
rect 3549 2777 3571 2783
rect 3485 2737 3507 2743
rect 3421 2684 3427 2716
rect 3405 2584 3411 2676
rect 3357 2544 3363 2556
rect 3277 2303 3283 2436
rect 3309 2424 3315 2516
rect 3325 2344 3331 2436
rect 3277 2297 3292 2303
rect 3277 2284 3283 2297
rect 3325 2264 3331 2276
rect 3261 2144 3267 2236
rect 3341 2184 3347 2496
rect 3373 2464 3379 2516
rect 3421 2503 3427 2576
rect 3437 2564 3443 2616
rect 3453 2584 3459 2636
rect 3469 2504 3475 2696
rect 3485 2684 3491 2716
rect 3501 2704 3507 2737
rect 3549 2524 3555 2777
rect 3565 2704 3571 2716
rect 3581 2704 3587 2897
rect 3597 2604 3603 2836
rect 3629 2564 3635 2756
rect 3645 2563 3651 3256
rect 3661 3004 3667 3216
rect 3693 3184 3699 3336
rect 3677 2944 3683 3136
rect 3709 3104 3715 3656
rect 3693 2984 3699 3056
rect 3709 2964 3715 3096
rect 3709 2944 3715 2956
rect 3677 2924 3683 2936
rect 3693 2924 3699 2936
rect 3661 2903 3667 2916
rect 3661 2897 3683 2903
rect 3661 2704 3667 2716
rect 3677 2684 3683 2897
rect 3693 2704 3699 2856
rect 3709 2784 3715 2856
rect 3645 2557 3660 2563
rect 3581 2524 3587 2536
rect 3412 2497 3427 2503
rect 3485 2484 3491 2516
rect 3389 2304 3395 2436
rect 3405 2304 3411 2356
rect 3421 2324 3427 2436
rect 3341 2164 3347 2176
rect 3373 2144 3379 2296
rect 3117 2124 3123 2136
rect 2989 1984 2995 1996
rect 2957 1784 2963 1876
rect 3005 1864 3011 1996
rect 3037 1984 3043 2096
rect 3005 1724 3011 1836
rect 3069 1724 3075 1916
rect 2989 1604 2995 1676
rect 2893 1557 2915 1563
rect 2829 1484 2835 1516
rect 2845 1484 2851 1496
rect 2829 1304 2835 1456
rect 2877 1344 2883 1376
rect 2893 1344 2899 1476
rect 2909 1384 2915 1557
rect 3005 1523 3011 1596
rect 3021 1584 3027 1696
rect 3069 1664 3075 1676
rect 3133 1624 3139 1676
rect 3149 1584 3155 2136
rect 3165 1904 3171 2036
rect 3181 1884 3187 2136
rect 3213 2104 3219 2118
rect 3277 1984 3283 2116
rect 3309 2084 3315 2116
rect 3357 2084 3363 2116
rect 3389 2044 3395 2296
rect 3421 2284 3427 2296
rect 3437 2144 3443 2456
rect 3469 2344 3475 2436
rect 3501 2323 3507 2516
rect 3485 2317 3507 2323
rect 3469 2284 3475 2316
rect 3437 2124 3443 2136
rect 3469 2126 3475 2136
rect 3405 2024 3411 2036
rect 3277 1897 3292 1903
rect 3181 1784 3187 1856
rect 3229 1784 3235 1876
rect 3021 1544 3027 1556
rect 3037 1544 3043 1556
rect 3053 1524 3059 1576
rect 3133 1524 3139 1536
rect 2996 1517 3011 1523
rect 2925 1363 2931 1516
rect 2941 1484 2947 1516
rect 3037 1504 3043 1516
rect 2941 1464 2947 1476
rect 3053 1403 3059 1516
rect 3069 1464 3075 1476
rect 3037 1397 3059 1403
rect 2909 1357 2931 1363
rect 2669 1257 2691 1263
rect 2589 984 2595 1016
rect 2621 1004 2627 1116
rect 2653 984 2659 1216
rect 2669 1184 2675 1257
rect 2717 1184 2723 1256
rect 2733 1184 2739 1276
rect 2733 1144 2739 1176
rect 2765 1164 2771 1276
rect 2797 1244 2803 1276
rect 2813 1264 2819 1296
rect 2877 1184 2883 1276
rect 2893 1184 2899 1236
rect 2765 1124 2771 1156
rect 2685 984 2691 996
rect 2733 984 2739 1116
rect 2461 944 2467 956
rect 2509 924 2515 976
rect 2749 964 2755 1076
rect 2765 1064 2771 1096
rect 2557 957 2572 963
rect 2557 924 2563 957
rect 2413 904 2419 916
rect 2429 784 2435 876
rect 2461 817 2499 823
rect 2461 784 2467 817
rect 2493 804 2499 817
rect 2477 784 2483 796
rect 2509 764 2515 916
rect 2525 804 2531 916
rect 2573 904 2579 936
rect 2637 924 2643 956
rect 2765 944 2771 956
rect 2781 944 2787 1076
rect 2797 1064 2803 1096
rect 2845 1044 2851 1076
rect 2893 1064 2899 1076
rect 2909 1064 2915 1357
rect 3021 1304 3027 1316
rect 3037 1304 3043 1397
rect 3069 1344 3075 1456
rect 3165 1384 3171 1476
rect 3181 1424 3187 1456
rect 3197 1384 3203 1736
rect 3213 1684 3219 1696
rect 3229 1624 3235 1756
rect 3261 1744 3267 1796
rect 3245 1623 3251 1736
rect 3261 1643 3267 1736
rect 3277 1724 3283 1897
rect 3309 1804 3315 1876
rect 3341 1764 3347 1956
rect 3357 1924 3363 1936
rect 3405 1903 3411 1976
rect 3421 1924 3427 1976
rect 3405 1897 3427 1903
rect 3373 1804 3379 1876
rect 3421 1864 3427 1897
rect 3437 1804 3443 1876
rect 3469 1764 3475 2036
rect 3485 1924 3491 2317
rect 3517 2284 3523 2376
rect 3549 2324 3555 2496
rect 3581 2484 3587 2516
rect 3581 2404 3587 2476
rect 3597 2304 3603 2416
rect 3629 2383 3635 2476
rect 3613 2377 3635 2383
rect 3533 2244 3539 2296
rect 3549 2284 3555 2296
rect 3549 2264 3555 2276
rect 3581 2244 3587 2256
rect 3565 2184 3571 2236
rect 3597 2203 3603 2296
rect 3581 2197 3603 2203
rect 3565 1923 3571 2096
rect 3581 2023 3587 2197
rect 3613 2183 3619 2377
rect 3636 2317 3644 2323
rect 3629 2284 3635 2316
rect 3597 2177 3619 2183
rect 3597 2063 3603 2177
rect 3629 2123 3635 2276
rect 3661 2164 3667 2536
rect 3677 2524 3683 2556
rect 3677 2304 3683 2356
rect 3693 2304 3699 2596
rect 3709 2484 3715 2676
rect 3725 2663 3731 3636
rect 3770 3614 3782 3616
rect 3755 3606 3757 3614
rect 3765 3606 3767 3614
rect 3775 3606 3777 3614
rect 3785 3606 3787 3614
rect 3795 3606 3797 3614
rect 3770 3604 3782 3606
rect 3757 3344 3763 3476
rect 3789 3326 3795 3336
rect 3821 3324 3827 3876
rect 3869 3864 3875 3876
rect 3901 3724 3907 3836
rect 3965 3764 3971 3876
rect 3869 3504 3875 3636
rect 3901 3583 3907 3716
rect 3892 3577 3907 3583
rect 3901 3484 3907 3496
rect 3917 3384 3923 3676
rect 3933 3504 3939 3516
rect 3949 3484 3955 3616
rect 3965 3484 3971 3496
rect 3981 3463 3987 3716
rect 4020 3517 4035 3523
rect 4013 3504 4019 3516
rect 3965 3457 3987 3463
rect 3965 3384 3971 3457
rect 3933 3324 3939 3336
rect 3949 3324 3955 3336
rect 3770 3214 3782 3216
rect 3755 3206 3757 3214
rect 3765 3206 3767 3214
rect 3775 3206 3777 3214
rect 3785 3206 3787 3214
rect 3795 3206 3797 3214
rect 3770 3204 3782 3206
rect 3741 3044 3747 3056
rect 3741 2964 3747 2976
rect 3757 2884 3763 3176
rect 3821 2984 3827 3096
rect 3837 3024 3843 3096
rect 3853 3084 3859 3316
rect 3770 2814 3782 2816
rect 3755 2806 3757 2814
rect 3765 2806 3767 2814
rect 3775 2806 3777 2814
rect 3785 2806 3787 2814
rect 3795 2806 3797 2814
rect 3770 2804 3782 2806
rect 3757 2664 3763 2716
rect 3837 2684 3843 2836
rect 3869 2664 3875 2694
rect 3725 2657 3747 2663
rect 3725 2564 3731 2636
rect 3741 2544 3747 2657
rect 3789 2464 3795 2536
rect 3821 2526 3827 2556
rect 3770 2414 3782 2416
rect 3755 2406 3757 2414
rect 3765 2406 3767 2414
rect 3775 2406 3777 2414
rect 3785 2406 3787 2414
rect 3795 2406 3797 2414
rect 3770 2404 3782 2406
rect 3725 2284 3731 2356
rect 3709 2264 3715 2276
rect 3693 2144 3699 2256
rect 3661 2124 3667 2136
rect 3613 2117 3635 2123
rect 3613 2104 3619 2117
rect 3677 2103 3683 2136
rect 3661 2097 3683 2103
rect 3597 2057 3619 2063
rect 3581 2017 3603 2023
rect 3581 1984 3587 1996
rect 3556 1917 3571 1923
rect 3533 1864 3539 1876
rect 3501 1784 3507 1836
rect 3277 1684 3283 1716
rect 3261 1637 3283 1643
rect 3245 1617 3267 1623
rect 3213 1384 3219 1496
rect 3245 1484 3251 1496
rect 3261 1384 3267 1617
rect 3277 1544 3283 1637
rect 3293 1344 3299 1436
rect 3309 1384 3315 1676
rect 3373 1524 3379 1756
rect 3469 1724 3475 1736
rect 3549 1724 3555 1816
rect 3565 1744 3571 1756
rect 3373 1503 3379 1516
rect 3469 1504 3475 1596
rect 3501 1504 3507 1676
rect 3364 1497 3379 1503
rect 3053 1284 3059 1296
rect 2973 1204 2979 1276
rect 3021 1264 3027 1276
rect 2973 1184 2979 1196
rect 2813 964 2819 1016
rect 2909 983 2915 1056
rect 2900 977 2915 983
rect 2877 944 2883 976
rect 2941 964 2947 1136
rect 3021 1104 3027 1116
rect 2765 924 2771 936
rect 2589 864 2595 916
rect 2605 784 2611 796
rect 2669 784 2675 916
rect 2397 644 2403 696
rect 2445 664 2451 696
rect 2461 644 2467 696
rect 2266 614 2278 616
rect 2251 606 2253 614
rect 2261 606 2263 614
rect 2271 606 2273 614
rect 2281 606 2283 614
rect 2291 606 2293 614
rect 2266 604 2278 606
rect 2173 597 2195 603
rect 2189 584 2195 597
rect 2196 577 2211 583
rect 2173 564 2179 576
rect 2205 564 2211 577
rect 2189 544 2195 556
rect 2141 537 2163 543
rect 2013 504 2019 516
rect 1965 364 1971 496
rect 2029 344 2035 496
rect 2045 424 2051 516
rect 1933 284 1939 294
rect 1949 284 1955 296
rect 1949 164 1955 276
rect 2045 204 2051 416
rect 2141 404 2147 537
rect 2173 424 2179 536
rect 2157 384 2163 416
rect 2077 324 2083 376
rect 2061 244 2067 296
rect 2141 284 2147 316
rect 2189 284 2195 536
rect 2221 444 2227 596
rect 2317 584 2323 616
rect 2461 584 2467 636
rect 2365 544 2371 556
rect 2061 164 2067 236
rect 2077 144 2083 176
rect 2093 163 2099 276
rect 2141 184 2147 276
rect 2205 264 2211 396
rect 2381 384 2387 416
rect 2365 304 2371 316
rect 2237 284 2243 296
rect 2365 244 2371 276
rect 2397 264 2403 396
rect 2461 344 2467 536
rect 2477 384 2483 516
rect 2493 384 2499 736
rect 2525 624 2531 716
rect 2557 624 2563 656
rect 2573 644 2579 656
rect 2557 384 2563 518
rect 2653 464 2659 656
rect 2701 564 2707 676
rect 2781 543 2787 936
rect 2909 924 2915 956
rect 2957 924 2963 1036
rect 2973 944 2979 1036
rect 3005 964 3011 1096
rect 3053 1044 3059 1056
rect 3060 1037 3075 1043
rect 3069 1024 3075 1037
rect 3069 964 3075 1016
rect 3101 984 3107 1276
rect 3117 1184 3123 1276
rect 3133 1264 3139 1336
rect 3245 1304 3251 1336
rect 3181 1124 3187 1276
rect 3245 1264 3251 1296
rect 3277 1184 3283 1336
rect 3309 1324 3315 1376
rect 3325 1264 3331 1476
rect 3341 1464 3347 1476
rect 3341 1304 3347 1376
rect 3389 1364 3395 1436
rect 3373 1343 3379 1356
rect 3373 1337 3411 1343
rect 3405 1323 3411 1337
rect 3405 1317 3427 1323
rect 3421 1303 3427 1317
rect 3421 1297 3436 1303
rect 3485 1303 3491 1316
rect 3476 1297 3491 1303
rect 3405 1284 3411 1296
rect 3277 1144 3283 1176
rect 3309 1124 3315 1176
rect 3133 1064 3139 1076
rect 3181 1063 3187 1116
rect 3197 1084 3203 1096
rect 3261 1077 3276 1083
rect 3181 1057 3196 1063
rect 3165 1024 3171 1056
rect 3085 964 3091 976
rect 2989 937 3004 943
rect 2861 844 2867 916
rect 2989 844 2995 937
rect 3101 943 3107 976
rect 3092 937 3107 943
rect 3005 917 3020 923
rect 3005 904 3011 917
rect 3069 903 3075 936
rect 3117 924 3123 956
rect 3149 944 3155 1016
rect 3197 964 3203 1036
rect 3229 1024 3235 1036
rect 3229 964 3235 976
rect 3028 897 3075 903
rect 3181 884 3187 896
rect 2909 704 2915 736
rect 2861 644 2867 656
rect 2829 544 2835 556
rect 2772 537 2787 543
rect 2877 524 2883 616
rect 2893 524 2899 696
rect 2957 684 2963 836
rect 3101 804 3107 836
rect 3229 784 3235 836
rect 3149 737 3164 743
rect 2989 544 2995 676
rect 3005 664 3011 696
rect 2509 304 2515 316
rect 2266 214 2278 216
rect 2251 206 2253 214
rect 2261 206 2263 214
rect 2271 206 2273 214
rect 2281 206 2283 214
rect 2291 206 2293 214
rect 2266 204 2278 206
rect 2148 177 2163 183
rect 2157 164 2163 177
rect 2093 157 2108 163
rect 2141 144 2147 156
rect 2173 144 2179 156
rect 2301 124 2307 156
rect 1757 84 1763 118
rect 2212 117 2236 123
rect 1965 84 1971 116
rect 2317 84 2323 236
rect 2413 184 2419 256
rect 2461 244 2467 276
rect 2509 184 2515 296
rect 2429 164 2435 176
rect 2461 144 2467 176
rect 2541 124 2547 256
rect 2557 223 2563 296
rect 2621 284 2627 336
rect 2637 264 2643 296
rect 2653 284 2659 316
rect 2685 304 2691 436
rect 2733 424 2739 516
rect 2797 484 2803 496
rect 2765 264 2771 336
rect 2813 284 2819 316
rect 2573 244 2579 256
rect 2589 244 2595 256
rect 2557 217 2579 223
rect 2557 144 2563 176
rect 2573 124 2579 217
rect 2589 184 2595 236
rect 2621 164 2627 196
rect 2669 144 2675 236
rect 2813 204 2819 276
rect 2877 264 2883 396
rect 2893 304 2899 516
rect 2829 184 2835 196
rect 2877 184 2883 216
rect 2893 184 2899 296
rect 2909 284 2915 416
rect 2925 184 2931 516
rect 2989 324 2995 436
rect 2973 284 2979 296
rect 2957 204 2963 276
rect 2989 264 2995 276
rect 3021 264 3027 676
rect 3037 564 3043 656
rect 3069 644 3075 676
rect 3085 664 3091 676
rect 3101 624 3107 696
rect 3117 684 3123 696
rect 3069 584 3075 596
rect 3117 544 3123 556
rect 3117 344 3123 356
rect 3133 344 3139 636
rect 3149 604 3155 737
rect 3229 704 3235 716
rect 3165 584 3171 636
rect 3181 584 3187 696
rect 3213 644 3219 696
rect 3149 524 3155 556
rect 3165 384 3171 516
rect 3181 504 3187 556
rect 3197 324 3203 576
rect 3229 544 3235 676
rect 3213 344 3219 476
rect 3213 324 3219 336
rect 2701 104 2707 156
rect 2733 104 2739 156
rect 2845 144 2851 156
rect 2925 144 2931 176
rect 2893 124 2899 136
rect 3005 124 3011 236
rect 3037 224 3043 316
rect 3124 297 3139 303
rect 3053 264 3059 296
rect 3117 184 3123 276
rect 3085 163 3091 176
rect 3133 164 3139 297
rect 3085 157 3100 163
rect 3213 104 3219 236
rect 3229 204 3235 536
rect 3245 404 3251 1036
rect 3261 944 3267 1077
rect 3325 1044 3331 1256
rect 3341 1097 3356 1103
rect 3277 924 3283 936
rect 3261 904 3267 916
rect 3293 884 3299 916
rect 3309 904 3315 1036
rect 3325 964 3331 976
rect 3341 964 3347 1097
rect 3373 1064 3379 1156
rect 3517 1143 3523 1676
rect 3533 1644 3539 1696
rect 3533 1584 3539 1636
rect 3549 1444 3555 1656
rect 3549 1324 3555 1376
rect 3565 1364 3571 1556
rect 3581 1464 3587 1816
rect 3597 1803 3603 2017
rect 3613 1924 3619 2057
rect 3661 1804 3667 2097
rect 3693 2044 3699 2136
rect 3677 1944 3683 2036
rect 3709 1984 3715 2156
rect 3725 1924 3731 2216
rect 3757 2124 3763 2296
rect 3789 2104 3795 2276
rect 3821 2084 3827 2396
rect 3885 2383 3891 2996
rect 3901 2764 3907 3236
rect 3933 3104 3939 3276
rect 3949 3104 3955 3316
rect 3981 3124 3987 3436
rect 3997 3124 4003 3296
rect 3949 3084 3955 3096
rect 3997 3084 4003 3116
rect 3933 2944 3939 3076
rect 3981 2924 3987 3076
rect 3901 2664 3907 2716
rect 3981 2564 3987 2756
rect 4029 2623 4035 3517
rect 4045 3464 4051 3616
rect 4061 3504 4067 3716
rect 4045 3344 4051 3416
rect 4061 3344 4067 3376
rect 4077 3343 4083 3897
rect 4141 3864 4147 3936
rect 4093 3784 4099 3816
rect 4157 3783 4163 3876
rect 4141 3777 4163 3783
rect 4141 3744 4147 3777
rect 4173 3764 4179 3936
rect 4237 3904 4243 3956
rect 4269 3884 4275 3996
rect 4365 3964 4371 4116
rect 4285 3884 4291 3956
rect 4269 3864 4275 3876
rect 4365 3784 4371 3836
rect 4381 3763 4387 4136
rect 4397 4004 4403 4156
rect 4509 4124 4515 4196
rect 4525 4164 4531 4256
rect 4541 4224 4547 4277
rect 4573 4264 4579 4276
rect 4557 4204 4563 4236
rect 4605 4164 4611 4276
rect 4621 4124 4627 4236
rect 4653 4124 4659 4296
rect 4708 4257 4723 4263
rect 4685 4123 4691 4236
rect 4685 4117 4700 4123
rect 4461 3964 4467 4036
rect 4477 3944 4483 4036
rect 4397 3904 4403 3916
rect 4413 3884 4419 3916
rect 4493 3897 4524 3903
rect 4397 3864 4403 3876
rect 4445 3863 4451 3896
rect 4461 3884 4467 3896
rect 4493 3883 4499 3897
rect 4477 3877 4499 3883
rect 4477 3863 4483 3877
rect 4445 3857 4483 3863
rect 4372 3757 4387 3763
rect 4157 3743 4163 3756
rect 4285 3744 4291 3756
rect 4157 3737 4179 3743
rect 4141 3724 4147 3736
rect 4173 3724 4179 3737
rect 4093 3464 4099 3536
rect 4109 3384 4115 3636
rect 4237 3524 4243 3596
rect 4301 3524 4307 3636
rect 4349 3523 4355 3756
rect 4365 3544 4371 3756
rect 4381 3724 4387 3736
rect 4397 3664 4403 3856
rect 4340 3517 4355 3523
rect 4141 3504 4147 3516
rect 4205 3444 4211 3496
rect 4253 3464 4259 3496
rect 4269 3484 4275 3496
rect 4317 3444 4323 3496
rect 4413 3484 4419 3536
rect 4429 3524 4435 3836
rect 4445 3584 4451 3736
rect 4477 3664 4483 3736
rect 4493 3724 4499 3756
rect 4509 3724 4515 3836
rect 4541 3744 4547 3876
rect 4573 3864 4579 3876
rect 4557 3763 4563 3836
rect 4605 3764 4611 4036
rect 4653 3964 4659 4116
rect 4621 3904 4627 3956
rect 4557 3757 4579 3763
rect 4365 3464 4371 3476
rect 4429 3464 4435 3496
rect 4445 3484 4451 3496
rect 4125 3364 4131 3436
rect 4141 3364 4147 3396
rect 4237 3383 4243 3436
rect 4237 3377 4259 3383
rect 4109 3344 4115 3356
rect 4077 3337 4099 3343
rect 4061 3184 4067 3316
rect 4077 3184 4083 3316
rect 4061 3103 4067 3176
rect 4093 3104 4099 3337
rect 4205 3324 4211 3336
rect 4052 3097 4067 3103
rect 4045 3064 4051 3076
rect 4093 2904 4099 3096
rect 4109 3064 4115 3116
rect 4173 3104 4179 3276
rect 4189 3104 4195 3316
rect 4221 3104 4227 3176
rect 4237 3124 4243 3356
rect 4253 3324 4259 3377
rect 4269 3324 4275 3356
rect 4333 3323 4339 3436
rect 4349 3364 4355 3396
rect 4365 3364 4371 3396
rect 4324 3317 4339 3323
rect 4269 3204 4275 3236
rect 4333 3144 4339 3236
rect 4301 3124 4307 3136
rect 4125 2944 4131 3036
rect 4141 3024 4147 3056
rect 4189 2924 4195 3096
rect 4221 2924 4227 3096
rect 4237 3084 4243 3096
rect 4253 3084 4259 3096
rect 4285 3064 4291 3096
rect 4317 3084 4323 3096
rect 4253 2984 4259 2996
rect 4317 2984 4323 3056
rect 4333 2964 4339 2996
rect 4285 2884 4291 2916
rect 4013 2617 4035 2623
rect 3997 2524 4003 2576
rect 3869 2377 3891 2383
rect 3869 2244 3875 2377
rect 3885 2304 3891 2356
rect 3917 2284 3923 2476
rect 3949 2302 3955 2336
rect 3917 2164 3923 2276
rect 3837 2044 3843 2116
rect 3853 2084 3859 2136
rect 3770 2014 3782 2016
rect 3755 2006 3757 2014
rect 3765 2006 3767 2014
rect 3775 2006 3777 2014
rect 3785 2006 3787 2014
rect 3795 2006 3797 2014
rect 3770 2004 3782 2006
rect 3741 1924 3747 1976
rect 3821 1944 3827 1996
rect 3837 1964 3843 2016
rect 3709 1824 3715 1876
rect 3597 1797 3619 1803
rect 3597 1764 3603 1776
rect 3613 1724 3619 1797
rect 3693 1784 3699 1796
rect 3741 1784 3747 1816
rect 3725 1744 3731 1756
rect 3821 1744 3827 1876
rect 3869 1764 3875 2036
rect 3869 1724 3875 1756
rect 3885 1744 3891 1836
rect 3661 1704 3667 1716
rect 3597 1604 3603 1636
rect 3661 1584 3667 1676
rect 3709 1624 3715 1716
rect 3725 1584 3731 1636
rect 3770 1614 3782 1616
rect 3755 1606 3757 1614
rect 3765 1606 3767 1614
rect 3775 1606 3777 1614
rect 3785 1606 3787 1614
rect 3795 1606 3797 1614
rect 3770 1604 3782 1606
rect 3805 1524 3811 1556
rect 3597 1504 3603 1516
rect 3725 1504 3731 1516
rect 3613 1437 3628 1443
rect 3581 1343 3587 1436
rect 3597 1364 3603 1376
rect 3565 1337 3587 1343
rect 3501 1137 3523 1143
rect 3501 1124 3507 1137
rect 3421 1104 3427 1116
rect 3405 1064 3411 1076
rect 3469 1064 3475 1076
rect 3517 1064 3523 1116
rect 3357 964 3363 996
rect 3373 984 3379 996
rect 3389 964 3395 1036
rect 3421 944 3427 1056
rect 3261 684 3267 876
rect 3389 724 3395 736
rect 3309 717 3324 723
rect 3261 564 3267 656
rect 3277 584 3283 696
rect 3293 684 3299 716
rect 3293 624 3299 636
rect 3277 524 3283 576
rect 3309 564 3315 717
rect 3325 704 3331 716
rect 3341 664 3347 676
rect 3357 663 3363 716
rect 3380 697 3395 703
rect 3348 657 3363 663
rect 3277 484 3283 516
rect 3373 504 3379 676
rect 3389 644 3395 697
rect 3277 304 3283 436
rect 3341 384 3347 476
rect 3373 464 3379 496
rect 3325 324 3331 356
rect 3357 304 3363 436
rect 3277 277 3292 283
rect 3261 144 3267 276
rect 3277 124 3283 277
rect 3357 264 3363 276
rect 3357 184 3363 256
rect 3373 224 3379 456
rect 3389 304 3395 636
rect 3405 263 3411 696
rect 3421 684 3427 716
rect 3421 664 3427 676
rect 3437 643 3443 696
rect 3421 637 3443 643
rect 3421 584 3427 637
rect 3437 304 3443 476
rect 3453 284 3459 1036
rect 3485 944 3491 1056
rect 3492 917 3507 923
rect 3485 584 3491 696
rect 3501 684 3507 917
rect 3533 904 3539 1036
rect 3565 943 3571 1337
rect 3613 1123 3619 1437
rect 3645 1344 3651 1456
rect 3677 1244 3683 1296
rect 3597 1117 3619 1123
rect 3597 1084 3603 1117
rect 3709 1123 3715 1496
rect 3725 1484 3731 1496
rect 3741 1344 3747 1456
rect 3757 1424 3763 1516
rect 3821 1444 3827 1696
rect 3773 1384 3779 1416
rect 3789 1284 3795 1376
rect 3770 1214 3782 1216
rect 3755 1206 3757 1214
rect 3765 1206 3767 1214
rect 3775 1206 3777 1214
rect 3785 1206 3787 1214
rect 3795 1206 3797 1214
rect 3770 1204 3782 1206
rect 3725 1124 3731 1196
rect 3700 1117 3715 1123
rect 3821 1104 3827 1356
rect 3837 1324 3843 1716
rect 3853 1584 3859 1716
rect 3869 1504 3875 1556
rect 3885 1504 3891 1736
rect 3885 1384 3891 1476
rect 3917 1364 3923 2136
rect 3933 2124 3939 2176
rect 3965 1984 3971 2436
rect 3949 1864 3955 1876
rect 3981 1823 3987 2276
rect 4013 2144 4019 2617
rect 4029 2584 4035 2596
rect 4045 2584 4051 2636
rect 4061 2364 4067 2536
rect 4077 2524 4083 2856
rect 4093 2584 4099 2696
rect 4109 2604 4115 2676
rect 4093 2544 4099 2576
rect 4109 2404 4115 2596
rect 4141 2504 4147 2716
rect 4093 2344 4099 2376
rect 4077 2304 4083 2336
rect 4141 2324 4147 2496
rect 4157 2463 4163 2856
rect 4173 2524 4179 2576
rect 4189 2544 4195 2576
rect 4221 2564 4227 2836
rect 4285 2824 4291 2876
rect 4317 2744 4323 2836
rect 4349 2784 4355 3116
rect 4365 3104 4371 3316
rect 4397 3164 4403 3436
rect 4413 3324 4419 3436
rect 4445 3344 4451 3476
rect 4461 3424 4467 3516
rect 4477 3464 4483 3476
rect 4477 3343 4483 3456
rect 4493 3444 4499 3496
rect 4509 3384 4515 3456
rect 4541 3384 4547 3476
rect 4557 3384 4563 3636
rect 4573 3524 4579 3757
rect 4621 3744 4627 3896
rect 4653 3884 4659 3936
rect 4669 3904 4675 3976
rect 4637 3764 4643 3776
rect 4685 3764 4691 4036
rect 4717 3884 4723 4257
rect 4749 4164 4755 4176
rect 4733 3944 4739 4116
rect 4733 3904 4739 3936
rect 4717 3764 4723 3876
rect 4733 3744 4739 3896
rect 4573 3383 4579 3436
rect 4573 3377 4595 3383
rect 4477 3337 4492 3343
rect 4413 3304 4419 3316
rect 4445 3304 4451 3316
rect 4461 3284 4467 3316
rect 4413 3044 4419 3116
rect 4365 2964 4371 2996
rect 4333 2724 4339 2756
rect 4381 2704 4387 3036
rect 4413 2924 4419 2936
rect 4429 2903 4435 3016
rect 4445 2984 4451 3056
rect 4461 2984 4467 3076
rect 4477 3044 4483 3096
rect 4493 3084 4499 3336
rect 4509 3324 4515 3376
rect 4557 3344 4563 3356
rect 4548 3337 4556 3343
rect 4541 3123 4547 3336
rect 4573 3324 4579 3356
rect 4589 3324 4595 3377
rect 4605 3344 4611 3436
rect 4621 3204 4627 3736
rect 4653 3484 4659 3536
rect 4669 3484 4675 3676
rect 4701 3564 4707 3636
rect 4685 3444 4691 3496
rect 4637 3364 4643 3396
rect 4653 3343 4659 3416
rect 4644 3337 4659 3343
rect 4525 3117 4547 3123
rect 4525 3084 4531 3117
rect 4493 3064 4499 3076
rect 4525 3064 4531 3076
rect 4541 3064 4547 3096
rect 4557 3084 4563 3136
rect 4477 2964 4483 3036
rect 4493 2984 4499 3036
rect 4525 2944 4531 2976
rect 4541 2944 4547 2976
rect 4477 2917 4524 2923
rect 4477 2904 4483 2917
rect 4573 2923 4579 3196
rect 4605 3104 4611 3156
rect 4589 2984 4595 3036
rect 4557 2917 4579 2923
rect 4413 2897 4435 2903
rect 4237 2684 4243 2696
rect 4365 2664 4371 2676
rect 4253 2564 4259 2656
rect 4317 2624 4323 2636
rect 4301 2504 4307 2516
rect 4365 2503 4371 2656
rect 4381 2584 4387 2636
rect 4413 2544 4419 2897
rect 4493 2702 4499 2756
rect 4429 2624 4435 2656
rect 4477 2564 4483 2596
rect 4493 2564 4499 2596
rect 4365 2497 4387 2503
rect 4157 2457 4179 2463
rect 4157 2384 4163 2416
rect 4173 2324 4179 2457
rect 4285 2324 4291 2376
rect 4141 2244 4147 2276
rect 4157 2264 4163 2276
rect 4061 2184 4067 2196
rect 4013 1884 4019 2076
rect 4109 1944 4115 2136
rect 4157 1984 4163 2256
rect 4141 1924 4147 1936
rect 4029 1824 4035 1896
rect 3981 1817 4003 1823
rect 3933 1724 3939 1756
rect 3949 1564 3955 1736
rect 3965 1483 3971 1796
rect 3981 1522 3987 1696
rect 3965 1477 3987 1483
rect 3917 1324 3923 1336
rect 3949 1326 3955 1476
rect 3837 1104 3843 1316
rect 3965 1264 3971 1456
rect 3581 964 3587 1036
rect 3613 944 3619 1096
rect 3725 1064 3731 1096
rect 3645 944 3651 956
rect 3565 937 3587 943
rect 3549 824 3555 916
rect 3565 884 3571 916
rect 3581 844 3587 937
rect 3629 924 3635 936
rect 3517 704 3523 716
rect 3581 704 3587 736
rect 3533 544 3539 676
rect 3549 584 3555 696
rect 3549 564 3555 576
rect 3469 484 3475 516
rect 3501 444 3507 536
rect 3597 504 3603 916
rect 3661 864 3667 916
rect 3677 903 3683 1036
rect 3757 964 3763 1036
rect 3709 944 3715 956
rect 3741 944 3747 956
rect 3693 924 3699 936
rect 3677 897 3692 903
rect 3709 783 3715 816
rect 3725 804 3731 896
rect 3741 864 3747 936
rect 3773 904 3779 1096
rect 3853 1084 3859 1196
rect 3869 1124 3875 1136
rect 3885 1104 3891 1236
rect 3981 1124 3987 1477
rect 3997 1124 4003 1817
rect 4061 1744 4067 1756
rect 4029 1684 4035 1716
rect 4077 1663 4083 1816
rect 4141 1784 4147 1896
rect 4157 1824 4163 1836
rect 4173 1783 4179 2316
rect 4237 2264 4243 2296
rect 4189 2224 4195 2256
rect 4189 1904 4195 2176
rect 4269 2164 4275 2236
rect 4301 2144 4307 2496
rect 4333 2284 4339 2336
rect 4317 2244 4323 2276
rect 4349 2244 4355 2256
rect 4333 2104 4339 2118
rect 4237 2044 4243 2056
rect 4205 1904 4211 1996
rect 4237 1984 4243 2036
rect 4157 1777 4179 1783
rect 4061 1657 4083 1663
rect 4013 1464 4019 1476
rect 4029 1464 4035 1496
rect 4045 1484 4051 1576
rect 3885 1064 3891 1076
rect 3901 1024 3907 1096
rect 3933 1084 3939 1116
rect 3949 1064 3955 1076
rect 3869 984 3875 996
rect 3837 924 3843 976
rect 3917 944 3923 1056
rect 3773 884 3779 896
rect 3770 814 3782 816
rect 3755 806 3757 814
rect 3765 806 3767 814
rect 3775 806 3777 814
rect 3785 806 3787 814
rect 3795 806 3797 814
rect 3770 804 3782 806
rect 3709 777 3747 783
rect 3741 764 3747 777
rect 3677 664 3683 676
rect 3709 664 3715 676
rect 3725 664 3731 756
rect 3821 724 3827 916
rect 3853 824 3859 896
rect 3613 584 3619 656
rect 3533 484 3539 496
rect 3613 444 3619 556
rect 3629 484 3635 516
rect 3645 323 3651 636
rect 3693 324 3699 636
rect 3821 564 3827 636
rect 3709 524 3715 556
rect 3725 544 3731 556
rect 3709 384 3715 436
rect 3770 414 3782 416
rect 3755 406 3757 414
rect 3765 406 3767 414
rect 3775 406 3777 414
rect 3785 406 3787 414
rect 3795 406 3797 414
rect 3770 404 3782 406
rect 3636 317 3651 323
rect 3501 284 3507 296
rect 3405 257 3420 263
rect 3405 203 3411 236
rect 3485 204 3491 276
rect 3533 264 3539 296
rect 3597 277 3612 283
rect 3549 264 3555 276
rect 3581 264 3587 276
rect 3389 197 3411 203
rect 3389 144 3395 197
rect 3549 184 3555 256
rect 3421 164 3427 176
rect 3421 126 3427 136
rect 3597 124 3603 277
rect 3821 283 3827 516
rect 3837 304 3843 736
rect 3853 624 3859 696
rect 3869 684 3875 856
rect 3885 724 3891 736
rect 3933 723 3939 1036
rect 3965 1024 3971 1116
rect 3949 824 3955 916
rect 3965 804 3971 916
rect 3981 904 3987 1036
rect 3997 924 4003 936
rect 3933 717 3955 723
rect 3917 644 3923 696
rect 3869 637 3884 643
rect 3869 544 3875 637
rect 3901 584 3907 596
rect 3949 564 3955 717
rect 3965 664 3971 676
rect 3933 524 3939 556
rect 3965 544 3971 656
rect 3949 537 3964 543
rect 3933 364 3939 516
rect 3869 324 3875 356
rect 3901 324 3907 336
rect 3933 304 3939 316
rect 3908 297 3923 303
rect 3853 284 3859 296
rect 3821 277 3836 283
rect 3645 264 3651 276
rect 3725 264 3731 276
rect 3613 124 3619 236
rect 3677 144 3683 176
rect 3741 124 3747 236
rect 3837 184 3843 276
rect 3885 264 3891 296
rect 3917 283 3923 297
rect 3917 277 3932 283
rect 3949 164 3955 537
rect 3981 504 3987 856
rect 4013 744 4019 1316
rect 4045 1104 4051 1296
rect 4061 1164 4067 1657
rect 4093 1563 4099 1756
rect 4093 1557 4115 1563
rect 4109 1524 4115 1557
rect 4125 1544 4131 1636
rect 4093 1364 4099 1476
rect 4141 1464 4147 1676
rect 4157 1584 4163 1777
rect 4189 1504 4195 1736
rect 4173 1464 4179 1496
rect 4109 1124 4115 1436
rect 4173 1384 4179 1396
rect 4189 1344 4195 1356
rect 4157 1304 4163 1336
rect 4205 1284 4211 1896
rect 4237 1724 4243 1856
rect 4253 1804 4259 1836
rect 4269 1684 4275 2036
rect 4285 1924 4291 1976
rect 4285 1904 4291 1916
rect 4333 1844 4339 1856
rect 4301 1784 4307 1836
rect 4317 1824 4323 1836
rect 4292 1757 4307 1763
rect 4244 1657 4259 1663
rect 4221 1624 4227 1636
rect 4221 1464 4227 1516
rect 4237 1503 4243 1636
rect 4253 1544 4259 1657
rect 4285 1584 4291 1696
rect 4301 1624 4307 1757
rect 4333 1723 4339 1836
rect 4324 1717 4339 1723
rect 4237 1497 4252 1503
rect 4285 1503 4291 1536
rect 4285 1497 4300 1503
rect 4221 1364 4227 1456
rect 4061 1084 4067 1096
rect 4029 984 4035 1076
rect 4029 944 4035 976
rect 4093 924 4099 1076
rect 4061 864 4067 916
rect 4093 702 4099 776
rect 4061 664 4067 696
rect 4109 684 4115 736
rect 3997 483 4003 516
rect 4013 504 4019 636
rect 4045 544 4051 596
rect 4061 563 4067 656
rect 4125 624 4131 1076
rect 4141 1064 4147 1096
rect 4157 1084 4163 1176
rect 4205 1124 4211 1176
rect 4221 1104 4227 1156
rect 4141 924 4147 976
rect 4173 944 4179 1076
rect 4189 624 4195 916
rect 4205 904 4211 1036
rect 4221 964 4227 1016
rect 4237 783 4243 1476
rect 4253 1144 4259 1476
rect 4269 1384 4275 1496
rect 4301 1464 4307 1476
rect 4301 1244 4307 1456
rect 4317 1404 4323 1716
rect 4349 1584 4355 2236
rect 4365 1984 4371 2476
rect 4365 1864 4371 1896
rect 4381 1524 4387 2497
rect 4397 2424 4403 2496
rect 4413 2204 4419 2236
rect 4429 1984 4435 2516
rect 4509 2504 4515 2676
rect 4541 2524 4547 2696
rect 4445 2264 4451 2336
rect 4477 2284 4483 2296
rect 4493 2284 4499 2336
rect 4500 2277 4524 2283
rect 4541 2244 4547 2516
rect 4493 2177 4531 2183
rect 4493 2164 4499 2177
rect 4525 2164 4531 2177
rect 4509 2124 4515 2156
rect 4509 2104 4515 2116
rect 4461 2084 4467 2096
rect 4525 1984 4531 2136
rect 4557 2104 4563 2917
rect 4573 2884 4579 2896
rect 4605 2884 4611 3056
rect 4573 2864 4579 2876
rect 4589 2724 4595 2836
rect 4621 2783 4627 3156
rect 4669 3103 4675 3336
rect 4701 3303 4707 3476
rect 4717 3324 4723 3436
rect 4733 3384 4739 3736
rect 4749 3544 4755 4116
rect 4781 3884 4787 4236
rect 4909 4184 4915 4256
rect 4829 4140 4835 4156
rect 4861 4064 4867 4136
rect 4909 3884 4915 3976
rect 4765 3724 4771 3836
rect 4797 3544 4803 3636
rect 4765 3424 4771 3456
rect 4781 3444 4787 3496
rect 4797 3464 4803 3476
rect 4813 3384 4819 3836
rect 4829 3604 4835 3836
rect 4845 3744 4851 3856
rect 4861 3684 4867 3696
rect 4861 3644 4867 3676
rect 4861 3524 4867 3536
rect 4877 3523 4883 3836
rect 4893 3684 4899 3716
rect 4909 3524 4915 3636
rect 4877 3517 4892 3523
rect 4829 3484 4835 3496
rect 4845 3464 4851 3496
rect 4893 3464 4899 3476
rect 4909 3464 4915 3516
rect 4781 3344 4787 3356
rect 4733 3303 4739 3316
rect 4701 3297 4739 3303
rect 4781 3303 4787 3316
rect 4781 3297 4796 3303
rect 4717 3144 4723 3236
rect 4660 3097 4675 3103
rect 4685 3064 4691 3116
rect 4637 3044 4643 3056
rect 4653 2903 4659 3056
rect 4701 3024 4707 3056
rect 4669 2964 4675 2996
rect 4701 2924 4707 2936
rect 4644 2897 4659 2903
rect 4637 2864 4643 2876
rect 4605 2777 4627 2783
rect 4573 2584 4579 2616
rect 4589 2384 4595 2496
rect 4605 2444 4611 2777
rect 4653 2704 4659 2776
rect 4701 2743 4707 2856
rect 4717 2763 4723 3016
rect 4733 2984 4739 3276
rect 4749 3044 4755 3096
rect 4749 2944 4755 2976
rect 4717 2757 4739 2763
rect 4701 2737 4723 2743
rect 4621 2544 4627 2576
rect 4637 2524 4643 2636
rect 4701 2584 4707 2716
rect 4717 2704 4723 2737
rect 4733 2664 4739 2757
rect 4717 2624 4723 2656
rect 4749 2643 4755 2856
rect 4765 2724 4771 3136
rect 4781 2944 4787 3116
rect 4797 2904 4803 3116
rect 4829 3044 4835 3076
rect 4845 3003 4851 3376
rect 4861 3324 4867 3436
rect 4893 3364 4899 3376
rect 4877 3184 4883 3336
rect 4909 3324 4915 3436
rect 4925 3343 4931 3836
rect 4941 3824 4947 3956
rect 4957 3903 4963 4396
rect 4973 4384 4979 4656
rect 4989 4524 4995 4776
rect 5037 4724 5043 4736
rect 5037 4564 5043 4576
rect 5037 4524 5043 4536
rect 4973 4184 4979 4236
rect 4989 4204 4995 4296
rect 5021 4284 5027 4496
rect 5037 4384 5043 4516
rect 5037 4144 5043 4236
rect 5053 4124 5059 4756
rect 5085 4344 5091 4836
rect 5197 4704 5203 4756
rect 5124 4657 5132 4663
rect 5133 4644 5139 4656
rect 5133 4524 5139 4596
rect 5149 4544 5155 4696
rect 5213 4684 5219 4816
rect 5309 4784 5315 4796
rect 5229 4664 5235 4696
rect 5213 4584 5219 4616
rect 5165 4524 5171 4576
rect 5229 4540 5235 4636
rect 5274 4614 5286 4616
rect 5259 4606 5261 4614
rect 5269 4606 5271 4614
rect 5279 4606 5281 4614
rect 5289 4606 5291 4614
rect 5299 4606 5301 4614
rect 5274 4604 5286 4606
rect 5181 4524 5187 4536
rect 5133 4424 5139 4436
rect 5069 4244 5075 4296
rect 5133 4284 5139 4296
rect 5005 4084 5011 4116
rect 5069 4103 5075 4236
rect 5101 4144 5107 4216
rect 5149 4184 5155 4256
rect 5165 4204 5171 4336
rect 5229 4297 5244 4303
rect 5213 4284 5219 4296
rect 5188 4257 5203 4263
rect 5101 4124 5107 4136
rect 5165 4124 5171 4196
rect 5197 4184 5203 4257
rect 5229 4184 5235 4297
rect 5245 4264 5251 4276
rect 5274 4214 5286 4216
rect 5259 4206 5261 4214
rect 5269 4206 5271 4214
rect 5279 4206 5281 4214
rect 5289 4206 5291 4214
rect 5299 4206 5301 4214
rect 5274 4204 5286 4206
rect 5325 4184 5331 4936
rect 5341 4924 5347 4936
rect 5389 4924 5395 5056
rect 5437 4956 5443 5036
rect 5485 4884 5491 4936
rect 5341 4484 5347 4696
rect 5389 4584 5395 4596
rect 5421 4584 5427 4636
rect 5373 4564 5379 4576
rect 5405 4524 5411 4536
rect 5357 4404 5363 4516
rect 5421 4504 5427 4516
rect 5229 4140 5235 4156
rect 5053 4097 5075 4103
rect 5005 3984 5011 4076
rect 5021 3944 5027 4036
rect 5037 3904 5043 3976
rect 4957 3897 4979 3903
rect 4973 3884 4979 3897
rect 4941 3724 4947 3816
rect 4973 3763 4979 3876
rect 4964 3757 4979 3763
rect 4989 3743 4995 3896
rect 5053 3844 5059 4097
rect 5069 3984 5075 4016
rect 5165 3984 5171 4096
rect 5213 4084 5219 4136
rect 5117 3897 5132 3903
rect 4980 3737 4995 3743
rect 5021 3724 5027 3836
rect 5037 3744 5043 3776
rect 5069 3744 5075 3856
rect 5101 3744 5107 3756
rect 5069 3723 5075 3736
rect 5053 3717 5075 3723
rect 5053 3644 5059 3717
rect 5037 3544 5043 3636
rect 5069 3524 5075 3696
rect 5037 3504 5043 3516
rect 5069 3504 5075 3516
rect 4989 3424 4995 3456
rect 5053 3444 5059 3476
rect 5101 3444 5107 3736
rect 5117 3684 5123 3897
rect 5181 3884 5187 4076
rect 5197 3984 5203 4036
rect 5213 3924 5219 3936
rect 5181 3864 5187 3876
rect 5165 3744 5171 3836
rect 5213 3744 5219 3916
rect 5293 3844 5299 4176
rect 5341 4164 5347 4296
rect 5357 4264 5363 4396
rect 5389 4304 5395 4476
rect 5437 4464 5443 4516
rect 5309 4124 5315 4136
rect 5357 3904 5363 4256
rect 5373 4184 5379 4256
rect 5373 4164 5379 4176
rect 5389 3884 5395 3976
rect 5405 3884 5411 4376
rect 5437 4364 5443 4456
rect 5453 4384 5459 4836
rect 5501 4824 5507 4936
rect 5517 4924 5523 5096
rect 5533 5084 5539 5096
rect 5725 5084 5731 5136
rect 5901 5104 5907 5136
rect 6029 5124 6035 5156
rect 6285 5117 6300 5123
rect 6077 5104 6083 5116
rect 5597 4964 5603 5036
rect 5645 4944 5651 5016
rect 5629 4924 5635 4936
rect 5549 4804 5555 4896
rect 5565 4884 5571 4916
rect 5629 4904 5635 4916
rect 5677 4824 5683 4836
rect 5693 4804 5699 5036
rect 5725 4944 5731 5056
rect 5741 5024 5747 5056
rect 5805 4944 5811 5096
rect 5917 5084 5923 5096
rect 5965 5064 5971 5076
rect 5837 5057 5852 5063
rect 5837 4944 5843 5057
rect 5869 4984 5875 5036
rect 5981 5004 5987 5096
rect 6061 5084 6067 5096
rect 5917 4950 5923 4996
rect 6013 4956 6019 5036
rect 6029 5024 6035 5036
rect 6061 4944 6067 5076
rect 6093 5004 6099 5056
rect 6093 4964 6099 4996
rect 6125 4984 6131 5076
rect 6221 5064 6227 5076
rect 6285 5064 6291 5117
rect 6333 5064 6339 5076
rect 6148 5057 6172 5063
rect 6157 4984 6163 5057
rect 6189 5004 6195 5036
rect 6365 5024 6371 5056
rect 6109 4964 6115 4976
rect 5773 4924 5779 4936
rect 5805 4904 5811 4916
rect 5997 4824 6003 4836
rect 5533 4704 5539 4716
rect 5668 4697 5699 4703
rect 5469 4484 5475 4676
rect 5501 4663 5507 4696
rect 5549 4684 5555 4696
rect 5629 4684 5635 4696
rect 5693 4684 5699 4697
rect 5661 4664 5667 4676
rect 5725 4664 5731 4716
rect 5741 4664 5747 4716
rect 5773 4704 5779 4736
rect 5805 4684 5811 4716
rect 5981 4684 5987 4716
rect 6029 4704 6035 4716
rect 6061 4684 6067 4836
rect 6077 4704 6083 4776
rect 6109 4723 6115 4956
rect 6189 4940 6195 4976
rect 6237 4904 6243 4956
rect 6285 4924 6291 4936
rect 6349 4924 6355 4976
rect 6397 4964 6403 5036
rect 6413 5024 6419 5096
rect 6429 4984 6435 5036
rect 6461 5024 6467 5080
rect 6477 5064 6483 5076
rect 6493 5024 6499 5076
rect 6589 5064 6595 5076
rect 6365 4944 6371 4956
rect 6413 4924 6419 4936
rect 6429 4904 6435 4936
rect 6109 4717 6131 4723
rect 6109 4684 6115 4696
rect 6125 4684 6131 4717
rect 6237 4703 6243 4896
rect 6317 4824 6323 4836
rect 6228 4697 6243 4703
rect 6221 4684 6227 4696
rect 6381 4684 6387 4736
rect 6404 4717 6419 4723
rect 5492 4657 5507 4663
rect 5501 4584 5507 4657
rect 5565 4564 5571 4596
rect 5549 4484 5555 4496
rect 5581 4484 5587 4656
rect 5613 4624 5619 4636
rect 5773 4604 5779 4636
rect 5613 4524 5619 4536
rect 5645 4484 5651 4556
rect 5709 4544 5715 4576
rect 5789 4564 5795 4676
rect 5805 4544 5811 4556
rect 5677 4524 5683 4536
rect 5661 4504 5667 4516
rect 5469 4384 5475 4476
rect 5565 4384 5571 4436
rect 5677 4384 5683 4416
rect 5549 4324 5555 4336
rect 5437 4244 5443 4296
rect 5421 4224 5427 4236
rect 5421 4104 5427 4216
rect 5437 4124 5443 4236
rect 5453 4084 5459 4316
rect 5485 4243 5491 4276
rect 5485 4237 5507 4243
rect 5501 4144 5507 4237
rect 5549 4164 5555 4264
rect 5581 4257 5596 4263
rect 5549 4144 5555 4156
rect 5421 3864 5427 4036
rect 5229 3764 5235 3836
rect 5274 3814 5286 3816
rect 5259 3806 5261 3814
rect 5269 3806 5271 3814
rect 5279 3806 5281 3814
rect 5289 3806 5291 3814
rect 5299 3806 5301 3814
rect 5274 3804 5286 3806
rect 5261 3744 5267 3756
rect 5229 3524 5235 3636
rect 5245 3504 5251 3556
rect 5181 3497 5196 3503
rect 5117 3464 5123 3476
rect 5149 3444 5155 3476
rect 5053 3384 5059 3396
rect 5165 3384 5171 3496
rect 5181 3444 5187 3497
rect 5204 3477 5228 3483
rect 5181 3384 5187 3416
rect 4957 3344 4963 3376
rect 4925 3337 4947 3343
rect 4877 3044 4883 3096
rect 4845 2997 4867 3003
rect 4829 2944 4835 2976
rect 4845 2924 4851 2976
rect 4781 2884 4787 2896
rect 4797 2863 4803 2896
rect 4861 2863 4867 2997
rect 4877 2964 4883 2976
rect 4893 2964 4899 2996
rect 4909 2884 4915 3116
rect 4941 3083 4947 3337
rect 4989 3184 4995 3336
rect 5021 3324 5027 3356
rect 5085 3344 5091 3376
rect 5037 3304 5043 3336
rect 5149 3324 5155 3356
rect 5069 3264 5075 3296
rect 5085 3104 5091 3316
rect 5165 3304 5171 3336
rect 5197 3323 5203 3456
rect 5245 3443 5251 3496
rect 5229 3437 5251 3443
rect 5229 3323 5235 3437
rect 5274 3414 5286 3416
rect 5259 3406 5261 3414
rect 5269 3406 5271 3414
rect 5279 3406 5281 3414
rect 5289 3406 5291 3414
rect 5299 3406 5301 3414
rect 5274 3404 5286 3406
rect 5293 3344 5299 3356
rect 5197 3317 5219 3323
rect 5229 3317 5244 3323
rect 5197 3284 5203 3296
rect 5197 3124 5203 3176
rect 5213 3164 5219 3317
rect 5213 3124 5219 3136
rect 4941 3077 4963 3083
rect 4925 3024 4931 3056
rect 4941 3024 4947 3056
rect 4925 2904 4931 2916
rect 4781 2857 4803 2863
rect 4845 2857 4867 2863
rect 4781 2724 4787 2857
rect 4829 2784 4835 2836
rect 4781 2683 4787 2716
rect 4733 2637 4755 2643
rect 4765 2677 4787 2683
rect 4733 2604 4739 2637
rect 4749 2584 4755 2616
rect 4685 2544 4691 2576
rect 4685 2524 4691 2536
rect 4621 2384 4627 2436
rect 4717 2424 4723 2516
rect 4765 2384 4771 2677
rect 4781 2584 4787 2636
rect 4573 2304 4579 2316
rect 4781 2304 4787 2336
rect 4797 2324 4803 2776
rect 4845 2723 4851 2857
rect 4845 2717 4860 2723
rect 4925 2704 4931 2896
rect 4941 2884 4947 2956
rect 4957 2903 4963 3077
rect 4973 2924 4979 2996
rect 4989 2944 4995 3096
rect 4957 2897 4972 2903
rect 4941 2704 4947 2836
rect 4964 2777 4988 2783
rect 5005 2744 5011 2836
rect 5021 2724 5027 3096
rect 5085 3084 5091 3096
rect 5069 3044 5075 3076
rect 5101 3044 5107 3076
rect 5149 3044 5155 3096
rect 5165 3064 5171 3076
rect 5037 2964 5043 2996
rect 5053 2943 5059 2956
rect 5101 2944 5107 2956
rect 5044 2937 5059 2943
rect 5101 2804 5107 2916
rect 5117 2904 5123 2956
rect 5165 2943 5171 3036
rect 5149 2937 5171 2943
rect 5149 2924 5155 2937
rect 5181 2923 5187 3056
rect 5197 3024 5203 3036
rect 5197 2924 5203 2976
rect 5213 2964 5219 3096
rect 5229 3077 5244 3083
rect 5229 2984 5235 3077
rect 5274 3014 5286 3016
rect 5259 3006 5261 3014
rect 5269 3006 5271 3014
rect 5279 3006 5281 3014
rect 5289 3006 5291 3014
rect 5299 3006 5301 3014
rect 5274 3004 5286 3006
rect 5165 2917 5187 2923
rect 5165 2884 5171 2917
rect 5149 2824 5155 2836
rect 5117 2764 5123 2796
rect 4957 2704 4963 2716
rect 4996 2697 5027 2703
rect 4845 2683 4851 2696
rect 4909 2684 4915 2696
rect 4845 2677 4860 2683
rect 4925 2683 4931 2696
rect 5021 2683 5027 2697
rect 4925 2677 4963 2683
rect 5021 2677 5036 2683
rect 4813 2644 4819 2676
rect 4893 2657 4924 2663
rect 4829 2624 4835 2656
rect 4893 2604 4899 2657
rect 4909 2584 4915 2596
rect 4829 2524 4835 2536
rect 4813 2424 4819 2516
rect 4845 2424 4851 2556
rect 4877 2544 4883 2576
rect 4861 2537 4876 2543
rect 4861 2524 4867 2537
rect 4909 2504 4915 2536
rect 4941 2524 4947 2576
rect 4605 2264 4611 2276
rect 4653 2264 4659 2276
rect 4573 2244 4579 2256
rect 4621 2244 4627 2256
rect 4685 2184 4691 2296
rect 4605 2157 4620 2163
rect 4605 2144 4611 2157
rect 4676 2137 4691 2143
rect 4621 2124 4627 2136
rect 4557 2004 4563 2036
rect 4573 1984 4579 2116
rect 4605 2064 4611 2096
rect 4621 2043 4627 2116
rect 4685 2103 4691 2137
rect 4701 2124 4707 2156
rect 4685 2097 4700 2103
rect 4717 2084 4723 2256
rect 4765 2224 4771 2276
rect 4893 2264 4899 2276
rect 4829 2177 4867 2183
rect 4733 2143 4739 2156
rect 4733 2137 4780 2143
rect 4829 2124 4835 2177
rect 4861 2164 4867 2177
rect 4893 2164 4899 2176
rect 4845 2144 4851 2156
rect 4621 2037 4643 2043
rect 4429 1884 4435 1976
rect 4637 1944 4643 2037
rect 4685 1924 4691 1996
rect 4701 1984 4707 2016
rect 4724 1937 4748 1943
rect 4733 1897 4748 1903
rect 4445 1884 4451 1896
rect 4413 1784 4419 1856
rect 4397 1664 4403 1716
rect 4445 1644 4451 1876
rect 4493 1824 4499 1876
rect 4541 1863 4547 1896
rect 4557 1884 4563 1896
rect 4573 1877 4588 1883
rect 4573 1863 4579 1877
rect 4541 1857 4579 1863
rect 4509 1844 4515 1856
rect 4253 1124 4259 1136
rect 4269 1124 4275 1236
rect 4317 1204 4323 1356
rect 4333 1344 4339 1436
rect 4301 1104 4307 1116
rect 4317 1084 4323 1096
rect 4333 1084 4339 1236
rect 4349 1144 4355 1516
rect 4365 1444 4371 1516
rect 4381 1497 4396 1503
rect 4381 1464 4387 1497
rect 4397 1477 4412 1483
rect 4365 1383 4371 1436
rect 4365 1377 4387 1383
rect 4365 1344 4371 1356
rect 4381 1304 4387 1377
rect 4365 1124 4371 1296
rect 4381 1124 4387 1296
rect 4397 1104 4403 1477
rect 4429 1424 4435 1456
rect 4445 1383 4451 1416
rect 4429 1377 4451 1383
rect 4429 1344 4435 1377
rect 4461 1344 4467 1796
rect 4493 1744 4499 1756
rect 4477 1504 4483 1676
rect 4477 1484 4483 1496
rect 4525 1344 4531 1836
rect 4541 1784 4547 1857
rect 4605 1784 4611 1896
rect 4637 1804 4643 1876
rect 4589 1664 4595 1716
rect 4653 1684 4659 1836
rect 4701 1824 4707 1896
rect 4733 1784 4739 1897
rect 4781 1864 4787 1996
rect 4797 1864 4803 1896
rect 4813 1884 4819 2096
rect 4845 2064 4851 2136
rect 4909 2124 4915 2136
rect 4845 1864 4851 1876
rect 4861 1844 4867 1896
rect 4701 1744 4707 1776
rect 4749 1744 4755 1836
rect 4877 1784 4883 1916
rect 4909 1904 4915 1916
rect 4909 1884 4915 1896
rect 4893 1864 4899 1876
rect 4925 1804 4931 2416
rect 4941 2324 4947 2476
rect 4957 2404 4963 2677
rect 5069 2664 5075 2716
rect 4989 2384 4995 2536
rect 5037 2504 5043 2576
rect 5053 2564 5059 2656
rect 5101 2543 5107 2736
rect 5117 2704 5123 2756
rect 5165 2744 5171 2816
rect 5181 2784 5187 2896
rect 5133 2704 5139 2716
rect 5117 2544 5123 2556
rect 5101 2537 5116 2543
rect 5005 2344 5011 2436
rect 4989 2264 4995 2296
rect 5005 2244 5011 2316
rect 5021 2284 5027 2296
rect 5037 2284 5043 2436
rect 5117 2304 5123 2396
rect 5149 2364 5155 2696
rect 5181 2624 5187 2756
rect 5213 2684 5219 2936
rect 5245 2784 5251 2936
rect 5261 2924 5267 2956
rect 5277 2684 5283 2956
rect 5197 2644 5203 2676
rect 5274 2614 5286 2616
rect 5259 2606 5261 2614
rect 5269 2606 5271 2614
rect 5279 2606 5281 2614
rect 5289 2606 5291 2614
rect 5299 2606 5301 2614
rect 5274 2604 5286 2606
rect 5229 2584 5235 2596
rect 5213 2504 5219 2536
rect 5229 2524 5235 2576
rect 5165 2324 5171 2396
rect 5197 2384 5203 2416
rect 4941 1884 4947 2236
rect 4957 2164 4963 2196
rect 4989 2124 4995 2156
rect 4957 1984 4963 2116
rect 5005 2084 5011 2136
rect 4973 1904 4979 2036
rect 5021 1924 5027 2156
rect 5037 2064 5043 2276
rect 5053 2184 5059 2236
rect 5069 2224 5075 2256
rect 5085 2224 5091 2256
rect 5117 2104 5123 2296
rect 5197 2223 5203 2336
rect 5277 2324 5283 2376
rect 5229 2284 5235 2316
rect 5245 2284 5251 2296
rect 5220 2257 5235 2263
rect 5197 2217 5219 2223
rect 5197 2184 5203 2196
rect 5213 2164 5219 2217
rect 5133 2124 5139 2136
rect 5181 2124 5187 2136
rect 4957 1824 4963 1856
rect 4989 1824 4995 1836
rect 4765 1744 4771 1776
rect 4813 1744 4819 1776
rect 4877 1744 4883 1756
rect 4669 1704 4675 1716
rect 4797 1704 4803 1736
rect 4845 1704 4851 1716
rect 4573 1504 4579 1536
rect 4621 1524 4627 1536
rect 4653 1504 4659 1576
rect 4685 1544 4691 1636
rect 4669 1517 4700 1523
rect 4621 1483 4627 1496
rect 4669 1483 4675 1517
rect 4621 1477 4675 1483
rect 4541 1404 4547 1456
rect 4685 1384 4691 1416
rect 4717 1384 4723 1696
rect 4733 1584 4739 1636
rect 4797 1504 4803 1516
rect 4877 1504 4883 1716
rect 4893 1584 4899 1716
rect 4925 1584 4931 1776
rect 4941 1764 4947 1796
rect 5005 1744 5011 1896
rect 5005 1703 5011 1716
rect 5005 1697 5020 1703
rect 5037 1683 5043 2016
rect 5053 1904 5059 2096
rect 5101 2084 5107 2096
rect 5229 2024 5235 2257
rect 5293 2244 5299 2516
rect 5325 2304 5331 3836
rect 5405 3764 5411 3856
rect 5421 3663 5427 3836
rect 5437 3704 5443 3876
rect 5453 3724 5459 4076
rect 5485 4044 5491 4136
rect 5581 4104 5587 4257
rect 5645 4164 5651 4256
rect 5693 4164 5699 4176
rect 5709 4164 5715 4436
rect 5773 4404 5779 4536
rect 5869 4484 5875 4556
rect 5933 4544 5939 4616
rect 5949 4564 5955 4596
rect 5885 4424 5891 4496
rect 5725 4324 5731 4376
rect 5725 4304 5731 4316
rect 5629 4104 5635 4116
rect 5501 3923 5507 4056
rect 5485 3917 5507 3923
rect 5485 3884 5491 3917
rect 5533 3904 5539 4096
rect 5581 4024 5587 4096
rect 5645 3984 5651 4116
rect 5661 3984 5667 4136
rect 5693 4124 5699 4156
rect 5741 4144 5747 4256
rect 5741 4124 5747 4136
rect 5757 4124 5763 4136
rect 5773 4124 5779 4356
rect 5860 4317 5875 4323
rect 5789 4184 5795 4256
rect 5805 4184 5811 4196
rect 5645 3904 5651 3976
rect 5693 3904 5699 3996
rect 5741 3904 5747 3996
rect 5805 3944 5811 4156
rect 5821 4144 5827 4276
rect 5853 4164 5859 4276
rect 5869 4264 5875 4317
rect 5853 4144 5859 4156
rect 5917 4144 5923 4396
rect 5949 4384 5955 4516
rect 5965 4504 5971 4636
rect 5981 4564 5987 4676
rect 6029 4564 6035 4576
rect 6125 4564 6131 4676
rect 6237 4644 6243 4676
rect 6237 4564 6243 4576
rect 5981 4384 5987 4516
rect 6077 4497 6108 4503
rect 6077 4484 6083 4497
rect 5949 4304 5955 4356
rect 5965 4344 5971 4376
rect 6029 4344 6035 4436
rect 6013 4244 6019 4276
rect 6013 4144 6019 4216
rect 6077 4184 6083 4296
rect 6093 4184 6099 4476
rect 6141 4304 6147 4316
rect 6109 4184 6115 4236
rect 6125 4144 6131 4196
rect 5821 3904 5827 3936
rect 5501 3864 5507 3896
rect 5501 3844 5507 3856
rect 5469 3764 5475 3836
rect 5517 3784 5523 3836
rect 5533 3764 5539 3896
rect 5581 3764 5587 3776
rect 5597 3744 5603 3876
rect 5773 3864 5779 3896
rect 5837 3864 5843 3916
rect 5629 3724 5635 3836
rect 5613 3664 5619 3716
rect 5645 3704 5651 3736
rect 5693 3724 5699 3856
rect 5837 3784 5843 3856
rect 5869 3763 5875 4016
rect 5901 4004 5907 4036
rect 5917 3944 5923 4136
rect 6029 4044 6035 4136
rect 5885 3924 5891 3936
rect 5965 3924 5971 4036
rect 5917 3844 5923 3896
rect 5933 3824 5939 3876
rect 5949 3844 5955 3916
rect 5965 3784 5971 3836
rect 5869 3757 5891 3763
rect 5725 3744 5731 3756
rect 5885 3744 5891 3757
rect 5948 3750 5956 3756
rect 5981 3744 5987 3876
rect 5997 3764 6003 3936
rect 6013 3884 6019 4036
rect 6125 3904 6131 4136
rect 6157 4123 6163 4336
rect 6221 4304 6227 4436
rect 6237 4283 6243 4436
rect 6221 4277 6243 4283
rect 6173 4264 6179 4276
rect 6189 4204 6195 4236
rect 6205 4184 6211 4276
rect 6157 4117 6172 4123
rect 6141 4104 6147 4116
rect 6189 4104 6195 4136
rect 6013 3803 6019 3876
rect 6013 3797 6035 3803
rect 5869 3724 5875 3736
rect 5981 3724 5987 3736
rect 6013 3704 6019 3776
rect 6029 3764 6035 3797
rect 6029 3744 6035 3756
rect 6061 3724 6067 3864
rect 6109 3763 6115 3876
rect 6125 3864 6131 3876
rect 6109 3757 6124 3763
rect 6109 3704 6115 3757
rect 5421 3657 5443 3663
rect 5357 3424 5363 3456
rect 5405 3383 5411 3496
rect 5421 3464 5427 3636
rect 5437 3524 5443 3657
rect 5501 3484 5507 3596
rect 5613 3504 5619 3636
rect 5757 3544 5763 3636
rect 5492 3457 5507 3463
rect 5421 3424 5427 3456
rect 5405 3377 5427 3383
rect 5341 3304 5347 3376
rect 5373 3344 5379 3356
rect 5389 3324 5395 3356
rect 5373 3124 5379 3136
rect 5421 3104 5427 3377
rect 5469 3323 5475 3436
rect 5501 3383 5507 3457
rect 5517 3404 5523 3496
rect 5549 3484 5555 3496
rect 5613 3484 5619 3496
rect 5725 3484 5731 3536
rect 5821 3524 5827 3656
rect 5949 3544 5955 3636
rect 5501 3377 5523 3383
rect 5469 3317 5484 3323
rect 5501 3284 5507 3356
rect 5421 3084 5427 3096
rect 5357 3044 5363 3056
rect 5357 2984 5363 3016
rect 5373 2964 5379 3036
rect 5453 3024 5459 3056
rect 5469 3044 5475 3076
rect 5485 3024 5491 3036
rect 5341 2924 5347 2956
rect 5389 2944 5395 2956
rect 5357 2704 5363 2936
rect 5405 2924 5411 2936
rect 5373 2764 5379 2916
rect 5437 2904 5443 3016
rect 5469 2964 5475 2996
rect 5501 2984 5507 3096
rect 5517 3084 5523 3377
rect 5533 3324 5539 3476
rect 5709 3464 5715 3476
rect 5757 3463 5763 3516
rect 5773 3484 5779 3496
rect 5789 3484 5795 3496
rect 5821 3464 5827 3516
rect 5949 3504 5955 3516
rect 5997 3464 6003 3516
rect 6045 3484 6051 3636
rect 6077 3524 6083 3676
rect 6141 3624 6147 3896
rect 6189 3883 6195 3896
rect 6173 3877 6195 3883
rect 6173 3844 6179 3877
rect 6189 3764 6195 3856
rect 6205 3844 6211 3856
rect 6221 3763 6227 4277
rect 6253 4264 6259 4636
rect 6269 4544 6275 4576
rect 6285 4524 6291 4556
rect 6285 4504 6291 4516
rect 6269 4304 6275 4316
rect 6301 4303 6307 4556
rect 6365 4544 6371 4556
rect 6381 4544 6387 4656
rect 6397 4584 6403 4636
rect 6413 4544 6419 4717
rect 6445 4684 6451 4976
rect 6541 4884 6547 5036
rect 6621 4984 6627 5076
rect 6653 5043 6659 5056
rect 6701 5044 6707 5096
rect 6653 5037 6675 5043
rect 6637 4984 6643 5036
rect 6669 4984 6675 5037
rect 6621 4964 6627 4976
rect 6557 4924 6563 4956
rect 6701 4924 6707 5036
rect 6733 4924 6739 5136
rect 7181 5097 7196 5103
rect 7181 5083 7187 5097
rect 7172 5077 7187 5083
rect 7085 5064 7091 5076
rect 7229 5064 7235 5076
rect 7277 5064 7283 5076
rect 6932 5057 6947 5063
rect 6845 4984 6851 5056
rect 6605 4904 6611 4916
rect 6557 4724 6563 4836
rect 6589 4784 6595 4896
rect 6493 4704 6499 4716
rect 6461 4664 6467 4696
rect 6605 4664 6611 4736
rect 6733 4724 6739 4916
rect 6861 4904 6867 5056
rect 6941 4984 6947 5057
rect 6941 4964 6947 4976
rect 6893 4944 6899 4956
rect 6778 4814 6790 4816
rect 6763 4806 6765 4814
rect 6773 4806 6775 4814
rect 6783 4806 6785 4814
rect 6793 4806 6795 4814
rect 6803 4806 6805 4814
rect 6778 4804 6790 4806
rect 6845 4724 6851 4836
rect 6669 4704 6675 4716
rect 6877 4704 6883 4836
rect 6957 4704 6963 4736
rect 6733 4684 6739 4696
rect 6381 4524 6387 4536
rect 6397 4524 6403 4536
rect 6365 4517 6380 4523
rect 6349 4344 6355 4436
rect 6292 4297 6307 4303
rect 6285 4264 6291 4296
rect 6365 4284 6371 4517
rect 6429 4504 6435 4576
rect 6445 4524 6451 4536
rect 6237 4244 6243 4256
rect 6253 4184 6259 4236
rect 6349 4224 6355 4276
rect 6285 4144 6291 4156
rect 6349 4124 6355 4176
rect 6381 4164 6387 4456
rect 6445 4384 6451 4496
rect 6461 4484 6467 4656
rect 6477 4564 6483 4636
rect 6621 4544 6627 4556
rect 6477 4504 6483 4536
rect 6525 4464 6531 4516
rect 6509 4457 6524 4463
rect 6493 4384 6499 4416
rect 6413 4264 6419 4276
rect 6429 4143 6435 4356
rect 6413 4137 6435 4143
rect 6237 3984 6243 4116
rect 6285 4104 6291 4116
rect 6397 4104 6403 4136
rect 6413 4124 6419 4137
rect 6301 3944 6307 4036
rect 6237 3824 6243 3876
rect 6253 3864 6259 3896
rect 6269 3864 6275 3896
rect 6253 3824 6259 3856
rect 6221 3757 6243 3763
rect 6189 3704 6195 3736
rect 6221 3724 6227 3736
rect 6205 3704 6211 3716
rect 5757 3457 5779 3463
rect 5597 3424 5603 3456
rect 5565 3304 5571 3356
rect 5581 3344 5587 3376
rect 5581 3224 5587 3316
rect 5597 3224 5603 3336
rect 5645 3324 5651 3436
rect 5549 3044 5555 3096
rect 5485 2944 5491 2976
rect 5533 2944 5539 2976
rect 5549 2944 5555 3036
rect 5581 3024 5587 3056
rect 5508 2917 5539 2923
rect 5533 2904 5539 2917
rect 5421 2784 5427 2816
rect 5357 2604 5363 2696
rect 5373 2624 5379 2656
rect 5357 2544 5363 2576
rect 5373 2503 5379 2556
rect 5389 2504 5395 2716
rect 5405 2703 5411 2776
rect 5437 2764 5443 2816
rect 5565 2784 5571 2976
rect 5581 2924 5587 2956
rect 5597 2944 5603 3216
rect 5661 3084 5667 3296
rect 5693 3284 5699 3316
rect 5725 3304 5731 3316
rect 5613 3044 5619 3076
rect 5629 2984 5635 3036
rect 5597 2903 5603 2916
rect 5645 2904 5651 3036
rect 5661 2984 5667 2996
rect 5677 2944 5683 2956
rect 5693 2924 5699 2956
rect 5588 2897 5603 2903
rect 5453 2703 5459 2776
rect 5485 2724 5491 2756
rect 5533 2704 5539 2756
rect 5405 2697 5427 2703
rect 5405 2644 5411 2676
rect 5364 2497 5379 2503
rect 5274 2214 5286 2216
rect 5259 2206 5261 2214
rect 5269 2206 5271 2214
rect 5279 2206 5281 2214
rect 5289 2206 5291 2214
rect 5299 2206 5301 2214
rect 5274 2204 5286 2206
rect 5325 2183 5331 2236
rect 5341 2224 5347 2316
rect 5357 2184 5363 2256
rect 5389 2184 5395 2396
rect 5405 2384 5411 2596
rect 5421 2444 5427 2697
rect 5437 2697 5459 2703
rect 5437 2604 5443 2697
rect 5453 2664 5459 2676
rect 5597 2664 5603 2736
rect 5725 2704 5731 3276
rect 5757 3204 5763 3436
rect 5773 3284 5779 3457
rect 6045 3463 6051 3476
rect 6077 3464 6083 3516
rect 6125 3504 6131 3556
rect 6036 3457 6051 3463
rect 5805 3324 5811 3376
rect 5821 3364 5827 3416
rect 5869 3384 5875 3436
rect 5837 3264 5843 3356
rect 5965 3344 5971 3416
rect 5853 3324 5859 3336
rect 5757 3084 5763 3176
rect 5869 3124 5875 3196
rect 5741 3024 5747 3056
rect 5757 2944 5763 2976
rect 5789 2963 5795 3076
rect 5853 3044 5859 3076
rect 5780 2957 5795 2963
rect 5837 2924 5843 2956
rect 5757 2844 5763 2916
rect 5853 2884 5859 2996
rect 5837 2824 5843 2836
rect 5757 2704 5763 2716
rect 5805 2704 5811 2756
rect 5853 2744 5859 2816
rect 5869 2764 5875 3036
rect 5885 2964 5891 3236
rect 5965 3124 5971 3136
rect 5901 3104 5907 3116
rect 5901 3084 5907 3096
rect 5949 3024 5955 3056
rect 5981 3044 5987 3136
rect 6013 3104 6019 3316
rect 5997 3044 6003 3076
rect 6013 3044 6019 3076
rect 5917 2944 5923 2956
rect 5949 2924 5955 2956
rect 5965 2904 5971 3036
rect 6061 2924 6067 3116
rect 6093 3104 6099 3376
rect 6141 3343 6147 3616
rect 6173 3484 6179 3536
rect 6205 3524 6211 3576
rect 6221 3384 6227 3436
rect 6237 3404 6243 3757
rect 6285 3743 6291 3936
rect 6317 3864 6323 3996
rect 6349 3864 6355 3916
rect 6429 3904 6435 4116
rect 6445 3864 6451 3916
rect 6461 3903 6467 4336
rect 6509 4284 6515 4457
rect 6541 4424 6547 4536
rect 6589 4484 6595 4496
rect 6573 4464 6579 4476
rect 6637 4464 6643 4536
rect 6589 4384 6595 4416
rect 6653 4384 6659 4476
rect 6685 4424 6691 4536
rect 6749 4524 6755 4636
rect 6765 4624 6771 4676
rect 6893 4664 6899 4676
rect 6909 4644 6915 4656
rect 6957 4644 6963 4676
rect 6925 4624 6931 4636
rect 6973 4544 6979 5036
rect 7021 4944 7027 5016
rect 7101 4964 7107 5056
rect 7133 5024 7139 5056
rect 7197 5024 7203 5056
rect 7245 4984 7251 5016
rect 7197 4964 7203 4976
rect 7101 4944 7107 4956
rect 7117 4944 7123 4956
rect 7133 4937 7148 4943
rect 7021 4904 7027 4936
rect 7053 4724 7059 4936
rect 7133 4923 7139 4937
rect 7124 4917 7139 4923
rect 7101 4744 7107 4776
rect 7133 4763 7139 4836
rect 7197 4764 7203 4836
rect 7133 4757 7155 4763
rect 7053 4704 7059 4716
rect 7069 4664 7075 4676
rect 6509 4264 6515 4276
rect 6477 4244 6483 4256
rect 6541 4244 6547 4316
rect 6493 4164 6499 4216
rect 6493 3904 6499 4096
rect 6461 3897 6476 3903
rect 6509 3884 6515 4196
rect 6541 4184 6547 4196
rect 6557 4144 6563 4256
rect 6573 4204 6579 4336
rect 6605 4284 6611 4316
rect 6605 4156 6611 4236
rect 6621 4204 6627 4296
rect 6637 4184 6643 4376
rect 6701 4324 6707 4516
rect 6778 4414 6790 4416
rect 6763 4406 6765 4414
rect 6773 4406 6775 4414
rect 6783 4406 6785 4414
rect 6793 4406 6795 4414
rect 6803 4406 6805 4414
rect 6778 4404 6790 4406
rect 6829 4384 6835 4496
rect 6845 4364 6851 4536
rect 6877 4384 6883 4536
rect 6909 4484 6915 4496
rect 6925 4304 6931 4316
rect 6813 4264 6819 4276
rect 6717 4184 6723 4256
rect 6717 4144 6723 4176
rect 6557 3864 6563 4116
rect 6285 3737 6300 3743
rect 6269 3704 6275 3716
rect 6317 3664 6323 3856
rect 6397 3724 6403 3836
rect 6445 3704 6451 3716
rect 6397 3564 6403 3636
rect 6253 3484 6259 3556
rect 6461 3544 6467 3836
rect 6477 3724 6483 3736
rect 6493 3704 6499 3816
rect 6573 3804 6579 3876
rect 6532 3677 6547 3683
rect 6340 3537 6355 3543
rect 6269 3464 6275 3536
rect 6301 3424 6307 3516
rect 6317 3504 6323 3536
rect 6349 3503 6355 3537
rect 6372 3517 6387 3523
rect 6349 3497 6364 3503
rect 6381 3444 6387 3517
rect 6381 3384 6387 3436
rect 6397 3404 6403 3496
rect 6413 3484 6419 3516
rect 6429 3444 6435 3456
rect 6253 3344 6259 3356
rect 6269 3344 6275 3376
rect 6141 3337 6156 3343
rect 6413 3324 6419 3416
rect 6461 3384 6467 3496
rect 6477 3364 6483 3496
rect 6493 3364 6499 3616
rect 6509 3383 6515 3636
rect 6525 3524 6531 3656
rect 6525 3504 6531 3516
rect 6525 3424 6531 3436
rect 6541 3384 6547 3677
rect 6557 3484 6563 3616
rect 6573 3544 6579 3596
rect 6589 3584 6595 3836
rect 6621 3743 6627 3876
rect 6621 3737 6636 3743
rect 6605 3724 6611 3736
rect 6557 3424 6563 3476
rect 6573 3464 6579 3516
rect 6589 3384 6595 3436
rect 6605 3384 6611 3696
rect 6637 3644 6643 3736
rect 6653 3504 6659 3936
rect 6669 3888 6675 4136
rect 6685 3984 6691 4116
rect 6733 4084 6739 4116
rect 6813 4104 6819 4256
rect 6829 4184 6835 4196
rect 6845 4144 6851 4296
rect 6909 4284 6915 4296
rect 6861 4264 6867 4276
rect 6893 4244 6899 4276
rect 6861 4124 6867 4176
rect 6877 4103 6883 4236
rect 6925 4104 6931 4276
rect 6941 4164 6947 4476
rect 6973 4384 6979 4496
rect 6989 4484 6995 4636
rect 7053 4544 7059 4636
rect 6989 4444 6995 4456
rect 6989 4323 6995 4436
rect 6973 4317 6995 4323
rect 6973 4284 6979 4317
rect 6989 4263 6995 4276
rect 6980 4257 6995 4263
rect 7005 4203 7011 4536
rect 7021 4444 7027 4516
rect 7053 4483 7059 4516
rect 7069 4484 7075 4576
rect 7085 4504 7091 4636
rect 7101 4524 7107 4736
rect 7117 4664 7123 4716
rect 7149 4704 7155 4757
rect 7213 4744 7219 4916
rect 7197 4684 7203 4716
rect 7181 4664 7187 4676
rect 7213 4664 7219 4696
rect 7124 4657 7139 4663
rect 7117 4644 7123 4656
rect 7133 4584 7139 4657
rect 7133 4524 7139 4576
rect 7149 4504 7155 4556
rect 7213 4524 7219 4536
rect 7037 4477 7059 4483
rect 7021 4324 7027 4436
rect 7037 4324 7043 4477
rect 7053 4344 7059 4436
rect 7181 4343 7187 4436
rect 7181 4337 7203 4343
rect 7037 4284 7043 4316
rect 7053 4264 7059 4296
rect 6989 4197 7011 4203
rect 6989 4164 6995 4197
rect 7021 4184 7027 4236
rect 7117 4204 7123 4256
rect 7149 4183 7155 4336
rect 7181 4304 7187 4316
rect 7165 4264 7171 4276
rect 7149 4177 7171 4183
rect 6941 4144 6947 4156
rect 6989 4104 6995 4156
rect 7005 4144 7011 4156
rect 7165 4144 7171 4177
rect 7181 4164 7187 4196
rect 6877 4097 6892 4103
rect 6733 3904 6739 4076
rect 6778 4014 6790 4016
rect 6763 4006 6765 4014
rect 6773 4006 6775 4014
rect 6783 4006 6785 4014
rect 6793 4006 6795 4014
rect 6803 4006 6805 4014
rect 6778 4004 6790 4006
rect 6861 3984 6867 4096
rect 6749 3904 6755 3976
rect 6909 3924 6915 4036
rect 6685 3864 6691 3876
rect 6669 3744 6675 3796
rect 6701 3724 6707 3736
rect 6717 3503 6723 3896
rect 6845 3764 6851 3836
rect 6749 3744 6755 3756
rect 6861 3744 6867 3876
rect 6925 3744 6931 3876
rect 6733 3724 6739 3736
rect 6925 3724 6931 3736
rect 6941 3704 6947 3896
rect 6989 3764 6995 3916
rect 7005 3864 7011 3916
rect 7021 3904 7027 4116
rect 7085 3937 7100 3943
rect 7037 3904 7043 3916
rect 7012 3857 7027 3863
rect 6989 3744 6995 3756
rect 7005 3724 7011 3736
rect 6778 3614 6790 3616
rect 6763 3606 6765 3614
rect 6773 3606 6775 3614
rect 6783 3606 6785 3614
rect 6793 3606 6795 3614
rect 6803 3606 6805 3614
rect 6778 3604 6790 3606
rect 6861 3524 6867 3576
rect 6957 3544 6963 3636
rect 6717 3497 6732 3503
rect 6621 3464 6627 3496
rect 6893 3484 6899 3496
rect 6717 3463 6723 3476
rect 6717 3457 6739 3463
rect 6653 3444 6659 3456
rect 6509 3377 6531 3383
rect 6477 3344 6483 3356
rect 6509 3344 6515 3356
rect 6525 3324 6531 3377
rect 6157 3303 6163 3316
rect 6148 3297 6163 3303
rect 6301 3284 6307 3296
rect 6125 3104 6131 3236
rect 6333 3184 6339 3216
rect 6221 3124 6227 3156
rect 6381 3104 6387 3156
rect 6397 3124 6403 3136
rect 6445 3104 6451 3296
rect 6541 3284 6547 3296
rect 6461 3124 6467 3136
rect 6237 3077 6252 3083
rect 6077 3064 6083 3076
rect 6109 3064 6115 3076
rect 6125 2904 6131 3036
rect 6157 2944 6163 2956
rect 6205 2924 6211 3036
rect 5901 2683 5907 2836
rect 6029 2784 6035 2896
rect 5933 2717 5948 2723
rect 5933 2704 5939 2717
rect 5981 2704 5987 2776
rect 6205 2764 6211 2876
rect 6237 2784 6243 3077
rect 6317 3044 6323 3076
rect 6365 3064 6371 3076
rect 6269 2963 6275 3036
rect 6285 2964 6291 2976
rect 6301 2964 6307 2996
rect 6260 2957 6275 2963
rect 6301 2904 6307 2916
rect 5901 2677 5916 2683
rect 5949 2683 5955 2696
rect 5997 2684 6003 2696
rect 6061 2684 6067 2736
rect 5933 2677 5955 2683
rect 5469 2564 5475 2636
rect 5485 2564 5491 2596
rect 5501 2564 5507 2596
rect 5444 2477 5459 2483
rect 5421 2343 5427 2416
rect 5437 2384 5443 2456
rect 5453 2424 5459 2477
rect 5453 2344 5459 2396
rect 5517 2364 5523 2636
rect 5549 2624 5555 2656
rect 5565 2604 5571 2636
rect 5581 2584 5587 2616
rect 5597 2564 5603 2596
rect 5613 2584 5619 2676
rect 5549 2524 5555 2536
rect 5549 2463 5555 2516
rect 5604 2497 5619 2503
rect 5549 2457 5571 2463
rect 5421 2337 5443 2343
rect 5437 2304 5443 2337
rect 5533 2343 5539 2356
rect 5517 2337 5539 2343
rect 5517 2304 5523 2337
rect 5533 2304 5539 2316
rect 5437 2264 5443 2276
rect 5325 2177 5347 2183
rect 5341 2156 5347 2177
rect 5405 2164 5411 2236
rect 5293 2144 5299 2156
rect 5405 2144 5411 2156
rect 5277 2104 5283 2136
rect 5341 2064 5347 2116
rect 5437 2104 5443 2256
rect 5485 2184 5491 2256
rect 5549 2224 5555 2276
rect 5517 2164 5523 2196
rect 5565 2124 5571 2457
rect 5581 2384 5587 2456
rect 5597 2244 5603 2296
rect 5613 2184 5619 2497
rect 5629 2164 5635 2576
rect 5645 2524 5651 2636
rect 5661 2564 5667 2664
rect 5725 2644 5731 2676
rect 5741 2584 5747 2636
rect 5757 2523 5763 2576
rect 5748 2517 5763 2523
rect 5645 2364 5651 2436
rect 5773 2424 5779 2656
rect 5789 2524 5795 2656
rect 5709 2324 5715 2336
rect 5677 2284 5683 2316
rect 5709 2264 5715 2276
rect 5757 2204 5763 2296
rect 5757 2184 5763 2196
rect 5645 2144 5651 2176
rect 5693 2144 5699 2176
rect 5709 2144 5715 2176
rect 5549 2117 5564 2123
rect 5501 2104 5507 2116
rect 5149 1984 5155 2016
rect 5053 1844 5059 1896
rect 5021 1677 5043 1683
rect 4973 1524 4979 1676
rect 4733 1384 4739 1496
rect 4925 1484 4931 1496
rect 4781 1424 4787 1476
rect 4852 1457 4867 1463
rect 4765 1384 4771 1396
rect 4589 1344 4595 1356
rect 4461 1324 4467 1336
rect 4429 1244 4435 1316
rect 4381 1084 4387 1096
rect 4413 1084 4419 1116
rect 4429 1104 4435 1236
rect 4461 1084 4467 1276
rect 4493 1102 4499 1336
rect 4573 1324 4579 1336
rect 4637 1324 4643 1336
rect 4605 1244 4611 1316
rect 4653 1304 4659 1316
rect 4701 1284 4707 1356
rect 4829 1344 4835 1436
rect 4861 1364 4867 1457
rect 4909 1364 4915 1416
rect 4845 1344 4851 1356
rect 4733 1184 4739 1316
rect 4813 1124 4819 1136
rect 4685 1102 4691 1116
rect 4829 1084 4835 1096
rect 4845 1084 4851 1336
rect 4861 1324 4867 1336
rect 4941 1324 4947 1516
rect 4973 1424 4979 1456
rect 4989 1364 4995 1436
rect 5021 1344 5027 1677
rect 5037 1504 5043 1516
rect 5053 1484 5059 1716
rect 5069 1524 5075 1916
rect 5341 1904 5347 1916
rect 5373 1884 5379 1916
rect 5085 1824 5091 1856
rect 5085 1764 5091 1816
rect 5069 1424 5075 1456
rect 5085 1404 5091 1456
rect 5101 1424 5107 1816
rect 5149 1744 5155 1776
rect 5117 1704 5123 1736
rect 5117 1524 5123 1576
rect 5149 1524 5155 1716
rect 5165 1704 5171 1836
rect 5213 1824 5219 1876
rect 5437 1864 5443 1916
rect 5229 1824 5235 1856
rect 5274 1814 5286 1816
rect 5259 1806 5261 1814
rect 5269 1806 5271 1814
rect 5279 1806 5281 1814
rect 5289 1806 5291 1814
rect 5299 1806 5301 1814
rect 5274 1804 5286 1806
rect 5405 1804 5411 1836
rect 5517 1824 5523 1856
rect 5197 1664 5203 1696
rect 5181 1584 5187 1636
rect 5149 1504 5155 1516
rect 5117 1483 5123 1496
rect 5117 1477 5164 1483
rect 5085 1364 5091 1396
rect 5101 1344 5107 1416
rect 5117 1364 5123 1436
rect 5181 1424 5187 1456
rect 5213 1423 5219 1796
rect 5325 1764 5331 1796
rect 5341 1764 5347 1796
rect 5229 1724 5235 1756
rect 5373 1724 5379 1776
rect 5405 1704 5411 1756
rect 5421 1744 5427 1756
rect 5437 1724 5443 1776
rect 5453 1704 5459 1736
rect 5469 1704 5475 1796
rect 5533 1704 5539 1916
rect 5549 1784 5555 2117
rect 5613 2104 5619 2116
rect 5661 2104 5667 2116
rect 5613 1924 5619 2096
rect 5565 1844 5571 1876
rect 5581 1844 5587 1876
rect 5613 1844 5619 1916
rect 5661 1844 5667 1876
rect 5677 1864 5683 1876
rect 5597 1824 5603 1836
rect 5629 1804 5635 1836
rect 5581 1764 5587 1776
rect 5629 1744 5635 1776
rect 5645 1744 5651 1776
rect 5677 1763 5683 1856
rect 5677 1757 5692 1763
rect 5677 1724 5683 1757
rect 5485 1684 5491 1696
rect 5245 1664 5251 1676
rect 5229 1604 5235 1636
rect 5501 1624 5507 1636
rect 5549 1624 5555 1716
rect 5261 1524 5267 1576
rect 5405 1544 5411 1576
rect 5380 1537 5395 1543
rect 5389 1523 5395 1537
rect 5389 1517 5420 1523
rect 5229 1504 5235 1516
rect 5373 1504 5379 1516
rect 5213 1417 5235 1423
rect 5213 1364 5219 1396
rect 4941 1304 4947 1316
rect 4989 1184 4995 1336
rect 5005 1224 5011 1296
rect 5021 1144 5027 1316
rect 5117 1304 5123 1316
rect 5053 1184 5059 1216
rect 4877 1104 4883 1116
rect 4884 1097 4899 1103
rect 4269 943 4275 1076
rect 4333 1064 4339 1076
rect 4260 937 4275 943
rect 4285 864 4291 916
rect 4301 904 4307 1036
rect 4317 944 4323 956
rect 4333 944 4339 976
rect 4509 964 4515 1076
rect 4621 1044 4627 1056
rect 4749 1024 4755 1076
rect 4861 1064 4867 1096
rect 4317 824 4323 916
rect 4365 823 4371 936
rect 4381 843 4387 916
rect 4397 864 4403 956
rect 4653 944 4659 976
rect 4717 944 4723 996
rect 4381 837 4403 843
rect 4365 817 4387 823
rect 4221 777 4243 783
rect 4205 564 4211 736
rect 4221 724 4227 777
rect 4237 704 4243 756
rect 4253 684 4259 816
rect 4221 604 4227 636
rect 4061 557 4076 563
rect 3997 477 4019 483
rect 3997 324 4003 336
rect 3981 284 3987 316
rect 3997 163 4003 236
rect 3981 157 4003 163
rect 3949 144 3955 156
rect 3981 103 3987 157
rect 4013 124 4019 477
rect 4029 444 4035 516
rect 4093 464 4099 496
rect 4109 484 4115 516
rect 4205 504 4211 518
rect 4093 324 4099 456
rect 4125 444 4131 476
rect 4173 384 4179 476
rect 4045 164 4051 236
rect 4061 124 4067 136
rect 4077 124 4083 296
rect 4125 244 4131 296
rect 4157 283 4163 316
rect 4173 304 4179 356
rect 4148 277 4163 283
rect 4189 244 4195 336
rect 4221 264 4227 276
rect 4237 204 4243 536
rect 4253 524 4259 676
rect 4301 464 4307 696
rect 4333 644 4339 676
rect 4349 544 4355 796
rect 4381 724 4387 817
rect 4397 784 4403 837
rect 4429 804 4435 936
rect 4445 924 4451 936
rect 4509 926 4515 936
rect 4413 684 4419 696
rect 4445 684 4451 736
rect 4477 664 4483 856
rect 4493 704 4499 756
rect 4573 744 4579 916
rect 4637 784 4643 836
rect 4653 824 4659 916
rect 4701 904 4707 936
rect 4797 924 4803 976
rect 4669 784 4675 796
rect 4605 704 4611 756
rect 4717 744 4723 916
rect 4733 824 4739 916
rect 4813 884 4819 916
rect 4829 804 4835 936
rect 4893 824 4899 1097
rect 5021 1084 5027 1136
rect 5069 1084 5075 1176
rect 5213 1144 5219 1216
rect 4925 964 4931 1016
rect 4909 784 4915 796
rect 4653 684 4659 716
rect 4477 564 4483 656
rect 4541 564 4547 676
rect 4404 557 4419 563
rect 4413 544 4419 557
rect 4269 384 4275 436
rect 4269 224 4275 296
rect 4173 124 4179 156
rect 4189 144 4195 196
rect 4285 124 4291 176
rect 4301 144 4307 416
rect 4317 123 4323 516
rect 4333 364 4339 436
rect 4413 384 4419 516
rect 4429 484 4435 516
rect 4541 504 4547 518
rect 4333 264 4339 356
rect 4477 324 4483 456
rect 4493 384 4499 476
rect 4445 164 4451 236
rect 4365 144 4371 156
rect 4308 117 4323 123
rect 3981 97 3996 103
rect 4413 84 4419 136
rect 4429 64 4435 116
rect 4461 84 4467 216
rect 4477 144 4483 316
rect 4557 264 4563 336
rect 4573 304 4579 376
rect 4541 144 4547 256
rect 4589 244 4595 316
rect 4605 184 4611 316
rect 4621 164 4627 376
rect 4653 324 4659 676
rect 4669 564 4675 736
rect 4685 644 4691 696
rect 4717 684 4723 696
rect 4765 664 4771 776
rect 4845 703 4851 776
rect 4925 763 4931 956
rect 5149 944 5155 1016
rect 5076 917 5091 923
rect 4909 757 4931 763
rect 4845 697 4860 703
rect 4836 677 4851 683
rect 4765 644 4771 656
rect 4685 544 4691 576
rect 4740 557 4755 563
rect 4749 544 4755 557
rect 4772 517 4787 523
rect 4669 384 4675 436
rect 4749 324 4755 516
rect 4781 384 4787 517
rect 4797 364 4803 636
rect 4813 564 4819 656
rect 4845 424 4851 677
rect 4893 624 4899 716
rect 4909 544 4915 757
rect 4941 704 4947 736
rect 4989 724 4995 736
rect 5021 724 5027 756
rect 5053 744 5059 836
rect 5085 784 5091 917
rect 5076 737 5091 743
rect 4877 504 4883 518
rect 4669 244 4675 256
rect 4733 184 4739 316
rect 4797 264 4803 316
rect 4669 164 4675 176
rect 4509 84 4515 116
rect 4525 104 4531 136
rect 4541 104 4547 136
rect 4781 124 4787 156
rect 4877 144 4883 416
rect 4893 304 4899 476
rect 4909 364 4915 536
rect 4925 404 4931 656
rect 4941 464 4947 696
rect 4957 684 4963 716
rect 4989 544 4995 716
rect 5005 644 5011 696
rect 5037 684 5043 716
rect 5053 624 5059 696
rect 5037 584 5043 616
rect 5021 544 5027 556
rect 4909 284 4915 296
rect 4909 264 4915 276
rect 4925 244 4931 256
rect 4941 144 4947 436
rect 4973 264 4979 536
rect 5053 484 5059 616
rect 5069 524 5075 556
rect 5085 544 5091 737
rect 5101 684 5107 716
rect 5117 644 5123 696
rect 5165 664 5171 676
rect 5213 664 5219 1056
rect 5229 764 5235 1417
rect 5274 1414 5286 1416
rect 5259 1406 5261 1414
rect 5269 1406 5271 1414
rect 5279 1406 5281 1414
rect 5289 1406 5291 1414
rect 5299 1406 5301 1414
rect 5274 1404 5286 1406
rect 5325 1324 5331 1476
rect 5357 1324 5363 1496
rect 5421 1464 5427 1496
rect 5501 1484 5507 1496
rect 5517 1463 5523 1616
rect 5597 1504 5603 1596
rect 5613 1524 5619 1636
rect 5645 1564 5651 1716
rect 5693 1644 5699 1736
rect 5501 1457 5523 1463
rect 5309 1303 5315 1316
rect 5309 1297 5324 1303
rect 5357 1184 5363 1276
rect 5373 1224 5379 1336
rect 5389 1304 5395 1376
rect 5421 1284 5427 1436
rect 5501 1384 5507 1457
rect 5565 1364 5571 1436
rect 5629 1424 5635 1456
rect 5581 1364 5587 1396
rect 5437 1337 5452 1343
rect 5437 1324 5443 1337
rect 5533 1324 5539 1336
rect 5629 1324 5635 1336
rect 5274 1014 5286 1016
rect 5259 1006 5261 1014
rect 5269 1006 5271 1014
rect 5279 1006 5281 1014
rect 5289 1006 5291 1014
rect 5299 1006 5301 1014
rect 5274 1004 5286 1006
rect 5245 964 5251 976
rect 5309 724 5315 736
rect 5325 704 5331 836
rect 5341 804 5347 836
rect 5341 704 5347 796
rect 5149 583 5155 636
rect 5165 584 5171 616
rect 5133 577 5155 583
rect 5133 564 5139 577
rect 5005 324 5011 436
rect 5021 324 5027 336
rect 5053 304 5059 336
rect 5085 304 5091 516
rect 5101 444 5107 496
rect 5133 484 5139 556
rect 5149 544 5155 556
rect 5149 504 5155 536
rect 5165 524 5171 536
rect 5181 524 5187 636
rect 5197 504 5203 636
rect 5213 564 5219 596
rect 5229 584 5235 676
rect 5274 614 5286 616
rect 5259 606 5261 614
rect 5269 606 5271 614
rect 5279 606 5281 614
rect 5289 606 5291 614
rect 5299 606 5301 614
rect 5274 604 5286 606
rect 5309 544 5315 576
rect 5325 544 5331 696
rect 5357 684 5363 756
rect 5405 724 5411 1236
rect 5437 1204 5443 1236
rect 5501 1144 5507 1296
rect 5581 1284 5587 1296
rect 5613 1204 5619 1256
rect 5613 1104 5619 1196
rect 5453 1004 5459 1096
rect 5469 924 5475 1076
rect 5501 964 5507 1096
rect 5517 1004 5523 1076
rect 5597 984 5603 1016
rect 5613 984 5619 1076
rect 5629 984 5635 1136
rect 5437 904 5443 918
rect 5453 724 5459 856
rect 5501 724 5507 776
rect 5565 744 5571 836
rect 5581 784 5587 936
rect 5629 904 5635 916
rect 5645 724 5651 1556
rect 5661 1524 5667 1636
rect 5709 1604 5715 2116
rect 5741 1924 5747 2096
rect 5789 2024 5795 2036
rect 5805 1944 5811 2656
rect 5821 2564 5827 2636
rect 5885 2624 5891 2656
rect 5901 2584 5907 2616
rect 5837 2544 5843 2556
rect 5933 2524 5939 2677
rect 5949 2564 5955 2656
rect 5981 2544 5987 2636
rect 6013 2624 6019 2676
rect 6077 2664 6083 2680
rect 6173 2664 6179 2736
rect 6205 2704 6211 2756
rect 6253 2704 6259 2736
rect 6317 2704 6323 2816
rect 6349 2704 6355 2716
rect 6381 2664 6387 2936
rect 6429 2784 6435 3096
rect 6445 3084 6451 3096
rect 6541 3084 6547 3096
rect 6557 3084 6563 3216
rect 6573 3123 6579 3336
rect 6573 3117 6595 3123
rect 6573 3084 6579 3096
rect 6477 2844 6483 3076
rect 6493 2944 6499 2956
rect 6525 2944 6531 2976
rect 6557 2904 6563 3056
rect 6500 2877 6556 2883
rect 6573 2844 6579 2936
rect 6589 2884 6595 3117
rect 6605 3084 6611 3316
rect 6621 3284 6627 3316
rect 6637 3224 6643 3236
rect 6685 3184 6691 3436
rect 6701 3344 6707 3416
rect 6733 3363 6739 3457
rect 6717 3357 6739 3363
rect 6717 3323 6723 3357
rect 6701 3317 6723 3323
rect 6621 3084 6627 3176
rect 6637 3104 6643 3176
rect 6653 3104 6659 3116
rect 6605 2983 6611 3036
rect 6621 3024 6627 3076
rect 6685 3024 6691 3036
rect 6605 2977 6627 2983
rect 6621 2944 6627 2977
rect 6397 2737 6451 2743
rect 6029 2524 6035 2536
rect 5901 2304 5907 2316
rect 5933 2297 5948 2303
rect 5853 2264 5859 2276
rect 5933 2263 5939 2297
rect 5908 2257 5939 2263
rect 5821 2244 5827 2256
rect 5837 2164 5843 2196
rect 5853 2144 5859 2256
rect 5869 2184 5875 2216
rect 5949 2184 5955 2256
rect 5965 2204 5971 2256
rect 5997 2144 6003 2236
rect 6013 2184 6019 2296
rect 6013 2144 6019 2156
rect 6029 2140 6035 2236
rect 5837 1923 5843 2036
rect 5853 1964 5859 2096
rect 5885 2064 5891 2136
rect 6045 2124 6051 2616
rect 6109 2584 6115 2636
rect 6125 2624 6131 2656
rect 6157 2584 6163 2636
rect 6157 2564 6163 2576
rect 6173 2524 6179 2656
rect 6205 2624 6211 2656
rect 6285 2644 6291 2656
rect 6221 2564 6227 2636
rect 6237 2537 6275 2543
rect 6237 2524 6243 2537
rect 6269 2524 6275 2537
rect 6301 2503 6307 2556
rect 6381 2544 6387 2656
rect 6397 2584 6403 2737
rect 6445 2704 6451 2737
rect 6413 2624 6419 2696
rect 6413 2524 6419 2576
rect 6429 2544 6435 2676
rect 6461 2624 6467 2680
rect 6461 2584 6467 2616
rect 6477 2584 6483 2836
rect 6541 2784 6547 2816
rect 6605 2784 6611 2936
rect 6653 2904 6659 3016
rect 6669 2924 6675 2956
rect 6685 2944 6691 2956
rect 6701 2944 6707 3317
rect 6733 3183 6739 3336
rect 6749 3324 6755 3376
rect 6845 3323 6851 3476
rect 6925 3464 6931 3536
rect 6957 3504 6963 3516
rect 6941 3464 6947 3496
rect 6836 3317 6851 3323
rect 6877 3304 6883 3416
rect 6909 3344 6915 3356
rect 6925 3324 6931 3356
rect 6941 3224 6947 3336
rect 6778 3214 6790 3216
rect 6763 3206 6765 3214
rect 6773 3206 6775 3214
rect 6783 3206 6785 3214
rect 6793 3206 6795 3214
rect 6803 3206 6805 3214
rect 6778 3204 6790 3206
rect 6733 3177 6755 3183
rect 6717 3064 6723 3076
rect 6733 3044 6739 3096
rect 6717 2944 6723 3036
rect 6749 3024 6755 3177
rect 6861 3104 6867 3136
rect 6909 3124 6915 3196
rect 6957 3184 6963 3476
rect 6973 3184 6979 3616
rect 7021 3584 7027 3857
rect 7053 3744 7059 3856
rect 7085 3756 7091 3937
rect 7165 3924 7171 4136
rect 7149 3644 7155 3896
rect 7197 3884 7203 4337
rect 7229 4324 7235 4956
rect 7309 4944 7315 5076
rect 7332 5057 7340 5063
rect 7389 5024 7395 5056
rect 7396 5017 7411 5023
rect 7405 4944 7411 5017
rect 7245 4724 7251 4736
rect 7261 4704 7267 4896
rect 7277 4744 7283 4836
rect 7261 4684 7267 4696
rect 7277 4684 7283 4696
rect 7293 4683 7299 4936
rect 7284 4677 7299 4683
rect 7325 4664 7331 4676
rect 7245 4584 7251 4636
rect 7309 4564 7315 4636
rect 7341 4564 7347 4656
rect 7373 4564 7379 4576
rect 7357 4544 7363 4556
rect 7293 4344 7299 4436
rect 7277 4284 7283 4316
rect 7293 4284 7299 4296
rect 7373 4284 7379 4296
rect 7229 4063 7235 4236
rect 7277 4204 7283 4276
rect 7341 4204 7347 4256
rect 7373 4184 7379 4276
rect 7341 4164 7347 4176
rect 7245 4144 7251 4156
rect 7309 4144 7315 4156
rect 7213 4057 7235 4063
rect 7213 3884 7219 4057
rect 7165 3864 7171 3876
rect 7181 3723 7187 3836
rect 7197 3803 7203 3876
rect 7197 3797 7219 3803
rect 7197 3764 7203 3776
rect 7213 3744 7219 3797
rect 7172 3717 7187 3723
rect 7213 3684 7219 3716
rect 7101 3524 7107 3636
rect 7117 3623 7123 3636
rect 7117 3617 7139 3623
rect 7069 3504 7075 3516
rect 7133 3504 7139 3617
rect 7005 3444 7011 3496
rect 7021 3444 7027 3496
rect 6989 3344 6995 3376
rect 6797 2984 6803 3076
rect 6445 2537 6460 2543
rect 6292 2497 6307 2503
rect 6061 2284 6067 2316
rect 6093 2204 6099 2316
rect 6109 2264 6115 2296
rect 6077 2124 6083 2136
rect 5885 1944 5891 2056
rect 5901 1984 5907 2116
rect 5965 1984 5971 2116
rect 6077 2104 6083 2116
rect 6061 2024 6067 2036
rect 5837 1917 5859 1923
rect 5853 1904 5859 1917
rect 5997 1904 6003 1956
rect 5725 1724 5731 1836
rect 5741 1644 5747 1896
rect 5853 1824 5859 1896
rect 6045 1884 6051 1936
rect 6061 1904 6067 1956
rect 5853 1764 5859 1796
rect 5869 1743 5875 1876
rect 6109 1864 6115 1896
rect 6125 1884 6131 2436
rect 6253 2364 6259 2436
rect 6349 2384 6355 2456
rect 6157 2284 6163 2336
rect 6173 2304 6179 2356
rect 6365 2344 6371 2516
rect 6445 2444 6451 2537
rect 6477 2524 6483 2556
rect 6493 2524 6499 2536
rect 6461 2504 6467 2516
rect 6509 2424 6515 2776
rect 6589 2703 6595 2736
rect 6580 2697 6595 2703
rect 6525 2604 6531 2696
rect 6589 2664 6595 2676
rect 6541 2503 6547 2616
rect 6573 2564 6579 2576
rect 6589 2544 6595 2576
rect 6573 2524 6579 2536
rect 6532 2497 6547 2503
rect 6605 2484 6611 2716
rect 6621 2563 6627 2896
rect 6685 2824 6691 2936
rect 6717 2903 6723 2936
rect 6733 2924 6739 2976
rect 6845 2944 6851 2976
rect 6717 2897 6739 2903
rect 6637 2744 6643 2796
rect 6717 2744 6723 2876
rect 6637 2704 6643 2736
rect 6733 2684 6739 2897
rect 6778 2814 6790 2816
rect 6763 2806 6765 2814
rect 6773 2806 6775 2814
rect 6783 2806 6785 2814
rect 6793 2806 6795 2814
rect 6803 2806 6805 2814
rect 6778 2804 6790 2806
rect 6653 2644 6659 2656
rect 6621 2557 6643 2563
rect 6637 2544 6643 2557
rect 6541 2404 6547 2436
rect 6253 2284 6259 2316
rect 6349 2284 6355 2316
rect 6445 2284 6451 2316
rect 6237 2244 6243 2256
rect 6157 2224 6163 2236
rect 6253 2224 6259 2276
rect 6237 2184 6243 2216
rect 6285 2164 6291 2276
rect 6317 2164 6323 2276
rect 6429 2264 6435 2276
rect 6445 2264 6451 2276
rect 6333 2184 6339 2256
rect 6188 2150 6196 2156
rect 6221 2064 6227 2136
rect 6221 1904 6227 2056
rect 6237 1904 6243 2156
rect 6381 2144 6387 2216
rect 6397 2184 6403 2196
rect 6413 2164 6419 2236
rect 6509 2184 6515 2276
rect 6525 2164 6531 2236
rect 6269 2124 6275 2136
rect 6253 1904 6259 2056
rect 6317 1984 6323 2116
rect 6333 2064 6339 2116
rect 6381 2104 6387 2136
rect 6349 1917 6364 1923
rect 6349 1904 6355 1917
rect 6397 1904 6403 2016
rect 6413 1904 6419 2156
rect 6461 2144 6467 2156
rect 6477 2124 6483 2136
rect 6557 2104 6563 2476
rect 6637 2324 6643 2536
rect 6653 2524 6659 2556
rect 6717 2544 6723 2576
rect 6781 2544 6787 2696
rect 6829 2584 6835 2936
rect 6861 2884 6867 2956
rect 6845 2704 6851 2856
rect 6877 2764 6883 2916
rect 6893 2884 6899 3076
rect 6925 3043 6931 3176
rect 6941 3084 6947 3136
rect 6989 3104 6995 3316
rect 7037 3304 7043 3476
rect 7085 3464 7091 3496
rect 7069 3324 7075 3356
rect 7101 3323 7107 3436
rect 7165 3424 7171 3436
rect 7181 3364 7187 3576
rect 7229 3504 7235 4036
rect 7245 3963 7251 4076
rect 7261 3984 7267 4096
rect 7245 3957 7267 3963
rect 7261 3924 7267 3957
rect 7261 3904 7267 3916
rect 7277 3884 7283 3916
rect 7261 3764 7267 3796
rect 7293 3783 7299 4036
rect 7309 3844 7315 3896
rect 7341 3884 7347 4156
rect 7357 3884 7363 3916
rect 7357 3864 7363 3876
rect 7373 3864 7379 4116
rect 7389 4084 7395 4876
rect 7421 4864 7427 5036
rect 7437 4884 7443 5076
rect 7453 5004 7459 5096
rect 7501 5024 7507 5096
rect 7533 4964 7539 5036
rect 7421 4724 7427 4836
rect 7421 4644 7427 4696
rect 7453 4664 7459 4916
rect 7469 4804 7475 4836
rect 7469 4664 7475 4696
rect 7405 4524 7411 4536
rect 7405 4384 7411 4516
rect 7405 4184 7411 4276
rect 7421 4164 7427 4596
rect 7453 4544 7459 4636
rect 7485 4604 7491 4656
rect 7501 4523 7507 4896
rect 7533 4883 7539 4936
rect 7533 4877 7555 4883
rect 7517 4764 7523 4836
rect 7517 4704 7523 4716
rect 7485 4517 7507 4523
rect 7437 4324 7443 4498
rect 7437 4284 7443 4296
rect 7453 4284 7459 4516
rect 7469 4384 7475 4496
rect 7405 4044 7411 4156
rect 7421 4144 7427 4156
rect 7437 3883 7443 4256
rect 7485 4243 7491 4517
rect 7517 4463 7523 4656
rect 7533 4524 7539 4676
rect 7517 4457 7539 4463
rect 7501 4304 7507 4436
rect 7469 4237 7491 4243
rect 7453 4144 7459 4156
rect 7453 4124 7459 4136
rect 7437 3877 7459 3883
rect 7309 3784 7315 3836
rect 7341 3804 7347 3836
rect 7277 3777 7299 3783
rect 7277 3744 7283 3777
rect 7373 3744 7379 3836
rect 7389 3704 7395 3736
rect 7405 3664 7411 3756
rect 7453 3744 7459 3877
rect 7421 3704 7427 3736
rect 7453 3704 7459 3716
rect 7421 3684 7427 3696
rect 7261 3524 7267 3636
rect 7309 3544 7315 3636
rect 7213 3483 7219 3496
rect 7197 3477 7219 3483
rect 7117 3344 7123 3356
rect 7133 3324 7139 3336
rect 7092 3317 7107 3323
rect 7197 3323 7203 3477
rect 7213 3344 7219 3376
rect 7245 3344 7251 3476
rect 7261 3364 7267 3436
rect 7277 3324 7283 3536
rect 7309 3484 7315 3516
rect 7293 3444 7299 3476
rect 7197 3317 7212 3323
rect 7053 3304 7059 3316
rect 7165 3304 7171 3316
rect 7085 3124 7091 3136
rect 6957 3064 6963 3096
rect 6925 3037 6947 3043
rect 6925 2984 6931 3016
rect 6909 2863 6915 2936
rect 6893 2857 6915 2863
rect 6701 2504 6707 2516
rect 6717 2504 6723 2516
rect 6829 2424 6835 2476
rect 6778 2414 6790 2416
rect 6763 2406 6765 2414
rect 6773 2406 6775 2414
rect 6783 2406 6785 2414
rect 6793 2406 6795 2414
rect 6803 2406 6805 2414
rect 6778 2404 6790 2406
rect 6845 2384 6851 2636
rect 6877 2564 6883 2676
rect 6829 2324 6835 2336
rect 6861 2324 6867 2336
rect 6676 2317 6691 2323
rect 6573 2163 6579 2216
rect 6589 2184 6595 2296
rect 6637 2264 6643 2276
rect 6685 2264 6691 2317
rect 6637 2224 6643 2256
rect 6685 2244 6691 2256
rect 6701 2224 6707 2276
rect 6573 2157 6588 2163
rect 6573 2084 6579 2116
rect 6429 1984 6435 2056
rect 6461 1904 6467 1976
rect 6509 1904 6515 1916
rect 6541 1904 6547 1916
rect 6125 1864 6131 1876
rect 5901 1764 5907 1856
rect 6125 1804 6131 1836
rect 5965 1744 5971 1776
rect 6013 1744 6019 1796
rect 6109 1764 6115 1776
rect 6061 1744 6067 1756
rect 5853 1737 5875 1743
rect 5661 1184 5667 1416
rect 5677 1364 5683 1396
rect 5693 1364 5699 1516
rect 5709 1504 5715 1596
rect 5709 1384 5715 1456
rect 5741 1424 5747 1456
rect 5757 1364 5763 1736
rect 5837 1684 5843 1716
rect 5821 1464 5827 1476
rect 5789 1424 5795 1456
rect 5805 1364 5811 1396
rect 5837 1384 5843 1496
rect 5773 1324 5779 1336
rect 5741 1264 5747 1296
rect 5837 1144 5843 1236
rect 5773 1084 5779 1136
rect 5789 1084 5795 1116
rect 5853 1103 5859 1737
rect 5885 1604 5891 1716
rect 5901 1384 5907 1736
rect 6125 1724 6131 1756
rect 6157 1743 6163 1876
rect 6173 1844 6179 1896
rect 6189 1864 6195 1896
rect 6237 1884 6243 1896
rect 6477 1864 6483 1896
rect 6525 1884 6531 1896
rect 6157 1737 6172 1743
rect 6141 1724 6147 1736
rect 6189 1724 6195 1776
rect 6205 1724 6211 1756
rect 6221 1744 6227 1856
rect 6221 1724 6227 1736
rect 6269 1724 6275 1776
rect 6285 1724 6291 1776
rect 6301 1704 6307 1856
rect 6333 1744 6339 1856
rect 6349 1744 6355 1756
rect 6333 1724 6339 1736
rect 6349 1724 6355 1736
rect 6365 1724 6371 1796
rect 5933 1384 5939 1676
rect 5981 1644 5987 1696
rect 6029 1684 6035 1696
rect 5997 1524 6003 1636
rect 5949 1504 5955 1516
rect 6093 1504 6099 1516
rect 6013 1484 6019 1496
rect 5949 1424 5955 1476
rect 5981 1464 5987 1476
rect 5997 1424 6003 1456
rect 5901 1344 5907 1376
rect 5997 1324 6003 1336
rect 5885 1304 5891 1316
rect 5885 1104 5891 1156
rect 5853 1097 5875 1103
rect 5684 957 5699 963
rect 5693 784 5699 957
rect 5709 924 5715 1036
rect 5741 984 5747 1016
rect 5789 944 5795 1076
rect 5837 1064 5843 1076
rect 5757 864 5763 936
rect 5805 924 5811 1036
rect 5853 964 5859 1036
rect 5869 984 5875 1097
rect 5885 964 5891 1096
rect 5997 1084 6003 1316
rect 6013 1104 6019 1356
rect 6029 1344 6035 1416
rect 6045 1324 6051 1496
rect 6125 1484 6131 1496
rect 6061 1404 6067 1476
rect 6061 1344 6067 1396
rect 6077 1384 6083 1476
rect 6109 1384 6115 1476
rect 6205 1463 6211 1696
rect 6221 1484 6227 1636
rect 6333 1564 6339 1636
rect 6237 1484 6243 1496
rect 6285 1484 6291 1556
rect 6333 1524 6339 1536
rect 6365 1524 6371 1716
rect 6413 1703 6419 1736
rect 6429 1724 6435 1756
rect 6509 1744 6515 1876
rect 6541 1864 6547 1896
rect 6589 1864 6595 1896
rect 6605 1864 6611 1876
rect 6557 1744 6563 1776
rect 6413 1697 6435 1703
rect 6317 1464 6323 1516
rect 6397 1504 6403 1516
rect 6365 1484 6371 1496
rect 6381 1464 6387 1496
rect 6429 1484 6435 1697
rect 6445 1684 6451 1736
rect 6573 1724 6579 1836
rect 6589 1744 6595 1776
rect 6621 1744 6627 2036
rect 6637 1903 6643 2176
rect 6701 2164 6707 2196
rect 6653 2144 6659 2156
rect 6669 2104 6675 2116
rect 6717 2084 6723 2096
rect 6717 1984 6723 1996
rect 6637 1897 6652 1903
rect 6685 1864 6691 1936
rect 6733 1923 6739 2316
rect 6781 2144 6787 2276
rect 6893 2264 6899 2857
rect 6941 2684 6947 3037
rect 6989 2924 6995 2956
rect 6973 2684 6979 2836
rect 6941 2664 6947 2676
rect 6941 2624 6947 2636
rect 6957 2564 6963 2576
rect 6909 2503 6915 2516
rect 6941 2503 6947 2516
rect 6989 2504 6995 2656
rect 7005 2504 7011 3116
rect 7021 3044 7027 3076
rect 7037 2984 7043 3076
rect 7021 2924 7027 2956
rect 7053 2924 7059 2976
rect 7069 2944 7075 3096
rect 7085 2964 7091 3036
rect 7101 2984 7107 3076
rect 7117 2944 7123 3276
rect 7021 2644 7027 2916
rect 7069 2704 7075 2756
rect 7117 2704 7123 2896
rect 7133 2884 7139 2956
rect 7149 2944 7155 2996
rect 7165 2964 7171 3056
rect 7181 3004 7187 3096
rect 7197 3084 7203 3236
rect 7213 3124 7219 3316
rect 7309 3264 7315 3376
rect 7325 3364 7331 3516
rect 7341 3363 7347 3576
rect 7357 3504 7363 3636
rect 7357 3384 7363 3496
rect 7373 3484 7379 3496
rect 7389 3464 7395 3656
rect 7405 3504 7411 3636
rect 7437 3504 7443 3516
rect 7453 3504 7459 3516
rect 7469 3503 7475 4237
rect 7501 4223 7507 4276
rect 7485 4217 7507 4223
rect 7485 4184 7491 4217
rect 7517 4184 7523 4256
rect 7485 3664 7491 4076
rect 7501 3903 7507 4136
rect 7517 4084 7523 4156
rect 7501 3897 7516 3903
rect 7501 3884 7507 3897
rect 7533 3883 7539 4457
rect 7549 4164 7555 4877
rect 7565 4784 7571 5096
rect 7549 4104 7555 4116
rect 7517 3877 7539 3883
rect 7485 3524 7491 3636
rect 7501 3584 7507 3696
rect 7517 3683 7523 3877
rect 7533 3704 7539 3856
rect 7517 3677 7539 3683
rect 7517 3584 7523 3616
rect 7469 3497 7491 3503
rect 7373 3424 7379 3456
rect 7437 3444 7443 3476
rect 7389 3404 7395 3436
rect 7453 3384 7459 3456
rect 7485 3364 7491 3497
rect 7501 3464 7507 3556
rect 7341 3357 7363 3363
rect 7325 3324 7331 3336
rect 7341 3324 7347 3336
rect 7341 3084 7347 3256
rect 7357 3104 7363 3357
rect 7453 3337 7468 3343
rect 7405 3304 7411 3336
rect 7421 3304 7427 3316
rect 7437 3104 7443 3116
rect 7341 3063 7347 3076
rect 7389 3063 7395 3076
rect 7341 3057 7363 3063
rect 7213 2944 7219 3036
rect 7229 3024 7235 3056
rect 7172 2897 7187 2903
rect 7133 2764 7139 2876
rect 7149 2704 7155 2716
rect 7117 2684 7123 2696
rect 7165 2683 7171 2716
rect 7181 2704 7187 2897
rect 7165 2677 7187 2683
rect 7037 2544 7043 2636
rect 7053 2564 7059 2676
rect 7053 2544 7059 2556
rect 7053 2524 7059 2536
rect 7085 2524 7091 2636
rect 7101 2544 7107 2616
rect 6909 2497 6947 2503
rect 7101 2503 7107 2516
rect 7085 2497 7107 2503
rect 7085 2484 7091 2497
rect 6909 2284 6915 2456
rect 6925 2304 6931 2456
rect 7053 2384 7059 2436
rect 7117 2384 7123 2416
rect 6941 2284 6947 2376
rect 7085 2284 7091 2336
rect 7101 2317 7132 2323
rect 7101 2304 7107 2317
rect 7149 2303 7155 2676
rect 7165 2504 7171 2636
rect 7181 2484 7187 2677
rect 7197 2584 7203 2716
rect 7213 2704 7219 2736
rect 7213 2524 7219 2596
rect 7165 2324 7171 2376
rect 7197 2304 7203 2316
rect 7149 2297 7171 2303
rect 6877 2184 6883 2256
rect 6900 2237 6915 2243
rect 6893 2184 6899 2216
rect 6749 2104 6755 2116
rect 6778 2014 6790 2016
rect 6763 2006 6765 2014
rect 6773 2006 6775 2014
rect 6783 2006 6785 2014
rect 6793 2006 6795 2014
rect 6803 2006 6805 2014
rect 6778 2004 6790 2006
rect 6733 1917 6755 1923
rect 6733 1884 6739 1896
rect 6749 1884 6755 1917
rect 6829 1904 6835 1916
rect 6909 1904 6915 2237
rect 6973 2164 6979 2176
rect 6989 2144 6995 2156
rect 6925 1984 6931 2116
rect 6989 1984 6995 2136
rect 7005 2124 7011 2216
rect 7037 2204 7043 2276
rect 7085 2264 7091 2276
rect 7053 2183 7059 2256
rect 7085 2184 7091 2216
rect 7037 2177 7059 2183
rect 6925 1904 6931 1956
rect 6861 1897 6876 1903
rect 6493 1683 6499 1716
rect 6557 1704 6563 1716
rect 6477 1677 6499 1683
rect 6445 1504 6451 1516
rect 6205 1457 6227 1463
rect 6221 1384 6227 1457
rect 6237 1424 6243 1456
rect 6269 1444 6275 1456
rect 6429 1384 6435 1456
rect 6445 1444 6451 1476
rect 6109 1344 6115 1376
rect 6445 1364 6451 1396
rect 6141 1323 6147 1356
rect 6205 1344 6211 1356
rect 6132 1317 6147 1323
rect 6157 1104 6163 1176
rect 6253 1124 6259 1136
rect 6285 1124 6291 1356
rect 6333 1344 6339 1356
rect 6445 1344 6451 1356
rect 6317 1144 6323 1316
rect 6333 1304 6339 1336
rect 6477 1284 6483 1677
rect 6493 1464 6499 1476
rect 6509 1464 6515 1496
rect 6573 1444 6579 1476
rect 6509 1324 6515 1336
rect 6525 1304 6531 1356
rect 6589 1344 6595 1736
rect 6621 1703 6627 1736
rect 6637 1724 6643 1836
rect 6733 1764 6739 1776
rect 6685 1744 6691 1756
rect 6605 1697 6627 1703
rect 6605 1364 6611 1697
rect 6653 1684 6659 1696
rect 6749 1684 6755 1876
rect 6813 1864 6819 1896
rect 6861 1804 6867 1897
rect 6941 1883 6947 1916
rect 6957 1904 6963 1976
rect 7005 1904 7011 2096
rect 7012 1897 7027 1903
rect 6925 1877 6947 1883
rect 6877 1844 6883 1876
rect 6893 1864 6899 1876
rect 6813 1724 6819 1756
rect 6877 1744 6883 1776
rect 6829 1724 6835 1736
rect 6877 1724 6883 1736
rect 6893 1724 6899 1796
rect 6861 1704 6867 1716
rect 6925 1704 6931 1877
rect 7005 1844 7011 1876
rect 7021 1803 7027 1897
rect 7005 1797 7027 1803
rect 6749 1644 6755 1676
rect 6637 1484 6643 1636
rect 6778 1614 6790 1616
rect 6763 1606 6765 1614
rect 6773 1606 6775 1614
rect 6783 1606 6785 1614
rect 6793 1606 6795 1614
rect 6803 1606 6805 1614
rect 6778 1604 6790 1606
rect 6701 1504 6707 1516
rect 6861 1504 6867 1696
rect 6941 1684 6947 1736
rect 6957 1724 6963 1756
rect 6973 1744 6979 1756
rect 7005 1724 7011 1797
rect 7021 1744 7027 1776
rect 7037 1704 7043 2177
rect 7101 2164 7107 2196
rect 7117 2143 7123 2296
rect 7165 2184 7171 2297
rect 7149 2144 7155 2176
rect 7181 2163 7187 2276
rect 7213 2244 7219 2316
rect 7229 2223 7235 2916
rect 7245 2664 7251 2756
rect 7261 2604 7267 2696
rect 7261 2303 7267 2536
rect 7277 2343 7283 2776
rect 7325 2744 7331 2936
rect 7357 2804 7363 3057
rect 7389 3057 7404 3063
rect 7373 3004 7379 3036
rect 7373 2784 7379 2976
rect 7389 2944 7395 3057
rect 7453 2984 7459 3337
rect 7469 3064 7475 3316
rect 7485 3184 7491 3356
rect 7501 3184 7507 3436
rect 7517 3364 7523 3556
rect 7533 3444 7539 3677
rect 7517 3303 7523 3336
rect 7517 3297 7539 3303
rect 7485 3063 7491 3116
rect 7533 3063 7539 3297
rect 7476 3057 7491 3063
rect 7485 2944 7491 3057
rect 7517 3057 7539 3063
rect 7389 2904 7395 2936
rect 7373 2704 7379 2716
rect 7293 2544 7299 2696
rect 7309 2644 7315 2696
rect 7389 2664 7395 2736
rect 7453 2664 7459 2756
rect 7469 2724 7475 2876
rect 7501 2863 7507 3036
rect 7517 2884 7523 3057
rect 7533 2864 7539 2916
rect 7501 2857 7523 2863
rect 7485 2703 7491 2856
rect 7501 2764 7507 2836
rect 7485 2697 7507 2703
rect 7357 2644 7363 2656
rect 7309 2544 7315 2576
rect 7341 2564 7347 2596
rect 7357 2544 7363 2556
rect 7389 2484 7395 2516
rect 7341 2384 7347 2436
rect 7277 2337 7299 2343
rect 7261 2297 7283 2303
rect 7245 2264 7251 2296
rect 7261 2264 7267 2276
rect 7213 2217 7235 2223
rect 7181 2157 7196 2163
rect 7101 2137 7123 2143
rect 7101 2084 7107 2137
rect 7181 2124 7187 2157
rect 7213 2084 7219 2217
rect 7229 2104 7235 2116
rect 7053 1743 7059 1876
rect 7069 1844 7075 1896
rect 7085 1884 7091 1896
rect 7181 1844 7187 2076
rect 7261 1863 7267 1896
rect 7252 1857 7267 1863
rect 7117 1784 7123 1816
rect 7053 1737 7068 1743
rect 7005 1684 7011 1696
rect 6973 1504 6979 1516
rect 6653 1464 6659 1496
rect 6669 1464 6675 1476
rect 6717 1463 6723 1496
rect 6717 1457 6739 1463
rect 6685 1424 6691 1436
rect 6733 1384 6739 1457
rect 6781 1444 6787 1476
rect 6861 1444 6867 1476
rect 6925 1424 6931 1496
rect 6989 1484 6995 1516
rect 7005 1504 7011 1536
rect 7053 1524 7059 1737
rect 7133 1664 7139 1736
rect 7021 1484 7027 1496
rect 7021 1464 7027 1476
rect 6957 1384 6963 1456
rect 7053 1424 7059 1436
rect 7053 1384 7059 1396
rect 6557 1304 6563 1336
rect 6429 1184 6435 1276
rect 6589 1144 6595 1256
rect 6605 1144 6611 1336
rect 6653 1144 6659 1316
rect 6909 1264 6915 1336
rect 6778 1214 6790 1216
rect 6763 1206 6765 1214
rect 6773 1206 6775 1214
rect 6783 1206 6785 1214
rect 6793 1206 6795 1214
rect 6803 1206 6805 1214
rect 6778 1204 6790 1206
rect 6477 1124 6483 1136
rect 6509 1104 6515 1116
rect 6013 1084 6019 1096
rect 6125 1084 6131 1096
rect 5917 984 5923 996
rect 5965 944 5971 1036
rect 6109 944 6115 1076
rect 6141 964 6147 1036
rect 6157 984 6163 1096
rect 6221 1064 6227 1096
rect 6365 1084 6371 1096
rect 6189 984 6195 1056
rect 6157 964 6163 976
rect 6253 944 6259 1036
rect 6269 984 6275 1076
rect 6301 940 6307 1036
rect 5821 884 5827 936
rect 5837 924 5843 936
rect 6013 924 6019 936
rect 6029 924 6035 936
rect 6333 924 6339 1056
rect 6381 964 6387 1036
rect 6429 984 6435 1036
rect 6541 1024 6547 1056
rect 6573 1044 6579 1096
rect 6621 1084 6627 1116
rect 6637 1064 6643 1096
rect 6653 1084 6659 1136
rect 6669 1064 6675 1096
rect 6685 1063 6691 1096
rect 6685 1057 6707 1063
rect 6509 984 6515 996
rect 6573 984 6579 1016
rect 6701 984 6707 1057
rect 6717 984 6723 1136
rect 6893 1124 6899 1236
rect 6957 1184 6963 1296
rect 6973 1264 6979 1356
rect 7037 1344 7043 1356
rect 7069 1344 7075 1356
rect 7085 1323 7091 1336
rect 7069 1317 7091 1323
rect 7053 1184 7059 1276
rect 6852 1097 6867 1103
rect 6733 1044 6739 1056
rect 6381 944 6387 956
rect 6445 944 6451 956
rect 6541 924 6547 936
rect 5389 684 5395 716
rect 5309 424 5315 536
rect 5373 504 5379 636
rect 5421 564 5427 636
rect 5453 564 5459 696
rect 5661 684 5667 716
rect 5789 703 5795 836
rect 5885 784 5891 916
rect 5949 904 5955 916
rect 6045 884 6051 916
rect 5933 784 5939 836
rect 6045 724 6051 876
rect 5789 697 5804 703
rect 5789 684 5795 697
rect 5533 663 5539 676
rect 5533 657 5555 663
rect 5405 504 5411 516
rect 5348 497 5356 503
rect 5421 484 5427 536
rect 5469 504 5475 636
rect 5517 544 5523 636
rect 5549 544 5555 657
rect 5645 624 5651 676
rect 5757 643 5763 676
rect 5773 644 5779 656
rect 5741 637 5763 643
rect 5565 564 5571 576
rect 4973 143 4979 256
rect 4973 137 4988 143
rect 4589 84 4595 116
rect 4685 84 4691 116
rect 4797 104 4803 136
rect 5005 124 5011 236
rect 4829 104 4835 116
rect 4861 104 4867 116
rect 5037 84 5043 276
rect 5085 224 5091 276
rect 5101 204 5107 356
rect 5149 284 5155 296
rect 5117 277 5132 283
rect 5117 264 5123 277
rect 5165 264 5171 396
rect 5197 284 5203 356
rect 5213 284 5219 296
rect 5053 84 5059 116
rect 5069 104 5075 176
rect 5133 164 5139 256
rect 5181 224 5187 236
rect 5197 164 5203 196
rect 5101 144 5107 156
rect 5085 124 5091 136
rect 5197 104 5203 118
rect 5213 104 5219 216
rect 5229 184 5235 316
rect 5341 304 5347 316
rect 5252 297 5267 303
rect 5261 284 5267 297
rect 5341 284 5347 296
rect 5274 214 5286 216
rect 5259 206 5261 214
rect 5269 206 5271 214
rect 5279 206 5281 214
rect 5289 206 5291 214
rect 5299 206 5301 214
rect 5274 204 5286 206
rect 5325 204 5331 236
rect 5357 224 5363 316
rect 5389 304 5395 456
rect 5469 444 5475 476
rect 5469 324 5475 436
rect 5517 404 5523 516
rect 5549 484 5555 536
rect 5597 504 5603 556
rect 5629 504 5635 516
rect 5645 504 5651 536
rect 5677 503 5683 636
rect 5709 524 5715 636
rect 5741 584 5747 637
rect 5789 584 5795 656
rect 5741 544 5747 576
rect 5805 556 5811 656
rect 5853 544 5859 636
rect 5869 624 5875 676
rect 5901 644 5907 716
rect 6013 704 6019 716
rect 5981 644 5987 696
rect 6029 684 6035 696
rect 5997 664 6003 676
rect 5901 584 5907 616
rect 5997 584 6003 656
rect 6029 584 6035 656
rect 5981 544 5987 556
rect 5661 497 5683 503
rect 5613 384 5619 476
rect 5645 424 5651 496
rect 5405 284 5411 316
rect 5469 264 5475 316
rect 5629 297 5644 303
rect 5597 264 5603 276
rect 5437 244 5443 256
rect 5597 244 5603 256
rect 5325 184 5331 196
rect 5405 104 5411 216
rect 5421 124 5427 196
rect 5437 84 5443 236
rect 5485 144 5491 156
rect 5629 124 5635 297
rect 5661 264 5667 497
rect 5709 444 5715 516
rect 5693 364 5699 436
rect 5645 184 5651 236
rect 5693 184 5699 236
rect 5661 124 5667 176
rect 5709 124 5715 396
rect 5725 284 5731 296
rect 5741 284 5747 496
rect 5805 384 5811 456
rect 5869 324 5875 536
rect 6045 504 6051 556
rect 6061 524 6067 796
rect 6077 704 6083 896
rect 6141 704 6147 876
rect 6333 824 6339 916
rect 6333 784 6339 816
rect 6509 784 6515 896
rect 6541 864 6547 916
rect 6557 904 6563 956
rect 6605 924 6611 976
rect 6653 924 6659 956
rect 6477 704 6483 736
rect 6285 664 6291 676
rect 6349 664 6355 676
rect 6269 604 6275 636
rect 5757 124 5763 176
rect 5789 164 5795 276
rect 5821 264 5827 276
rect 5885 264 5891 276
rect 5933 264 5939 276
rect 5853 164 5859 196
rect 5885 144 5891 156
rect 5805 124 5811 136
rect 5517 104 5523 118
rect 5917 103 5923 236
rect 5949 164 5955 376
rect 5965 304 5971 316
rect 6077 284 6083 536
rect 6093 324 6099 596
rect 6109 464 6115 516
rect 6141 484 6147 556
rect 6157 504 6163 556
rect 6141 384 6147 456
rect 6237 384 6243 516
rect 6253 484 6259 536
rect 6253 364 6259 476
rect 6269 444 6275 536
rect 6173 284 6179 316
rect 6269 284 6275 436
rect 6285 324 6291 656
rect 6301 524 6307 616
rect 6333 384 6339 636
rect 6349 324 6355 656
rect 6413 584 6419 636
rect 6509 584 6515 756
rect 6541 664 6547 856
rect 6557 704 6563 776
rect 6381 544 6387 556
rect 6477 524 6483 576
rect 6525 563 6531 636
rect 6541 563 6547 656
rect 6573 584 6579 676
rect 6525 557 6547 563
rect 6541 544 6547 557
rect 6557 524 6563 556
rect 6365 504 6371 516
rect 6397 503 6403 516
rect 6429 503 6435 516
rect 6397 497 6435 503
rect 6285 304 6291 316
rect 6397 284 6403 356
rect 6445 344 6451 436
rect 6573 384 6579 556
rect 6413 284 6419 316
rect 6589 304 6595 776
rect 6605 704 6611 916
rect 6653 664 6659 916
rect 6733 904 6739 956
rect 6861 944 6867 1097
rect 6877 984 6883 1036
rect 6829 924 6835 936
rect 6861 904 6867 936
rect 6717 704 6723 716
rect 6733 684 6739 896
rect 6893 884 6899 1096
rect 6941 1064 6947 1076
rect 6925 944 6931 1056
rect 6957 984 6963 1056
rect 6941 944 6947 956
rect 6957 904 6963 976
rect 6973 864 6979 956
rect 6989 944 6995 1096
rect 7005 1004 7011 1136
rect 7069 1103 7075 1317
rect 7101 1104 7107 1436
rect 7117 1384 7123 1456
rect 7133 1364 7139 1436
rect 7149 1364 7155 1836
rect 7229 1783 7235 1836
rect 7245 1804 7251 1856
rect 7213 1777 7235 1783
rect 7213 1756 7219 1777
rect 7277 1723 7283 2297
rect 7293 2264 7299 2337
rect 7437 2304 7443 2356
rect 7309 2144 7315 2156
rect 7309 1924 7315 2136
rect 7293 1724 7299 1896
rect 7261 1717 7283 1723
rect 7165 1684 7171 1716
rect 7197 1684 7203 1716
rect 7165 1524 7171 1676
rect 7181 1504 7187 1656
rect 7261 1644 7267 1717
rect 7309 1684 7315 1736
rect 7293 1664 7299 1676
rect 7325 1624 7331 2216
rect 7357 2184 7363 2236
rect 7389 2203 7395 2264
rect 7389 2197 7411 2203
rect 7341 2144 7347 2176
rect 7373 2124 7379 2156
rect 7405 1963 7411 2197
rect 7421 2144 7427 2276
rect 7453 2244 7459 2516
rect 7469 2484 7475 2616
rect 7485 2524 7491 2676
rect 7469 2184 7475 2316
rect 7485 2304 7491 2516
rect 7501 2184 7507 2697
rect 7517 2683 7523 2857
rect 7533 2704 7539 2836
rect 7517 2677 7539 2683
rect 7517 2344 7523 2516
rect 7533 2504 7539 2677
rect 7533 2384 7539 2476
rect 7549 2404 7555 4076
rect 7565 3924 7571 4296
rect 7565 3884 7571 3896
rect 7565 3724 7571 3736
rect 7533 2144 7539 2156
rect 7389 1957 7411 1963
rect 7389 1924 7395 1957
rect 7341 1884 7347 1916
rect 7389 1904 7395 1916
rect 7405 1884 7411 1936
rect 7341 1864 7347 1876
rect 7357 1744 7363 1836
rect 7373 1764 7379 1776
rect 7389 1744 7395 1756
rect 7421 1744 7427 1796
rect 7437 1743 7443 2116
rect 7469 1984 7475 2096
rect 7453 1904 7459 1916
rect 7485 1864 7491 1916
rect 7533 1903 7539 2136
rect 7524 1897 7539 1903
rect 7453 1784 7459 1856
rect 7453 1764 7459 1776
rect 7437 1737 7459 1743
rect 7357 1723 7363 1736
rect 7348 1717 7363 1723
rect 7181 1443 7187 1476
rect 7245 1444 7251 1464
rect 7181 1437 7203 1443
rect 7133 1184 7139 1336
rect 7197 1304 7203 1437
rect 7229 1344 7235 1356
rect 7069 1097 7091 1103
rect 7069 1044 7075 1056
rect 6778 814 6790 816
rect 6763 806 6765 814
rect 6773 806 6775 814
rect 6783 806 6785 814
rect 6793 806 6795 814
rect 6803 806 6805 814
rect 6778 804 6790 806
rect 6925 704 6931 716
rect 6653 604 6659 656
rect 6621 564 6627 596
rect 6701 584 6707 676
rect 6829 664 6835 696
rect 6941 683 6947 716
rect 6941 677 6956 683
rect 6852 577 6883 583
rect 6877 564 6883 577
rect 6509 284 6515 296
rect 6157 277 6172 283
rect 6013 264 6019 276
rect 6125 264 6131 276
rect 6157 264 6163 277
rect 6276 277 6284 283
rect 6205 264 6211 276
rect 6221 264 6227 276
rect 6253 264 6259 276
rect 6260 257 6275 263
rect 6029 164 6035 236
rect 5933 124 5939 136
rect 6109 104 6115 236
rect 6173 104 6179 236
rect 6237 164 6243 216
rect 6269 144 6275 257
rect 6285 124 6291 236
rect 6381 124 6387 136
rect 6413 123 6419 276
rect 6477 144 6483 236
rect 6541 184 6547 296
rect 6621 263 6627 556
rect 6653 523 6659 556
rect 6701 544 6707 556
rect 6812 550 6820 556
rect 6941 544 6947 596
rect 6957 584 6963 676
rect 6973 563 6979 836
rect 7005 743 7011 956
rect 6989 737 7011 743
rect 6989 664 6995 737
rect 6989 564 6995 576
rect 6957 557 6979 563
rect 6781 524 6787 536
rect 6653 517 6668 523
rect 6669 384 6675 516
rect 6877 483 6883 536
rect 6893 524 6899 536
rect 6877 477 6899 483
rect 6778 414 6790 416
rect 6763 406 6765 414
rect 6773 406 6775 414
rect 6783 406 6785 414
rect 6793 406 6795 414
rect 6803 406 6805 414
rect 6778 404 6790 406
rect 6669 364 6675 376
rect 6877 304 6883 316
rect 6685 264 6691 276
rect 6829 264 6835 276
rect 6861 264 6867 276
rect 6621 257 6636 263
rect 6589 124 6595 236
rect 6637 164 6643 256
rect 6717 244 6723 256
rect 6637 144 6643 156
rect 6669 144 6675 236
rect 6413 117 6428 123
rect 6189 104 6195 116
rect 6317 104 6323 116
rect 6333 104 6339 116
rect 6701 104 6707 136
rect 6717 124 6723 236
rect 6749 184 6755 216
rect 6781 124 6787 156
rect 6877 123 6883 276
rect 6893 204 6899 477
rect 6925 444 6931 516
rect 6868 117 6883 123
rect 5917 97 5932 103
rect 6909 103 6915 236
rect 6957 223 6963 557
rect 6989 343 6995 556
rect 7005 384 7011 716
rect 7037 657 7052 663
rect 7037 584 7043 657
rect 7069 583 7075 636
rect 7085 584 7091 1097
rect 7101 964 7107 1056
rect 7117 1044 7123 1096
rect 7133 944 7139 1076
rect 7133 904 7139 916
rect 7101 704 7107 876
rect 7133 784 7139 876
rect 7149 763 7155 1096
rect 7165 923 7171 1296
rect 7181 1284 7187 1296
rect 7245 1104 7251 1356
rect 7277 1344 7283 1616
rect 7293 1364 7299 1476
rect 7309 1324 7315 1456
rect 7357 1384 7363 1476
rect 7405 1344 7411 1376
rect 7453 1344 7459 1737
rect 7469 1543 7475 1836
rect 7485 1584 7491 1696
rect 7501 1684 7507 1856
rect 7517 1784 7523 1896
rect 7533 1784 7539 1876
rect 7549 1864 7555 2236
rect 7549 1804 7555 1836
rect 7565 1743 7571 3696
rect 7549 1737 7571 1743
rect 7469 1537 7491 1543
rect 7469 1464 7475 1476
rect 7485 1383 7491 1537
rect 7469 1377 7491 1383
rect 7293 1304 7299 1316
rect 7181 1084 7187 1096
rect 7197 984 7203 1096
rect 7245 1004 7251 1096
rect 7197 944 7203 976
rect 7261 924 7267 1276
rect 7293 1104 7299 1296
rect 7277 984 7283 1056
rect 7309 984 7315 996
rect 7165 917 7187 923
rect 7181 784 7187 917
rect 7197 864 7203 916
rect 7133 757 7155 763
rect 7053 577 7075 583
rect 7053 564 7059 577
rect 7053 544 7059 556
rect 7133 444 7139 757
rect 7213 743 7219 916
rect 7197 737 7219 743
rect 7149 503 7155 696
rect 7165 524 7171 536
rect 7181 504 7187 556
rect 7149 497 7171 503
rect 7165 344 7171 497
rect 6973 337 6995 343
rect 6973 284 6979 337
rect 7197 343 7203 737
rect 7309 704 7315 736
rect 7229 624 7235 696
rect 7325 644 7331 1336
rect 7405 1104 7411 1336
rect 7469 1264 7475 1377
rect 7485 1284 7491 1356
rect 7501 1324 7507 1456
rect 7469 1104 7475 1236
rect 7373 1084 7379 1096
rect 7469 1064 7475 1076
rect 7501 1064 7507 1316
rect 7517 1064 7523 1076
rect 7341 944 7347 1036
rect 7373 984 7379 1036
rect 7405 963 7411 1036
rect 7517 984 7523 1016
rect 7533 1004 7539 1636
rect 7549 1104 7555 1737
rect 7565 1484 7571 1496
rect 7565 1284 7571 1296
rect 7389 957 7411 963
rect 7357 944 7363 956
rect 7341 704 7347 716
rect 7357 684 7363 936
rect 7389 903 7395 957
rect 7380 897 7395 903
rect 7405 784 7411 936
rect 7421 924 7427 956
rect 7389 724 7395 736
rect 7229 524 7235 616
rect 7437 584 7443 696
rect 7533 684 7539 916
rect 7549 784 7555 916
rect 7197 337 7219 343
rect 6989 284 6995 316
rect 6973 264 6979 276
rect 7005 264 7011 296
rect 6941 217 6963 223
rect 6941 184 6947 217
rect 6973 164 6979 196
rect 7005 164 7011 256
rect 7021 224 7027 336
rect 7149 284 7155 316
rect 7053 164 7059 276
rect 7149 204 7155 276
rect 7197 244 7203 316
rect 7213 304 7219 337
rect 7293 324 7299 476
rect 7373 444 7379 516
rect 7405 323 7411 436
rect 7396 317 7411 323
rect 7197 157 7212 163
rect 6925 144 6931 156
rect 6957 144 6963 156
rect 7037 144 7043 156
rect 7197 124 7203 157
rect 7229 144 7235 316
rect 7373 304 7379 316
rect 7405 304 7411 317
rect 7245 164 7251 236
rect 7261 184 7267 296
rect 7309 144 7315 156
rect 7357 144 7363 296
rect 7421 284 7427 556
rect 7453 384 7459 636
rect 7501 564 7507 576
rect 7469 304 7475 336
rect 7421 264 7427 276
rect 7437 264 7443 276
rect 7389 184 7395 236
rect 7421 156 7427 256
rect 7388 150 7396 156
rect 7485 144 7491 276
rect 7501 184 7507 536
rect 7517 284 7523 296
rect 7533 284 7539 436
rect 7565 344 7571 1256
rect 6900 97 6915 103
rect 7101 103 7107 116
rect 7101 97 7123 103
rect 7117 84 7123 97
rect 5421 64 5427 76
rect 2509 -17 2515 36
rect 3261 -17 3267 36
rect 3309 -17 3315 36
rect 2509 -23 2531 -17
rect 3245 -23 3267 -17
rect 3293 -23 3315 -17
rect 3565 -17 3571 36
rect 3645 -17 3651 36
rect 3770 14 3782 16
rect 3755 6 3757 14
rect 3765 6 3767 14
rect 3775 6 3777 14
rect 3785 6 3787 14
rect 3795 6 3797 14
rect 3770 4 3782 6
rect 4045 -17 4051 36
rect 4093 -17 4099 36
rect 4925 -17 4931 36
rect 3565 -23 3587 -17
rect 3629 -23 3651 -17
rect 4029 -23 4051 -17
rect 4077 -23 4099 -17
rect 4909 -23 4931 -17
rect 5677 -23 5683 16
rect 5693 -17 5699 36
rect 5693 -23 5715 -17
rect 5741 -23 5747 36
rect 5789 -17 5795 36
rect 5837 -17 5843 36
rect 6013 -17 6019 36
rect 5773 -23 5795 -17
rect 5821 -23 5843 -17
rect 5997 -23 6019 -17
rect 6061 -17 6067 36
rect 6365 -17 6371 36
rect 6413 -17 6419 36
rect 6461 -17 6467 36
rect 6621 -17 6627 36
rect 6778 14 6790 16
rect 6763 6 6765 14
rect 6773 6 6775 14
rect 6783 6 6785 14
rect 6793 6 6795 14
rect 6803 6 6805 14
rect 6778 4 6790 6
rect 6061 -23 6083 -17
rect 6349 -23 6371 -17
rect 6397 -23 6419 -17
rect 6445 -23 6467 -17
rect 6605 -23 6627 -17
rect 7165 -17 7171 36
rect 7165 -23 7187 -17
<< m3contact >>
rect 3852 5216 3860 5224
rect 3884 5216 3892 5224
rect 739 5206 747 5214
rect 749 5206 757 5214
rect 759 5206 767 5214
rect 769 5206 777 5214
rect 779 5206 787 5214
rect 789 5206 797 5214
rect 3747 5206 3755 5214
rect 3757 5206 3765 5214
rect 3767 5206 3775 5214
rect 3777 5206 3785 5214
rect 3787 5206 3795 5214
rect 3797 5206 3805 5214
rect 380 5116 388 5124
rect 476 5116 484 5124
rect 1020 5116 1028 5124
rect 1100 5116 1108 5124
rect 2732 5116 2740 5124
rect 2892 5116 2900 5124
rect 3420 5116 3428 5124
rect 3580 5116 3588 5124
rect 204 5096 212 5104
rect 124 5076 132 5084
rect 76 5036 84 5044
rect 76 4956 84 4964
rect 188 5016 196 5024
rect 188 4936 196 4944
rect 220 5056 228 5064
rect 268 5056 276 5064
rect 316 5056 324 5064
rect 396 5056 404 5064
rect 236 5036 244 5044
rect 348 5036 356 5044
rect 300 5016 308 5024
rect 236 4956 244 4964
rect 268 4936 276 4944
rect 380 4936 388 4944
rect 220 4916 228 4924
rect 300 4916 308 4924
rect 316 4916 324 4924
rect 108 4756 116 4764
rect 12 4556 20 4564
rect 204 4756 212 4764
rect 124 4676 132 4684
rect 44 4516 52 4524
rect 92 4516 100 4524
rect 188 4656 196 4664
rect 156 4576 164 4584
rect 188 4556 196 4564
rect 300 4856 308 4864
rect 348 4736 356 4744
rect 268 4676 276 4684
rect 220 4536 228 4544
rect 300 4536 308 4544
rect 332 4536 340 4544
rect 236 4516 244 4524
rect 284 4516 292 4524
rect 76 4276 84 4284
rect 76 4116 84 4124
rect 76 3916 84 3924
rect 124 3876 132 3884
rect 76 3716 84 3724
rect 844 5096 852 5104
rect 444 5076 452 5084
rect 684 5076 692 5084
rect 412 4976 420 4984
rect 604 5036 612 5044
rect 748 5036 756 5044
rect 476 4936 484 4944
rect 428 4916 436 4924
rect 412 4736 420 4744
rect 572 4896 580 4904
rect 492 4816 500 4824
rect 556 4816 564 4824
rect 492 4756 500 4764
rect 460 4716 468 4724
rect 364 4696 372 4704
rect 460 4696 468 4704
rect 444 4676 452 4684
rect 396 4636 404 4644
rect 428 4636 436 4644
rect 620 4936 628 4944
rect 716 4936 724 4944
rect 764 4916 772 4924
rect 652 4836 660 4844
rect 684 4836 692 4844
rect 604 4796 612 4804
rect 572 4736 580 4744
rect 556 4696 564 4704
rect 604 4696 612 4704
rect 636 4696 644 4704
rect 524 4676 532 4684
rect 380 4536 388 4544
rect 396 4536 404 4544
rect 460 4536 468 4544
rect 412 4516 420 4524
rect 508 4516 516 4524
rect 380 4496 388 4504
rect 348 4456 356 4464
rect 396 4456 404 4464
rect 220 4296 228 4304
rect 300 4296 308 4304
rect 188 4256 196 4264
rect 188 4156 196 4164
rect 236 4276 244 4284
rect 268 4256 276 4264
rect 268 4156 276 4164
rect 220 4136 228 4144
rect 396 4336 404 4344
rect 444 4456 452 4464
rect 460 4356 468 4364
rect 428 4316 436 4324
rect 380 4296 388 4304
rect 428 4296 436 4304
rect 364 4276 372 4284
rect 380 4256 388 4264
rect 412 4256 420 4264
rect 428 4256 436 4264
rect 348 4236 356 4244
rect 332 4216 340 4224
rect 348 4176 356 4184
rect 332 4156 340 4164
rect 364 4156 372 4164
rect 204 4076 212 4084
rect 236 4116 244 4124
rect 300 4116 308 4124
rect 252 3916 260 3924
rect 332 3916 340 3924
rect 236 3896 244 3904
rect 284 3896 292 3904
rect 412 3896 420 3904
rect 332 3876 340 3884
rect 220 3856 228 3864
rect 316 3796 324 3804
rect 204 3756 212 3764
rect 236 3736 244 3744
rect 284 3736 292 3744
rect 300 3736 308 3744
rect 364 3776 372 3784
rect 476 4216 484 4224
rect 620 4676 628 4684
rect 572 4656 580 4664
rect 556 4556 564 4564
rect 812 4896 820 4904
rect 748 4876 756 4884
rect 700 4816 708 4824
rect 684 4796 692 4804
rect 668 4676 676 4684
rect 668 4556 676 4564
rect 604 4536 612 4544
rect 540 4516 548 4524
rect 588 4516 596 4524
rect 508 4496 516 4504
rect 524 4496 532 4504
rect 524 4276 532 4284
rect 556 4376 564 4384
rect 572 4236 580 4244
rect 540 4216 548 4224
rect 492 4196 500 4204
rect 588 4196 596 4204
rect 492 4176 500 4184
rect 476 4096 484 4104
rect 636 4516 644 4524
rect 739 4806 747 4814
rect 749 4806 757 4814
rect 759 4806 767 4814
rect 769 4806 777 4814
rect 779 4806 787 4814
rect 789 4806 797 4814
rect 828 4876 836 4884
rect 700 4776 708 4784
rect 700 4716 708 4724
rect 812 4716 820 4724
rect 716 4696 724 4704
rect 732 4696 740 4704
rect 892 5056 900 5064
rect 972 5056 980 5064
rect 876 4936 884 4944
rect 908 5036 916 5044
rect 924 4996 932 5004
rect 1036 5096 1044 5104
rect 1292 5102 1300 5104
rect 1004 4956 1012 4964
rect 940 4936 948 4944
rect 924 4916 932 4924
rect 860 4816 868 4824
rect 860 4736 868 4744
rect 860 4716 868 4724
rect 844 4696 852 4704
rect 700 4636 708 4644
rect 700 4476 708 4484
rect 636 4336 644 4344
rect 684 4336 692 4344
rect 620 4216 628 4224
rect 668 4256 676 4264
rect 652 4176 660 4184
rect 604 4156 612 4164
rect 652 4156 660 4164
rect 684 4176 692 4184
rect 572 4116 580 4124
rect 620 4116 628 4124
rect 572 4096 580 4104
rect 556 4036 564 4044
rect 540 3916 548 3924
rect 524 3896 532 3904
rect 508 3856 516 3864
rect 684 4096 692 4104
rect 668 4056 676 4064
rect 636 3916 644 3924
rect 620 3896 628 3904
rect 588 3876 596 3884
rect 556 3836 564 3844
rect 524 3776 532 3784
rect 428 3736 436 3744
rect 252 3716 260 3724
rect 236 3696 244 3704
rect 172 3516 180 3524
rect 12 3476 20 3484
rect 124 3476 132 3484
rect 172 3476 180 3484
rect 12 3436 20 3444
rect 188 3356 196 3364
rect 332 3696 340 3704
rect 428 3696 436 3704
rect 300 3636 308 3644
rect 348 3636 356 3644
rect 380 3636 388 3644
rect 332 3516 340 3524
rect 316 3476 324 3484
rect 364 3496 372 3504
rect 332 3356 340 3364
rect 124 3316 132 3324
rect 156 3316 164 3324
rect 236 3316 244 3324
rect 492 3716 500 3724
rect 492 3696 500 3704
rect 508 3696 516 3704
rect 492 3676 500 3684
rect 412 3496 420 3504
rect 460 3496 468 3504
rect 476 3496 484 3504
rect 380 3456 388 3464
rect 444 3456 452 3464
rect 460 3356 468 3364
rect 412 3336 420 3344
rect 588 3718 596 3724
rect 588 3716 596 3718
rect 604 3716 612 3724
rect 796 4536 804 4544
rect 828 4656 836 4664
rect 860 4536 868 4544
rect 860 4516 868 4524
rect 828 4476 836 4484
rect 739 4406 747 4414
rect 749 4406 757 4414
rect 759 4406 767 4414
rect 769 4406 777 4414
rect 779 4406 787 4414
rect 789 4406 797 4414
rect 812 4356 820 4364
rect 732 4336 740 4344
rect 780 4296 788 4304
rect 764 4276 772 4284
rect 844 4416 852 4424
rect 860 4336 868 4344
rect 860 4316 868 4324
rect 892 4836 900 4844
rect 1292 5096 1300 5102
rect 1516 5096 1524 5104
rect 1740 5096 1748 5104
rect 1804 5096 1812 5104
rect 1836 5096 1844 5104
rect 1964 5096 1972 5104
rect 2108 5096 2116 5104
rect 2236 5096 2244 5104
rect 2412 5096 2420 5104
rect 2492 5096 2500 5104
rect 2508 5096 2516 5104
rect 1068 5076 1076 5084
rect 1500 5076 1508 5084
rect 1468 5056 1476 5064
rect 1516 5056 1524 5064
rect 1100 5036 1108 5044
rect 1052 5016 1060 5024
rect 1276 5016 1284 5024
rect 1228 4996 1236 5004
rect 1164 4976 1172 4984
rect 1116 4936 1124 4944
rect 1180 4936 1188 4944
rect 1212 4936 1220 4944
rect 1020 4916 1028 4924
rect 1132 4916 1140 4924
rect 1068 4896 1076 4904
rect 1148 4896 1156 4904
rect 1020 4816 1028 4824
rect 1004 4796 1012 4804
rect 908 4736 916 4744
rect 892 4696 900 4704
rect 1004 4696 1012 4704
rect 908 4676 916 4684
rect 924 4656 932 4664
rect 972 4656 980 4664
rect 924 4636 932 4644
rect 956 4616 964 4624
rect 988 4596 996 4604
rect 988 4556 996 4564
rect 1052 4656 1060 4664
rect 1020 4516 1028 4524
rect 908 4356 916 4364
rect 908 4336 916 4344
rect 1196 4816 1204 4824
rect 1212 4756 1220 4764
rect 1116 4736 1124 4744
rect 1148 4696 1156 4704
rect 1132 4656 1140 4664
rect 1084 4636 1092 4644
rect 1116 4636 1124 4644
rect 1164 4636 1172 4644
rect 1052 4496 1060 4504
rect 956 4436 964 4444
rect 1020 4396 1028 4404
rect 1068 4476 1076 4484
rect 1068 4356 1076 4364
rect 1020 4296 1028 4304
rect 876 4276 884 4284
rect 796 4256 804 4264
rect 828 4256 836 4264
rect 860 4236 868 4244
rect 828 4216 836 4224
rect 796 4176 804 4184
rect 796 4156 804 4164
rect 812 4136 820 4144
rect 764 4096 772 4104
rect 812 4076 820 4084
rect 716 4036 724 4044
rect 739 4006 747 4014
rect 749 4006 757 4014
rect 759 4006 767 4014
rect 769 4006 777 4014
rect 779 4006 787 4014
rect 789 4006 797 4014
rect 908 4236 916 4244
rect 876 4216 884 4224
rect 876 4176 884 4184
rect 892 4156 900 4164
rect 972 4256 980 4264
rect 1052 4256 1060 4264
rect 1068 4256 1076 4264
rect 1052 4216 1060 4224
rect 956 4196 964 4204
rect 1148 4596 1156 4604
rect 1228 4556 1236 4564
rect 1420 5036 1428 5044
rect 1436 5036 1444 5044
rect 1404 4936 1412 4944
rect 1292 4916 1300 4924
rect 1340 4896 1348 4904
rect 1340 4776 1348 4784
rect 1308 4716 1316 4724
rect 1116 4536 1124 4544
rect 1244 4536 1252 4544
rect 1116 4516 1124 4524
rect 1148 4516 1156 4524
rect 1164 4516 1172 4524
rect 1164 4476 1172 4484
rect 1244 4516 1252 4524
rect 1212 4496 1220 4504
rect 1276 4496 1284 4504
rect 1196 4436 1204 4444
rect 1180 4336 1188 4344
rect 1100 4216 1108 4224
rect 924 4136 932 4144
rect 940 4136 948 4144
rect 1004 4136 1012 4144
rect 876 4116 884 4124
rect 956 4116 964 4124
rect 1004 4116 1012 4124
rect 844 4096 852 4104
rect 924 4096 932 4104
rect 988 4096 996 4104
rect 924 4076 932 4084
rect 1036 4056 1044 4064
rect 860 3976 868 3984
rect 956 3976 964 3984
rect 844 3836 852 3844
rect 1164 4276 1172 4284
rect 1324 4596 1332 4604
rect 1356 4716 1364 4724
rect 1356 4696 1364 4704
rect 1372 4676 1380 4684
rect 1356 4576 1364 4584
rect 1308 4516 1316 4524
rect 1356 4516 1364 4524
rect 1292 4456 1300 4464
rect 1196 4276 1204 4284
rect 1212 4276 1220 4284
rect 1196 4176 1204 4184
rect 1196 4118 1204 4124
rect 1196 4116 1204 4118
rect 1180 4056 1188 4064
rect 1148 3956 1156 3964
rect 1116 3936 1124 3944
rect 1052 3916 1060 3924
rect 1148 3916 1156 3924
rect 908 3896 916 3904
rect 972 3896 980 3904
rect 908 3876 916 3884
rect 860 3816 868 3824
rect 716 3776 724 3784
rect 876 3776 884 3784
rect 796 3756 804 3764
rect 796 3736 804 3744
rect 924 3776 932 3784
rect 940 3756 948 3764
rect 908 3716 916 3724
rect 739 3606 747 3614
rect 749 3606 757 3614
rect 759 3606 767 3614
rect 769 3606 777 3614
rect 779 3606 787 3614
rect 789 3606 797 3614
rect 796 3556 804 3564
rect 844 3676 852 3684
rect 924 3676 932 3684
rect 876 3616 884 3624
rect 636 3536 644 3544
rect 812 3536 820 3544
rect 844 3536 852 3544
rect 620 3496 628 3504
rect 700 3496 708 3504
rect 748 3496 756 3504
rect 556 3476 564 3484
rect 524 3456 532 3464
rect 652 3416 660 3424
rect 524 3336 532 3344
rect 44 3096 52 3104
rect 92 3096 100 3104
rect 156 3096 164 3104
rect 252 3096 260 3104
rect 348 3096 356 3104
rect 12 2976 20 2984
rect 12 2656 20 2664
rect 12 2596 20 2604
rect 92 2936 100 2944
rect 428 3116 436 3124
rect 572 3316 580 3324
rect 604 3136 612 3144
rect 636 3136 644 3144
rect 572 3116 580 3124
rect 620 3116 628 3124
rect 556 3096 564 3104
rect 364 3036 372 3044
rect 476 3036 484 3044
rect 540 3036 548 3044
rect 252 2956 260 2964
rect 300 2956 308 2964
rect 348 2956 356 2964
rect 108 2856 116 2864
rect 220 2916 228 2924
rect 236 2916 244 2924
rect 204 2856 212 2864
rect 284 2936 292 2944
rect 268 2916 276 2924
rect 124 2676 132 2684
rect 204 2656 212 2664
rect 140 2576 148 2584
rect 220 2576 228 2584
rect 172 2536 180 2544
rect 140 2518 148 2524
rect 140 2516 148 2518
rect 236 2436 244 2444
rect 428 2976 436 2984
rect 428 2936 436 2944
rect 524 2936 532 2944
rect 300 2916 308 2924
rect 348 2916 356 2924
rect 380 2916 388 2924
rect 476 2916 484 2924
rect 300 2876 308 2884
rect 300 2856 308 2864
rect 444 2896 452 2904
rect 412 2756 420 2764
rect 364 2716 372 2724
rect 316 2696 324 2704
rect 364 2696 372 2704
rect 428 2696 436 2704
rect 300 2576 308 2584
rect 300 2556 308 2564
rect 284 2516 292 2524
rect 252 2376 260 2384
rect 268 2356 276 2364
rect 428 2656 436 2664
rect 364 2616 372 2624
rect 364 2596 372 2604
rect 540 2856 548 2864
rect 460 2836 468 2844
rect 460 2736 468 2744
rect 444 2636 452 2644
rect 396 2576 404 2584
rect 364 2556 372 2564
rect 332 2516 340 2524
rect 348 2516 356 2524
rect 428 2518 436 2524
rect 428 2516 436 2518
rect 508 2716 516 2724
rect 556 2776 564 2784
rect 636 3076 644 3084
rect 620 2956 628 2964
rect 572 2736 580 2744
rect 524 2696 532 2704
rect 540 2696 548 2704
rect 588 2696 596 2704
rect 476 2656 484 2664
rect 636 2916 644 2924
rect 812 3456 820 3464
rect 684 3376 692 3384
rect 764 3376 772 3384
rect 716 3296 724 3304
rect 700 3276 708 3284
rect 684 3236 692 3244
rect 668 3136 676 3144
rect 700 3136 708 3144
rect 684 3096 692 3104
rect 739 3206 747 3214
rect 749 3206 757 3214
rect 759 3206 767 3214
rect 769 3206 777 3214
rect 779 3206 787 3214
rect 789 3206 797 3214
rect 716 3096 724 3104
rect 748 3096 756 3104
rect 668 3036 676 3044
rect 668 2976 676 2984
rect 796 3036 804 3044
rect 796 2996 804 3004
rect 860 3516 868 3524
rect 860 3496 868 3504
rect 892 3516 900 3524
rect 956 3696 964 3704
rect 940 3616 948 3624
rect 940 3576 948 3584
rect 908 3496 916 3504
rect 924 3496 932 3504
rect 860 3396 868 3404
rect 1036 3876 1044 3884
rect 1052 3876 1060 3884
rect 988 3756 996 3764
rect 1004 3756 1012 3764
rect 1052 3756 1060 3764
rect 1020 3736 1028 3744
rect 1036 3716 1044 3724
rect 1116 3856 1124 3864
rect 1132 3836 1140 3844
rect 1260 4316 1268 4324
rect 1324 4336 1332 4344
rect 1276 4276 1284 4284
rect 1388 4636 1396 4644
rect 1388 4576 1396 4584
rect 1404 4536 1412 4544
rect 1388 4436 1396 4444
rect 1372 4296 1380 4304
rect 1324 4256 1332 4264
rect 1292 4136 1300 4144
rect 1292 4116 1300 4124
rect 1260 4036 1268 4044
rect 1356 4236 1364 4244
rect 1660 5076 1668 5084
rect 1772 5076 1780 5084
rect 1548 5036 1556 5044
rect 1580 5036 1588 5044
rect 1532 4956 1540 4964
rect 1532 4936 1540 4944
rect 1484 4916 1492 4924
rect 1452 4702 1460 4704
rect 1452 4696 1460 4702
rect 1468 4676 1476 4684
rect 1468 4596 1476 4604
rect 1436 4576 1444 4584
rect 1420 4496 1428 4504
rect 1388 4256 1396 4264
rect 1356 4116 1364 4124
rect 1404 4136 1412 4144
rect 1388 4116 1396 4124
rect 1516 4896 1524 4904
rect 1516 4716 1524 4724
rect 1772 5036 1780 5044
rect 1708 4996 1716 5004
rect 1612 4976 1620 4984
rect 1660 4956 1668 4964
rect 1580 4916 1588 4924
rect 1596 4776 1604 4784
rect 1564 4736 1572 4744
rect 1564 4696 1572 4704
rect 1580 4636 1588 4644
rect 1548 4596 1556 4604
rect 1564 4576 1572 4584
rect 1548 4556 1556 4564
rect 1484 4536 1492 4544
rect 1500 4536 1508 4544
rect 1660 4916 1668 4924
rect 1628 4856 1636 4864
rect 1676 4796 1684 4804
rect 1836 5076 1844 5084
rect 1884 5076 1892 5084
rect 2012 5076 2020 5084
rect 1852 5036 1860 5044
rect 1884 4996 1892 5004
rect 1788 4976 1796 4984
rect 1724 4956 1732 4964
rect 1724 4936 1732 4944
rect 2060 5056 2068 5064
rect 2044 4976 2052 4984
rect 2172 5076 2180 5084
rect 2252 5076 2260 5084
rect 2140 5036 2148 5044
rect 2140 5016 2148 5024
rect 2348 5056 2356 5064
rect 2243 5006 2251 5014
rect 2253 5006 2261 5014
rect 2263 5006 2271 5014
rect 2273 5006 2281 5014
rect 2283 5006 2291 5014
rect 2293 5006 2301 5014
rect 1820 4918 1828 4924
rect 1820 4916 1828 4918
rect 2044 4916 2052 4924
rect 2108 4916 2116 4924
rect 2124 4916 2132 4924
rect 2156 4916 2164 4924
rect 1756 4896 1764 4904
rect 1948 4896 1956 4904
rect 1980 4896 1988 4904
rect 1964 4876 1972 4884
rect 1804 4776 1812 4784
rect 1948 4776 1956 4784
rect 1708 4716 1716 4724
rect 1868 4736 1876 4744
rect 1900 4736 1908 4744
rect 1836 4716 1844 4724
rect 1644 4702 1652 4704
rect 1644 4696 1652 4702
rect 1820 4696 1828 4704
rect 1772 4676 1780 4684
rect 1660 4656 1668 4664
rect 1644 4616 1652 4624
rect 1612 4556 1620 4564
rect 1788 4656 1796 4664
rect 1772 4616 1780 4624
rect 1740 4576 1748 4584
rect 1820 4576 1828 4584
rect 1708 4556 1716 4564
rect 1772 4556 1780 4564
rect 1676 4536 1684 4544
rect 1500 4516 1508 4524
rect 1532 4516 1540 4524
rect 1612 4516 1620 4524
rect 1468 4496 1476 4504
rect 1452 4336 1460 4344
rect 1548 4456 1556 4464
rect 1660 4396 1668 4404
rect 1644 4356 1652 4364
rect 1484 4336 1492 4344
rect 1516 4336 1524 4344
rect 1612 4336 1620 4344
rect 1516 4316 1524 4324
rect 1452 4276 1460 4284
rect 1500 4256 1508 4264
rect 1468 4116 1476 4124
rect 1452 4076 1460 4084
rect 1388 4056 1396 4064
rect 1436 4056 1444 4064
rect 1372 4016 1380 4024
rect 1276 3996 1284 4004
rect 1292 3936 1300 3944
rect 1356 3936 1364 3944
rect 1260 3916 1268 3924
rect 1324 3896 1332 3904
rect 1228 3796 1236 3804
rect 1228 3776 1236 3784
rect 988 3616 996 3624
rect 1180 3716 1188 3724
rect 1196 3716 1204 3724
rect 1132 3696 1140 3704
rect 1196 3696 1204 3704
rect 1100 3656 1108 3664
rect 1068 3616 1076 3624
rect 1084 3536 1092 3544
rect 1052 3496 1060 3504
rect 1116 3496 1124 3504
rect 1100 3476 1108 3484
rect 988 3456 996 3464
rect 1036 3456 1044 3464
rect 1020 3396 1028 3404
rect 1052 3396 1060 3404
rect 940 3376 948 3384
rect 924 3336 932 3344
rect 1036 3376 1044 3384
rect 956 3336 964 3344
rect 1052 3316 1060 3324
rect 1068 3316 1076 3324
rect 876 3296 884 3304
rect 908 3296 916 3304
rect 972 3296 980 3304
rect 892 3276 900 3284
rect 956 3176 964 3184
rect 940 3116 948 3124
rect 860 3096 868 3104
rect 844 3056 852 3064
rect 908 3056 916 3064
rect 988 3056 996 3064
rect 1004 3056 1012 3064
rect 828 2956 836 2964
rect 860 2956 868 2964
rect 716 2916 724 2924
rect 739 2806 747 2814
rect 749 2806 757 2814
rect 759 2806 767 2814
rect 769 2806 777 2814
rect 779 2806 787 2814
rect 789 2806 797 2814
rect 652 2702 660 2704
rect 652 2696 660 2702
rect 620 2676 628 2684
rect 572 2656 580 2664
rect 652 2656 660 2664
rect 524 2636 532 2644
rect 604 2636 612 2644
rect 476 2556 484 2564
rect 492 2536 500 2544
rect 460 2496 468 2504
rect 316 2456 324 2464
rect 412 2436 420 2444
rect 364 2396 372 2404
rect 156 2296 164 2304
rect 204 2296 212 2304
rect 220 2296 228 2304
rect 252 2296 260 2304
rect 268 2296 276 2304
rect 12 2156 20 2164
rect 12 1936 20 1944
rect 12 1796 20 1804
rect 12 1356 20 1364
rect 188 2276 196 2284
rect 236 2280 244 2284
rect 236 2276 244 2280
rect 44 2156 52 2164
rect 156 2156 164 2164
rect 204 2156 212 2164
rect 44 2136 52 2144
rect 92 2136 100 2144
rect 172 2136 180 2144
rect 76 2116 84 2124
rect 124 2116 132 2124
rect 188 2116 196 2124
rect 76 2096 84 2104
rect 108 2076 116 2084
rect 332 2276 340 2284
rect 428 2256 436 2264
rect 508 2416 516 2424
rect 492 2316 500 2324
rect 588 2616 596 2624
rect 556 2576 564 2584
rect 636 2616 644 2624
rect 572 2356 580 2364
rect 604 2356 612 2364
rect 316 2156 324 2164
rect 444 2156 452 2164
rect 476 2156 484 2164
rect 284 2136 292 2144
rect 252 2116 260 2124
rect 268 2116 276 2124
rect 380 2136 388 2144
rect 332 2116 340 2124
rect 348 2096 356 2104
rect 396 2096 404 2104
rect 476 2076 484 2084
rect 204 2016 212 2024
rect 412 1976 420 1984
rect 492 1956 500 1964
rect 300 1936 308 1944
rect 220 1916 228 1924
rect 268 1916 276 1924
rect 140 1902 148 1904
rect 140 1896 148 1902
rect 236 1896 244 1904
rect 540 2256 548 2264
rect 572 2256 580 2264
rect 556 2236 564 2244
rect 556 2196 564 2204
rect 620 2316 628 2324
rect 524 2116 532 2124
rect 540 2116 548 2124
rect 556 2096 564 2104
rect 540 2076 548 2084
rect 572 2076 580 2084
rect 604 2076 612 2084
rect 524 1956 532 1964
rect 556 1916 564 1924
rect 508 1896 516 1904
rect 172 1876 180 1884
rect 332 1876 340 1884
rect 204 1856 212 1864
rect 140 1736 148 1744
rect 108 1716 116 1724
rect 316 1836 324 1844
rect 300 1796 308 1804
rect 236 1736 244 1744
rect 220 1716 228 1724
rect 268 1716 276 1724
rect 220 1696 228 1704
rect 364 1836 372 1844
rect 524 1856 532 1864
rect 476 1756 484 1764
rect 716 2636 724 2644
rect 780 2636 788 2644
rect 780 2596 788 2604
rect 764 2536 772 2544
rect 812 2536 820 2544
rect 739 2406 747 2414
rect 749 2406 757 2414
rect 759 2406 767 2414
rect 769 2406 777 2414
rect 779 2406 787 2414
rect 789 2406 797 2414
rect 812 2356 820 2364
rect 860 2936 868 2944
rect 844 2796 852 2804
rect 828 2316 836 2324
rect 828 2296 836 2304
rect 684 2216 692 2224
rect 732 2216 740 2224
rect 924 2956 932 2964
rect 972 2956 980 2964
rect 908 2916 916 2924
rect 892 2856 900 2864
rect 876 2836 884 2844
rect 892 2836 900 2844
rect 860 2756 868 2764
rect 860 2716 868 2724
rect 1004 2996 1012 3004
rect 1068 3176 1076 3184
rect 1180 3476 1188 3484
rect 1116 3456 1124 3464
rect 1116 3316 1124 3324
rect 1116 3136 1124 3144
rect 1068 2976 1076 2984
rect 1164 3316 1172 3324
rect 1292 3718 1300 3724
rect 1292 3716 1300 3718
rect 1308 3496 1316 3504
rect 1436 4036 1444 4044
rect 1484 3996 1492 4004
rect 1420 3956 1428 3964
rect 1356 3836 1364 3844
rect 1340 3796 1348 3804
rect 1468 3856 1476 3864
rect 1420 3776 1428 3784
rect 1404 3736 1412 3744
rect 1388 3636 1396 3644
rect 1340 3556 1348 3564
rect 1532 4276 1540 4284
rect 1580 4276 1588 4284
rect 1548 4256 1556 4264
rect 1532 4236 1540 4244
rect 1564 4236 1572 4244
rect 1532 4136 1540 4144
rect 1628 4276 1636 4284
rect 1596 4216 1604 4224
rect 1708 4496 1716 4504
rect 1740 4516 1748 4524
rect 1772 4516 1780 4524
rect 1740 4396 1748 4404
rect 1756 4376 1764 4384
rect 1692 4216 1700 4224
rect 1628 4196 1636 4204
rect 1676 4196 1684 4204
rect 1596 4176 1604 4184
rect 1612 4156 1620 4164
rect 1580 4136 1588 4144
rect 1532 4016 1540 4024
rect 1516 3976 1524 3984
rect 1516 3936 1524 3944
rect 1660 4156 1668 4164
rect 1804 4416 1812 4424
rect 1916 4696 1924 4704
rect 1964 4696 1972 4704
rect 1852 4656 1860 4664
rect 1932 4676 1940 4684
rect 1916 4656 1924 4664
rect 1900 4616 1908 4624
rect 1868 4576 1876 4584
rect 1900 4496 1908 4504
rect 1852 4436 1860 4444
rect 1868 4296 1876 4304
rect 1788 4216 1796 4224
rect 1788 4196 1796 4204
rect 1676 4136 1684 4144
rect 1756 4136 1764 4144
rect 1884 4216 1892 4224
rect 1836 4176 1844 4184
rect 1820 4156 1828 4164
rect 1804 4136 1812 4144
rect 1740 4116 1748 4124
rect 1740 4096 1748 4104
rect 1724 4076 1732 4084
rect 1628 3976 1636 3984
rect 1548 3936 1556 3944
rect 1580 3936 1588 3944
rect 1612 3936 1620 3944
rect 1548 3896 1556 3904
rect 1516 3876 1524 3884
rect 1644 3876 1652 3884
rect 1484 3736 1492 3744
rect 1468 3696 1476 3704
rect 1468 3616 1476 3624
rect 1500 3616 1508 3624
rect 1452 3536 1460 3544
rect 1244 3456 1252 3464
rect 1244 3376 1252 3384
rect 1212 3316 1220 3324
rect 1196 3296 1204 3304
rect 1308 3296 1316 3304
rect 1148 3276 1156 3284
rect 1148 3236 1156 3244
rect 1196 3216 1204 3224
rect 1276 3196 1284 3204
rect 1324 3196 1332 3204
rect 1196 3116 1204 3124
rect 1244 3116 1252 3124
rect 1132 3056 1140 3064
rect 956 2896 964 2904
rect 956 2856 964 2864
rect 1036 2916 1044 2924
rect 988 2896 996 2904
rect 972 2796 980 2804
rect 1052 2796 1060 2804
rect 1052 2756 1060 2764
rect 1020 2716 1028 2724
rect 892 2676 900 2684
rect 1068 2716 1076 2724
rect 1036 2696 1044 2704
rect 1084 2696 1092 2704
rect 940 2676 948 2684
rect 1004 2676 1012 2684
rect 908 2656 916 2664
rect 940 2636 948 2644
rect 1020 2636 1028 2644
rect 972 2616 980 2624
rect 1020 2616 1028 2624
rect 956 2596 964 2604
rect 988 2536 996 2544
rect 940 2436 948 2444
rect 1052 2576 1060 2584
rect 1228 2936 1236 2944
rect 1116 2916 1124 2924
rect 1260 2916 1268 2924
rect 1116 2776 1124 2784
rect 1148 2696 1156 2704
rect 1132 2676 1140 2684
rect 1212 2856 1220 2864
rect 1244 2836 1252 2844
rect 1292 3116 1300 3124
rect 1436 3496 1444 3504
rect 1452 3496 1460 3504
rect 1356 3456 1364 3464
rect 1500 3476 1508 3484
rect 1388 3396 1396 3404
rect 1356 3336 1364 3344
rect 1404 3276 1412 3284
rect 1692 3856 1700 3864
rect 1692 3816 1700 3824
rect 1612 3696 1620 3704
rect 1788 3976 1796 3984
rect 1772 3936 1780 3944
rect 1900 4156 1908 4164
rect 1836 4076 1844 4084
rect 1852 4076 1860 4084
rect 1820 3896 1828 3904
rect 1964 4676 1972 4684
rect 2076 4896 2084 4904
rect 2220 4856 2228 4864
rect 2060 4776 2068 4784
rect 2092 4776 2100 4784
rect 2044 4696 2052 4704
rect 2236 4776 2244 4784
rect 2188 4736 2196 4744
rect 2172 4696 2180 4704
rect 1996 4676 2004 4684
rect 2028 4676 2036 4684
rect 1980 4656 1988 4664
rect 1980 4576 1988 4584
rect 1932 4536 1940 4544
rect 2604 5096 2612 5104
rect 2764 5096 2772 5104
rect 2860 5096 2868 5104
rect 3036 5096 3044 5104
rect 3052 5096 3060 5104
rect 3212 5102 3220 5104
rect 3212 5096 3220 5102
rect 3276 5096 3284 5104
rect 3532 5096 3540 5104
rect 3708 5096 3716 5104
rect 2476 5076 2484 5084
rect 2572 5076 2580 5084
rect 2412 5036 2420 5044
rect 2476 5036 2484 5044
rect 2444 5016 2452 5024
rect 2380 4956 2388 4964
rect 2540 5056 2548 5064
rect 2492 4996 2500 5004
rect 2460 4956 2468 4964
rect 2572 4956 2580 4964
rect 2492 4936 2500 4944
rect 2636 5076 2644 5084
rect 2716 5036 2724 5044
rect 2700 5016 2708 5024
rect 2716 5016 2724 5024
rect 2780 4976 2788 4984
rect 2764 4956 2772 4964
rect 2364 4916 2372 4924
rect 2444 4916 2452 4924
rect 2524 4916 2532 4924
rect 2620 4916 2628 4924
rect 2668 4916 2676 4924
rect 2588 4876 2596 4884
rect 2156 4676 2164 4684
rect 2220 4676 2228 4684
rect 2284 4676 2292 4684
rect 2108 4656 2116 4664
rect 2012 4616 2020 4624
rect 2060 4616 2068 4624
rect 2060 4556 2068 4564
rect 1996 4536 2004 4544
rect 2044 4536 2052 4544
rect 1964 4516 1972 4524
rect 2012 4516 2020 4524
rect 2076 4516 2084 4524
rect 1932 4496 1940 4504
rect 2028 4496 2036 4504
rect 2140 4616 2148 4624
rect 2124 4576 2132 4584
rect 2156 4556 2164 4564
rect 2124 4536 2132 4544
rect 2108 4496 2116 4504
rect 2092 4416 2100 4424
rect 2092 4296 2100 4304
rect 1980 4236 1988 4244
rect 1996 4216 2004 4224
rect 1948 4136 1956 4144
rect 1932 4116 1940 4124
rect 1852 3996 1860 4004
rect 1868 3996 1876 4004
rect 1900 3896 1908 3904
rect 1820 3876 1828 3884
rect 1964 3996 1972 4004
rect 1884 3816 1892 3824
rect 1852 3776 1860 3784
rect 1804 3736 1812 3744
rect 1836 3736 1844 3744
rect 1884 3716 1892 3724
rect 1724 3676 1732 3684
rect 1660 3576 1668 3584
rect 1660 3556 1668 3564
rect 1676 3556 1684 3564
rect 1628 3496 1636 3504
rect 1548 3476 1556 3484
rect 1532 3456 1540 3464
rect 1436 3376 1444 3384
rect 1532 3376 1540 3384
rect 1564 3376 1572 3384
rect 1516 3356 1524 3364
rect 1436 3316 1444 3324
rect 1420 3136 1428 3144
rect 1308 3056 1316 3064
rect 1308 3016 1316 3024
rect 1292 2996 1300 3004
rect 1388 3036 1396 3044
rect 1404 3016 1412 3024
rect 1388 2976 1396 2984
rect 1340 2936 1348 2944
rect 1356 2936 1364 2944
rect 1388 2936 1396 2944
rect 1356 2916 1364 2924
rect 1308 2836 1316 2844
rect 1292 2796 1300 2804
rect 1276 2716 1284 2724
rect 1212 2696 1220 2704
rect 1180 2676 1188 2684
rect 1244 2676 1252 2684
rect 1164 2656 1172 2664
rect 1196 2656 1204 2664
rect 1164 2616 1172 2624
rect 1116 2596 1124 2604
rect 1132 2516 1140 2524
rect 1260 2616 1268 2624
rect 1260 2576 1268 2584
rect 1068 2496 1076 2504
rect 1116 2496 1124 2504
rect 988 2336 996 2344
rect 1100 2476 1108 2484
rect 1132 2476 1140 2484
rect 1100 2376 1108 2384
rect 1068 2316 1076 2324
rect 1228 2496 1236 2504
rect 1420 2936 1428 2944
rect 1404 2896 1412 2904
rect 1340 2816 1348 2824
rect 1356 2816 1364 2824
rect 1420 2816 1428 2824
rect 1356 2776 1364 2784
rect 1340 2756 1348 2764
rect 1340 2736 1348 2744
rect 1404 2696 1412 2704
rect 1372 2676 1380 2684
rect 1388 2656 1396 2664
rect 1356 2616 1364 2624
rect 1356 2576 1364 2584
rect 1372 2556 1380 2564
rect 1340 2536 1348 2544
rect 1468 3216 1476 3224
rect 1468 2876 1476 2884
rect 1452 2856 1460 2864
rect 1468 2836 1476 2844
rect 1436 2736 1444 2744
rect 1436 2676 1444 2684
rect 1436 2616 1444 2624
rect 1420 2596 1428 2604
rect 1452 2576 1460 2584
rect 1404 2556 1412 2564
rect 1452 2516 1460 2524
rect 1308 2356 1316 2364
rect 1196 2336 1204 2344
rect 1292 2336 1300 2344
rect 1180 2316 1188 2324
rect 860 2296 868 2304
rect 924 2302 932 2304
rect 924 2296 932 2302
rect 1324 2316 1332 2324
rect 1324 2296 1332 2304
rect 1372 2336 1380 2344
rect 1452 2496 1460 2504
rect 1420 2396 1428 2404
rect 1500 2956 1508 2964
rect 1564 3236 1572 3244
rect 1628 3256 1636 3264
rect 1612 3216 1620 3224
rect 1772 3596 1780 3604
rect 1740 3576 1748 3584
rect 1724 3536 1732 3544
rect 1724 3516 1732 3524
rect 1676 3496 1684 3504
rect 1692 3496 1700 3504
rect 1756 3496 1764 3504
rect 1708 3476 1716 3484
rect 1676 3356 1684 3364
rect 1724 3356 1732 3364
rect 1756 3356 1764 3364
rect 1820 3576 1828 3584
rect 1836 3496 1844 3504
rect 1852 3496 1860 3504
rect 1868 3476 1876 3484
rect 1868 3436 1876 3444
rect 1932 3876 1940 3884
rect 1948 3776 1956 3784
rect 2044 4276 2052 4284
rect 2076 4256 2084 4264
rect 2012 4196 2020 4204
rect 2108 4196 2116 4204
rect 2204 4516 2212 4524
rect 2172 4476 2180 4484
rect 2156 4456 2164 4464
rect 2140 4216 2148 4224
rect 2092 4176 2100 4184
rect 2124 4176 2132 4184
rect 2028 4116 2036 4124
rect 2044 3996 2052 4004
rect 2172 4296 2180 4304
rect 2124 4116 2132 4124
rect 2140 4076 2148 4084
rect 2140 3976 2148 3984
rect 2060 3916 2068 3924
rect 1996 3896 2004 3904
rect 2012 3876 2020 3884
rect 2124 3836 2132 3844
rect 1948 3756 1956 3764
rect 1980 3756 1988 3764
rect 1996 3756 2004 3764
rect 1916 3716 1924 3724
rect 2188 4236 2196 4244
rect 2243 4606 2251 4614
rect 2253 4606 2261 4614
rect 2263 4606 2271 4614
rect 2273 4606 2281 4614
rect 2283 4606 2291 4614
rect 2293 4606 2301 4614
rect 2396 4596 2404 4604
rect 2316 4576 2324 4584
rect 2268 4556 2276 4564
rect 2236 4476 2244 4484
rect 2252 4456 2260 4464
rect 2556 4796 2564 4804
rect 2572 4736 2580 4744
rect 2508 4656 2516 4664
rect 2508 4616 2516 4624
rect 2620 4796 2628 4804
rect 2652 4796 2660 4804
rect 2604 4756 2612 4764
rect 2556 4656 2564 4664
rect 2588 4656 2596 4664
rect 2540 4596 2548 4604
rect 2524 4556 2532 4564
rect 2604 4616 2612 4624
rect 2636 4616 2644 4624
rect 2620 4596 2628 4604
rect 2556 4556 2564 4564
rect 2604 4556 2612 4564
rect 2412 4536 2420 4544
rect 2428 4516 2436 4524
rect 2508 4516 2516 4524
rect 2540 4516 2548 4524
rect 2396 4496 2404 4504
rect 2524 4496 2532 4504
rect 2332 4456 2340 4464
rect 2332 4416 2340 4424
rect 2348 4376 2356 4384
rect 2243 4206 2251 4214
rect 2253 4206 2261 4214
rect 2263 4206 2271 4214
rect 2273 4206 2281 4214
rect 2283 4206 2291 4214
rect 2293 4206 2301 4214
rect 2236 4176 2244 4184
rect 2188 4156 2196 4164
rect 2220 4156 2228 4164
rect 2172 4036 2180 4044
rect 2156 3876 2164 3884
rect 2140 3816 2148 3824
rect 2156 3776 2164 3784
rect 2076 3756 2084 3764
rect 2220 3936 2228 3944
rect 2252 3856 2260 3864
rect 2243 3806 2251 3814
rect 2253 3806 2261 3814
rect 2263 3806 2271 3814
rect 2273 3806 2281 3814
rect 2283 3806 2291 3814
rect 2293 3806 2301 3814
rect 2252 3776 2260 3784
rect 2220 3756 2228 3764
rect 2028 3736 2036 3744
rect 2140 3736 2148 3744
rect 2188 3736 2196 3744
rect 2252 3736 2260 3744
rect 1996 3716 2004 3724
rect 2044 3716 2052 3724
rect 1932 3696 1940 3704
rect 1996 3596 2004 3604
rect 1900 3556 1908 3564
rect 1980 3536 1988 3544
rect 1948 3516 1956 3524
rect 2028 3596 2036 3604
rect 2028 3576 2036 3584
rect 2044 3576 2052 3584
rect 2012 3536 2020 3544
rect 2012 3516 2020 3524
rect 2140 3676 2148 3684
rect 2172 3636 2180 3644
rect 2092 3556 2100 3564
rect 2092 3536 2100 3544
rect 2092 3516 2100 3524
rect 2156 3516 2164 3524
rect 2124 3496 2132 3504
rect 2172 3496 2180 3504
rect 1932 3476 1940 3484
rect 1916 3416 1924 3424
rect 1884 3396 1892 3404
rect 2012 3456 2020 3464
rect 1996 3436 2004 3444
rect 1948 3356 1956 3364
rect 1964 3356 1972 3364
rect 1852 3336 1860 3344
rect 1916 3336 1924 3344
rect 1788 3296 1796 3304
rect 1852 3296 1860 3304
rect 1740 3256 1748 3264
rect 1724 3236 1732 3244
rect 1660 3156 1668 3164
rect 1596 3116 1604 3124
rect 1644 3056 1652 3064
rect 1548 2956 1556 2964
rect 1516 2936 1524 2944
rect 1532 2916 1540 2924
rect 1500 2856 1508 2864
rect 1580 2956 1588 2964
rect 1676 2956 1684 2964
rect 1756 3036 1764 3044
rect 1724 2996 1732 3004
rect 1740 2996 1748 3004
rect 1772 2976 1780 2984
rect 1820 3196 1828 3204
rect 1740 2956 1748 2964
rect 1788 2956 1796 2964
rect 1708 2936 1716 2944
rect 1788 2936 1796 2944
rect 1676 2916 1684 2924
rect 1772 2916 1780 2924
rect 1980 3316 1988 3324
rect 1884 3216 1892 3224
rect 1868 3176 1876 3184
rect 1948 3096 1956 3104
rect 1884 3036 1892 3044
rect 1868 2996 1876 3004
rect 1484 2776 1492 2784
rect 1532 2776 1540 2784
rect 1564 2836 1572 2844
rect 1660 2816 1668 2824
rect 1628 2756 1636 2764
rect 1564 2716 1572 2724
rect 1596 2696 1604 2704
rect 1660 2696 1668 2704
rect 1644 2676 1652 2684
rect 1484 2636 1492 2644
rect 1516 2636 1524 2644
rect 1804 2896 1812 2904
rect 1852 2896 1860 2904
rect 1724 2836 1732 2844
rect 1692 2796 1700 2804
rect 1708 2736 1716 2744
rect 1756 2776 1764 2784
rect 1788 2736 1796 2744
rect 1772 2696 1780 2704
rect 1708 2676 1716 2684
rect 1740 2676 1748 2684
rect 1676 2656 1684 2664
rect 1500 2596 1508 2604
rect 1484 2536 1492 2544
rect 1500 2536 1508 2544
rect 1532 2616 1540 2624
rect 1548 2616 1556 2624
rect 1580 2556 1588 2564
rect 1532 2516 1540 2524
rect 1564 2516 1572 2524
rect 1500 2476 1508 2484
rect 1564 2476 1572 2484
rect 1484 2416 1492 2424
rect 1468 2376 1476 2384
rect 1388 2316 1396 2324
rect 1484 2316 1492 2324
rect 860 2276 868 2284
rect 1340 2276 1348 2284
rect 1404 2276 1412 2284
rect 668 2136 676 2144
rect 812 2136 820 2144
rect 1100 2176 1108 2184
rect 1372 2256 1380 2264
rect 1068 2136 1076 2144
rect 1132 2136 1140 2144
rect 1180 2136 1188 2144
rect 1228 2136 1236 2144
rect 652 2116 660 2124
rect 684 2116 692 2124
rect 924 2116 932 2124
rect 652 2076 660 2084
rect 732 2076 740 2084
rect 732 2036 740 2044
rect 739 2006 747 2014
rect 749 2006 757 2014
rect 759 2006 767 2014
rect 769 2006 777 2014
rect 779 2006 787 2014
rect 789 2006 797 2014
rect 652 1956 660 1964
rect 828 1896 836 1904
rect 620 1876 628 1884
rect 668 1856 676 1864
rect 572 1796 580 1804
rect 588 1796 596 1804
rect 572 1776 580 1784
rect 652 1776 660 1784
rect 588 1756 596 1764
rect 380 1716 388 1724
rect 428 1716 436 1724
rect 412 1536 420 1544
rect 540 1716 548 1724
rect 508 1696 516 1704
rect 556 1696 564 1704
rect 508 1636 516 1644
rect 44 1496 52 1504
rect 108 1496 116 1504
rect 140 1496 148 1504
rect 220 1496 228 1504
rect 444 1496 452 1504
rect 492 1496 500 1504
rect 124 1416 132 1424
rect 300 1456 308 1464
rect 188 1376 196 1384
rect 380 1436 388 1444
rect 428 1416 436 1424
rect 380 1376 388 1384
rect 284 1336 292 1344
rect 412 1336 420 1344
rect 172 1316 180 1324
rect 252 1318 260 1324
rect 252 1316 260 1318
rect 364 1236 372 1244
rect 380 1176 388 1184
rect 460 1156 468 1164
rect 156 1036 164 1044
rect 268 996 276 1004
rect 220 936 228 944
rect 12 776 20 784
rect 188 876 196 884
rect 252 936 260 944
rect 316 1036 324 1044
rect 284 956 292 964
rect 300 936 308 944
rect 636 1536 644 1544
rect 604 1516 612 1524
rect 524 1496 532 1504
rect 540 1496 548 1504
rect 780 1876 788 1884
rect 844 1816 852 1824
rect 844 1756 852 1764
rect 684 1736 692 1744
rect 652 1496 660 1504
rect 668 1476 676 1484
rect 572 1456 580 1464
rect 700 1716 708 1724
rect 748 1676 756 1684
rect 739 1606 747 1614
rect 749 1606 757 1614
rect 759 1606 767 1614
rect 769 1606 777 1614
rect 779 1606 787 1614
rect 789 1606 797 1614
rect 908 2076 916 2084
rect 988 2116 996 2124
rect 1068 2116 1076 2124
rect 1164 2116 1172 2124
rect 972 2096 980 2104
rect 876 2056 884 2064
rect 924 2056 932 2064
rect 956 2056 964 2064
rect 892 1716 900 1724
rect 972 2036 980 2044
rect 1036 2056 1044 2064
rect 1004 1996 1012 2004
rect 972 1916 980 1924
rect 988 1896 996 1904
rect 940 1856 948 1864
rect 988 1856 996 1864
rect 1020 1856 1028 1864
rect 956 1836 964 1844
rect 972 1816 980 1824
rect 1052 1916 1060 1924
rect 1132 1916 1140 1924
rect 1116 1876 1124 1884
rect 1036 1816 1044 1824
rect 988 1756 996 1764
rect 1004 1736 1012 1744
rect 1068 1736 1076 1744
rect 972 1716 980 1724
rect 908 1696 916 1704
rect 892 1676 900 1684
rect 860 1636 868 1644
rect 812 1496 820 1504
rect 716 1476 724 1484
rect 524 1396 532 1404
rect 572 1376 580 1384
rect 652 1356 660 1364
rect 604 1336 612 1344
rect 748 1396 756 1404
rect 748 1356 756 1364
rect 684 1336 692 1344
rect 700 1336 708 1344
rect 956 1656 964 1664
rect 1036 1696 1044 1704
rect 1260 2118 1268 2124
rect 1260 2116 1268 2118
rect 1180 1856 1188 1864
rect 1324 2036 1332 2044
rect 1276 1956 1284 1964
rect 1260 1896 1268 1904
rect 1212 1836 1220 1844
rect 1244 1836 1252 1844
rect 1196 1816 1204 1824
rect 1068 1676 1076 1684
rect 1084 1676 1092 1684
rect 1116 1696 1124 1704
rect 1052 1656 1060 1664
rect 1100 1656 1108 1664
rect 1020 1636 1028 1644
rect 1004 1556 1012 1564
rect 1004 1516 1012 1524
rect 1068 1616 1076 1624
rect 1020 1496 1028 1504
rect 1036 1496 1044 1504
rect 1148 1676 1156 1684
rect 1148 1656 1156 1664
rect 1420 2256 1428 2264
rect 1404 2196 1412 2204
rect 1388 2176 1396 2184
rect 1404 2156 1412 2164
rect 1372 2016 1380 2024
rect 1292 1916 1300 1924
rect 1388 1916 1396 1924
rect 1340 1896 1348 1904
rect 1372 1876 1380 1884
rect 1228 1756 1236 1764
rect 1260 1736 1268 1744
rect 1228 1676 1236 1684
rect 1244 1676 1252 1684
rect 1212 1616 1220 1624
rect 1180 1596 1188 1604
rect 1132 1576 1140 1584
rect 1116 1556 1124 1564
rect 1116 1516 1124 1524
rect 1356 1836 1364 1844
rect 1388 1816 1396 1824
rect 1356 1796 1364 1804
rect 1388 1756 1396 1764
rect 1324 1736 1332 1744
rect 1484 2236 1492 2244
rect 1484 2216 1492 2224
rect 1468 2176 1476 2184
rect 1436 2156 1444 2164
rect 1420 1896 1428 1904
rect 1548 2396 1556 2404
rect 1564 2376 1572 2384
rect 1564 2336 1572 2344
rect 1532 2196 1540 2204
rect 1532 2136 1540 2144
rect 1500 2096 1508 2104
rect 1564 2216 1572 2224
rect 1548 2056 1556 2064
rect 1452 2036 1460 2044
rect 1516 1996 1524 2004
rect 1468 1956 1476 1964
rect 1484 1936 1492 1944
rect 1452 1916 1460 1924
rect 1468 1896 1476 1904
rect 1420 1796 1428 1804
rect 1676 2636 1684 2644
rect 1660 2616 1668 2624
rect 1660 2576 1668 2584
rect 1644 2536 1652 2544
rect 1628 2396 1636 2404
rect 1628 2316 1636 2324
rect 1660 2316 1668 2324
rect 1724 2536 1732 2544
rect 1708 2376 1716 2384
rect 1996 3216 2004 3224
rect 2140 3436 2148 3444
rect 2060 3416 2068 3424
rect 2028 3316 2036 3324
rect 2044 3316 2052 3324
rect 2044 3256 2052 3264
rect 2220 3496 2228 3504
rect 2188 3476 2196 3484
rect 2156 3316 2164 3324
rect 2060 3216 2068 3224
rect 2108 3176 2116 3184
rect 2044 3136 2052 3144
rect 2076 3136 2084 3144
rect 1996 3096 2004 3104
rect 1932 3016 1940 3024
rect 1900 2936 1908 2944
rect 2060 3036 2068 3044
rect 2060 3016 2068 3024
rect 2252 3436 2260 3444
rect 2243 3406 2251 3414
rect 2253 3406 2261 3414
rect 2263 3406 2271 3414
rect 2273 3406 2281 3414
rect 2283 3406 2291 3414
rect 2293 3406 2301 3414
rect 2220 3336 2228 3344
rect 2508 4476 2516 4484
rect 2508 4436 2516 4444
rect 2524 4416 2532 4424
rect 2396 4336 2404 4344
rect 2460 4336 2468 4344
rect 2428 4296 2436 4304
rect 2364 4276 2372 4284
rect 2508 4296 2516 4304
rect 2412 4276 2420 4284
rect 2476 4276 2484 4284
rect 2428 4256 2436 4264
rect 2460 4256 2468 4264
rect 2524 4256 2532 4264
rect 2492 4216 2500 4224
rect 2444 4176 2452 4184
rect 2476 4176 2484 4184
rect 2572 4496 2580 4504
rect 2620 4416 2628 4424
rect 2556 4296 2564 4304
rect 2572 4276 2580 4284
rect 2588 4256 2596 4264
rect 2572 4196 2580 4204
rect 2588 4176 2596 4184
rect 2540 4156 2548 4164
rect 2572 4156 2580 4164
rect 2348 4116 2356 4124
rect 2396 4116 2404 4124
rect 2332 3976 2340 3984
rect 2460 4096 2468 4104
rect 2508 4096 2516 4104
rect 2556 4096 2564 4104
rect 2428 4076 2436 4084
rect 2396 3956 2404 3964
rect 2396 3936 2404 3944
rect 2364 3916 2372 3924
rect 2364 3856 2372 3864
rect 2332 3816 2340 3824
rect 2348 3756 2356 3764
rect 2380 3756 2388 3764
rect 2364 3716 2372 3724
rect 2348 3596 2356 3604
rect 2332 3456 2340 3464
rect 2220 3276 2228 3284
rect 2204 3156 2212 3164
rect 2108 3116 2116 3124
rect 2172 3116 2180 3124
rect 2092 2976 2100 2984
rect 1980 2936 1988 2944
rect 1996 2936 2004 2944
rect 2060 2936 2068 2944
rect 1948 2916 1956 2924
rect 1964 2916 1972 2924
rect 1884 2856 1892 2864
rect 1836 2836 1844 2844
rect 1884 2796 1892 2804
rect 1868 2776 1876 2784
rect 1916 2736 1924 2744
rect 1980 2896 1988 2904
rect 1964 2816 1972 2824
rect 1948 2716 1956 2724
rect 1820 2676 1828 2684
rect 1852 2676 1860 2684
rect 1900 2676 1908 2684
rect 1932 2676 1940 2684
rect 1836 2596 1844 2604
rect 1900 2636 1908 2644
rect 1852 2576 1860 2584
rect 1916 2576 1924 2584
rect 1964 2556 1972 2564
rect 1820 2536 1828 2544
rect 1852 2536 1860 2544
rect 1788 2476 1796 2484
rect 1852 2516 1860 2524
rect 1772 2376 1780 2384
rect 1740 2316 1748 2324
rect 1756 2296 1764 2304
rect 1772 2296 1780 2304
rect 1692 2276 1700 2284
rect 1708 2276 1716 2284
rect 1612 2196 1620 2204
rect 1628 2196 1636 2204
rect 1596 2176 1604 2184
rect 1580 2016 1588 2024
rect 1740 2256 1748 2264
rect 1724 2236 1732 2244
rect 1740 2236 1748 2244
rect 1708 2216 1716 2224
rect 1724 2176 1732 2184
rect 1708 2156 1716 2164
rect 1692 2136 1700 2144
rect 1692 2096 1700 2104
rect 1740 2116 1748 2124
rect 1756 2116 1764 2124
rect 1724 2096 1732 2104
rect 1740 2096 1748 2104
rect 1724 2076 1732 2084
rect 1580 1996 1588 2004
rect 1628 1996 1636 2004
rect 1564 1916 1572 1924
rect 1660 1956 1668 1964
rect 1580 1896 1588 1904
rect 1516 1856 1524 1864
rect 1468 1756 1476 1764
rect 1484 1756 1492 1764
rect 1340 1696 1348 1704
rect 1356 1636 1364 1644
rect 1308 1576 1316 1584
rect 1308 1536 1316 1544
rect 1260 1516 1268 1524
rect 1276 1516 1284 1524
rect 1132 1496 1140 1504
rect 1148 1496 1156 1504
rect 1084 1476 1092 1484
rect 1036 1436 1044 1444
rect 1068 1436 1076 1444
rect 1084 1436 1092 1444
rect 988 1416 996 1424
rect 908 1376 916 1384
rect 892 1336 900 1344
rect 508 1316 516 1324
rect 636 1276 644 1284
rect 716 1296 724 1304
rect 739 1206 747 1214
rect 749 1206 757 1214
rect 759 1206 767 1214
rect 769 1206 777 1214
rect 779 1206 787 1214
rect 789 1206 797 1214
rect 460 1016 468 1024
rect 396 996 404 1004
rect 380 976 388 984
rect 444 976 452 984
rect 396 956 404 964
rect 412 956 420 964
rect 268 916 276 924
rect 348 916 356 924
rect 380 916 388 924
rect 268 876 276 884
rect 348 876 356 884
rect 236 816 244 824
rect 156 776 164 784
rect 316 816 324 824
rect 140 702 148 704
rect 140 696 148 702
rect 252 696 260 704
rect 76 596 84 604
rect 220 676 228 684
rect 252 656 260 664
rect 364 696 372 704
rect 428 936 436 944
rect 428 916 436 924
rect 476 956 484 964
rect 508 956 516 964
rect 476 916 484 924
rect 460 856 468 864
rect 412 816 420 824
rect 412 796 420 804
rect 428 716 436 724
rect 412 696 420 704
rect 348 676 356 684
rect 316 656 324 664
rect 204 636 212 644
rect 268 636 276 644
rect 300 636 308 644
rect 236 596 244 604
rect 284 596 292 604
rect 188 576 196 584
rect 124 536 132 544
rect 220 536 228 544
rect 108 356 116 364
rect 60 176 68 184
rect 188 356 196 364
rect 188 316 196 324
rect 140 216 148 224
rect 124 176 132 184
rect 28 136 36 144
rect 156 136 164 144
rect 12 116 20 124
rect 76 116 84 124
rect 332 596 340 604
rect 300 576 308 584
rect 396 676 404 684
rect 380 596 388 604
rect 396 576 404 584
rect 780 1136 788 1144
rect 636 1116 644 1124
rect 700 1116 708 1124
rect 684 1096 692 1104
rect 588 1056 596 1064
rect 620 956 628 964
rect 1020 1396 1028 1404
rect 1068 1376 1076 1384
rect 1052 1336 1060 1344
rect 1180 1476 1188 1484
rect 1148 1396 1156 1404
rect 1100 1336 1108 1344
rect 1148 1336 1156 1344
rect 1212 1456 1220 1464
rect 1260 1376 1268 1384
rect 1244 1356 1252 1364
rect 1164 1276 1172 1284
rect 1196 1276 1204 1284
rect 1180 1256 1188 1264
rect 1196 1236 1204 1244
rect 1244 1296 1252 1304
rect 1260 1296 1268 1304
rect 1276 1276 1284 1284
rect 1292 1256 1300 1264
rect 1372 1516 1380 1524
rect 1340 1496 1348 1504
rect 1324 1416 1332 1424
rect 1340 1396 1348 1404
rect 1324 1356 1332 1364
rect 1356 1336 1364 1344
rect 1452 1736 1460 1744
rect 1500 1736 1508 1744
rect 1404 1676 1412 1684
rect 1404 1656 1412 1664
rect 1468 1656 1476 1664
rect 1500 1616 1508 1624
rect 1436 1496 1444 1504
rect 1596 1876 1604 1884
rect 1676 1876 1684 1884
rect 1548 1796 1556 1804
rect 1564 1796 1572 1804
rect 1676 1816 1684 1824
rect 1644 1796 1652 1804
rect 1580 1756 1588 1764
rect 1628 1756 1636 1764
rect 1644 1736 1652 1744
rect 1612 1716 1620 1724
rect 1548 1696 1556 1704
rect 1612 1696 1620 1704
rect 1532 1676 1540 1684
rect 1516 1576 1524 1584
rect 1532 1556 1540 1564
rect 1516 1496 1524 1504
rect 1452 1476 1460 1484
rect 1484 1456 1492 1464
rect 1564 1476 1572 1484
rect 1548 1456 1556 1464
rect 1548 1436 1556 1444
rect 1644 1636 1652 1644
rect 1596 1456 1604 1464
rect 1420 1376 1428 1384
rect 1452 1376 1460 1384
rect 1532 1376 1540 1384
rect 1356 1296 1364 1304
rect 1324 1256 1332 1264
rect 1308 1216 1316 1224
rect 1340 1216 1348 1224
rect 1164 1176 1172 1184
rect 1212 1176 1220 1184
rect 1004 1116 1012 1124
rect 1052 1116 1060 1124
rect 1084 1116 1092 1124
rect 1100 1116 1108 1124
rect 972 1096 980 1104
rect 860 1076 868 1084
rect 812 1016 820 1024
rect 652 956 660 964
rect 604 936 612 944
rect 604 916 612 924
rect 540 876 548 884
rect 684 716 692 724
rect 476 636 484 644
rect 508 636 516 644
rect 460 596 468 604
rect 460 536 468 544
rect 668 656 676 664
rect 652 576 660 584
rect 860 1016 868 1024
rect 748 916 756 924
rect 812 918 820 924
rect 812 916 820 918
rect 739 806 747 814
rect 749 806 757 814
rect 759 806 767 814
rect 769 806 777 814
rect 779 806 787 814
rect 789 806 797 814
rect 1212 1116 1220 1124
rect 1116 1096 1124 1104
rect 988 1076 996 1084
rect 1100 1076 1108 1084
rect 1164 1076 1172 1084
rect 908 996 916 1004
rect 1116 996 1124 1004
rect 940 976 948 984
rect 956 976 964 984
rect 1148 936 1156 944
rect 1084 918 1092 924
rect 1084 916 1092 918
rect 1116 776 1124 784
rect 860 736 868 744
rect 828 716 836 724
rect 1052 716 1060 724
rect 1212 1016 1220 1024
rect 1196 956 1204 964
rect 1180 936 1188 944
rect 1180 916 1188 924
rect 1180 896 1188 904
rect 1244 996 1252 1004
rect 1356 996 1364 1004
rect 1260 956 1268 964
rect 1516 1356 1524 1364
rect 1404 1276 1412 1284
rect 1452 1296 1460 1304
rect 1580 1396 1588 1404
rect 1596 1396 1604 1404
rect 1580 1376 1588 1384
rect 1564 1356 1572 1364
rect 1628 1416 1636 1424
rect 1436 1076 1444 1084
rect 1404 1036 1412 1044
rect 1388 976 1396 984
rect 1516 1296 1524 1304
rect 1564 1296 1572 1304
rect 1612 1236 1620 1244
rect 1532 1216 1540 1224
rect 1516 1116 1524 1124
rect 1516 1076 1524 1084
rect 1452 996 1460 1004
rect 1516 996 1524 1004
rect 1420 956 1428 964
rect 1708 1876 1716 1884
rect 1692 1776 1700 1784
rect 1692 1756 1700 1764
rect 1708 1736 1716 1744
rect 1724 1656 1732 1664
rect 1868 2496 1876 2504
rect 1948 2496 1956 2504
rect 1996 2856 2004 2864
rect 2076 2876 2084 2884
rect 2028 2836 2036 2844
rect 2060 2836 2068 2844
rect 2012 2736 2020 2744
rect 2060 2736 2068 2744
rect 2012 2616 2020 2624
rect 1868 2476 1876 2484
rect 1916 2476 1924 2484
rect 1948 2416 1956 2424
rect 1852 2296 1860 2304
rect 1820 2276 1828 2284
rect 1884 2276 1892 2284
rect 1836 2216 1844 2224
rect 1836 2196 1844 2204
rect 1804 2096 1812 2104
rect 1932 2236 1940 2244
rect 1900 2136 1908 2144
rect 1884 2096 1892 2104
rect 1932 2076 1940 2084
rect 1852 2056 1860 2064
rect 1820 2036 1828 2044
rect 1772 1996 1780 2004
rect 1836 1976 1844 1984
rect 1820 1876 1828 1884
rect 1804 1816 1812 1824
rect 1868 1916 1876 1924
rect 1916 1916 1924 1924
rect 1868 1896 1876 1904
rect 1900 1896 1908 1904
rect 1932 1876 1940 1884
rect 1916 1796 1924 1804
rect 1900 1776 1908 1784
rect 1852 1756 1860 1764
rect 1932 1756 1940 1764
rect 1788 1716 1796 1724
rect 1804 1676 1812 1684
rect 1868 1676 1876 1684
rect 1772 1656 1780 1664
rect 1756 1636 1764 1644
rect 1740 1576 1748 1584
rect 1836 1656 1844 1664
rect 1820 1596 1828 1604
rect 1836 1596 1844 1604
rect 1932 1596 1940 1604
rect 1964 2396 1972 2404
rect 1964 2316 1972 2324
rect 2012 2496 2020 2504
rect 2044 2656 2052 2664
rect 2044 2636 2052 2644
rect 2076 2716 2084 2724
rect 2172 3056 2180 3064
rect 2188 3056 2196 3064
rect 2140 3036 2148 3044
rect 2156 3016 2164 3024
rect 2124 2956 2132 2964
rect 2156 2956 2164 2964
rect 2124 2936 2132 2944
rect 2124 2876 2132 2884
rect 2316 3196 2324 3204
rect 2364 3536 2372 3544
rect 2412 3716 2420 3724
rect 2396 3696 2404 3704
rect 2508 4076 2516 4084
rect 2556 4076 2564 4084
rect 2508 3916 2516 3924
rect 2460 3896 2468 3904
rect 2764 4936 2772 4944
rect 2780 4936 2788 4944
rect 2700 4796 2708 4804
rect 2972 5016 2980 5024
rect 3084 5076 3092 5084
rect 3356 5076 3364 5084
rect 3436 5076 3444 5084
rect 3452 5076 3460 5084
rect 3660 5076 3668 5084
rect 2892 4976 2900 4984
rect 3004 4976 3012 4984
rect 3036 4956 3044 4964
rect 2940 4936 2948 4944
rect 2892 4916 2900 4924
rect 2972 4916 2980 4924
rect 2684 4736 2692 4744
rect 2908 4796 2916 4804
rect 3020 4796 3028 4804
rect 2956 4756 2964 4764
rect 3148 5036 3156 5044
rect 3244 5036 3252 5044
rect 3340 5036 3348 5044
rect 3116 4976 3124 4984
rect 3148 4976 3156 4984
rect 3084 4956 3092 4964
rect 3196 4936 3204 4944
rect 3340 4976 3348 4984
rect 3292 4936 3300 4944
rect 3388 5056 3396 5064
rect 3468 5056 3476 5064
rect 3356 4956 3364 4964
rect 3420 4976 3428 4984
rect 3548 4996 3556 5004
rect 3596 4996 3604 5004
rect 3516 4936 3524 4944
rect 3628 4936 3636 4944
rect 3228 4916 3236 4924
rect 3500 4916 3508 4924
rect 3580 4916 3588 4924
rect 3132 4876 3140 4884
rect 3228 4876 3236 4884
rect 3164 4736 3172 4744
rect 2716 4676 2724 4684
rect 2684 4656 2692 4664
rect 2700 4656 2708 4664
rect 2668 4576 2676 4584
rect 2668 4556 2676 4564
rect 2860 4656 2868 4664
rect 2892 4636 2900 4644
rect 2940 4636 2948 4644
rect 2716 4556 2724 4564
rect 2732 4536 2740 4544
rect 2652 4416 2660 4424
rect 2684 4516 2692 4524
rect 2764 4516 2772 4524
rect 2844 4516 2852 4524
rect 3052 4536 3060 4544
rect 2716 4496 2724 4504
rect 2780 4496 2788 4504
rect 2796 4496 2804 4504
rect 2700 4456 2708 4464
rect 2764 4336 2772 4344
rect 2828 4456 2836 4464
rect 2828 4356 2836 4364
rect 2684 4316 2692 4324
rect 3164 4676 3172 4684
rect 3148 4656 3156 4664
rect 3196 4656 3204 4664
rect 3212 4576 3220 4584
rect 2924 4496 2932 4504
rect 3052 4496 3060 4504
rect 3116 4496 3124 4504
rect 2924 4456 2932 4464
rect 2748 4296 2756 4304
rect 2812 4296 2820 4304
rect 2844 4296 2852 4304
rect 2876 4296 2884 4304
rect 2636 4276 2644 4284
rect 2668 4276 2676 4284
rect 2668 3956 2676 3964
rect 2604 3936 2612 3944
rect 2668 3936 2676 3944
rect 2620 3916 2628 3924
rect 2556 3856 2564 3864
rect 2444 3776 2452 3784
rect 2476 3736 2484 3744
rect 2508 3696 2516 3704
rect 2428 3676 2436 3684
rect 2636 3896 2644 3904
rect 2652 3896 2660 3904
rect 2636 3776 2644 3784
rect 2620 3716 2628 3724
rect 2572 3656 2580 3664
rect 2620 3596 2628 3604
rect 2428 3536 2436 3544
rect 2444 3536 2452 3544
rect 2476 3536 2484 3544
rect 2380 3516 2388 3524
rect 2444 3496 2452 3504
rect 2364 3476 2372 3484
rect 2348 3436 2356 3444
rect 2348 3356 2356 3364
rect 2380 3416 2388 3424
rect 2540 3502 2548 3504
rect 2540 3496 2548 3502
rect 2636 3456 2644 3464
rect 2396 3376 2404 3384
rect 2380 3356 2388 3364
rect 2348 3316 2356 3324
rect 2508 3376 2516 3384
rect 2492 3336 2500 3344
rect 2796 4276 2804 4284
rect 2844 4276 2852 4284
rect 2732 4256 2740 4264
rect 2812 4256 2820 4264
rect 2892 4276 2900 4284
rect 2796 4196 2804 4204
rect 2828 4196 2836 4204
rect 2988 4416 2996 4424
rect 3020 4296 3028 4304
rect 2748 4136 2756 4144
rect 2908 4136 2916 4144
rect 2780 4116 2788 4124
rect 2700 4076 2708 4084
rect 2716 3916 2724 3924
rect 2684 3896 2692 3904
rect 2748 3896 2756 3904
rect 2700 3876 2708 3884
rect 2668 3536 2676 3544
rect 2716 3796 2724 3804
rect 2748 3776 2756 3784
rect 2732 3716 2740 3724
rect 2684 3516 2692 3524
rect 2748 3516 2756 3524
rect 2732 3496 2740 3504
rect 2812 3976 2820 3984
rect 2780 3916 2788 3924
rect 2780 3856 2788 3864
rect 2780 3816 2788 3824
rect 2956 4276 2964 4284
rect 3004 4256 3012 4264
rect 3036 4276 3044 4284
rect 3116 4436 3124 4444
rect 3132 4436 3140 4444
rect 3084 4336 3092 4344
rect 3180 4496 3188 4504
rect 3228 4516 3236 4524
rect 3404 4876 3412 4884
rect 3308 4836 3316 4844
rect 3260 4616 3268 4624
rect 3196 4416 3204 4424
rect 3148 4356 3156 4364
rect 3196 4356 3204 4364
rect 3180 4336 3188 4344
rect 3260 4456 3268 4464
rect 3260 4416 3268 4424
rect 3228 4316 3236 4324
rect 3052 4236 3060 4244
rect 3148 4256 3156 4264
rect 3196 4256 3204 4264
rect 3116 4216 3124 4224
rect 3084 4196 3092 4204
rect 3020 4176 3028 4184
rect 3020 4156 3028 4164
rect 3020 4116 3028 4124
rect 2956 4096 2964 4104
rect 2988 3976 2996 3984
rect 2940 3936 2948 3944
rect 2972 3936 2980 3944
rect 2844 3902 2852 3904
rect 2844 3896 2852 3902
rect 2908 3896 2916 3904
rect 2988 3876 2996 3884
rect 2844 3836 2852 3844
rect 2700 3476 2708 3484
rect 2764 3476 2772 3484
rect 2684 3396 2692 3404
rect 2572 3316 2580 3324
rect 2380 3296 2388 3304
rect 2364 3196 2372 3204
rect 2380 3156 2388 3164
rect 2236 3116 2244 3124
rect 2252 3096 2260 3104
rect 2243 3006 2251 3014
rect 2253 3006 2261 3014
rect 2263 3006 2271 3014
rect 2273 3006 2281 3014
rect 2283 3006 2291 3014
rect 2293 3006 2301 3014
rect 2444 3116 2452 3124
rect 2476 3116 2484 3124
rect 2620 3296 2628 3304
rect 2604 3276 2612 3284
rect 2540 3136 2548 3144
rect 2572 3136 2580 3144
rect 2380 2976 2388 2984
rect 2268 2876 2276 2884
rect 2172 2856 2180 2864
rect 2220 2856 2228 2864
rect 2172 2836 2180 2844
rect 2156 2756 2164 2764
rect 2140 2696 2148 2704
rect 2108 2676 2116 2684
rect 2124 2676 2132 2684
rect 2076 2616 2084 2624
rect 2060 2596 2068 2604
rect 2092 2496 2100 2504
rect 2028 2376 2036 2384
rect 2012 2316 2020 2324
rect 1964 2256 1972 2264
rect 2076 2256 2084 2264
rect 1980 2196 1988 2204
rect 1980 2116 1988 2124
rect 1996 2116 2004 2124
rect 2012 2116 2020 2124
rect 2012 2076 2020 2084
rect 2028 2036 2036 2044
rect 2028 1976 2036 1984
rect 1964 1896 1972 1904
rect 1964 1876 1972 1884
rect 1996 1856 2004 1864
rect 2060 1916 2068 1924
rect 2060 1816 2068 1824
rect 1980 1756 1988 1764
rect 2044 1756 2052 1764
rect 2060 1736 2068 1744
rect 2044 1716 2052 1724
rect 2092 2236 2100 2244
rect 2204 2796 2212 2804
rect 2300 2736 2308 2744
rect 2220 2696 2228 2704
rect 2172 2576 2180 2584
rect 2140 2536 2148 2544
rect 2140 2496 2148 2504
rect 2156 2456 2164 2464
rect 2243 2606 2251 2614
rect 2253 2606 2261 2614
rect 2263 2606 2271 2614
rect 2273 2606 2281 2614
rect 2283 2606 2291 2614
rect 2293 2606 2301 2614
rect 2348 2916 2356 2924
rect 2364 2856 2372 2864
rect 2204 2556 2212 2564
rect 2332 2556 2340 2564
rect 2300 2496 2308 2504
rect 2316 2496 2324 2504
rect 2188 2396 2196 2404
rect 2124 2336 2132 2344
rect 2188 2336 2196 2344
rect 2172 2316 2180 2324
rect 2156 2296 2164 2304
rect 2252 2296 2260 2304
rect 2268 2256 2276 2264
rect 2204 2236 2212 2244
rect 2220 2216 2228 2224
rect 2243 2206 2251 2214
rect 2253 2206 2261 2214
rect 2263 2206 2271 2214
rect 2273 2206 2281 2214
rect 2283 2206 2291 2214
rect 2293 2206 2301 2214
rect 2188 2196 2196 2204
rect 2508 3056 2516 3064
rect 2460 2936 2468 2944
rect 2492 2936 2500 2944
rect 2428 2916 2436 2924
rect 2476 2916 2484 2924
rect 2412 2676 2420 2684
rect 2540 3036 2548 3044
rect 2540 2956 2548 2964
rect 2604 2956 2612 2964
rect 2636 3256 2644 3264
rect 2652 3196 2660 3204
rect 2636 3176 2644 3184
rect 2652 3176 2660 3184
rect 2652 3136 2660 3144
rect 2668 3116 2676 3124
rect 2652 3036 2660 3044
rect 2636 3016 2644 3024
rect 2636 2996 2644 3004
rect 2572 2916 2580 2924
rect 2620 2896 2628 2904
rect 2556 2876 2564 2884
rect 2588 2836 2596 2844
rect 2524 2776 2532 2784
rect 2540 2702 2548 2704
rect 2540 2696 2548 2702
rect 2508 2676 2516 2684
rect 2428 2656 2436 2664
rect 2572 2596 2580 2604
rect 2380 2496 2388 2504
rect 2396 2376 2404 2384
rect 2380 2316 2388 2324
rect 2428 2316 2436 2324
rect 2588 2516 2596 2524
rect 2492 2496 2500 2504
rect 2492 2456 2500 2464
rect 2460 2376 2468 2384
rect 2476 2316 2484 2324
rect 2668 2996 2676 3004
rect 2668 2956 2676 2964
rect 2652 2936 2660 2944
rect 2748 3456 2756 3464
rect 2812 3796 2820 3804
rect 3036 4096 3044 4104
rect 3244 4116 3252 4124
rect 3148 4096 3156 4104
rect 3132 3996 3140 4004
rect 3052 3976 3060 3984
rect 3196 3976 3204 3984
rect 3036 3956 3044 3964
rect 3180 3936 3188 3944
rect 3244 3936 3252 3944
rect 3036 3916 3044 3924
rect 3116 3896 3124 3904
rect 3244 3916 3252 3924
rect 3292 4736 3300 4744
rect 3324 4716 3332 4724
rect 3356 4716 3364 4724
rect 3388 4716 3396 4724
rect 3324 4656 3332 4664
rect 3372 4656 3380 4664
rect 3452 4836 3460 4844
rect 3564 4836 3572 4844
rect 3516 4776 3524 4784
rect 3452 4716 3460 4724
rect 3500 4716 3508 4724
rect 3436 4696 3444 4704
rect 3340 4616 3348 4624
rect 3388 4616 3396 4624
rect 3404 4616 3412 4624
rect 3356 4536 3364 4544
rect 3292 4496 3300 4504
rect 3340 4456 3348 4464
rect 3628 4876 3636 4884
rect 3612 4796 3620 4804
rect 3644 4776 3652 4784
rect 3580 4736 3588 4744
rect 3468 4676 3476 4684
rect 3548 4676 3556 4684
rect 3596 4676 3604 4684
rect 3676 4996 3684 5004
rect 3724 4996 3732 5004
rect 3756 4976 3764 4984
rect 3788 4956 3796 4964
rect 3724 4936 3732 4944
rect 4764 5216 4772 5224
rect 6755 5206 6763 5214
rect 6765 5206 6773 5214
rect 6775 5206 6783 5214
rect 6785 5206 6793 5214
rect 6795 5206 6803 5214
rect 6805 5206 6813 5214
rect 4204 5156 4212 5164
rect 6028 5156 6036 5164
rect 6156 5156 6164 5164
rect 4444 5136 4452 5144
rect 4636 5136 4644 5144
rect 4924 5136 4932 5144
rect 4956 5136 4964 5144
rect 5436 5136 5444 5144
rect 5532 5136 5540 5144
rect 5548 5136 5556 5144
rect 5724 5136 5732 5144
rect 5900 5136 5908 5144
rect 4732 5116 4740 5124
rect 4780 5116 4788 5124
rect 4796 5116 4804 5124
rect 4828 5116 4836 5124
rect 4876 5116 4884 5124
rect 4972 5116 4980 5124
rect 5036 5116 5044 5124
rect 5068 5116 5076 5124
rect 3948 5096 3956 5104
rect 4076 5102 4084 5104
rect 4076 5096 4084 5102
rect 4092 5056 4100 5064
rect 3900 4956 3908 4964
rect 3964 4956 3972 4964
rect 4492 5096 4500 5104
rect 4604 5096 4612 5104
rect 4252 5076 4260 5084
rect 4172 4976 4180 4984
rect 4060 4936 4068 4944
rect 4140 4936 4148 4944
rect 3740 4916 3748 4924
rect 3948 4916 3956 4924
rect 4028 4916 4036 4924
rect 3836 4896 3844 4904
rect 3724 4816 3732 4824
rect 3747 4806 3755 4814
rect 3757 4806 3765 4814
rect 3767 4806 3775 4814
rect 3777 4806 3785 4814
rect 3787 4806 3795 4814
rect 3797 4806 3805 4814
rect 3836 4776 3844 4784
rect 3708 4756 3716 4764
rect 3692 4736 3700 4744
rect 3820 4736 3828 4744
rect 3724 4696 3732 4704
rect 3916 4896 3924 4904
rect 3996 4896 4004 4904
rect 4076 4916 4084 4924
rect 4172 4916 4180 4924
rect 4044 4876 4052 4884
rect 3932 4856 3940 4864
rect 3996 4856 4004 4864
rect 3948 4716 3956 4724
rect 3676 4676 3684 4684
rect 3772 4676 3780 4684
rect 3596 4656 3604 4664
rect 3660 4656 3668 4664
rect 3500 4636 3508 4644
rect 3580 4636 3588 4644
rect 3468 4616 3476 4624
rect 3452 4596 3460 4604
rect 3436 4536 3444 4544
rect 3404 4516 3412 4524
rect 3436 4516 3444 4524
rect 3388 4496 3396 4504
rect 3420 4496 3428 4504
rect 3372 4436 3380 4444
rect 3324 4416 3332 4424
rect 3404 4356 3412 4364
rect 3276 4176 3284 4184
rect 3276 4156 3284 4164
rect 3388 4276 3396 4284
rect 3420 4276 3428 4284
rect 3404 4196 3412 4204
rect 3324 4136 3332 4144
rect 3292 4116 3300 4124
rect 3148 3876 3156 3884
rect 3212 3876 3220 3884
rect 3036 3856 3044 3864
rect 3020 3816 3028 3824
rect 2876 3776 2884 3784
rect 3132 3776 3140 3784
rect 2940 3756 2948 3764
rect 3260 3816 3268 3824
rect 3212 3776 3220 3784
rect 2972 3736 2980 3744
rect 3212 3736 3220 3744
rect 3260 3736 3268 3744
rect 2892 3716 2900 3724
rect 2908 3716 2916 3724
rect 2844 3696 2852 3704
rect 2876 3576 2884 3584
rect 2796 3536 2804 3544
rect 2860 3516 2868 3524
rect 2860 3496 2868 3504
rect 2796 3476 2804 3484
rect 2748 3416 2756 3424
rect 2732 3396 2740 3404
rect 2732 3376 2740 3384
rect 2732 3296 2740 3304
rect 2812 3456 2820 3464
rect 2860 3476 2868 3484
rect 2844 3436 2852 3444
rect 2828 3336 2836 3344
rect 2796 3316 2804 3324
rect 2860 3318 2868 3324
rect 2860 3316 2868 3318
rect 2796 3296 2804 3304
rect 2860 3296 2868 3304
rect 2764 3196 2772 3204
rect 2780 3156 2788 3164
rect 2748 3136 2756 3144
rect 2764 3116 2772 3124
rect 2716 3096 2724 3104
rect 2780 3096 2788 3104
rect 2732 3076 2740 3084
rect 2796 3076 2804 3084
rect 2796 3056 2804 3064
rect 2700 2976 2708 2984
rect 2796 2956 2804 2964
rect 2684 2936 2692 2944
rect 2700 2936 2708 2944
rect 2732 2916 2740 2924
rect 2716 2896 2724 2904
rect 2700 2876 2708 2884
rect 2844 2976 2852 2984
rect 2844 2956 2852 2964
rect 2924 3696 2932 3704
rect 2908 3556 2916 3564
rect 3004 3718 3012 3724
rect 3004 3716 3012 3718
rect 3164 3716 3172 3724
rect 3196 3716 3204 3724
rect 3148 3696 3156 3704
rect 2956 3576 2964 3584
rect 3052 3556 3060 3564
rect 2988 3536 2996 3544
rect 2972 3496 2980 3504
rect 3180 3636 3188 3644
rect 3100 3536 3108 3544
rect 3100 3496 3108 3504
rect 2956 3476 2964 3484
rect 3020 3476 3028 3484
rect 3036 3476 3044 3484
rect 2924 3456 2932 3464
rect 2940 3456 2948 3464
rect 2892 3376 2900 3384
rect 2940 3196 2948 3204
rect 3084 3476 3092 3484
rect 3004 3316 3012 3324
rect 2972 3176 2980 3184
rect 2956 3136 2964 3144
rect 2988 3116 2996 3124
rect 2940 3096 2948 3104
rect 2860 2936 2868 2944
rect 2796 2896 2804 2904
rect 2828 2896 2836 2904
rect 2764 2876 2772 2884
rect 2764 2856 2772 2864
rect 2716 2716 2724 2724
rect 2684 2696 2692 2704
rect 2780 2696 2788 2704
rect 2684 2636 2692 2644
rect 2652 2616 2660 2624
rect 2652 2556 2660 2564
rect 2684 2536 2692 2544
rect 2716 2516 2724 2524
rect 2636 2496 2644 2504
rect 2700 2496 2708 2504
rect 2620 2436 2628 2444
rect 2524 2416 2532 2424
rect 2508 2376 2516 2384
rect 2460 2276 2468 2284
rect 2108 2136 2116 2144
rect 2380 2156 2388 2164
rect 2332 2136 2340 2144
rect 2124 2116 2132 2124
rect 2172 2056 2180 2064
rect 2156 1816 2164 1824
rect 2092 1736 2100 1744
rect 1964 1696 1972 1704
rect 1964 1616 1972 1624
rect 1868 1576 1876 1584
rect 1916 1576 1924 1584
rect 1948 1576 1956 1584
rect 1756 1496 1764 1504
rect 1788 1496 1796 1504
rect 1804 1496 1812 1504
rect 1884 1496 1892 1504
rect 1660 1436 1668 1444
rect 1660 1296 1668 1304
rect 1644 1276 1652 1284
rect 1756 1456 1764 1464
rect 1788 1456 1796 1464
rect 1724 1396 1732 1404
rect 1692 1376 1700 1384
rect 1756 1376 1764 1384
rect 1708 1356 1716 1364
rect 1740 1356 1748 1364
rect 1756 1336 1764 1344
rect 1788 1356 1796 1364
rect 1916 1476 1924 1484
rect 1804 1336 1812 1344
rect 1692 1296 1700 1304
rect 1756 1296 1764 1304
rect 1692 1276 1700 1284
rect 1676 1216 1684 1224
rect 1644 1116 1652 1124
rect 1548 1096 1556 1104
rect 1596 1096 1604 1104
rect 1580 976 1588 984
rect 1612 956 1620 964
rect 1228 936 1236 944
rect 1292 936 1300 944
rect 1308 936 1316 944
rect 1372 936 1380 944
rect 1468 936 1476 944
rect 1244 916 1252 924
rect 1324 916 1332 924
rect 1436 916 1444 924
rect 1212 896 1220 904
rect 1324 896 1332 904
rect 1372 896 1380 904
rect 1228 876 1236 884
rect 1260 816 1268 824
rect 1484 916 1492 924
rect 1468 876 1476 884
rect 1484 876 1492 884
rect 1532 876 1540 884
rect 1580 876 1588 884
rect 1596 876 1604 884
rect 1324 776 1332 784
rect 1164 736 1172 744
rect 1308 736 1316 744
rect 1276 716 1284 724
rect 892 696 900 704
rect 924 702 932 704
rect 924 696 932 702
rect 1164 696 1172 704
rect 732 636 740 644
rect 732 616 740 624
rect 700 556 708 564
rect 524 516 532 524
rect 588 516 596 524
rect 620 516 628 524
rect 428 496 436 504
rect 364 476 372 484
rect 444 416 452 424
rect 764 556 772 564
rect 812 536 820 544
rect 588 496 596 504
rect 684 496 692 504
rect 796 496 804 504
rect 652 456 660 464
rect 460 376 468 384
rect 220 236 228 244
rect 268 276 276 284
rect 252 216 260 224
rect 380 236 388 244
rect 588 316 596 324
rect 620 316 628 324
rect 556 296 564 304
rect 636 296 644 304
rect 540 276 548 284
rect 668 316 676 324
rect 940 616 948 624
rect 908 596 916 604
rect 892 556 900 564
rect 860 536 868 544
rect 924 536 932 544
rect 716 476 724 484
rect 828 476 836 484
rect 739 406 747 414
rect 749 406 757 414
rect 759 406 767 414
rect 769 406 777 414
rect 779 406 787 414
rect 789 406 797 414
rect 716 316 724 324
rect 668 276 676 284
rect 684 276 692 284
rect 700 276 708 284
rect 588 256 596 264
rect 556 176 564 184
rect 236 136 244 144
rect 300 136 308 144
rect 492 136 500 144
rect 684 256 692 264
rect 348 116 356 124
rect 76 96 84 104
rect 188 96 196 104
rect 252 56 260 64
rect 812 296 820 304
rect 812 256 820 264
rect 796 136 804 144
rect 764 96 772 104
rect 876 296 884 304
rect 924 276 932 284
rect 860 236 868 244
rect 892 256 900 264
rect 844 116 852 124
rect 956 556 964 564
rect 956 496 964 504
rect 956 316 964 324
rect 972 236 980 244
rect 1292 676 1300 684
rect 1340 676 1348 684
rect 1388 676 1396 684
rect 1164 656 1172 664
rect 1148 636 1156 644
rect 1116 596 1124 604
rect 1244 616 1252 624
rect 1212 576 1220 584
rect 1196 556 1204 564
rect 1404 656 1412 664
rect 1356 596 1364 604
rect 1196 536 1204 544
rect 1052 516 1060 524
rect 1068 516 1076 524
rect 1020 496 1028 504
rect 1036 376 1044 384
rect 1004 336 1012 344
rect 1004 296 1012 304
rect 1132 416 1140 424
rect 1084 336 1092 344
rect 1276 516 1284 524
rect 1164 396 1172 404
rect 1196 396 1204 404
rect 1020 276 1028 284
rect 988 216 996 224
rect 1324 416 1332 424
rect 1388 576 1396 584
rect 1436 556 1444 564
rect 1404 536 1412 544
rect 1404 516 1412 524
rect 1420 516 1428 524
rect 1500 836 1508 844
rect 1548 796 1556 804
rect 1516 676 1524 684
rect 1516 656 1524 664
rect 1500 576 1508 584
rect 1532 556 1540 564
rect 1516 536 1524 544
rect 1388 456 1396 464
rect 1468 396 1476 404
rect 1580 716 1588 724
rect 1580 676 1588 684
rect 1612 836 1620 844
rect 1724 1116 1732 1124
rect 1644 1076 1652 1084
rect 1708 996 1716 1004
rect 1836 1316 1844 1324
rect 1820 1296 1828 1304
rect 1804 1276 1812 1284
rect 1804 1256 1812 1264
rect 1852 1256 1860 1264
rect 1900 1236 1908 1244
rect 1852 1216 1860 1224
rect 1836 956 1844 964
rect 1868 936 1876 944
rect 1724 896 1732 904
rect 1660 776 1668 784
rect 1628 756 1636 764
rect 1820 776 1828 784
rect 1740 696 1748 704
rect 1820 696 1828 704
rect 1852 702 1860 704
rect 1852 696 1860 702
rect 1692 676 1700 684
rect 1660 656 1668 664
rect 1708 656 1716 664
rect 1596 576 1604 584
rect 1564 536 1572 544
rect 1612 536 1620 544
rect 1676 616 1684 624
rect 1644 556 1652 564
rect 1692 556 1700 564
rect 1772 556 1780 564
rect 1644 536 1652 544
rect 1676 536 1684 544
rect 1708 536 1716 544
rect 1628 496 1636 504
rect 1532 476 1540 484
rect 1516 396 1524 404
rect 1484 336 1492 344
rect 1196 302 1204 304
rect 1196 296 1204 302
rect 1260 276 1268 284
rect 1164 256 1172 264
rect 1148 236 1156 244
rect 988 136 996 144
rect 1004 136 1012 144
rect 1052 136 1060 144
rect 1100 136 1108 144
rect 1196 216 1204 224
rect 1212 196 1220 204
rect 1132 156 1140 164
rect 1196 156 1204 164
rect 1180 136 1188 144
rect 1276 216 1284 224
rect 1228 136 1236 144
rect 1068 96 1076 104
rect 1276 96 1284 104
rect 844 36 852 44
rect 940 36 948 44
rect 684 16 692 24
rect 716 16 724 24
rect 828 16 836 24
rect 739 6 747 14
rect 749 6 757 14
rect 759 6 767 14
rect 769 6 777 14
rect 779 6 787 14
rect 789 6 797 14
rect 860 16 868 24
rect 1036 76 1044 84
rect 988 16 996 24
rect 1164 36 1172 44
rect 1388 156 1396 164
rect 1372 76 1380 84
rect 1260 36 1268 44
rect 1340 36 1348 44
rect 1596 396 1604 404
rect 1612 336 1620 344
rect 1564 296 1572 304
rect 1548 256 1556 264
rect 1436 216 1444 224
rect 1516 236 1524 244
rect 1484 196 1492 204
rect 1468 176 1476 184
rect 1516 176 1524 184
rect 1468 156 1476 164
rect 1532 156 1540 164
rect 1436 136 1444 144
rect 1468 116 1476 124
rect 1500 96 1508 104
rect 1404 16 1412 24
rect 1580 276 1588 284
rect 1644 276 1652 284
rect 1644 236 1652 244
rect 1628 196 1636 204
rect 1596 156 1604 164
rect 1660 156 1668 164
rect 1644 36 1652 44
rect 1564 16 1572 24
rect 1596 16 1604 24
rect 1708 516 1716 524
rect 1788 516 1796 524
rect 1708 356 1716 364
rect 1724 336 1732 344
rect 1820 616 1828 624
rect 1852 616 1860 624
rect 1820 576 1828 584
rect 1948 1456 1956 1464
rect 1980 1576 1988 1584
rect 2380 1956 2388 1964
rect 2300 1916 2308 1924
rect 2204 1876 2212 1884
rect 2220 1876 2228 1884
rect 2188 1856 2196 1864
rect 2268 1856 2276 1864
rect 2188 1816 2196 1824
rect 2332 1816 2340 1824
rect 2243 1806 2251 1814
rect 2253 1806 2261 1814
rect 2263 1806 2271 1814
rect 2273 1806 2281 1814
rect 2283 1806 2291 1814
rect 2293 1806 2301 1814
rect 2220 1796 2228 1804
rect 2172 1736 2180 1744
rect 2188 1736 2196 1744
rect 2108 1716 2116 1724
rect 2188 1716 2196 1724
rect 2108 1696 2116 1704
rect 2156 1696 2164 1704
rect 2204 1696 2212 1704
rect 2220 1696 2228 1704
rect 2076 1676 2084 1684
rect 2012 1596 2020 1604
rect 1996 1556 2004 1564
rect 1980 1536 1988 1544
rect 1996 1536 2004 1544
rect 2028 1576 2036 1584
rect 2092 1576 2100 1584
rect 2140 1576 2148 1584
rect 2076 1556 2084 1564
rect 2060 1536 2068 1544
rect 2012 1496 2020 1504
rect 2044 1496 2052 1504
rect 1932 1396 1940 1404
rect 1964 1356 1972 1364
rect 1948 1336 1956 1344
rect 1980 1336 1988 1344
rect 1996 1336 2004 1344
rect 1964 1096 1972 1104
rect 2028 1436 2036 1444
rect 2012 1316 2020 1324
rect 2060 1376 2068 1384
rect 2044 1336 2052 1344
rect 2028 1276 2036 1284
rect 2044 1256 2052 1264
rect 2012 1136 2020 1144
rect 2204 1536 2212 1544
rect 2172 1516 2180 1524
rect 2188 1516 2196 1524
rect 2172 1456 2180 1464
rect 2156 1436 2164 1444
rect 2172 1436 2180 1444
rect 2124 1376 2132 1384
rect 2140 1376 2148 1384
rect 2188 1376 2196 1384
rect 2156 1296 2164 1304
rect 2092 1216 2100 1224
rect 2076 1136 2084 1144
rect 1980 1076 1988 1084
rect 1996 1076 2004 1084
rect 1964 1016 1972 1024
rect 1996 956 2004 964
rect 2060 1076 2068 1084
rect 2060 1016 2068 1024
rect 2108 1196 2116 1204
rect 2172 1236 2180 1244
rect 2188 1236 2196 1244
rect 2172 1196 2180 1204
rect 2188 1176 2196 1184
rect 2268 1656 2276 1664
rect 2300 1656 2308 1664
rect 2252 1616 2260 1624
rect 2268 1596 2276 1604
rect 2252 1576 2260 1584
rect 2284 1576 2292 1584
rect 2236 1536 2244 1544
rect 2220 1496 2228 1504
rect 2284 1476 2292 1484
rect 2300 1476 2308 1484
rect 2236 1456 2244 1464
rect 2252 1456 2260 1464
rect 2348 1736 2356 1744
rect 2444 2256 2452 2264
rect 2828 2776 2836 2784
rect 2844 2776 2852 2784
rect 2812 2676 2820 2684
rect 2748 2656 2756 2664
rect 2812 2636 2820 2644
rect 2796 2556 2804 2564
rect 2764 2536 2772 2544
rect 2764 2516 2772 2524
rect 2732 2376 2740 2384
rect 2604 2356 2612 2364
rect 2636 2356 2644 2364
rect 2492 2236 2500 2244
rect 2540 2236 2548 2244
rect 2556 2156 2564 2164
rect 2588 2156 2596 2164
rect 2620 2276 2628 2284
rect 2668 2276 2676 2284
rect 2700 2276 2708 2284
rect 2620 2256 2628 2264
rect 2652 2216 2660 2224
rect 2540 2116 2548 2124
rect 2588 2116 2596 2124
rect 2524 2076 2532 2084
rect 2716 2196 2724 2204
rect 2668 2136 2676 2144
rect 2700 2136 2708 2144
rect 2748 2156 2756 2164
rect 2796 2316 2804 2324
rect 2764 2136 2772 2144
rect 2780 2116 2788 2124
rect 2668 2096 2676 2104
rect 2604 2056 2612 2064
rect 2524 2016 2532 2024
rect 2540 2016 2548 2024
rect 2492 1896 2500 1904
rect 2540 1896 2548 1904
rect 2588 1896 2596 1904
rect 2620 1902 2628 1904
rect 2620 1896 2628 1902
rect 2428 1876 2436 1884
rect 2460 1876 2468 1884
rect 2524 1856 2532 1864
rect 2412 1836 2420 1844
rect 2588 1856 2596 1864
rect 2620 1856 2628 1864
rect 2588 1836 2596 1844
rect 2556 1796 2564 1804
rect 2556 1776 2564 1784
rect 2460 1756 2468 1764
rect 2444 1736 2452 1744
rect 2396 1716 2404 1724
rect 2428 1696 2436 1704
rect 2364 1676 2372 1684
rect 2380 1676 2388 1684
rect 2332 1636 2340 1644
rect 2380 1536 2388 1544
rect 2412 1676 2420 1684
rect 2412 1576 2420 1584
rect 2396 1516 2404 1524
rect 2476 1676 2484 1684
rect 2892 2976 2900 2984
rect 2972 2976 2980 2984
rect 2940 2956 2948 2964
rect 2924 2916 2932 2924
rect 2908 2896 2916 2904
rect 2940 2796 2948 2804
rect 2892 2756 2900 2764
rect 2844 2696 2852 2704
rect 2876 2656 2884 2664
rect 3036 3196 3044 3204
rect 3084 3456 3092 3464
rect 3068 3216 3076 3224
rect 3052 3176 3060 3184
rect 3068 3116 3076 3124
rect 3100 3436 3108 3444
rect 3164 3476 3172 3484
rect 3196 3516 3204 3524
rect 3212 3516 3220 3524
rect 3180 3416 3188 3424
rect 3116 3356 3124 3364
rect 3148 3356 3156 3364
rect 3100 3136 3108 3144
rect 3100 3096 3108 3104
rect 3052 3036 3060 3044
rect 3004 2836 3012 2844
rect 3036 2756 3044 2764
rect 3020 2736 3028 2744
rect 3084 2996 3092 3004
rect 3068 2916 3076 2924
rect 2956 2696 2964 2704
rect 2924 2656 2932 2664
rect 2924 2596 2932 2604
rect 2860 2536 2868 2544
rect 3052 2676 3060 2684
rect 2988 2656 2996 2664
rect 3052 2656 3060 2664
rect 2972 2636 2980 2644
rect 3068 2636 3076 2644
rect 3004 2576 3012 2584
rect 2972 2556 2980 2564
rect 2988 2556 2996 2564
rect 3004 2536 3012 2544
rect 2956 2496 2964 2504
rect 3004 2496 3012 2504
rect 3068 2496 3076 2504
rect 2860 2336 2868 2344
rect 2924 2336 2932 2344
rect 2844 2296 2852 2304
rect 2828 2216 2836 2224
rect 2812 1976 2820 1984
rect 2844 2196 2852 2204
rect 2908 2276 2916 2284
rect 2892 2196 2900 2204
rect 2908 2156 2916 2164
rect 2892 2136 2900 2144
rect 2860 2036 2868 2044
rect 2828 1936 2836 1944
rect 2796 1896 2804 1904
rect 2844 1896 2852 1904
rect 2748 1876 2756 1884
rect 2796 1876 2804 1884
rect 2876 1876 2884 1884
rect 2892 1876 2900 1884
rect 2732 1856 2740 1864
rect 2700 1776 2708 1784
rect 2620 1736 2628 1744
rect 2572 1716 2580 1724
rect 2556 1576 2564 1584
rect 2508 1556 2516 1564
rect 2444 1536 2452 1544
rect 2524 1536 2532 1544
rect 2556 1536 2564 1544
rect 2540 1516 2548 1524
rect 2620 1516 2628 1524
rect 2380 1496 2388 1504
rect 2444 1496 2452 1504
rect 2524 1496 2532 1504
rect 2508 1476 2516 1484
rect 2380 1456 2388 1464
rect 2300 1436 2308 1444
rect 2316 1436 2324 1444
rect 2243 1406 2251 1414
rect 2253 1406 2261 1414
rect 2263 1406 2271 1414
rect 2273 1406 2281 1414
rect 2283 1406 2291 1414
rect 2293 1406 2301 1414
rect 2220 1396 2228 1404
rect 2396 1416 2404 1424
rect 2332 1336 2340 1344
rect 2364 1336 2372 1344
rect 2220 1256 2228 1264
rect 2140 1136 2148 1144
rect 2204 1136 2212 1144
rect 2140 1096 2148 1104
rect 2156 1096 2164 1104
rect 2124 1076 2132 1084
rect 2092 1016 2100 1024
rect 2124 1016 2132 1024
rect 2140 1016 2148 1024
rect 2076 996 2084 1004
rect 1964 936 1972 944
rect 2012 916 2020 924
rect 2028 916 2036 924
rect 1964 896 1972 904
rect 1932 796 1940 804
rect 1916 676 1924 684
rect 1948 676 1956 684
rect 1916 616 1924 624
rect 1884 596 1892 604
rect 1868 556 1876 564
rect 1932 556 1940 564
rect 1836 536 1844 544
rect 1820 516 1828 524
rect 1884 456 1892 464
rect 1932 436 1940 444
rect 1884 416 1892 424
rect 1804 316 1812 324
rect 1868 316 1876 324
rect 1708 302 1716 304
rect 1708 296 1716 302
rect 1772 296 1780 304
rect 1804 276 1812 284
rect 1852 276 1860 284
rect 1772 136 1780 144
rect 1692 116 1700 124
rect 2076 916 2084 924
rect 2012 796 2020 804
rect 2092 816 2100 824
rect 2076 756 2084 764
rect 2028 736 2036 744
rect 2060 736 2068 744
rect 2044 696 2052 704
rect 1996 656 2004 664
rect 2012 656 2020 664
rect 2012 616 2020 624
rect 2092 716 2100 724
rect 2188 1076 2196 1084
rect 2172 996 2180 1004
rect 2188 916 2196 924
rect 2124 736 2132 744
rect 2108 696 2116 704
rect 2140 616 2148 624
rect 1996 556 2004 564
rect 2076 556 2084 564
rect 1980 536 1988 544
rect 2268 1176 2276 1184
rect 2236 1096 2244 1104
rect 2300 1316 2308 1324
rect 2332 1316 2340 1324
rect 2316 1296 2324 1304
rect 2348 1296 2356 1304
rect 2300 1156 2308 1164
rect 2348 1196 2356 1204
rect 2444 1396 2452 1404
rect 2476 1336 2484 1344
rect 2460 1296 2468 1304
rect 2636 1456 2644 1464
rect 2684 1616 2692 1624
rect 2812 1836 2820 1844
rect 2860 1796 2868 1804
rect 2780 1776 2788 1784
rect 2764 1756 2772 1764
rect 2764 1716 2772 1724
rect 2732 1696 2740 1704
rect 2748 1696 2756 1704
rect 2700 1596 2708 1604
rect 2684 1536 2692 1544
rect 2588 1376 2596 1384
rect 2540 1356 2548 1364
rect 2556 1356 2564 1364
rect 2700 1516 2708 1524
rect 2684 1456 2692 1464
rect 2700 1456 2708 1464
rect 2732 1596 2740 1604
rect 2732 1576 2740 1584
rect 2764 1616 2772 1624
rect 2764 1576 2772 1584
rect 2748 1516 2756 1524
rect 2844 1716 2852 1724
rect 2860 1696 2868 1704
rect 2828 1656 2836 1664
rect 2796 1616 2804 1624
rect 2764 1476 2772 1484
rect 2716 1416 2724 1424
rect 2764 1416 2772 1424
rect 2700 1376 2708 1384
rect 2748 1376 2756 1384
rect 2668 1336 2676 1344
rect 2684 1336 2692 1344
rect 2556 1316 2564 1324
rect 2620 1316 2628 1324
rect 2524 1296 2532 1304
rect 2556 1296 2564 1304
rect 2428 1236 2436 1244
rect 2492 1276 2500 1284
rect 2508 1276 2516 1284
rect 2540 1276 2548 1284
rect 2524 1176 2532 1184
rect 2364 1136 2372 1144
rect 2444 1136 2452 1144
rect 2508 1136 2516 1144
rect 2476 1116 2484 1124
rect 2412 1096 2420 1104
rect 2540 1096 2548 1104
rect 2364 1076 2372 1084
rect 2428 1076 2436 1084
rect 2492 1076 2500 1084
rect 2508 1076 2516 1084
rect 2243 1006 2251 1014
rect 2253 1006 2261 1014
rect 2263 1006 2271 1014
rect 2273 1006 2281 1014
rect 2283 1006 2291 1014
rect 2293 1006 2301 1014
rect 2220 956 2228 964
rect 2204 736 2212 744
rect 2204 696 2212 704
rect 2252 956 2260 964
rect 2412 1016 2420 1024
rect 2444 1016 2452 1024
rect 2396 996 2404 1004
rect 2380 956 2388 964
rect 2348 916 2356 924
rect 2268 796 2276 804
rect 2364 896 2372 904
rect 2332 776 2340 784
rect 2364 776 2372 784
rect 2348 736 2356 744
rect 2332 696 2340 704
rect 2572 1196 2580 1204
rect 2732 1316 2740 1324
rect 2860 1576 2868 1584
rect 2876 1576 2884 1584
rect 3004 2316 3012 2324
rect 3132 3336 3140 3344
rect 3212 3476 3220 3484
rect 3228 3436 3236 3444
rect 3292 4036 3300 4044
rect 3308 3896 3316 3904
rect 3532 4576 3540 4584
rect 3612 4576 3620 4584
rect 3676 4536 3684 4544
rect 3564 4516 3572 4524
rect 3724 4516 3732 4524
rect 3484 4436 3492 4444
rect 3580 4436 3588 4444
rect 3468 4356 3476 4364
rect 3500 4316 3508 4324
rect 3468 4276 3476 4284
rect 3564 4276 3572 4284
rect 3516 4256 3524 4264
rect 3548 4256 3556 4264
rect 3484 4236 3492 4244
rect 3484 4156 3492 4164
rect 3340 4116 3348 4124
rect 3548 4116 3556 4124
rect 3644 4456 3652 4464
rect 3747 4406 3755 4414
rect 3757 4406 3765 4414
rect 3767 4406 3775 4414
rect 3777 4406 3785 4414
rect 3787 4406 3795 4414
rect 3797 4406 3805 4414
rect 3724 4336 3732 4344
rect 3612 4316 3620 4324
rect 3708 4316 3716 4324
rect 3820 4316 3828 4324
rect 3804 4296 3812 4304
rect 3676 4276 3684 4284
rect 3644 4256 3652 4264
rect 3724 4256 3732 4264
rect 3596 4236 3604 4244
rect 3580 4176 3588 4184
rect 3772 4176 3780 4184
rect 3612 4136 3620 4144
rect 3868 4696 3876 4704
rect 3980 4676 3988 4684
rect 3884 4656 3892 4664
rect 4108 4896 4116 4904
rect 4092 4756 4100 4764
rect 4076 4736 4084 4744
rect 4092 4696 4100 4704
rect 4060 4636 4068 4644
rect 3868 4556 3876 4564
rect 3980 4536 3988 4544
rect 4028 4536 4036 4544
rect 3932 4516 3940 4524
rect 3852 4456 3860 4464
rect 3868 4436 3876 4444
rect 4124 4856 4132 4864
rect 4124 4756 4132 4764
rect 4156 4716 4164 4724
rect 4188 4776 4196 4784
rect 4172 4696 4180 4704
rect 4236 4956 4244 4964
rect 4316 5056 4324 5064
rect 4492 4976 4500 4984
rect 4300 4936 4308 4944
rect 4348 4936 4356 4944
rect 4396 4936 4404 4944
rect 4252 4776 4260 4784
rect 4204 4756 4212 4764
rect 4428 4896 4436 4904
rect 4364 4796 4372 4804
rect 4252 4716 4260 4724
rect 4220 4676 4228 4684
rect 4188 4556 4196 4564
rect 4284 4556 4292 4564
rect 4316 4556 4324 4564
rect 4156 4536 4164 4544
rect 4220 4536 4228 4544
rect 4092 4516 4100 4524
rect 4268 4516 4276 4524
rect 4028 4496 4036 4504
rect 4060 4496 4068 4504
rect 4140 4476 4148 4484
rect 4076 4456 4084 4464
rect 4044 4396 4052 4404
rect 4012 4376 4020 4384
rect 3900 4196 3908 4204
rect 3948 4196 3956 4204
rect 3964 4176 3972 4184
rect 3916 4136 3924 4144
rect 3644 4118 3652 4124
rect 3644 4116 3652 4118
rect 3836 4116 3844 4124
rect 3852 4116 3860 4124
rect 3500 4096 3508 4104
rect 3548 4096 3556 4104
rect 3564 4096 3572 4104
rect 3884 4096 3892 4104
rect 3388 4036 3396 4044
rect 3356 3896 3364 3904
rect 3436 3896 3444 3904
rect 3516 3896 3524 3904
rect 3324 3876 3332 3884
rect 3308 3856 3316 3864
rect 3324 3836 3332 3844
rect 3324 3796 3332 3804
rect 3388 3876 3396 3884
rect 3532 3876 3540 3884
rect 3452 3836 3460 3844
rect 3340 3776 3348 3784
rect 3500 3776 3508 3784
rect 3308 3736 3316 3744
rect 3324 3716 3332 3724
rect 3404 3716 3412 3724
rect 3292 3696 3300 3704
rect 3292 3596 3300 3604
rect 3276 3476 3284 3484
rect 3260 3456 3268 3464
rect 3260 3436 3268 3444
rect 3244 3376 3252 3384
rect 3212 3356 3220 3364
rect 3196 3296 3204 3304
rect 3244 3296 3252 3304
rect 3228 3256 3236 3264
rect 3196 3156 3204 3164
rect 3212 3156 3220 3164
rect 3340 3596 3348 3604
rect 3388 3636 3396 3644
rect 3356 3576 3364 3584
rect 3372 3576 3380 3584
rect 3324 3516 3332 3524
rect 3324 3336 3332 3344
rect 3404 3536 3412 3544
rect 3436 3516 3444 3524
rect 3372 3476 3380 3484
rect 3372 3456 3380 3464
rect 3404 3456 3412 3464
rect 4028 4296 4036 4304
rect 4236 4456 4244 4464
rect 4204 4356 4212 4364
rect 4172 4316 4180 4324
rect 4444 4702 4452 4704
rect 4444 4696 4452 4702
rect 4300 4536 4308 4544
rect 3996 4176 4004 4184
rect 4060 4236 4068 4244
rect 4108 4236 4116 4244
rect 4092 4196 4100 4204
rect 4044 4156 4052 4164
rect 4076 4156 4084 4164
rect 3996 4136 4004 4144
rect 4044 4136 4052 4144
rect 3964 4096 3972 4104
rect 3900 4036 3908 4044
rect 3747 4006 3755 4014
rect 3757 4006 3765 4014
rect 3767 4006 3775 4014
rect 3777 4006 3785 4014
rect 3787 4006 3795 4014
rect 3797 4006 3805 4014
rect 3756 3936 3764 3944
rect 3564 3896 3572 3904
rect 3628 3902 3636 3904
rect 3628 3896 3636 3902
rect 4140 4156 4148 4164
rect 4188 4136 4196 4144
rect 4124 4116 4132 4124
rect 4172 4116 4180 4124
rect 4076 4076 4084 4084
rect 4028 4056 4036 4064
rect 4012 3956 4020 3964
rect 4140 4096 4148 4104
rect 4396 4556 4404 4564
rect 4380 4476 4388 4484
rect 4284 4296 4292 4304
rect 4300 4296 4308 4304
rect 4332 4296 4340 4304
rect 4364 4296 4372 4304
rect 4300 4256 4308 4264
rect 4300 4236 4308 4244
rect 4316 4216 4324 4224
rect 4284 4136 4292 4144
rect 4364 4236 4372 4244
rect 4380 4176 4388 4184
rect 4556 5076 4564 5084
rect 4748 5076 4756 5084
rect 4796 5076 4804 5084
rect 4812 5076 4820 5084
rect 4876 5076 4884 5084
rect 4652 5056 4660 5064
rect 4700 5056 4708 5064
rect 4764 5056 4772 5064
rect 4812 5056 4820 5064
rect 4828 5056 4836 5064
rect 4924 5056 4932 5064
rect 4556 5036 4564 5044
rect 4588 5036 4596 5044
rect 4588 4936 4596 4944
rect 4796 4936 4804 4944
rect 4620 4876 4628 4884
rect 4588 4796 4596 4804
rect 4748 4776 4756 4784
rect 4748 4756 4756 4764
rect 4732 4696 4740 4704
rect 4588 4636 4596 4644
rect 4620 4636 4628 4644
rect 4540 4556 4548 4564
rect 4556 4556 4564 4564
rect 4412 4516 4420 4524
rect 4444 4316 4452 4324
rect 4428 4302 4436 4304
rect 4428 4296 4436 4302
rect 4572 4516 4580 4524
rect 4556 4436 4564 4444
rect 4652 4616 4660 4624
rect 4796 4716 4804 4724
rect 4956 4996 4964 5004
rect 4988 4996 4996 5004
rect 4892 4976 4900 4984
rect 4972 4976 4980 4984
rect 4860 4956 4868 4964
rect 5116 5076 5124 5084
rect 5148 5116 5156 5124
rect 5180 5116 5188 5124
rect 5516 5116 5524 5124
rect 5612 5116 5620 5124
rect 5340 5096 5348 5104
rect 5180 5076 5188 5084
rect 5228 5076 5236 5084
rect 5356 5076 5364 5084
rect 5404 5096 5412 5104
rect 5468 5096 5476 5104
rect 5068 5056 5076 5064
rect 5148 5056 5156 5064
rect 5212 5056 5220 5064
rect 5388 5056 5396 5064
rect 5452 5056 5460 5064
rect 5004 4976 5012 4984
rect 5251 5006 5259 5014
rect 5261 5006 5269 5014
rect 5271 5006 5279 5014
rect 5281 5006 5289 5014
rect 5291 5006 5299 5014
rect 5301 5006 5309 5014
rect 5372 4976 5380 4984
rect 5020 4956 5028 4964
rect 5164 4956 5172 4964
rect 5196 4936 5204 4944
rect 5228 4936 5236 4944
rect 5340 4936 5348 4944
rect 5052 4916 5060 4924
rect 4876 4896 4884 4904
rect 4780 4696 4788 4704
rect 4796 4616 4804 4624
rect 4668 4576 4676 4584
rect 4764 4576 4772 4584
rect 4780 4576 4788 4584
rect 4796 4576 4804 4584
rect 4764 4556 4772 4564
rect 4636 4536 4644 4544
rect 4844 4596 4852 4604
rect 4908 4676 4916 4684
rect 4908 4636 4916 4644
rect 4828 4556 4836 4564
rect 4812 4516 4820 4524
rect 4876 4536 4884 4544
rect 4748 4476 4756 4484
rect 4844 4476 4852 4484
rect 4620 4456 4628 4464
rect 4700 4416 4708 4424
rect 4812 4356 4820 4364
rect 4828 4336 4836 4344
rect 4972 4796 4980 4804
rect 5148 4896 5156 4904
rect 5068 4876 5076 4884
rect 4988 4776 4996 4784
rect 4972 4756 4980 4764
rect 4972 4676 4980 4684
rect 4972 4656 4980 4664
rect 4956 4616 4964 4624
rect 4940 4496 4948 4504
rect 4940 4436 4948 4444
rect 4924 4376 4932 4384
rect 4908 4336 4916 4344
rect 4956 4396 4964 4404
rect 4604 4296 4612 4304
rect 4652 4296 4660 4304
rect 4780 4296 4788 4304
rect 4860 4296 4868 4304
rect 4892 4296 4900 4304
rect 4524 4256 4532 4264
rect 4508 4196 4516 4204
rect 4348 4156 4356 4164
rect 4476 4156 4484 4164
rect 4380 4136 4388 4144
rect 4332 4116 4340 4124
rect 4268 4096 4276 4104
rect 4300 4096 4308 4104
rect 4236 4076 4244 4084
rect 4124 3976 4132 3984
rect 4268 3996 4276 4004
rect 4204 3956 4212 3964
rect 4236 3956 4244 3964
rect 4124 3936 4132 3944
rect 4140 3936 4148 3944
rect 4172 3936 4180 3944
rect 3820 3876 3828 3884
rect 3836 3876 3844 3884
rect 3564 3856 3572 3864
rect 3564 3796 3572 3804
rect 3500 3716 3508 3724
rect 3532 3716 3540 3724
rect 3548 3716 3556 3724
rect 3532 3676 3540 3684
rect 3500 3656 3508 3664
rect 3612 3776 3620 3784
rect 3596 3756 3604 3764
rect 3580 3716 3588 3724
rect 3580 3696 3588 3704
rect 3724 3696 3732 3704
rect 3708 3656 3716 3664
rect 3580 3616 3588 3624
rect 3500 3496 3508 3504
rect 3372 3416 3380 3424
rect 3484 3416 3492 3424
rect 3468 3376 3476 3384
rect 3356 3296 3364 3304
rect 3340 3256 3348 3264
rect 3276 3216 3284 3224
rect 3132 3116 3140 3124
rect 3148 3116 3156 3124
rect 3244 3116 3252 3124
rect 3180 3076 3188 3084
rect 3324 3116 3332 3124
rect 3260 3056 3268 3064
rect 3308 3056 3316 3064
rect 3244 3036 3252 3044
rect 3116 2996 3124 3004
rect 3164 2996 3172 3004
rect 3228 2956 3236 2964
rect 3212 2936 3220 2944
rect 3276 2956 3284 2964
rect 3324 3016 3332 3024
rect 3324 2956 3332 2964
rect 3372 3196 3380 3204
rect 3404 3296 3412 3304
rect 3420 3296 3428 3304
rect 3388 3176 3396 3184
rect 3420 3156 3428 3164
rect 3436 3156 3444 3164
rect 3356 3096 3364 3104
rect 3388 3096 3396 3104
rect 3372 3076 3380 3084
rect 3340 2936 3348 2944
rect 3372 2956 3380 2964
rect 3260 2916 3268 2924
rect 3212 2896 3220 2904
rect 3196 2836 3204 2844
rect 3228 2816 3236 2824
rect 3132 2776 3140 2784
rect 3116 2736 3124 2744
rect 3244 2776 3252 2784
rect 3228 2756 3236 2764
rect 3148 2736 3156 2744
rect 3308 2896 3316 2904
rect 3116 2676 3124 2684
rect 3260 2676 3268 2684
rect 3276 2676 3284 2684
rect 3260 2596 3268 2604
rect 3148 2536 3156 2544
rect 3276 2536 3284 2544
rect 3180 2516 3188 2524
rect 3228 2516 3236 2524
rect 3228 2456 3236 2464
rect 3228 2396 3236 2404
rect 3116 2376 3124 2384
rect 3180 2376 3188 2384
rect 3212 2376 3220 2384
rect 2988 2156 2996 2164
rect 3036 2156 3044 2164
rect 3084 2156 3092 2164
rect 3148 2156 3156 2164
rect 2956 2136 2964 2144
rect 2988 2136 2996 2144
rect 2940 2056 2948 2064
rect 3324 2876 3332 2884
rect 3372 2836 3380 2844
rect 3340 2736 3348 2744
rect 3356 2736 3364 2744
rect 3372 2716 3380 2724
rect 3372 2676 3380 2684
rect 3356 2616 3364 2624
rect 3420 2856 3428 2864
rect 3404 2776 3412 2784
rect 3628 3516 3636 3524
rect 3612 3496 3620 3504
rect 3564 3476 3572 3484
rect 3484 3336 3492 3344
rect 3532 3336 3540 3344
rect 3452 3076 3460 3084
rect 3692 3516 3700 3524
rect 3660 3456 3668 3464
rect 3612 3396 3620 3404
rect 3596 3356 3604 3364
rect 3692 3336 3700 3344
rect 3516 3316 3524 3324
rect 3580 3316 3588 3324
rect 3628 3316 3636 3324
rect 3500 3296 3508 3304
rect 3500 3136 3508 3144
rect 3500 3096 3508 3104
rect 3468 3036 3476 3044
rect 3468 2996 3476 3004
rect 3436 2736 3444 2744
rect 3660 3296 3668 3304
rect 3644 3256 3652 3264
rect 3580 3196 3588 3204
rect 3564 3176 3572 3184
rect 3548 3116 3556 3124
rect 3548 3096 3556 3104
rect 3628 3096 3636 3104
rect 3516 2936 3524 2944
rect 3612 3056 3620 3064
rect 3628 2936 3636 2944
rect 3548 2916 3556 2924
rect 3596 2916 3604 2924
rect 3532 2876 3540 2884
rect 3500 2856 3508 2864
rect 3564 2876 3572 2884
rect 3548 2796 3556 2804
rect 3420 2716 3428 2724
rect 3452 2716 3460 2724
rect 3484 2716 3492 2724
rect 3436 2696 3444 2704
rect 3468 2696 3476 2704
rect 3404 2676 3412 2684
rect 3388 2596 3396 2604
rect 3436 2616 3444 2624
rect 3420 2576 3428 2584
rect 3356 2556 3364 2564
rect 3260 2376 3268 2384
rect 3340 2496 3348 2504
rect 3308 2416 3316 2424
rect 3324 2336 3332 2344
rect 3292 2296 3300 2304
rect 3244 2276 3252 2284
rect 3276 2276 3284 2284
rect 3292 2276 3300 2284
rect 3276 2256 3284 2264
rect 3324 2256 3332 2264
rect 3452 2576 3460 2584
rect 3452 2556 3460 2564
rect 3516 2696 3524 2704
rect 3500 2536 3508 2544
rect 3564 2716 3572 2724
rect 3596 2836 3604 2844
rect 3628 2756 3636 2764
rect 3612 2696 3620 2704
rect 3596 2596 3604 2604
rect 3660 3216 3668 3224
rect 3692 3176 3700 3184
rect 3676 3136 3684 3144
rect 3660 2996 3668 3004
rect 3724 3636 3732 3644
rect 3692 2976 3700 2984
rect 3708 2956 3716 2964
rect 3692 2936 3700 2944
rect 3676 2916 3684 2924
rect 3660 2716 3668 2724
rect 3692 2856 3700 2864
rect 3708 2856 3716 2864
rect 3708 2776 3716 2784
rect 3692 2596 3700 2604
rect 3580 2536 3588 2544
rect 3596 2536 3604 2544
rect 3660 2536 3668 2544
rect 3500 2516 3508 2524
rect 3596 2516 3604 2524
rect 3468 2496 3476 2504
rect 3484 2476 3492 2484
rect 3372 2456 3380 2464
rect 3436 2456 3444 2464
rect 3388 2436 3396 2444
rect 3404 2356 3412 2364
rect 3420 2316 3428 2324
rect 3372 2296 3380 2304
rect 3420 2296 3428 2304
rect 3356 2276 3364 2284
rect 3340 2156 3348 2164
rect 3068 2136 3076 2144
rect 3116 2136 3124 2144
rect 3148 2136 3156 2144
rect 3260 2136 3268 2144
rect 3052 2116 3060 2124
rect 3036 2096 3044 2104
rect 3100 2096 3108 2104
rect 2956 2016 2964 2024
rect 2988 1996 2996 2004
rect 3004 1996 3012 2004
rect 2972 1876 2980 1884
rect 3068 1976 3076 1984
rect 3068 1916 3076 1924
rect 3052 1876 3060 1884
rect 3004 1856 3012 1864
rect 3004 1836 3012 1844
rect 3116 1716 3124 1724
rect 3020 1696 3028 1704
rect 3084 1696 3092 1704
rect 2988 1596 2996 1604
rect 3004 1596 3012 1604
rect 2924 1576 2932 1584
rect 2828 1516 2836 1524
rect 2860 1496 2868 1504
rect 2844 1476 2852 1484
rect 2828 1456 2836 1464
rect 2812 1316 2820 1324
rect 2844 1376 2852 1384
rect 2876 1376 2884 1384
rect 2956 1536 2964 1544
rect 2940 1516 2948 1524
rect 3052 1676 3060 1684
rect 3068 1676 3076 1684
rect 3132 1616 3140 1624
rect 3164 2036 3172 2044
rect 3276 2116 3284 2124
rect 3308 2116 3316 2124
rect 3212 2096 3220 2104
rect 3356 2076 3364 2084
rect 3404 2156 3412 2164
rect 3468 2336 3476 2344
rect 3452 2316 3460 2324
rect 3516 2376 3524 2384
rect 3468 2276 3476 2284
rect 3468 2136 3476 2144
rect 3436 2116 3444 2124
rect 3388 2036 3396 2044
rect 3468 2036 3476 2044
rect 3404 2016 3412 2024
rect 3404 1976 3412 1984
rect 3420 1976 3428 1984
rect 3340 1956 3348 1964
rect 3324 1916 3332 1924
rect 3228 1876 3236 1884
rect 3260 1876 3268 1884
rect 3180 1856 3188 1864
rect 3260 1796 3268 1804
rect 3228 1756 3236 1764
rect 3020 1576 3028 1584
rect 3052 1576 3060 1584
rect 3020 1556 3028 1564
rect 3036 1536 3044 1544
rect 3132 1536 3140 1544
rect 3036 1516 3044 1524
rect 3084 1516 3092 1524
rect 3116 1516 3124 1524
rect 2956 1496 2964 1504
rect 2940 1456 2948 1464
rect 3084 1496 3092 1504
rect 3068 1456 3076 1464
rect 2956 1376 2964 1384
rect 2892 1336 2900 1344
rect 2796 1296 2804 1304
rect 2812 1296 2820 1304
rect 2844 1296 2852 1304
rect 2652 1216 2660 1224
rect 2620 1196 2628 1204
rect 2604 1076 2612 1084
rect 2588 1016 2596 1024
rect 2556 996 2564 1004
rect 2636 1096 2644 1104
rect 2620 996 2628 1004
rect 2716 1256 2724 1264
rect 2796 1236 2804 1244
rect 2892 1236 2900 1244
rect 2892 1176 2900 1184
rect 2764 1156 2772 1164
rect 2732 1136 2740 1144
rect 2732 1116 2740 1124
rect 2764 1116 2772 1124
rect 2828 1116 2836 1124
rect 2684 1096 2692 1104
rect 2684 996 2692 1004
rect 2764 1096 2772 1104
rect 2796 1096 2804 1104
rect 2748 1076 2756 1084
rect 2508 976 2516 984
rect 2540 976 2548 984
rect 2588 976 2596 984
rect 2620 976 2628 984
rect 2652 976 2660 984
rect 2460 956 2468 964
rect 2780 1076 2788 1084
rect 2764 1056 2772 1064
rect 2540 956 2548 964
rect 2572 956 2580 964
rect 2700 956 2708 964
rect 2748 956 2756 964
rect 2764 956 2772 964
rect 2412 916 2420 924
rect 2556 916 2564 924
rect 2476 796 2484 804
rect 2492 796 2500 804
rect 2396 776 2404 784
rect 2428 776 2436 784
rect 2828 1076 2836 1084
rect 2844 1080 2852 1084
rect 2844 1076 2852 1080
rect 2892 1076 2900 1084
rect 2924 1336 2932 1344
rect 3052 1376 3060 1384
rect 3180 1416 3188 1424
rect 3212 1676 3220 1684
rect 3228 1616 3236 1624
rect 3292 1896 3300 1904
rect 3308 1796 3316 1804
rect 3324 1776 3332 1784
rect 3356 1936 3364 1944
rect 3388 1896 3396 1904
rect 3404 1876 3412 1884
rect 3452 1896 3460 1904
rect 3436 1876 3444 1884
rect 3420 1856 3428 1864
rect 3372 1796 3380 1804
rect 3436 1796 3444 1804
rect 3500 2296 3508 2304
rect 3580 2476 3588 2484
rect 3596 2416 3604 2424
rect 3580 2396 3588 2404
rect 3548 2316 3556 2324
rect 3548 2296 3556 2304
rect 3548 2256 3556 2264
rect 3532 2236 3540 2244
rect 3580 2236 3588 2244
rect 3564 2176 3572 2184
rect 3564 2096 3572 2104
rect 3628 2356 3636 2364
rect 3628 2316 3636 2324
rect 3628 2276 3636 2284
rect 3612 2156 3620 2164
rect 3644 2236 3652 2244
rect 3676 2516 3684 2524
rect 3676 2496 3684 2504
rect 3676 2356 3684 2364
rect 3747 3606 3755 3614
rect 3757 3606 3765 3614
rect 3767 3606 3775 3614
rect 3777 3606 3785 3614
rect 3787 3606 3795 3614
rect 3797 3606 3805 3614
rect 3788 3336 3796 3344
rect 3868 3856 3876 3864
rect 3900 3836 3908 3844
rect 3852 3736 3860 3744
rect 3932 3736 3940 3744
rect 4060 3716 4068 3724
rect 3916 3676 3924 3684
rect 3868 3496 3876 3504
rect 3900 3476 3908 3484
rect 3948 3616 3956 3624
rect 3932 3516 3940 3524
rect 3964 3476 3972 3484
rect 4044 3616 4052 3624
rect 4012 3516 4020 3524
rect 3932 3336 3940 3344
rect 3820 3316 3828 3324
rect 3948 3316 3956 3324
rect 3747 3206 3755 3214
rect 3757 3206 3765 3214
rect 3767 3206 3775 3214
rect 3777 3206 3785 3214
rect 3787 3206 3795 3214
rect 3797 3206 3805 3214
rect 3756 3176 3764 3184
rect 3740 3056 3748 3064
rect 3740 2976 3748 2984
rect 3820 3096 3828 3104
rect 3932 3276 3940 3284
rect 3900 3236 3908 3244
rect 3836 3016 3844 3024
rect 3884 2996 3892 3004
rect 3804 2916 3812 2924
rect 3756 2876 3764 2884
rect 3836 2836 3844 2844
rect 3747 2806 3755 2814
rect 3757 2806 3765 2814
rect 3767 2806 3775 2814
rect 3777 2806 3785 2814
rect 3787 2806 3795 2814
rect 3797 2806 3805 2814
rect 3756 2716 3764 2724
rect 3724 2556 3732 2564
rect 3868 2656 3876 2664
rect 3820 2556 3828 2564
rect 3740 2536 3748 2544
rect 3708 2476 3716 2484
rect 3788 2456 3796 2464
rect 3747 2406 3755 2414
rect 3757 2406 3765 2414
rect 3767 2406 3775 2414
rect 3777 2406 3785 2414
rect 3787 2406 3795 2414
rect 3797 2406 3805 2414
rect 3820 2396 3828 2404
rect 3724 2356 3732 2364
rect 3692 2256 3700 2264
rect 3708 2256 3716 2264
rect 3660 2156 3668 2164
rect 3724 2216 3732 2224
rect 3708 2156 3716 2164
rect 3660 2136 3668 2144
rect 3644 2116 3652 2124
rect 3596 2036 3604 2044
rect 3580 1996 3588 2004
rect 3516 1896 3524 1904
rect 3580 1896 3588 1904
rect 3500 1876 3508 1884
rect 3564 1876 3572 1884
rect 3532 1856 3540 1864
rect 3484 1836 3492 1844
rect 3500 1836 3508 1844
rect 3548 1816 3556 1824
rect 3580 1816 3588 1824
rect 3500 1776 3508 1784
rect 3372 1756 3380 1764
rect 3468 1756 3476 1764
rect 3292 1716 3300 1724
rect 3308 1696 3316 1704
rect 3276 1676 3284 1684
rect 3308 1676 3316 1684
rect 3244 1516 3252 1524
rect 3212 1496 3220 1504
rect 3244 1496 3252 1504
rect 3276 1456 3284 1464
rect 3212 1376 3220 1384
rect 3468 1736 3476 1744
rect 3564 1756 3572 1764
rect 3404 1718 3412 1724
rect 3404 1716 3412 1718
rect 3532 1696 3540 1704
rect 3516 1676 3524 1684
rect 3468 1596 3476 1604
rect 3372 1516 3380 1524
rect 3340 1476 3348 1484
rect 3308 1376 3316 1384
rect 3068 1336 3076 1344
rect 3292 1336 3300 1344
rect 3020 1296 3028 1304
rect 3004 1276 3012 1284
rect 3020 1276 3028 1284
rect 3052 1276 3060 1284
rect 3116 1276 3124 1284
rect 2972 1196 2980 1204
rect 2924 1176 2932 1184
rect 2972 1176 2980 1184
rect 2940 1136 2948 1144
rect 2908 1056 2916 1064
rect 2844 1036 2852 1044
rect 2876 1036 2884 1044
rect 2812 1016 2820 1024
rect 2876 976 2884 984
rect 3020 1116 3028 1124
rect 3036 1116 3044 1124
rect 2956 1036 2964 1044
rect 2972 1036 2980 1044
rect 2764 936 2772 944
rect 2780 936 2788 944
rect 2812 936 2820 944
rect 2844 936 2852 944
rect 2876 936 2884 944
rect 2588 916 2596 924
rect 2636 916 2644 924
rect 2668 916 2676 924
rect 2716 916 2724 924
rect 2572 896 2580 904
rect 2588 856 2596 864
rect 2524 796 2532 804
rect 2604 796 2612 804
rect 2636 776 2644 784
rect 2508 756 2516 764
rect 2492 736 2500 744
rect 2396 696 2404 704
rect 2444 696 2452 704
rect 2460 696 2468 704
rect 2220 656 2228 664
rect 2396 636 2404 644
rect 2460 636 2468 644
rect 2316 616 2324 624
rect 2243 606 2251 614
rect 2253 606 2261 614
rect 2263 606 2271 614
rect 2273 606 2281 614
rect 2283 606 2291 614
rect 2293 606 2301 614
rect 2220 596 2228 604
rect 2188 576 2196 584
rect 2172 556 2180 564
rect 2076 516 2084 524
rect 2012 496 2020 504
rect 1964 356 1972 364
rect 2044 416 2052 424
rect 2028 336 2036 344
rect 1948 296 1956 304
rect 1932 276 1940 284
rect 1884 176 1892 184
rect 2188 536 2196 544
rect 2156 516 2164 524
rect 2156 416 2164 424
rect 2172 416 2180 424
rect 2140 396 2148 404
rect 2076 376 2084 384
rect 2076 316 2084 324
rect 2140 316 2148 324
rect 2060 296 2068 304
rect 2108 296 2116 304
rect 2156 296 2164 304
rect 2364 556 2372 564
rect 2460 556 2468 564
rect 2300 536 2308 544
rect 2364 516 2372 524
rect 2316 496 2324 504
rect 2220 436 2228 444
rect 2380 416 2388 424
rect 2204 396 2212 404
rect 2188 276 2196 284
rect 2044 196 2052 204
rect 2060 156 2068 164
rect 2396 396 2404 404
rect 2300 316 2308 324
rect 2364 316 2372 324
rect 2236 276 2244 284
rect 2476 516 2484 524
rect 2508 696 2516 704
rect 2572 696 2580 704
rect 2604 696 2612 704
rect 2748 696 2756 704
rect 2620 656 2628 664
rect 2572 636 2580 644
rect 2524 616 2532 624
rect 2556 616 2564 624
rect 2556 556 2564 564
rect 2700 556 2708 564
rect 2700 536 2708 544
rect 2764 536 2772 544
rect 3084 1080 3092 1084
rect 3084 1076 3092 1080
rect 3052 1036 3060 1044
rect 3068 1016 3076 1024
rect 3196 1276 3204 1284
rect 3132 1256 3140 1264
rect 3244 1256 3252 1264
rect 3308 1316 3316 1324
rect 3340 1376 3348 1384
rect 3372 1356 3380 1364
rect 3388 1356 3396 1364
rect 3356 1336 3364 1344
rect 3372 1316 3380 1324
rect 3420 1336 3428 1344
rect 3484 1336 3492 1344
rect 3436 1316 3444 1324
rect 3468 1316 3476 1324
rect 3484 1316 3492 1324
rect 3500 1296 3508 1304
rect 3372 1276 3380 1284
rect 3404 1276 3412 1284
rect 3308 1256 3316 1264
rect 3324 1256 3332 1264
rect 3196 1176 3204 1184
rect 3276 1176 3284 1184
rect 3308 1176 3316 1184
rect 3276 1136 3284 1144
rect 3180 1116 3188 1124
rect 3276 1116 3284 1124
rect 3132 1076 3140 1084
rect 3164 1076 3172 1084
rect 3196 1076 3204 1084
rect 3244 1056 3252 1064
rect 3116 1036 3124 1044
rect 3196 1036 3204 1044
rect 3244 1036 3252 1044
rect 3148 1016 3156 1024
rect 3164 1016 3172 1024
rect 3084 976 3092 984
rect 3100 976 3108 984
rect 3004 956 3012 964
rect 2860 916 2868 924
rect 2908 916 2916 924
rect 2956 916 2964 924
rect 2828 856 2836 864
rect 2940 896 2948 904
rect 3068 936 3076 944
rect 3004 896 3012 904
rect 3228 1016 3236 1024
rect 3228 976 3236 984
rect 3164 936 3172 944
rect 3116 916 3124 924
rect 3148 916 3156 924
rect 3228 916 3236 924
rect 3180 876 3188 884
rect 2860 836 2868 844
rect 2956 836 2964 844
rect 2988 836 2996 844
rect 3228 836 3236 844
rect 2908 736 2916 744
rect 2876 696 2884 704
rect 2892 696 2900 704
rect 2940 696 2948 704
rect 2860 656 2868 664
rect 2876 616 2884 624
rect 2828 556 2836 564
rect 3100 796 3108 804
rect 3228 776 3236 784
rect 2988 716 2996 724
rect 3020 716 3028 724
rect 3084 716 3092 724
rect 3020 696 3028 704
rect 3052 696 3060 704
rect 3100 696 3108 704
rect 3116 696 3124 704
rect 2940 676 2948 684
rect 3020 676 3028 684
rect 3084 676 3092 684
rect 3004 656 3012 664
rect 2988 536 2996 544
rect 2716 516 2724 524
rect 2892 516 2900 524
rect 2652 456 2660 464
rect 2492 376 2500 384
rect 2460 336 2468 344
rect 2620 336 2628 344
rect 2428 316 2436 324
rect 2508 296 2516 304
rect 2604 296 2612 304
rect 2444 276 2452 284
rect 2412 256 2420 264
rect 2364 236 2372 244
rect 2243 206 2251 214
rect 2253 206 2261 214
rect 2263 206 2271 214
rect 2273 206 2281 214
rect 2283 206 2291 214
rect 2293 206 2301 214
rect 2140 176 2148 184
rect 2172 156 2180 164
rect 2300 156 2308 164
rect 2076 136 2084 144
rect 2140 136 2148 144
rect 2284 136 2292 144
rect 1852 116 1860 124
rect 2140 96 2148 104
rect 2220 96 2228 104
rect 2460 236 2468 244
rect 2524 256 2532 264
rect 2540 256 2548 264
rect 2428 176 2436 184
rect 2460 176 2468 184
rect 2508 176 2516 184
rect 2396 156 2404 164
rect 2492 136 2500 144
rect 2652 316 2660 324
rect 2796 476 2804 484
rect 2732 416 2740 424
rect 2876 396 2884 404
rect 2700 336 2708 344
rect 2764 336 2772 344
rect 2684 296 2692 304
rect 2700 296 2708 304
rect 2812 316 2820 324
rect 2780 296 2788 304
rect 2860 276 2868 284
rect 2572 256 2580 264
rect 2588 256 2596 264
rect 2636 256 2644 264
rect 2684 256 2692 264
rect 2732 256 2740 264
rect 2588 236 2596 244
rect 2556 176 2564 184
rect 2620 196 2628 204
rect 2908 416 2916 424
rect 2828 256 2836 264
rect 2876 216 2884 224
rect 2812 196 2820 204
rect 2828 196 2836 204
rect 2988 316 2996 324
rect 2956 296 2964 304
rect 2972 276 2980 284
rect 2940 256 2948 264
rect 3036 656 3044 664
rect 3068 636 3076 644
rect 3132 636 3140 644
rect 3100 616 3108 624
rect 3068 596 3076 604
rect 3052 556 3060 564
rect 3116 556 3124 564
rect 3036 496 3044 504
rect 3068 496 3076 504
rect 3196 716 3204 724
rect 3228 696 3236 704
rect 3164 636 3172 644
rect 3148 596 3156 604
rect 3212 636 3220 644
rect 3180 576 3188 584
rect 3196 576 3204 584
rect 3148 556 3156 564
rect 3180 496 3188 504
rect 3164 376 3172 384
rect 3068 336 3076 344
rect 3116 336 3124 344
rect 3228 536 3236 544
rect 3212 476 3220 484
rect 3212 336 3220 344
rect 3116 316 3124 324
rect 2988 256 2996 264
rect 2956 196 2964 204
rect 2748 176 2756 184
rect 2892 176 2900 184
rect 2924 176 2932 184
rect 2796 156 2804 164
rect 2860 156 2868 164
rect 2636 136 2644 144
rect 2668 136 2676 144
rect 2572 116 2580 124
rect 2652 116 2660 124
rect 2684 116 2692 124
rect 2716 136 2724 144
rect 2844 136 2852 144
rect 2892 136 2900 144
rect 3116 296 3124 304
rect 3068 276 3076 284
rect 3116 276 3124 284
rect 3052 256 3060 264
rect 3036 216 3044 224
rect 3164 276 3172 284
rect 3180 256 3188 264
rect 3100 156 3108 164
rect 3132 156 3140 164
rect 3164 136 3172 144
rect 3276 1076 3284 1084
rect 3308 1076 3316 1084
rect 3372 1156 3380 1164
rect 3324 1036 3332 1044
rect 3276 936 3284 944
rect 3260 896 3268 904
rect 3324 976 3332 984
rect 3548 1656 3556 1664
rect 3532 1576 3540 1584
rect 3564 1556 3572 1564
rect 3548 1436 3556 1444
rect 3548 1376 3556 1384
rect 3644 1916 3652 1924
rect 3644 1896 3652 1904
rect 3628 1876 3636 1884
rect 3676 2036 3684 2044
rect 3692 2036 3700 2044
rect 3708 1976 3716 1984
rect 3676 1936 3684 1944
rect 3788 2276 3796 2284
rect 3756 2116 3764 2124
rect 3772 2096 3780 2104
rect 3996 3296 4004 3304
rect 3980 3116 3988 3124
rect 3948 3096 3956 3104
rect 3996 3076 4004 3084
rect 3916 2916 3924 2924
rect 3980 2916 3988 2924
rect 3996 2776 4004 2784
rect 3900 2756 3908 2764
rect 3980 2756 3988 2764
rect 3900 2716 3908 2724
rect 3900 2656 3908 2664
rect 3948 2576 3956 2584
rect 4012 2696 4020 2704
rect 4060 3496 4068 3504
rect 4044 3416 4052 3424
rect 4060 3376 4068 3384
rect 4092 3876 4100 3884
rect 4156 3876 4164 3884
rect 4092 3816 4100 3824
rect 4124 3756 4132 3764
rect 4204 3916 4212 3924
rect 4188 3896 4196 3904
rect 4284 3956 4292 3964
rect 4364 3956 4372 3964
rect 4348 3876 4356 3884
rect 4364 3776 4372 3784
rect 4156 3756 4164 3764
rect 4172 3756 4180 3764
rect 4284 3756 4292 3764
rect 4348 3756 4356 3764
rect 4412 4136 4420 4144
rect 4428 4140 4436 4144
rect 4428 4136 4436 4140
rect 4604 4276 4612 4284
rect 4636 4276 4644 4284
rect 4572 4256 4580 4264
rect 4540 4216 4548 4224
rect 4556 4196 4564 4204
rect 4748 4276 4756 4284
rect 4780 4276 4788 4284
rect 4700 4256 4708 4264
rect 4556 4116 4564 4124
rect 4396 3996 4404 4004
rect 4460 3956 4468 3964
rect 4476 3936 4484 3944
rect 4396 3916 4404 3924
rect 4412 3916 4420 3924
rect 4444 3916 4452 3924
rect 4444 3896 4452 3904
rect 4460 3896 4468 3904
rect 4476 3896 4484 3904
rect 4396 3856 4404 3864
rect 4540 3876 4548 3884
rect 4140 3736 4148 3744
rect 4268 3740 4276 3744
rect 4268 3736 4276 3740
rect 4332 3716 4340 3724
rect 4092 3536 4100 3544
rect 4236 3596 4244 3604
rect 4140 3516 4148 3524
rect 4300 3516 4308 3524
rect 4380 3716 4388 3724
rect 4396 3656 4404 3664
rect 4364 3536 4372 3544
rect 4412 3536 4420 3544
rect 4380 3516 4388 3524
rect 4268 3496 4276 3504
rect 4300 3476 4308 3484
rect 4284 3456 4292 3464
rect 4444 3756 4452 3764
rect 4492 3756 4500 3764
rect 4444 3736 4452 3744
rect 4572 3856 4580 3864
rect 4668 3976 4676 3984
rect 4620 3956 4628 3964
rect 4652 3956 4660 3964
rect 4652 3936 4660 3944
rect 4620 3896 4628 3904
rect 4540 3736 4548 3744
rect 4556 3736 4564 3744
rect 4476 3656 4484 3664
rect 4444 3576 4452 3584
rect 4444 3536 4452 3544
rect 4428 3516 4436 3524
rect 4460 3516 4468 3524
rect 4444 3496 4452 3504
rect 4364 3456 4372 3464
rect 4204 3436 4212 3444
rect 4412 3436 4420 3444
rect 4108 3376 4116 3384
rect 4124 3356 4132 3364
rect 4172 3356 4180 3364
rect 4076 3176 4084 3184
rect 4044 3096 4052 3104
rect 4108 3336 4116 3344
rect 4204 3336 4212 3344
rect 4108 3316 4116 3324
rect 4188 3316 4196 3324
rect 4108 3116 4116 3124
rect 4044 3056 4052 3064
rect 4060 2918 4068 2924
rect 4060 2916 4068 2918
rect 4220 3296 4228 3304
rect 4220 3176 4228 3184
rect 4268 3356 4276 3364
rect 4252 3316 4260 3324
rect 4348 3396 4356 3404
rect 4364 3316 4372 3324
rect 4252 3296 4260 3304
rect 4284 3276 4292 3284
rect 4268 3196 4276 3204
rect 4316 3156 4324 3164
rect 4268 3136 4276 3144
rect 4300 3136 4308 3144
rect 4236 3116 4244 3124
rect 4348 3116 4356 3124
rect 4172 3096 4180 3104
rect 4236 3096 4244 3104
rect 4284 3096 4292 3104
rect 4124 2936 4132 2944
rect 4204 3076 4212 3084
rect 4204 2936 4212 2944
rect 4252 3076 4260 3084
rect 4316 3076 4324 3084
rect 4316 3056 4324 3064
rect 4252 2996 4260 3004
rect 4268 2936 4276 2944
rect 4332 2936 4340 2944
rect 4188 2916 4196 2924
rect 4252 2916 4260 2924
rect 4092 2896 4100 2904
rect 4188 2876 4196 2884
rect 4284 2876 4292 2884
rect 4076 2856 4084 2864
rect 4156 2856 4164 2864
rect 4060 2716 4068 2724
rect 4060 2656 4068 2664
rect 4044 2636 4052 2644
rect 3996 2576 4004 2584
rect 3996 2516 4004 2524
rect 3836 2316 3844 2324
rect 3884 2356 3892 2364
rect 3948 2336 3956 2344
rect 3884 2276 3892 2284
rect 3868 2236 3876 2244
rect 3932 2176 3940 2184
rect 3916 2136 3924 2144
rect 3820 2076 3828 2084
rect 3852 2076 3860 2084
rect 3836 2036 3844 2044
rect 3868 2036 3876 2044
rect 3836 2016 3844 2024
rect 3747 2006 3755 2014
rect 3757 2006 3765 2014
rect 3767 2006 3775 2014
rect 3777 2006 3785 2014
rect 3787 2006 3795 2014
rect 3797 2006 3805 2014
rect 3820 1996 3828 2004
rect 3740 1976 3748 1984
rect 3836 1956 3844 1964
rect 3820 1936 3828 1944
rect 3676 1916 3684 1924
rect 3724 1916 3732 1924
rect 3708 1896 3716 1904
rect 3692 1876 3700 1884
rect 3708 1876 3716 1884
rect 3740 1836 3748 1844
rect 3708 1816 3716 1824
rect 3740 1816 3748 1824
rect 3596 1776 3604 1784
rect 3660 1796 3668 1804
rect 3692 1796 3700 1804
rect 3644 1756 3652 1764
rect 3724 1756 3732 1764
rect 3884 1836 3892 1844
rect 3868 1756 3876 1764
rect 3820 1736 3828 1744
rect 3900 1776 3908 1784
rect 3612 1716 3620 1724
rect 3836 1716 3844 1724
rect 3852 1716 3860 1724
rect 3660 1696 3668 1704
rect 3660 1676 3668 1684
rect 3596 1596 3604 1604
rect 3820 1696 3828 1704
rect 3724 1636 3732 1644
rect 3708 1616 3716 1624
rect 3747 1606 3755 1614
rect 3757 1606 3765 1614
rect 3767 1606 3775 1614
rect 3777 1606 3785 1614
rect 3787 1606 3795 1614
rect 3797 1606 3805 1614
rect 3804 1556 3812 1564
rect 3596 1516 3604 1524
rect 3676 1516 3684 1524
rect 3724 1516 3732 1524
rect 3756 1516 3764 1524
rect 3708 1496 3716 1504
rect 3644 1476 3652 1484
rect 3580 1456 3588 1464
rect 3644 1456 3652 1464
rect 3692 1456 3700 1464
rect 3596 1376 3604 1384
rect 3532 1316 3540 1324
rect 3548 1316 3556 1324
rect 3532 1296 3540 1304
rect 3420 1116 3428 1124
rect 3500 1116 3508 1124
rect 3388 1076 3396 1084
rect 3548 1076 3556 1084
rect 3404 1056 3412 1064
rect 3420 1056 3428 1064
rect 3468 1056 3476 1064
rect 3484 1056 3492 1064
rect 3516 1056 3524 1064
rect 3388 1036 3396 1044
rect 3356 996 3364 1004
rect 3372 996 3380 1004
rect 3340 956 3348 964
rect 3260 876 3268 884
rect 3292 876 3300 884
rect 3356 876 3364 884
rect 3372 776 3380 784
rect 3292 716 3300 724
rect 3260 656 3268 664
rect 3292 676 3300 684
rect 3292 616 3300 624
rect 3276 576 3284 584
rect 3324 716 3332 724
rect 3388 716 3396 724
rect 3420 716 3428 724
rect 3340 656 3348 664
rect 3372 676 3380 684
rect 3292 556 3300 564
rect 3276 516 3284 524
rect 3356 516 3364 524
rect 3404 696 3412 704
rect 3388 636 3396 644
rect 3276 476 3284 484
rect 3244 396 3252 404
rect 3372 456 3380 464
rect 3340 376 3348 384
rect 3324 356 3332 364
rect 3260 276 3268 284
rect 3228 196 3236 204
rect 3260 136 3268 144
rect 3356 276 3364 284
rect 3356 256 3364 264
rect 3388 296 3396 304
rect 3388 276 3396 284
rect 3420 656 3428 664
rect 3436 496 3444 504
rect 3436 476 3444 484
rect 3468 716 3476 724
rect 3468 676 3476 684
rect 3580 1316 3588 1324
rect 3596 1296 3604 1304
rect 3628 1436 3636 1444
rect 3628 1356 3636 1364
rect 3676 1296 3684 1304
rect 3676 1236 3684 1244
rect 3724 1476 3732 1484
rect 3740 1456 3748 1464
rect 3820 1436 3828 1444
rect 3756 1416 3764 1424
rect 3772 1416 3780 1424
rect 3772 1376 3780 1384
rect 3788 1376 3796 1384
rect 3740 1336 3748 1344
rect 3772 1316 3780 1324
rect 3820 1356 3828 1364
rect 3788 1276 3796 1284
rect 3747 1206 3755 1214
rect 3757 1206 3765 1214
rect 3767 1206 3775 1214
rect 3777 1206 3785 1214
rect 3787 1206 3795 1214
rect 3797 1206 3805 1214
rect 3724 1196 3732 1204
rect 3724 1116 3732 1124
rect 3868 1556 3876 1564
rect 3900 1696 3908 1704
rect 3884 1496 3892 1504
rect 3868 1476 3876 1484
rect 3980 2276 3988 2284
rect 3964 1976 3972 1984
rect 3948 1856 3956 1864
rect 4028 2596 4036 2604
rect 4060 2556 4068 2564
rect 4124 2736 4132 2744
rect 4140 2716 4148 2724
rect 4092 2696 4100 2704
rect 4108 2596 4116 2604
rect 4092 2576 4100 2584
rect 4124 2516 4132 2524
rect 4108 2396 4116 2404
rect 4092 2376 4100 2384
rect 4060 2356 4068 2364
rect 4092 2336 4100 2344
rect 4220 2836 4228 2844
rect 4172 2576 4180 2584
rect 4188 2576 4196 2584
rect 4284 2816 4292 2824
rect 4476 3476 4484 3484
rect 4476 3456 4484 3464
rect 4460 3416 4468 3424
rect 4460 3356 4468 3364
rect 4444 3336 4452 3344
rect 4524 3476 4532 3484
rect 4604 3756 4612 3764
rect 4636 3880 4644 3884
rect 4636 3876 4644 3880
rect 4636 3776 4644 3784
rect 4748 4176 4756 4184
rect 4732 4116 4740 4124
rect 4732 3936 4740 3944
rect 4700 3876 4708 3884
rect 4668 3756 4676 3764
rect 4604 3496 4612 3504
rect 4588 3476 4596 3484
rect 4556 3376 4564 3384
rect 4492 3356 4500 3364
rect 4444 3316 4452 3324
rect 4460 3316 4468 3324
rect 4412 3296 4420 3304
rect 4460 3276 4468 3284
rect 4396 3156 4404 3164
rect 4396 3096 4404 3104
rect 4364 3076 4372 3084
rect 4396 3056 4404 3064
rect 4444 3096 4452 3104
rect 4444 3056 4452 3064
rect 4380 3036 4388 3044
rect 4412 3036 4420 3044
rect 4348 2776 4356 2784
rect 4332 2756 4340 2764
rect 4316 2736 4324 2744
rect 4316 2716 4324 2724
rect 4332 2716 4340 2724
rect 4428 3016 4436 3024
rect 4412 2936 4420 2944
rect 4556 3356 4564 3364
rect 4540 3336 4548 3344
rect 4524 3136 4532 3144
rect 4604 3336 4612 3344
rect 4604 3316 4612 3324
rect 4652 3536 4660 3544
rect 4700 3556 4708 3564
rect 4716 3496 4724 3504
rect 4684 3436 4692 3444
rect 4652 3416 4660 3424
rect 4668 3336 4676 3344
rect 4572 3196 4580 3204
rect 4620 3196 4628 3204
rect 4556 3136 4564 3144
rect 4492 3056 4500 3064
rect 4524 3056 4532 3064
rect 4492 3036 4500 3044
rect 4604 3156 4612 3164
rect 4620 3156 4628 3164
rect 4588 3116 4596 3124
rect 4588 2976 4596 2984
rect 4348 2696 4356 2704
rect 4236 2676 4244 2684
rect 4396 2676 4404 2684
rect 4364 2656 4372 2664
rect 4316 2616 4324 2624
rect 4220 2556 4228 2564
rect 4252 2518 4260 2524
rect 4252 2516 4260 2518
rect 4300 2496 4308 2504
rect 4380 2636 4388 2644
rect 4444 2896 4452 2904
rect 4476 2896 4484 2904
rect 4492 2896 4500 2904
rect 4428 2756 4436 2764
rect 4492 2756 4500 2764
rect 4540 2696 4548 2704
rect 4428 2616 4436 2624
rect 4428 2516 4436 2524
rect 4156 2416 4164 2424
rect 4284 2376 4292 2384
rect 4140 2316 4148 2324
rect 4284 2316 4292 2324
rect 4076 2296 4084 2304
rect 4124 2296 4132 2304
rect 4156 2276 4164 2284
rect 4156 2256 4164 2264
rect 4060 2196 4068 2204
rect 4044 2176 4052 2184
rect 4076 2156 4084 2164
rect 4012 2136 4020 2144
rect 4108 2136 4116 2144
rect 4140 2118 4148 2124
rect 4140 2116 4148 2118
rect 4140 1916 4148 1924
rect 4140 1896 4148 1904
rect 3964 1796 3972 1804
rect 3932 1756 3940 1764
rect 3948 1556 3956 1564
rect 3980 1696 3988 1704
rect 3916 1356 3924 1364
rect 3916 1316 3924 1324
rect 3964 1256 3972 1264
rect 3852 1196 3860 1204
rect 3836 1096 3844 1104
rect 3580 956 3588 964
rect 3596 956 3604 964
rect 3660 1076 3668 1084
rect 3708 1076 3716 1084
rect 3724 1056 3732 1064
rect 3644 956 3652 964
rect 3516 896 3524 904
rect 3564 876 3572 884
rect 3612 936 3620 944
rect 3628 936 3636 944
rect 3596 916 3604 924
rect 3580 836 3588 844
rect 3548 816 3556 824
rect 3580 736 3588 744
rect 3516 716 3524 724
rect 3484 576 3492 584
rect 3564 676 3572 684
rect 3548 576 3556 584
rect 3532 536 3540 544
rect 3484 516 3492 524
rect 3468 476 3476 484
rect 3708 956 3716 964
rect 3740 956 3748 964
rect 3756 956 3764 964
rect 3692 916 3700 924
rect 3724 896 3732 904
rect 3660 856 3668 864
rect 3708 816 3716 824
rect 3612 776 3620 784
rect 3868 1136 3876 1144
rect 4028 1816 4036 1824
rect 4076 1816 4084 1824
rect 4044 1776 4052 1784
rect 4060 1736 4068 1744
rect 4028 1676 4036 1684
rect 4156 1816 4164 1824
rect 4236 2256 4244 2264
rect 4188 2176 4196 2184
rect 4268 2156 4276 2164
rect 4364 2476 4372 2484
rect 4332 2336 4340 2344
rect 4348 2280 4356 2284
rect 4348 2276 4356 2280
rect 4348 2256 4356 2264
rect 4348 2236 4356 2244
rect 4300 2136 4308 2144
rect 4332 2096 4340 2104
rect 4236 2056 4244 2064
rect 4236 2036 4244 2044
rect 4204 1996 4212 2004
rect 4092 1756 4100 1764
rect 4044 1576 4052 1584
rect 4012 1476 4020 1484
rect 4028 1456 4036 1464
rect 3964 1116 3972 1124
rect 3996 1116 4004 1124
rect 3884 1096 3892 1104
rect 3820 1076 3828 1084
rect 3852 1076 3860 1084
rect 3884 1056 3892 1064
rect 3932 1076 3940 1084
rect 3916 1056 3924 1064
rect 3948 1056 3956 1064
rect 3900 1016 3908 1024
rect 3868 996 3876 1004
rect 3836 976 3844 984
rect 3772 876 3780 884
rect 3740 856 3748 864
rect 3747 806 3755 814
rect 3757 806 3765 814
rect 3767 806 3775 814
rect 3777 806 3785 814
rect 3787 806 3795 814
rect 3797 806 3805 814
rect 3724 796 3732 804
rect 3724 756 3732 764
rect 3740 756 3748 764
rect 3628 716 3636 724
rect 3676 716 3684 724
rect 3852 896 3860 904
rect 3884 896 3892 904
rect 3868 856 3876 864
rect 3852 816 3860 824
rect 3836 736 3844 744
rect 3612 656 3620 664
rect 3676 656 3684 664
rect 3708 656 3716 664
rect 3804 636 3812 644
rect 3548 496 3556 504
rect 3596 496 3604 504
rect 3532 476 3540 484
rect 3628 476 3636 484
rect 3500 436 3508 444
rect 3612 436 3620 444
rect 3708 556 3716 564
rect 3724 556 3732 564
rect 3820 556 3828 564
rect 3756 536 3764 544
rect 3708 516 3716 524
rect 3708 436 3716 444
rect 3756 436 3764 444
rect 3747 406 3755 414
rect 3757 406 3765 414
rect 3767 406 3775 414
rect 3777 406 3785 414
rect 3787 406 3795 414
rect 3797 406 3805 414
rect 3532 296 3540 304
rect 3548 296 3556 304
rect 3660 296 3668 304
rect 3468 276 3476 284
rect 3500 276 3508 284
rect 3372 216 3380 224
rect 3548 276 3556 284
rect 3580 256 3588 264
rect 3484 196 3492 204
rect 3420 176 3428 184
rect 3388 136 3396 144
rect 3420 136 3428 144
rect 3324 116 3332 124
rect 3724 276 3732 284
rect 3884 736 3892 744
rect 3980 1076 3988 1084
rect 3964 1016 3972 1024
rect 3948 816 3956 824
rect 3996 936 4004 944
rect 3980 856 3988 864
rect 3964 796 3972 804
rect 3948 736 3956 744
rect 3868 676 3876 684
rect 3932 676 3940 684
rect 3852 616 3860 624
rect 3916 636 3924 644
rect 3900 596 3908 604
rect 3964 676 3972 684
rect 3964 656 3972 664
rect 3948 556 3956 564
rect 3900 536 3908 544
rect 3852 516 3860 524
rect 3884 376 3892 384
rect 3868 356 3876 364
rect 3932 356 3940 364
rect 3900 316 3908 324
rect 3852 296 3860 304
rect 3900 296 3908 304
rect 3836 276 3844 284
rect 3644 256 3652 264
rect 3724 256 3732 264
rect 3612 236 3620 244
rect 3692 236 3700 244
rect 3676 176 3684 184
rect 3932 296 3940 304
rect 3884 256 3892 264
rect 4044 1296 4052 1304
rect 4140 1676 4148 1684
rect 4124 1636 4132 1644
rect 4108 1576 4116 1584
rect 4108 1516 4116 1524
rect 4108 1496 4116 1504
rect 4092 1476 4100 1484
rect 4172 1756 4180 1764
rect 4188 1736 4196 1744
rect 4188 1496 4196 1504
rect 4172 1456 4180 1464
rect 4108 1436 4116 1444
rect 4076 1236 4084 1244
rect 4060 1156 4068 1164
rect 4172 1396 4180 1404
rect 4124 1336 4132 1344
rect 4188 1336 4196 1344
rect 4124 1296 4132 1304
rect 4156 1296 4164 1304
rect 4236 1856 4244 1864
rect 4252 1836 4260 1844
rect 4252 1796 4260 1804
rect 4236 1716 4244 1724
rect 4284 1976 4292 1984
rect 4284 1916 4292 1924
rect 4300 1856 4308 1864
rect 4300 1836 4308 1844
rect 4332 1836 4340 1844
rect 4316 1816 4324 1824
rect 4284 1716 4292 1724
rect 4284 1696 4292 1704
rect 4268 1676 4276 1684
rect 4236 1656 4244 1664
rect 4236 1636 4244 1644
rect 4220 1616 4228 1624
rect 4220 1516 4228 1524
rect 4300 1616 4308 1624
rect 4252 1536 4260 1544
rect 4284 1536 4292 1544
rect 4268 1496 4276 1504
rect 4236 1476 4244 1484
rect 4252 1476 4260 1484
rect 4220 1356 4228 1364
rect 4220 1316 4228 1324
rect 4204 1276 4212 1284
rect 4156 1176 4164 1184
rect 4204 1176 4212 1184
rect 4060 1096 4068 1104
rect 4140 1096 4148 1104
rect 4124 1076 4132 1084
rect 4028 936 4036 944
rect 4108 936 4116 944
rect 4076 916 4084 924
rect 4092 916 4100 924
rect 4060 856 4068 864
rect 4092 776 4100 784
rect 4012 736 4020 744
rect 3996 716 4004 724
rect 4060 696 4068 704
rect 4108 736 4116 744
rect 4028 676 4036 684
rect 4060 656 4068 664
rect 3980 496 3988 504
rect 4044 596 4052 604
rect 4220 1156 4228 1164
rect 4140 1056 4148 1064
rect 4140 976 4148 984
rect 4156 936 4164 944
rect 4172 936 4180 944
rect 4140 896 4148 904
rect 4220 1016 4228 1024
rect 4300 1456 4308 1464
rect 4284 1376 4292 1384
rect 4364 1896 4372 1904
rect 4348 1576 4356 1584
rect 4396 2416 4404 2424
rect 4412 2196 4420 2204
rect 4508 2496 4516 2504
rect 4444 2336 4452 2344
rect 4492 2336 4500 2344
rect 4524 2316 4532 2324
rect 4476 2276 4484 2284
rect 4524 2256 4532 2264
rect 4540 2236 4548 2244
rect 4492 2156 4500 2164
rect 4508 2156 4516 2164
rect 4524 2136 4532 2144
rect 4460 2096 4468 2104
rect 4508 2096 4516 2104
rect 4476 2076 4484 2084
rect 4572 2876 4580 2884
rect 4572 2856 4580 2864
rect 4684 3316 4692 3324
rect 4716 3436 4724 3444
rect 4828 4156 4836 4164
rect 4860 4056 4868 4064
rect 4908 3976 4916 3984
rect 4828 3916 4836 3924
rect 4876 3916 4884 3924
rect 4940 3956 4948 3964
rect 4924 3916 4932 3924
rect 4860 3876 4868 3884
rect 4844 3856 4852 3864
rect 4796 3736 4804 3744
rect 4764 3716 4772 3724
rect 4748 3536 4756 3544
rect 4796 3536 4804 3544
rect 4796 3456 4804 3464
rect 4844 3716 4852 3724
rect 4860 3696 4868 3704
rect 4860 3636 4868 3644
rect 4828 3596 4836 3604
rect 4860 3536 4868 3544
rect 4892 3676 4900 3684
rect 4908 3516 4916 3524
rect 4828 3496 4836 3504
rect 4828 3456 4836 3464
rect 4892 3456 4900 3464
rect 4908 3456 4916 3464
rect 4732 3376 4740 3384
rect 4812 3376 4820 3384
rect 4844 3376 4852 3384
rect 4732 3336 4740 3344
rect 4780 3336 4788 3344
rect 4716 3316 4724 3324
rect 4812 3316 4820 3324
rect 4732 3276 4740 3284
rect 4828 3276 4836 3284
rect 4716 3136 4724 3144
rect 4684 3116 4692 3124
rect 4636 3036 4644 3044
rect 4716 3016 4724 3024
rect 4700 2936 4708 2944
rect 4636 2856 4644 2864
rect 4700 2856 4708 2864
rect 4588 2716 4596 2724
rect 4572 2616 4580 2624
rect 4652 2776 4660 2784
rect 4620 2756 4628 2764
rect 4636 2716 4644 2724
rect 4812 3256 4820 3264
rect 4764 3136 4772 3144
rect 4748 3116 4756 3124
rect 4748 3096 4756 3104
rect 4748 3036 4756 3044
rect 4748 2856 4756 2864
rect 4700 2716 4708 2724
rect 4668 2696 4676 2704
rect 4636 2636 4644 2644
rect 4892 3376 4900 3384
rect 4876 3336 4884 3344
rect 4860 3276 4868 3284
rect 5052 4756 5060 4764
rect 5036 4716 5044 4724
rect 5036 4656 5044 4664
rect 5036 4576 5044 4584
rect 5020 4536 5028 4544
rect 5004 4516 5012 4524
rect 5036 4516 5044 4524
rect 5020 4496 5028 4504
rect 5020 4276 5028 4284
rect 4988 4196 4996 4204
rect 4972 4176 4980 4184
rect 4972 4156 4980 4164
rect 5036 4136 5044 4144
rect 5212 4816 5220 4824
rect 5196 4756 5204 4764
rect 5148 4696 5156 4704
rect 5164 4696 5172 4704
rect 5100 4676 5108 4684
rect 5132 4656 5140 4664
rect 5132 4596 5140 4604
rect 5116 4536 5124 4544
rect 5308 4796 5316 4804
rect 5228 4696 5236 4704
rect 5212 4676 5220 4684
rect 5244 4656 5252 4664
rect 5228 4636 5236 4644
rect 5212 4616 5220 4624
rect 5164 4576 5172 4584
rect 5196 4576 5204 4584
rect 5212 4576 5220 4584
rect 5148 4536 5156 4544
rect 5251 4606 5259 4614
rect 5261 4606 5269 4614
rect 5271 4606 5279 4614
rect 5281 4606 5289 4614
rect 5291 4606 5299 4614
rect 5301 4606 5309 4614
rect 5244 4536 5252 4544
rect 5180 4516 5188 4524
rect 5260 4516 5268 4524
rect 5100 4496 5108 4504
rect 5132 4416 5140 4424
rect 5084 4336 5092 4344
rect 5164 4336 5172 4344
rect 5100 4296 5108 4304
rect 5148 4296 5156 4304
rect 5084 4276 5092 4284
rect 5132 4276 5140 4284
rect 5148 4256 5156 4264
rect 5068 4236 5076 4244
rect 5052 4116 5060 4124
rect 5100 4216 5108 4224
rect 5212 4276 5220 4284
rect 5164 4196 5172 4204
rect 5100 4136 5108 4144
rect 5244 4276 5252 4284
rect 5251 4206 5259 4214
rect 5261 4206 5269 4214
rect 5271 4206 5279 4214
rect 5281 4206 5289 4214
rect 5291 4206 5299 4214
rect 5301 4206 5309 4214
rect 5388 4916 5396 4924
rect 5484 4876 5492 4884
rect 5420 4716 5428 4724
rect 5388 4676 5396 4684
rect 5436 4656 5444 4664
rect 5388 4596 5396 4604
rect 5372 4576 5380 4584
rect 5420 4576 5428 4584
rect 5404 4516 5412 4524
rect 5340 4476 5348 4484
rect 5420 4496 5428 4504
rect 5388 4476 5396 4484
rect 5356 4396 5364 4404
rect 5228 4176 5236 4184
rect 5260 4176 5268 4184
rect 5292 4176 5300 4184
rect 5324 4176 5332 4184
rect 5228 4156 5236 4164
rect 5116 4116 5124 4124
rect 5004 4076 5012 4084
rect 5004 3976 5012 3984
rect 5036 3976 5044 3984
rect 5020 3936 5028 3944
rect 4988 3896 4996 3904
rect 5036 3896 5044 3904
rect 4956 3876 4964 3884
rect 4940 3816 4948 3824
rect 5164 4096 5172 4104
rect 5068 4076 5076 4084
rect 5068 4016 5076 4024
rect 5180 4076 5188 4084
rect 5212 4076 5220 4084
rect 5116 3936 5124 3944
rect 5084 3896 5092 3904
rect 5068 3856 5076 3864
rect 5052 3836 5060 3844
rect 5036 3776 5044 3784
rect 5100 3756 5108 3764
rect 5036 3736 5044 3744
rect 5020 3716 5028 3724
rect 5084 3716 5092 3724
rect 5068 3696 5076 3704
rect 5052 3636 5060 3644
rect 5036 3536 5044 3544
rect 5036 3516 5044 3524
rect 5068 3516 5076 3524
rect 4940 3496 4948 3504
rect 5004 3456 5012 3464
rect 5036 3456 5044 3464
rect 5196 3976 5204 3984
rect 5212 3936 5220 3944
rect 5180 3856 5188 3864
rect 5148 3756 5156 3764
rect 5228 3876 5236 3884
rect 5436 4456 5444 4464
rect 5404 4376 5412 4384
rect 5356 4256 5364 4264
rect 5340 4156 5348 4164
rect 5308 4136 5316 4144
rect 5308 4116 5316 4124
rect 5340 3936 5348 3944
rect 5372 4156 5380 4164
rect 5388 4116 5396 4124
rect 5388 3976 5396 3984
rect 5356 3896 5364 3904
rect 6732 5136 6740 5144
rect 6012 5116 6020 5124
rect 6076 5116 6084 5124
rect 6188 5116 6196 5124
rect 6220 5116 6228 5124
rect 6060 5096 6068 5104
rect 6092 5096 6100 5104
rect 5532 5076 5540 5084
rect 5580 5076 5588 5084
rect 5724 5076 5732 5084
rect 5772 5076 5780 5084
rect 5724 5056 5732 5064
rect 5644 5016 5652 5024
rect 5564 4956 5572 4964
rect 5612 4956 5620 4964
rect 5628 4936 5636 4944
rect 5596 4916 5604 4924
rect 5660 4916 5668 4924
rect 5500 4816 5508 4824
rect 5628 4896 5636 4904
rect 5564 4876 5572 4884
rect 5676 4816 5684 4824
rect 5740 5016 5748 5024
rect 5916 5076 5924 5084
rect 5852 5056 5860 5064
rect 5916 5056 5924 5064
rect 5964 5056 5972 5064
rect 6060 5076 6068 5084
rect 6076 5076 6084 5084
rect 6124 5076 6132 5084
rect 6268 5076 6276 5084
rect 5916 4996 5924 5004
rect 5980 4996 5988 5004
rect 5868 4976 5876 4984
rect 6028 5016 6036 5024
rect 6092 5056 6100 5064
rect 6092 4996 6100 5004
rect 6300 5116 6308 5124
rect 6332 5116 6340 5124
rect 6604 5096 6612 5104
rect 6332 5076 6340 5084
rect 6220 5056 6228 5064
rect 6300 5056 6308 5064
rect 6332 5056 6340 5064
rect 6380 5056 6388 5064
rect 6364 5016 6372 5024
rect 6188 4996 6196 5004
rect 6108 4976 6116 4984
rect 6188 4976 6196 4984
rect 6348 4976 6356 4984
rect 5740 4936 5748 4944
rect 5772 4936 5780 4944
rect 5804 4936 5812 4944
rect 5852 4936 5860 4944
rect 5948 4936 5956 4944
rect 6076 4936 6084 4944
rect 5708 4916 5716 4924
rect 5804 4916 5812 4924
rect 5740 4896 5748 4904
rect 5884 4856 5892 4864
rect 6060 4836 6068 4844
rect 5996 4816 6004 4824
rect 5548 4796 5556 4804
rect 5692 4796 5700 4804
rect 5996 4756 6004 4764
rect 5724 4716 5732 4724
rect 5500 4696 5508 4704
rect 5532 4696 5540 4704
rect 5548 4696 5556 4704
rect 5628 4696 5636 4704
rect 5660 4676 5668 4684
rect 5804 4716 5812 4724
rect 5980 4716 5988 4724
rect 6028 4716 6036 4724
rect 5756 4696 5764 4704
rect 5772 4696 5780 4704
rect 5836 4696 5844 4704
rect 6076 4776 6084 4784
rect 6140 4916 6148 4924
rect 6204 4916 6212 4924
rect 6284 4936 6292 4944
rect 6412 5016 6420 5024
rect 6476 5056 6484 5064
rect 6588 5056 6596 5064
rect 6460 5016 6468 5024
rect 6492 5016 6500 5024
rect 6428 4976 6436 4984
rect 6444 4976 6452 4984
rect 6364 4956 6372 4964
rect 6396 4956 6404 4964
rect 6412 4936 6420 4944
rect 6316 4916 6324 4924
rect 6364 4916 6372 4924
rect 6236 4896 6244 4904
rect 6428 4896 6436 4904
rect 6108 4696 6116 4704
rect 6220 4696 6228 4704
rect 6316 4816 6324 4824
rect 6380 4736 6388 4744
rect 5788 4676 5796 4684
rect 5900 4676 5908 4684
rect 6060 4676 6068 4684
rect 6284 4676 6292 4684
rect 5740 4656 5748 4664
rect 5564 4596 5572 4604
rect 5484 4536 5492 4544
rect 5516 4536 5524 4544
rect 5516 4516 5524 4524
rect 5612 4616 5620 4624
rect 5772 4596 5780 4604
rect 5708 4576 5716 4584
rect 5612 4536 5620 4544
rect 5932 4616 5940 4624
rect 5852 4576 5860 4584
rect 5804 4536 5812 4544
rect 5676 4516 5684 4524
rect 5660 4496 5668 4504
rect 5468 4476 5476 4484
rect 5548 4476 5556 4484
rect 5580 4476 5588 4484
rect 5644 4476 5652 4484
rect 5676 4416 5684 4424
rect 5452 4376 5460 4384
rect 5564 4376 5572 4384
rect 5436 4356 5444 4364
rect 5452 4316 5460 4324
rect 5548 4316 5556 4324
rect 5436 4236 5444 4244
rect 5420 4216 5428 4224
rect 5420 4096 5428 4104
rect 5484 4156 5492 4164
rect 5548 4156 5556 4164
rect 5500 4136 5508 4144
rect 5532 4136 5540 4144
rect 5452 4076 5460 4084
rect 5436 3916 5444 3924
rect 5404 3856 5412 3864
rect 5420 3856 5428 3864
rect 5292 3836 5300 3844
rect 5324 3836 5332 3844
rect 5251 3806 5259 3814
rect 5261 3806 5269 3814
rect 5271 3806 5279 3814
rect 5281 3806 5289 3814
rect 5291 3806 5299 3814
rect 5301 3806 5309 3814
rect 5228 3756 5236 3764
rect 5260 3756 5268 3764
rect 5212 3736 5220 3744
rect 5132 3716 5140 3724
rect 5212 3716 5220 3724
rect 5132 3696 5140 3704
rect 5116 3676 5124 3684
rect 5244 3556 5252 3564
rect 5228 3516 5236 3524
rect 5116 3456 5124 3464
rect 5052 3436 5060 3444
rect 5100 3436 5108 3444
rect 5148 3436 5156 3444
rect 5052 3396 5060 3404
rect 5228 3456 5236 3464
rect 5180 3436 5188 3444
rect 5180 3416 5188 3424
rect 5164 3376 5172 3384
rect 4940 3356 4948 3364
rect 4924 3316 4932 3324
rect 4908 3116 4916 3124
rect 4876 3036 4884 3044
rect 4844 2976 4852 2984
rect 4796 2896 4804 2904
rect 4780 2876 4788 2884
rect 4876 2976 4884 2984
rect 4988 3336 4996 3344
rect 5004 3336 5012 3344
rect 4956 3316 4964 3324
rect 5132 3336 5140 3344
rect 5084 3316 5092 3324
rect 5004 3296 5012 3304
rect 5036 3296 5044 3304
rect 5068 3256 5076 3264
rect 5036 3116 5044 3124
rect 5212 3376 5220 3384
rect 5251 3406 5259 3414
rect 5261 3406 5269 3414
rect 5271 3406 5279 3414
rect 5281 3406 5289 3414
rect 5291 3406 5299 3414
rect 5301 3406 5309 3414
rect 5276 3356 5284 3364
rect 5292 3356 5300 3364
rect 5132 3296 5140 3304
rect 5164 3296 5172 3304
rect 5196 3276 5204 3284
rect 5196 3176 5204 3184
rect 5212 3156 5220 3164
rect 5212 3136 5220 3144
rect 5020 3096 5028 3104
rect 5212 3096 5220 3104
rect 4940 2956 4948 2964
rect 4924 2896 4932 2904
rect 4908 2876 4916 2884
rect 4828 2836 4836 2844
rect 4796 2776 4804 2784
rect 4828 2776 4836 2784
rect 4764 2716 4772 2724
rect 4764 2696 4772 2704
rect 4748 2616 4756 2624
rect 4732 2596 4740 2604
rect 4684 2576 4692 2584
rect 4700 2576 4708 2584
rect 4684 2516 4692 2524
rect 4604 2436 4612 2444
rect 4620 2436 4628 2444
rect 4716 2416 4724 2424
rect 4780 2576 4788 2584
rect 4588 2376 4596 2384
rect 4764 2376 4772 2384
rect 4780 2336 4788 2344
rect 4572 2316 4580 2324
rect 4860 2836 4868 2844
rect 4972 2996 4980 3004
rect 4988 2936 4996 2944
rect 5004 2896 5012 2904
rect 4940 2876 4948 2884
rect 5004 2836 5012 2844
rect 4956 2776 4964 2784
rect 5084 3076 5092 3084
rect 5132 3076 5140 3084
rect 5132 3056 5140 3064
rect 5164 3056 5172 3064
rect 5180 3056 5188 3064
rect 5100 3036 5108 3044
rect 5148 3036 5156 3044
rect 5164 3036 5172 3044
rect 5052 2956 5060 2964
rect 5100 2956 5108 2964
rect 5116 2956 5124 2964
rect 5084 2916 5092 2924
rect 5100 2916 5108 2924
rect 5196 3016 5204 3024
rect 5260 3056 5268 3064
rect 5251 3006 5259 3014
rect 5261 3006 5269 3014
rect 5271 3006 5279 3014
rect 5281 3006 5289 3014
rect 5291 3006 5299 3014
rect 5301 3006 5309 3014
rect 5212 2956 5220 2964
rect 5276 2956 5284 2964
rect 5132 2896 5140 2904
rect 5180 2896 5188 2904
rect 5148 2816 5156 2824
rect 5164 2816 5172 2824
rect 5100 2796 5108 2804
rect 5116 2796 5124 2804
rect 5116 2756 5124 2764
rect 5100 2736 5108 2744
rect 4956 2716 4964 2724
rect 5020 2716 5028 2724
rect 5068 2716 5076 2724
rect 4844 2696 4852 2704
rect 4860 2696 4868 2704
rect 4908 2696 4916 2704
rect 4940 2696 4948 2704
rect 5036 2696 5044 2704
rect 4892 2596 4900 2604
rect 4908 2596 4916 2604
rect 4876 2576 4884 2584
rect 4940 2576 4948 2584
rect 4828 2516 4836 2524
rect 4860 2516 4868 2524
rect 4876 2496 4884 2504
rect 4908 2496 4916 2504
rect 4940 2476 4948 2484
rect 4812 2416 4820 2424
rect 4844 2416 4852 2424
rect 4924 2416 4932 2424
rect 4796 2316 4804 2324
rect 4604 2276 4612 2284
rect 4652 2256 4660 2264
rect 4572 2236 4580 2244
rect 4620 2236 4628 2244
rect 4748 2276 4756 2284
rect 4796 2276 4804 2284
rect 4572 2136 4580 2144
rect 4604 2136 4612 2144
rect 4620 2136 4628 2144
rect 4572 2116 4580 2124
rect 4652 2116 4660 2124
rect 4556 2096 4564 2104
rect 4556 1996 4564 2004
rect 4604 2096 4612 2104
rect 4604 2056 4612 2064
rect 4700 2116 4708 2124
rect 4892 2256 4900 2264
rect 4764 2216 4772 2224
rect 4748 2156 4756 2164
rect 4844 2156 4852 2164
rect 4860 2156 4868 2164
rect 4892 2156 4900 2164
rect 4780 2116 4788 2124
rect 4812 2096 4820 2104
rect 4716 2076 4724 2084
rect 4412 1916 4420 1924
rect 4700 2016 4708 2024
rect 4684 1996 4692 2004
rect 4780 1996 4788 2004
rect 4460 1916 4468 1924
rect 4492 1916 4500 1924
rect 4636 1916 4644 1924
rect 4668 1916 4676 1924
rect 4444 1896 4452 1904
rect 4556 1896 4564 1904
rect 4604 1896 4612 1904
rect 4428 1876 4436 1884
rect 4412 1856 4420 1864
rect 4428 1756 4436 1764
rect 4396 1736 4404 1744
rect 4396 1656 4404 1664
rect 4508 1836 4516 1844
rect 4492 1816 4500 1824
rect 4460 1796 4468 1804
rect 4444 1636 4452 1644
rect 4348 1516 4356 1524
rect 4380 1516 4388 1524
rect 4316 1396 4324 1404
rect 4268 1236 4276 1244
rect 4300 1236 4308 1244
rect 4332 1336 4340 1344
rect 4332 1316 4340 1324
rect 4332 1296 4340 1304
rect 4332 1236 4340 1244
rect 4316 1196 4324 1204
rect 4252 1116 4260 1124
rect 4268 1116 4276 1124
rect 4300 1096 4308 1104
rect 4380 1456 4388 1464
rect 4364 1436 4372 1444
rect 4364 1356 4372 1364
rect 4364 1296 4372 1304
rect 4348 1136 4356 1144
rect 4364 1116 4372 1124
rect 4444 1416 4452 1424
rect 4444 1356 4452 1364
rect 4492 1756 4500 1764
rect 4476 1736 4484 1744
rect 4476 1676 4484 1684
rect 4508 1536 4516 1544
rect 4508 1496 4516 1504
rect 4476 1476 4484 1484
rect 4572 1836 4580 1844
rect 4636 1796 4644 1804
rect 4540 1756 4548 1764
rect 4572 1736 4580 1744
rect 4700 1816 4708 1824
rect 4860 2116 4868 2124
rect 4908 2116 4916 2124
rect 4844 2056 4852 2064
rect 4908 1916 4916 1924
rect 4844 1856 4852 1864
rect 4748 1836 4756 1844
rect 4812 1836 4820 1844
rect 4908 1876 4916 1884
rect 4892 1856 4900 1864
rect 5052 2656 5060 2664
rect 5084 2656 5092 2664
rect 5036 2576 5044 2584
rect 4956 2396 4964 2404
rect 5180 2756 5188 2764
rect 5132 2696 5140 2704
rect 5116 2556 5124 2564
rect 5084 2516 5092 2524
rect 5132 2516 5140 2524
rect 5116 2496 5124 2504
rect 5036 2436 5044 2444
rect 4988 2376 4996 2384
rect 5004 2336 5012 2344
rect 4940 2316 4948 2324
rect 4972 2276 4980 2284
rect 4988 2256 4996 2264
rect 5116 2396 5124 2404
rect 5244 2776 5252 2784
rect 5228 2716 5236 2724
rect 5212 2676 5220 2684
rect 5180 2616 5188 2624
rect 5251 2606 5259 2614
rect 5261 2606 5269 2614
rect 5271 2606 5279 2614
rect 5281 2606 5289 2614
rect 5291 2606 5299 2614
rect 5301 2606 5309 2614
rect 5228 2596 5236 2604
rect 5228 2576 5236 2584
rect 5164 2556 5172 2564
rect 5196 2516 5204 2524
rect 5292 2516 5300 2524
rect 5212 2496 5220 2504
rect 5196 2416 5204 2424
rect 5164 2396 5172 2404
rect 5148 2356 5156 2364
rect 5276 2376 5284 2384
rect 5196 2336 5204 2344
rect 5020 2276 5028 2284
rect 5084 2276 5092 2284
rect 5004 2236 5012 2244
rect 4956 2196 4964 2204
rect 5020 2156 5028 2164
rect 4988 2116 4996 2124
rect 5004 2076 5012 2084
rect 4956 1976 4964 1984
rect 5052 2236 5060 2244
rect 5068 2216 5076 2224
rect 5228 2316 5236 2324
rect 5244 2276 5252 2284
rect 5196 2196 5204 2204
rect 5148 2156 5156 2164
rect 5132 2116 5140 2124
rect 5180 2116 5188 2124
rect 5212 2116 5220 2124
rect 5052 2096 5060 2104
rect 5116 2096 5124 2104
rect 5148 2096 5156 2104
rect 5036 2056 5044 2064
rect 5036 2016 5044 2024
rect 4972 1896 4980 1904
rect 5004 1896 5012 1904
rect 4940 1876 4948 1884
rect 4972 1856 4980 1864
rect 4988 1816 4996 1824
rect 4924 1796 4932 1804
rect 4796 1776 4804 1784
rect 4876 1776 4884 1784
rect 4924 1776 4932 1784
rect 4876 1756 4884 1764
rect 4796 1736 4804 1744
rect 4668 1716 4676 1724
rect 4844 1716 4852 1724
rect 4876 1716 4884 1724
rect 4844 1696 4852 1704
rect 4652 1676 4660 1684
rect 4588 1656 4596 1664
rect 4652 1576 4660 1584
rect 4572 1536 4580 1544
rect 4620 1536 4628 1544
rect 4684 1536 4692 1544
rect 4684 1416 4692 1424
rect 4540 1396 4548 1404
rect 4732 1636 4740 1644
rect 4748 1536 4756 1544
rect 4796 1516 4804 1524
rect 4956 1756 4964 1764
rect 5020 1716 5028 1724
rect 4972 1676 4980 1684
rect 5100 2076 5108 2084
rect 5388 3736 5396 3744
rect 5628 4256 5636 4264
rect 5676 4256 5684 4264
rect 5692 4176 5700 4184
rect 5948 4596 5956 4604
rect 5900 4516 5908 4524
rect 5868 4476 5876 4484
rect 5884 4416 5892 4424
rect 5772 4396 5780 4404
rect 5916 4396 5924 4404
rect 5724 4376 5732 4384
rect 5772 4356 5780 4364
rect 5836 4356 5844 4364
rect 5724 4316 5732 4324
rect 5644 4156 5652 4164
rect 5708 4156 5716 4164
rect 5612 4136 5620 4144
rect 5660 4136 5668 4144
rect 5644 4116 5652 4124
rect 5532 4096 5540 4104
rect 5628 4096 5636 4104
rect 5500 4056 5508 4064
rect 5484 4036 5492 4044
rect 5580 4016 5588 4024
rect 5740 4136 5748 4144
rect 5820 4316 5828 4324
rect 5852 4316 5860 4324
rect 5804 4196 5812 4204
rect 5788 4176 5796 4184
rect 5804 4156 5812 4164
rect 5692 4116 5700 4124
rect 5708 4116 5716 4124
rect 5756 4116 5764 4124
rect 5708 4096 5716 4104
rect 5740 4096 5748 4104
rect 5692 3996 5700 4004
rect 5740 3996 5748 4004
rect 5644 3976 5652 3984
rect 5836 4176 5844 4184
rect 6012 4656 6020 4664
rect 6028 4576 6036 4584
rect 6380 4656 6388 4664
rect 6188 4636 6196 4644
rect 6236 4636 6244 4644
rect 6236 4576 6244 4584
rect 6124 4556 6132 4564
rect 5996 4536 6004 4544
rect 6156 4536 6164 4544
rect 6076 4516 6084 4524
rect 6156 4516 6164 4524
rect 6188 4516 6196 4524
rect 5964 4496 5972 4504
rect 6172 4496 6180 4504
rect 6012 4476 6020 4484
rect 6076 4476 6084 4484
rect 6092 4476 6100 4484
rect 6204 4476 6212 4484
rect 5964 4376 5972 4384
rect 5948 4356 5956 4364
rect 6028 4336 6036 4344
rect 6028 4316 6036 4324
rect 6060 4316 6068 4324
rect 6012 4276 6020 4284
rect 6028 4276 6036 4284
rect 5996 4256 6004 4264
rect 6012 4236 6020 4244
rect 6012 4216 6020 4224
rect 6220 4456 6228 4464
rect 6220 4436 6228 4444
rect 6156 4336 6164 4344
rect 6140 4316 6148 4324
rect 6124 4196 6132 4204
rect 6076 4176 6084 4184
rect 6108 4176 6116 4184
rect 5820 4136 5828 4144
rect 5852 4136 5860 4144
rect 6140 4136 6148 4144
rect 5820 4116 5828 4124
rect 5868 4116 5876 4124
rect 5868 4016 5876 4024
rect 5820 3936 5828 3944
rect 5788 3916 5796 3924
rect 5500 3896 5508 3904
rect 5772 3896 5780 3904
rect 5468 3836 5476 3844
rect 5500 3836 5508 3844
rect 5516 3776 5524 3784
rect 5628 3876 5636 3884
rect 5708 3876 5716 3884
rect 5548 3856 5556 3864
rect 5580 3776 5588 3784
rect 5532 3756 5540 3764
rect 5564 3756 5572 3764
rect 5692 3856 5700 3864
rect 5724 3856 5732 3864
rect 5772 3856 5780 3864
rect 5836 3856 5844 3864
rect 5596 3736 5604 3744
rect 5660 3756 5668 3764
rect 5516 3716 5524 3724
rect 5612 3716 5620 3724
rect 5436 3696 5444 3704
rect 5740 3756 5748 3764
rect 5900 3996 5908 4004
rect 6012 4036 6020 4044
rect 6028 4036 6036 4044
rect 5884 3936 5892 3944
rect 5916 3936 5924 3944
rect 5996 3936 6004 3944
rect 5916 3836 5924 3844
rect 5980 3876 5988 3884
rect 5948 3836 5956 3844
rect 5932 3816 5940 3824
rect 5964 3776 5972 3784
rect 5948 3756 5956 3764
rect 6140 4116 6148 4124
rect 6172 4276 6180 4284
rect 6204 4276 6212 4284
rect 6188 4196 6196 4204
rect 6188 4096 6196 4104
rect 6140 3896 6148 3904
rect 6124 3876 6132 3884
rect 6012 3776 6020 3784
rect 5724 3736 5732 3744
rect 5772 3736 5780 3744
rect 5692 3716 5700 3724
rect 5868 3716 5876 3724
rect 5980 3716 5988 3724
rect 6028 3736 6036 3744
rect 6076 3736 6084 3744
rect 6028 3716 6036 3724
rect 5644 3696 5652 3704
rect 6012 3696 6020 3704
rect 5404 3496 5412 3504
rect 5340 3456 5348 3464
rect 5340 3376 5348 3384
rect 5612 3656 5620 3664
rect 5820 3656 5828 3664
rect 5500 3596 5508 3604
rect 5724 3536 5732 3544
rect 5756 3536 5764 3544
rect 5612 3496 5620 3504
rect 5420 3456 5428 3464
rect 5420 3416 5428 3424
rect 5372 3356 5380 3364
rect 5404 3356 5412 3364
rect 5404 3336 5412 3344
rect 5372 3136 5380 3144
rect 5452 3316 5460 3324
rect 6012 3556 6020 3564
rect 5948 3536 5956 3544
rect 5756 3516 5764 3524
rect 5820 3516 5828 3524
rect 5996 3516 6004 3524
rect 5548 3476 5556 3484
rect 5516 3396 5524 3404
rect 5500 3356 5508 3364
rect 5468 3296 5476 3304
rect 5484 3236 5492 3244
rect 5500 3116 5508 3124
rect 5420 3076 5428 3084
rect 5356 3036 5364 3044
rect 5356 3016 5364 3024
rect 5436 3016 5444 3024
rect 5484 3016 5492 3024
rect 5340 2956 5348 2964
rect 5372 2956 5380 2964
rect 5388 2956 5396 2964
rect 5356 2936 5364 2944
rect 5404 2936 5412 2944
rect 5372 2916 5380 2924
rect 5388 2916 5396 2924
rect 5420 2916 5428 2924
rect 5708 3456 5716 3464
rect 5788 3496 5796 3504
rect 5772 3476 5780 3484
rect 5948 3496 5956 3504
rect 5980 3496 5988 3504
rect 5932 3476 5940 3484
rect 5980 3476 5988 3484
rect 6172 3836 6180 3844
rect 6204 3836 6212 3844
rect 6188 3756 6196 3764
rect 6268 4576 6276 4584
rect 6284 4556 6292 4564
rect 6364 4556 6372 4564
rect 6284 4496 6292 4504
rect 6268 4316 6276 4324
rect 6284 4296 6292 4304
rect 6396 4576 6404 4584
rect 6492 4936 6500 4944
rect 6460 4916 6468 4924
rect 6668 5056 6676 5064
rect 6716 5056 6724 5064
rect 6700 5036 6708 5044
rect 6636 4976 6644 4984
rect 6556 4956 6564 4964
rect 6620 4956 6628 4964
rect 6636 4936 6644 4944
rect 6684 4936 6692 4944
rect 7052 5116 7060 5124
rect 7180 5116 7188 5124
rect 6828 5096 6836 5104
rect 6876 5096 6884 5104
rect 6940 5096 6948 5104
rect 7132 5096 7140 5104
rect 7164 5096 7172 5104
rect 6956 5076 6964 5084
rect 7036 5076 7044 5084
rect 7084 5076 7092 5084
rect 7308 5096 7316 5104
rect 7356 5096 7364 5104
rect 7276 5076 7284 5084
rect 7308 5076 7316 5084
rect 7324 5076 7332 5084
rect 6844 5056 6852 5064
rect 6604 4916 6612 4924
rect 6652 4916 6660 4924
rect 6700 4916 6708 4924
rect 6588 4896 6596 4904
rect 6604 4736 6612 4744
rect 6492 4716 6500 4724
rect 6556 4716 6564 4724
rect 6508 4696 6516 4704
rect 6556 4696 6564 4704
rect 6540 4676 6548 4684
rect 7004 5056 7012 5064
rect 7084 5056 7092 5064
rect 7228 5056 7236 5064
rect 6892 4956 6900 4964
rect 6940 4956 6948 4964
rect 6908 4916 6916 4924
rect 6956 4916 6964 4924
rect 6860 4896 6868 4904
rect 6755 4806 6763 4814
rect 6765 4806 6773 4814
rect 6775 4806 6783 4814
rect 6785 4806 6793 4814
rect 6795 4806 6803 4814
rect 6805 4806 6813 4814
rect 6668 4716 6676 4724
rect 6732 4716 6740 4724
rect 6844 4716 6852 4724
rect 6956 4736 6964 4744
rect 6924 4716 6932 4724
rect 6652 4696 6660 4704
rect 6716 4696 6724 4704
rect 6732 4696 6740 4704
rect 6876 4696 6884 4704
rect 6956 4696 6964 4704
rect 6620 4676 6628 4684
rect 6700 4656 6708 4664
rect 6428 4576 6436 4584
rect 6332 4536 6340 4544
rect 6396 4536 6404 4544
rect 6332 4496 6340 4504
rect 6348 4336 6356 4344
rect 6348 4316 6356 4324
rect 6380 4516 6388 4524
rect 6444 4516 6452 4524
rect 6444 4496 6452 4504
rect 6380 4456 6388 4464
rect 6348 4276 6356 4284
rect 6252 4256 6260 4264
rect 6236 4236 6244 4244
rect 6348 4216 6356 4224
rect 6252 4176 6260 4184
rect 6348 4176 6356 4184
rect 6252 4156 6260 4164
rect 6284 4136 6292 4144
rect 6300 4136 6308 4144
rect 6332 4136 6340 4144
rect 6492 4576 6500 4584
rect 6476 4556 6484 4564
rect 6476 4536 6484 4544
rect 6540 4536 6548 4544
rect 6620 4536 6628 4544
rect 6492 4496 6500 4504
rect 6460 4476 6468 4484
rect 6492 4416 6500 4424
rect 6428 4356 6436 4364
rect 6412 4256 6420 4264
rect 6380 4156 6388 4164
rect 6460 4336 6468 4344
rect 6444 4276 6452 4284
rect 6428 4116 6436 4124
rect 6284 4096 6292 4104
rect 6396 4096 6404 4104
rect 6236 3976 6244 3984
rect 6316 3996 6324 4004
rect 6284 3936 6292 3944
rect 6300 3936 6308 3944
rect 6268 3896 6276 3904
rect 6236 3876 6244 3884
rect 6252 3856 6260 3864
rect 6236 3816 6244 3824
rect 6252 3816 6260 3824
rect 6156 3736 6164 3744
rect 6220 3736 6228 3744
rect 6156 3696 6164 3704
rect 6188 3696 6196 3704
rect 6204 3696 6212 3704
rect 6140 3616 6148 3624
rect 6124 3556 6132 3564
rect 6076 3516 6084 3524
rect 6028 3476 6036 3484
rect 6044 3476 6052 3484
rect 5612 3376 5620 3384
rect 5596 3336 5604 3344
rect 5628 3336 5636 3344
rect 5580 3316 5588 3324
rect 5548 3296 5556 3304
rect 5564 3296 5572 3304
rect 5708 3336 5716 3344
rect 5660 3316 5668 3324
rect 5740 3316 5748 3324
rect 5660 3296 5668 3304
rect 5580 3216 5588 3224
rect 5596 3216 5604 3224
rect 5548 3036 5556 3044
rect 5532 2976 5540 2984
rect 5452 2956 5460 2964
rect 5564 2976 5572 2984
rect 5548 2936 5556 2944
rect 5500 2916 5508 2924
rect 5548 2916 5556 2924
rect 5516 2896 5524 2904
rect 5532 2896 5540 2904
rect 5420 2816 5428 2824
rect 5436 2816 5444 2824
rect 5404 2776 5412 2784
rect 5372 2756 5380 2764
rect 5388 2716 5396 2724
rect 5356 2596 5364 2604
rect 5372 2556 5380 2564
rect 5340 2536 5348 2544
rect 5580 2956 5588 2964
rect 5644 3116 5652 3124
rect 5724 3296 5732 3304
rect 5692 3276 5700 3284
rect 5724 3276 5732 3284
rect 5692 3096 5700 3104
rect 5628 3036 5636 3044
rect 5644 3036 5652 3044
rect 5628 2976 5636 2984
rect 5596 2936 5604 2944
rect 5580 2916 5588 2924
rect 5596 2916 5604 2924
rect 5660 2996 5668 3004
rect 5676 2956 5684 2964
rect 5708 2956 5716 2964
rect 5708 2936 5716 2944
rect 5452 2776 5460 2784
rect 5436 2756 5444 2764
rect 5436 2716 5444 2724
rect 5484 2756 5492 2764
rect 5532 2756 5540 2764
rect 5580 2756 5588 2764
rect 5596 2736 5604 2744
rect 5404 2596 5412 2604
rect 5388 2496 5396 2504
rect 5388 2396 5396 2404
rect 5340 2316 5348 2324
rect 5251 2206 5259 2214
rect 5261 2206 5269 2214
rect 5271 2206 5279 2214
rect 5281 2206 5289 2214
rect 5291 2206 5299 2214
rect 5301 2206 5309 2214
rect 5372 2276 5380 2284
rect 5340 2216 5348 2224
rect 6108 3476 6116 3484
rect 5820 3416 5828 3424
rect 5804 3376 5812 3384
rect 5788 3336 5796 3344
rect 5964 3416 5972 3424
rect 5868 3376 5876 3384
rect 5836 3356 5844 3364
rect 5772 3276 5780 3284
rect 6092 3376 6100 3384
rect 5852 3336 5860 3344
rect 5948 3340 5956 3344
rect 5948 3336 5956 3340
rect 6076 3336 6084 3344
rect 6012 3316 6020 3324
rect 6076 3316 6084 3324
rect 5788 3256 5796 3264
rect 5836 3256 5844 3264
rect 5756 3196 5764 3204
rect 5868 3196 5876 3204
rect 5756 3176 5764 3184
rect 5820 3116 5828 3124
rect 5772 3096 5780 3104
rect 5852 2996 5860 3004
rect 5836 2956 5844 2964
rect 5804 2916 5812 2924
rect 5756 2836 5764 2844
rect 5836 2816 5844 2824
rect 5852 2816 5860 2824
rect 5804 2756 5812 2764
rect 5756 2716 5764 2724
rect 5964 3136 5972 3144
rect 5980 3136 5988 3144
rect 5900 3116 5908 3124
rect 5900 3076 5908 3084
rect 6060 3176 6068 3184
rect 6060 3116 6068 3124
rect 6012 3096 6020 3104
rect 5980 3036 5988 3044
rect 5996 3036 6004 3044
rect 5932 2956 5940 2964
rect 5948 2956 5956 2964
rect 5916 2936 5924 2944
rect 6028 2956 6036 2964
rect 5980 2936 5988 2944
rect 6012 2936 6020 2944
rect 6204 3576 6212 3584
rect 6172 3536 6180 3544
rect 6156 3516 6164 3524
rect 6156 3476 6164 3484
rect 6252 3756 6260 3764
rect 6348 3916 6356 3924
rect 6444 3916 6452 3924
rect 6380 3876 6388 3884
rect 6412 3876 6420 3884
rect 6524 4456 6532 4464
rect 6572 4516 6580 4524
rect 6556 4496 6564 4504
rect 6588 4496 6596 4504
rect 6572 4476 6580 4484
rect 6668 4496 6676 4504
rect 6652 4476 6660 4484
rect 6636 4456 6644 4464
rect 6540 4416 6548 4424
rect 6588 4416 6596 4424
rect 6892 4656 6900 4664
rect 6908 4636 6916 4644
rect 6956 4636 6964 4644
rect 6764 4616 6772 4624
rect 6924 4616 6932 4624
rect 7020 5016 7028 5024
rect 7004 4956 7012 4964
rect 7244 5036 7252 5044
rect 7132 5016 7140 5024
rect 7196 5016 7204 5024
rect 7244 5016 7252 5024
rect 7196 4976 7204 4984
rect 7100 4956 7108 4964
rect 7228 4956 7236 4964
rect 7004 4936 7012 4944
rect 7052 4936 7060 4944
rect 7116 4936 7124 4944
rect 7020 4896 7028 4904
rect 7068 4916 7076 4924
rect 7148 4916 7156 4924
rect 7068 4896 7076 4904
rect 7100 4776 7108 4784
rect 7100 4736 7108 4744
rect 7052 4696 7060 4704
rect 7020 4676 7028 4684
rect 7068 4656 7076 4664
rect 6908 4536 6916 4544
rect 6748 4516 6756 4524
rect 6828 4516 6836 4524
rect 6684 4416 6692 4424
rect 6636 4376 6644 4384
rect 6524 4296 6532 4304
rect 6508 4276 6516 4284
rect 6556 4296 6564 4304
rect 6556 4256 6564 4264
rect 6476 4236 6484 4244
rect 6540 4236 6548 4244
rect 6492 4216 6500 4224
rect 6508 4196 6516 4204
rect 6540 4196 6548 4204
rect 6492 3896 6500 3904
rect 6604 4316 6612 4324
rect 6604 4236 6612 4244
rect 6572 4196 6580 4204
rect 6620 4196 6628 4204
rect 6796 4496 6804 4504
rect 6796 4476 6804 4484
rect 6755 4406 6763 4414
rect 6765 4406 6773 4414
rect 6775 4406 6783 4414
rect 6785 4406 6793 4414
rect 6795 4406 6803 4414
rect 6805 4406 6813 4414
rect 6828 4376 6836 4384
rect 6924 4516 6932 4524
rect 6956 4516 6964 4524
rect 6924 4496 6932 4504
rect 6972 4496 6980 4504
rect 6908 4476 6916 4484
rect 6940 4476 6948 4484
rect 6876 4376 6884 4384
rect 6844 4356 6852 4364
rect 6700 4316 6708 4324
rect 6764 4316 6772 4324
rect 6844 4316 6852 4324
rect 6924 4316 6932 4324
rect 6844 4296 6852 4304
rect 6716 4276 6724 4284
rect 6668 4256 6676 4264
rect 6812 4256 6820 4264
rect 6716 4136 6724 4144
rect 6508 3876 6516 3884
rect 6652 3936 6660 3944
rect 6380 3856 6388 3864
rect 6492 3856 6500 3864
rect 6556 3856 6564 3864
rect 6268 3716 6276 3724
rect 6412 3756 6420 3764
rect 6332 3716 6340 3724
rect 6396 3716 6404 3724
rect 6364 3696 6372 3704
rect 6444 3696 6452 3704
rect 6316 3656 6324 3664
rect 6252 3556 6260 3564
rect 6316 3556 6324 3564
rect 6396 3556 6404 3564
rect 6492 3816 6500 3824
rect 6476 3736 6484 3744
rect 6572 3796 6580 3804
rect 6556 3736 6564 3744
rect 6508 3716 6516 3724
rect 6572 3716 6580 3724
rect 6524 3656 6532 3664
rect 6492 3616 6500 3624
rect 6476 3576 6484 3584
rect 6268 3536 6276 3544
rect 6460 3536 6468 3544
rect 6412 3516 6420 3524
rect 6380 3436 6388 3444
rect 6300 3416 6308 3424
rect 6236 3396 6244 3404
rect 6476 3496 6484 3504
rect 6412 3476 6420 3484
rect 6428 3436 6436 3444
rect 6412 3416 6420 3424
rect 6396 3396 6404 3404
rect 6220 3376 6228 3384
rect 6268 3376 6276 3384
rect 6252 3356 6260 3364
rect 6460 3376 6468 3384
rect 6524 3496 6532 3504
rect 6524 3416 6532 3424
rect 6556 3616 6564 3624
rect 6572 3596 6580 3604
rect 6604 3776 6612 3784
rect 6604 3736 6612 3744
rect 6588 3576 6596 3584
rect 6572 3536 6580 3544
rect 6572 3516 6580 3524
rect 6556 3416 6564 3424
rect 6636 3636 6644 3644
rect 6828 4236 6836 4244
rect 6828 4196 6836 4204
rect 6860 4276 6868 4284
rect 6908 4276 6916 4284
rect 6860 4256 6868 4264
rect 6892 4236 6900 4244
rect 6860 4176 6868 4184
rect 6812 4096 6820 4104
rect 6860 4096 6868 4104
rect 6892 4116 6900 4124
rect 7068 4576 7076 4584
rect 7004 4536 7012 4544
rect 7052 4536 7060 4544
rect 6988 4476 6996 4484
rect 6988 4456 6996 4464
rect 6988 4296 6996 4304
rect 7036 4496 7044 4504
rect 7132 4716 7140 4724
rect 7196 4756 7204 4764
rect 7212 4736 7220 4744
rect 7196 4716 7204 4724
rect 7148 4696 7156 4704
rect 7180 4676 7188 4684
rect 7116 4636 7124 4644
rect 7212 4656 7220 4664
rect 7164 4636 7172 4644
rect 7148 4556 7156 4564
rect 7212 4556 7220 4564
rect 7132 4516 7140 4524
rect 7196 4536 7204 4544
rect 7212 4536 7220 4544
rect 7084 4496 7092 4504
rect 7148 4496 7156 4504
rect 7020 4436 7028 4444
rect 7052 4336 7060 4344
rect 7148 4336 7156 4344
rect 7020 4316 7028 4324
rect 7084 4296 7092 4304
rect 7052 4256 7060 4264
rect 7084 4256 7092 4264
rect 7132 4256 7140 4264
rect 7116 4196 7124 4204
rect 7020 4176 7028 4184
rect 7180 4316 7188 4324
rect 7164 4276 7172 4284
rect 7180 4196 7188 4204
rect 6940 4156 6948 4164
rect 7004 4156 7012 4164
rect 6924 4096 6932 4104
rect 6988 4096 6996 4104
rect 6732 4076 6740 4084
rect 6684 3976 6692 3984
rect 6755 4006 6763 4014
rect 6765 4006 6773 4014
rect 6775 4006 6783 4014
rect 6785 4006 6793 4014
rect 6795 4006 6803 4014
rect 6805 4006 6813 4014
rect 6748 3976 6756 3984
rect 6908 3916 6916 3924
rect 7004 3916 7012 3924
rect 6716 3896 6724 3904
rect 6892 3896 6900 3904
rect 6940 3896 6948 3904
rect 6668 3880 6676 3884
rect 6668 3876 6676 3880
rect 6684 3856 6692 3864
rect 6668 3796 6676 3804
rect 6700 3736 6708 3744
rect 6684 3716 6692 3724
rect 6668 3636 6676 3644
rect 6860 3876 6868 3884
rect 6908 3876 6916 3884
rect 6924 3876 6932 3884
rect 6748 3756 6756 3764
rect 6844 3756 6852 3764
rect 6876 3756 6884 3764
rect 6732 3736 6740 3744
rect 6924 3736 6932 3744
rect 6764 3716 6772 3724
rect 6956 3876 6964 3884
rect 6972 3856 6980 3864
rect 7052 4096 7060 4104
rect 7132 4036 7140 4044
rect 7036 3916 7044 3924
rect 7020 3896 7028 3904
rect 6988 3756 6996 3764
rect 7004 3736 7012 3744
rect 6972 3716 6980 3724
rect 6940 3696 6948 3704
rect 6755 3606 6763 3614
rect 6765 3606 6773 3614
rect 6775 3606 6783 3614
rect 6785 3606 6793 3614
rect 6795 3606 6803 3614
rect 6805 3606 6813 3614
rect 6860 3576 6868 3584
rect 6972 3616 6980 3624
rect 6892 3536 6900 3544
rect 6924 3536 6932 3544
rect 6956 3536 6964 3544
rect 6844 3516 6852 3524
rect 6892 3496 6900 3504
rect 6684 3476 6692 3484
rect 6828 3476 6836 3484
rect 6620 3456 6628 3464
rect 6652 3436 6660 3444
rect 6476 3356 6484 3364
rect 6508 3336 6516 3344
rect 6588 3376 6596 3384
rect 6604 3376 6612 3384
rect 6652 3356 6660 3364
rect 6572 3336 6580 3344
rect 6124 3316 6132 3324
rect 6524 3316 6532 3324
rect 6300 3296 6308 3304
rect 6444 3296 6452 3304
rect 6524 3296 6532 3304
rect 6108 3276 6116 3284
rect 6332 3216 6340 3224
rect 6332 3176 6340 3184
rect 6220 3156 6228 3164
rect 6364 3156 6372 3164
rect 6380 3156 6388 3164
rect 6268 3116 6276 3124
rect 6396 3136 6404 3144
rect 6428 3136 6436 3144
rect 6540 3276 6548 3284
rect 6556 3216 6564 3224
rect 6460 3136 6468 3144
rect 6316 3096 6324 3104
rect 6444 3096 6452 3104
rect 6540 3096 6548 3104
rect 6108 3076 6116 3084
rect 6124 3076 6132 3084
rect 6076 3056 6084 3064
rect 5996 2916 6004 2924
rect 6156 2956 6164 2964
rect 6172 2936 6180 2944
rect 5868 2756 5876 2764
rect 5724 2696 5732 2704
rect 5756 2696 5764 2704
rect 5788 2696 5796 2704
rect 5852 2696 5860 2704
rect 6204 2876 6212 2884
rect 5980 2776 5988 2784
rect 6300 3076 6308 3084
rect 6364 3056 6372 3064
rect 6300 2996 6308 3004
rect 6284 2956 6292 2964
rect 6284 2936 6292 2944
rect 6300 2896 6308 2904
rect 6316 2816 6324 2824
rect 6204 2756 6212 2764
rect 6060 2736 6068 2744
rect 6172 2736 6180 2744
rect 6044 2716 6052 2724
rect 5996 2696 6004 2704
rect 6124 2696 6132 2704
rect 5452 2656 5460 2664
rect 5500 2656 5508 2664
rect 5436 2596 5444 2604
rect 5468 2556 5476 2564
rect 5436 2516 5444 2524
rect 5436 2456 5444 2464
rect 5420 2436 5428 2444
rect 5420 2416 5428 2424
rect 5404 2376 5412 2384
rect 5404 2336 5412 2344
rect 5452 2416 5460 2424
rect 5452 2396 5460 2404
rect 5564 2636 5572 2644
rect 5548 2616 5556 2624
rect 5580 2616 5588 2624
rect 5564 2596 5572 2604
rect 5644 2636 5652 2644
rect 5612 2576 5620 2584
rect 5628 2576 5636 2584
rect 5548 2536 5556 2544
rect 5516 2356 5524 2364
rect 5532 2356 5540 2364
rect 5420 2316 5428 2324
rect 5500 2316 5508 2324
rect 5532 2316 5540 2324
rect 5436 2276 5444 2284
rect 5436 2256 5444 2264
rect 5404 2236 5412 2244
rect 5292 2156 5300 2164
rect 5356 2176 5364 2184
rect 5388 2176 5396 2184
rect 5404 2156 5412 2164
rect 5276 2136 5284 2144
rect 5388 2136 5396 2144
rect 5340 2116 5348 2124
rect 5276 2096 5284 2104
rect 5548 2216 5556 2224
rect 5484 2176 5492 2184
rect 5452 2136 5460 2144
rect 5580 2456 5588 2464
rect 5596 2236 5604 2244
rect 5596 2176 5604 2184
rect 5612 2176 5620 2184
rect 5788 2656 5796 2664
rect 5676 2636 5684 2644
rect 5724 2636 5732 2644
rect 5740 2576 5748 2584
rect 5756 2576 5764 2584
rect 5660 2556 5668 2564
rect 5676 2516 5684 2524
rect 5772 2416 5780 2424
rect 5644 2356 5652 2364
rect 5676 2316 5684 2324
rect 5708 2316 5716 2324
rect 5660 2256 5668 2264
rect 5708 2256 5716 2264
rect 5676 2236 5684 2244
rect 5724 2236 5732 2244
rect 5772 2256 5780 2264
rect 5756 2196 5764 2204
rect 5660 2176 5668 2184
rect 5756 2176 5764 2184
rect 5628 2156 5636 2164
rect 5500 2116 5508 2124
rect 5340 2056 5348 2064
rect 5468 2036 5476 2044
rect 5148 2016 5156 2024
rect 5228 2016 5236 2024
rect 5068 1916 5076 1924
rect 5340 1916 5348 1924
rect 5532 1916 5540 1924
rect 5052 1896 5060 1904
rect 5052 1836 5060 1844
rect 4892 1576 4900 1584
rect 4988 1656 4996 1664
rect 4940 1516 4948 1524
rect 4876 1496 4884 1504
rect 4924 1476 4932 1484
rect 4780 1416 4788 1424
rect 4764 1396 4772 1404
rect 4540 1376 4548 1384
rect 4716 1376 4724 1384
rect 4732 1376 4740 1384
rect 4588 1356 4596 1364
rect 4700 1356 4708 1364
rect 4492 1336 4500 1344
rect 4556 1336 4564 1344
rect 4572 1336 4580 1344
rect 4636 1336 4644 1344
rect 4460 1316 4468 1324
rect 4412 1256 4420 1264
rect 4460 1276 4468 1284
rect 4428 1236 4436 1244
rect 4412 1116 4420 1124
rect 4396 1096 4404 1104
rect 4604 1316 4612 1324
rect 4652 1296 4660 1304
rect 4908 1416 4916 1424
rect 4844 1356 4852 1364
rect 4828 1336 4836 1344
rect 4860 1336 4868 1344
rect 4732 1316 4740 1324
rect 4828 1316 4836 1324
rect 4700 1276 4708 1284
rect 4604 1236 4612 1244
rect 4732 1176 4740 1184
rect 4684 1116 4692 1124
rect 4812 1116 4820 1124
rect 4828 1096 4836 1104
rect 4972 1376 4980 1384
rect 4956 1356 4964 1364
rect 4988 1356 4996 1364
rect 5036 1516 5044 1524
rect 5116 1876 5124 1884
rect 5372 1876 5380 1884
rect 5164 1836 5172 1844
rect 5100 1816 5108 1824
rect 5068 1516 5076 1524
rect 5052 1476 5060 1484
rect 5116 1736 5124 1744
rect 5148 1716 5156 1724
rect 5132 1676 5140 1684
rect 5116 1576 5124 1584
rect 5468 1896 5476 1904
rect 5516 1876 5524 1884
rect 5436 1856 5444 1864
rect 5212 1816 5220 1824
rect 5251 1806 5259 1814
rect 5261 1806 5269 1814
rect 5271 1806 5279 1814
rect 5281 1806 5289 1814
rect 5291 1806 5299 1814
rect 5301 1806 5309 1814
rect 5212 1796 5220 1804
rect 5324 1796 5332 1804
rect 5404 1796 5412 1804
rect 5468 1796 5476 1804
rect 5164 1696 5172 1704
rect 5196 1656 5204 1664
rect 5180 1576 5188 1584
rect 5148 1516 5156 1524
rect 5100 1416 5108 1424
rect 5372 1776 5380 1784
rect 5436 1776 5444 1784
rect 5228 1756 5236 1764
rect 5324 1756 5332 1764
rect 5356 1756 5364 1764
rect 5420 1756 5428 1764
rect 5452 1736 5460 1744
rect 5436 1716 5444 1724
rect 5500 1716 5508 1724
rect 5612 2116 5620 2124
rect 5660 2116 5668 2124
rect 5708 2116 5716 2124
rect 5788 2116 5796 2124
rect 5692 1896 5700 1904
rect 5676 1856 5684 1864
rect 5612 1836 5620 1844
rect 5596 1816 5604 1824
rect 5628 1796 5636 1804
rect 5548 1776 5556 1784
rect 5580 1776 5588 1784
rect 5564 1716 5572 1724
rect 5644 1716 5652 1724
rect 5676 1716 5684 1724
rect 5404 1696 5412 1704
rect 5436 1696 5444 1704
rect 5452 1696 5460 1704
rect 5532 1696 5540 1704
rect 5388 1676 5396 1684
rect 5484 1676 5492 1684
rect 5516 1676 5524 1684
rect 5244 1656 5252 1664
rect 5596 1696 5604 1704
rect 5500 1616 5508 1624
rect 5516 1616 5524 1624
rect 5548 1616 5556 1624
rect 5228 1596 5236 1604
rect 5260 1576 5268 1584
rect 5404 1576 5412 1584
rect 5228 1516 5236 1524
rect 5372 1516 5380 1524
rect 5500 1516 5508 1524
rect 5356 1496 5364 1504
rect 5324 1476 5332 1484
rect 5180 1376 5188 1384
rect 5116 1356 5124 1364
rect 5196 1356 5204 1364
rect 4988 1336 4996 1344
rect 5020 1336 5028 1344
rect 4940 1296 4948 1304
rect 5020 1316 5028 1324
rect 5036 1316 5044 1324
rect 5164 1316 5172 1324
rect 5004 1216 5012 1224
rect 5116 1296 5124 1304
rect 5148 1296 5156 1304
rect 5052 1216 5060 1224
rect 5212 1216 5220 1224
rect 5068 1176 5076 1184
rect 5020 1136 5028 1144
rect 4876 1116 4884 1124
rect 4316 1076 4324 1084
rect 4380 1076 4388 1084
rect 4412 1076 4420 1084
rect 4428 1076 4436 1084
rect 4460 1076 4468 1084
rect 4508 1076 4516 1084
rect 4652 1076 4660 1084
rect 4844 1076 4852 1084
rect 4252 936 4260 944
rect 4332 1056 4340 1064
rect 4332 976 4340 984
rect 4316 956 4324 964
rect 4620 1056 4628 1064
rect 4860 1056 4868 1064
rect 4748 1016 4756 1024
rect 4716 996 4724 1004
rect 4652 976 4660 984
rect 4364 956 4372 964
rect 4412 956 4420 964
rect 4332 936 4340 944
rect 4284 856 4292 864
rect 4252 816 4260 824
rect 4316 816 4324 824
rect 4796 976 4804 984
rect 4780 956 4788 964
rect 4444 936 4452 944
rect 4508 936 4516 944
rect 4700 936 4708 944
rect 4780 936 4788 944
rect 4396 856 4404 864
rect 4204 736 4212 744
rect 4124 616 4132 624
rect 4188 616 4196 624
rect 4236 756 4244 764
rect 4220 716 4228 724
rect 4348 796 4356 804
rect 4268 696 4276 704
rect 4316 696 4324 704
rect 4284 676 4292 684
rect 4220 596 4228 604
rect 3996 336 4004 344
rect 3980 316 3988 324
rect 3964 296 3972 304
rect 3948 156 3956 164
rect 2332 96 2340 104
rect 2700 96 2708 104
rect 2732 96 2740 104
rect 3996 136 4004 144
rect 4076 496 4084 504
rect 4204 496 4212 504
rect 4108 476 4116 484
rect 4172 476 4180 484
rect 4092 456 4100 464
rect 4028 436 4036 444
rect 4108 436 4116 444
rect 4124 436 4132 444
rect 4172 356 4180 364
rect 4092 296 4100 304
rect 4044 156 4052 164
rect 4060 136 4068 144
rect 4140 276 4148 284
rect 4220 276 4228 284
rect 4124 236 4132 244
rect 4188 236 4196 244
rect 4252 516 4260 524
rect 4332 636 4340 644
rect 4364 756 4372 764
rect 4476 856 4484 864
rect 4428 796 4436 804
rect 4396 776 4404 784
rect 4444 736 4452 744
rect 4380 716 4388 724
rect 4412 696 4420 704
rect 4492 756 4500 764
rect 4860 956 4868 964
rect 4700 896 4708 904
rect 4700 876 4708 884
rect 4652 816 4660 824
rect 4668 796 4676 804
rect 4636 776 4644 784
rect 4604 756 4612 764
rect 4812 876 4820 884
rect 4732 816 4740 824
rect 4860 916 4868 924
rect 5036 1116 5044 1124
rect 5196 1136 5204 1144
rect 5212 1136 5220 1144
rect 5132 1096 5140 1104
rect 4924 1076 4932 1084
rect 5084 1076 5092 1084
rect 5212 1056 5220 1064
rect 4924 1016 4932 1024
rect 5148 1016 5156 1024
rect 5116 956 5124 964
rect 4892 816 4900 824
rect 4828 796 4836 804
rect 4908 796 4916 804
rect 4764 776 4772 784
rect 4780 776 4788 784
rect 4844 776 4852 784
rect 4716 736 4724 744
rect 4604 696 4612 704
rect 4636 696 4644 704
rect 4652 676 4660 684
rect 4364 656 4372 664
rect 4476 656 4484 664
rect 4380 636 4388 644
rect 4396 536 4404 544
rect 4316 516 4324 524
rect 4348 516 4356 524
rect 4300 456 4308 464
rect 4268 436 4276 444
rect 4300 416 4308 424
rect 4252 276 4260 284
rect 4268 216 4276 224
rect 4188 196 4196 204
rect 4236 196 4244 204
rect 4172 156 4180 164
rect 4076 116 4084 124
rect 4284 116 4292 124
rect 4476 496 4484 504
rect 4540 496 4548 504
rect 4428 476 4436 484
rect 4492 476 4500 484
rect 4476 456 4484 464
rect 4412 376 4420 384
rect 4332 356 4340 364
rect 4572 376 4580 384
rect 4620 376 4628 384
rect 4508 336 4516 344
rect 4428 322 4436 324
rect 4428 316 4436 322
rect 4476 316 4484 324
rect 4396 296 4404 304
rect 4380 276 4388 284
rect 4380 256 4388 264
rect 4444 236 4452 244
rect 4460 216 4468 224
rect 4364 156 4372 164
rect 4380 156 4388 164
rect 4444 156 4452 164
rect 4348 136 4356 144
rect 4364 116 4372 124
rect 1692 76 1700 84
rect 1756 76 1764 84
rect 1964 76 1972 84
rect 2092 76 2100 84
rect 2252 76 2260 84
rect 2316 76 2324 84
rect 4348 76 4356 84
rect 4412 76 4420 84
rect 4492 296 4500 304
rect 4540 296 4548 304
rect 4540 256 4548 264
rect 4556 256 4564 264
rect 4588 236 4596 244
rect 4636 336 4644 344
rect 4716 696 4724 704
rect 4796 716 4804 724
rect 4828 696 4836 704
rect 5084 936 5092 944
rect 5148 936 5156 944
rect 4940 916 4948 924
rect 4860 736 4868 744
rect 4812 656 4820 664
rect 4684 636 4692 644
rect 4732 636 4740 644
rect 4764 636 4772 644
rect 4684 576 4692 584
rect 4668 556 4676 564
rect 4732 536 4740 544
rect 4684 516 4692 524
rect 4668 376 4676 384
rect 4700 336 4708 344
rect 4812 496 4820 504
rect 4892 616 4900 624
rect 5020 756 5028 764
rect 4924 736 4932 744
rect 5116 916 5124 924
rect 5180 918 5188 924
rect 5180 916 5188 918
rect 4988 716 4996 724
rect 5020 716 5028 724
rect 4924 656 4932 664
rect 4876 496 4884 504
rect 4892 476 4900 484
rect 4844 416 4852 424
rect 4876 416 4884 424
rect 4796 356 4804 364
rect 4652 316 4660 324
rect 4732 316 4740 324
rect 4748 316 4756 324
rect 4796 316 4804 324
rect 4636 296 4644 304
rect 4700 296 4708 304
rect 4700 256 4708 264
rect 4668 236 4676 244
rect 4748 296 4756 304
rect 4828 296 4836 304
rect 4812 276 4820 284
rect 4732 176 4740 184
rect 4668 156 4676 164
rect 4476 136 4484 144
rect 4524 136 4532 144
rect 4540 136 4548 144
rect 4668 136 4676 144
rect 4732 136 4740 144
rect 4956 676 4964 684
rect 5036 676 5044 684
rect 5004 636 5012 644
rect 5036 616 5044 624
rect 5052 616 5060 624
rect 4972 536 4980 544
rect 4988 536 4996 544
rect 5020 536 5028 544
rect 4940 456 4948 464
rect 4940 436 4948 444
rect 4924 396 4932 404
rect 4908 356 4916 364
rect 4908 296 4916 304
rect 4924 276 4932 284
rect 4924 256 4932 264
rect 5068 556 5076 564
rect 5100 716 5108 724
rect 5196 716 5204 724
rect 5100 676 5108 684
rect 5164 676 5172 684
rect 5251 1406 5259 1414
rect 5261 1406 5269 1414
rect 5271 1406 5279 1414
rect 5281 1406 5289 1414
rect 5291 1406 5299 1414
rect 5301 1406 5309 1414
rect 5500 1476 5508 1484
rect 5420 1456 5428 1464
rect 5596 1596 5604 1604
rect 5564 1516 5572 1524
rect 5676 1696 5684 1704
rect 5692 1636 5700 1644
rect 5644 1556 5652 1564
rect 5612 1516 5620 1524
rect 5532 1496 5540 1504
rect 5548 1476 5556 1484
rect 5388 1436 5396 1444
rect 5420 1436 5428 1444
rect 5388 1376 5396 1384
rect 5308 1316 5316 1324
rect 5356 1276 5364 1284
rect 5404 1316 5412 1324
rect 5484 1356 5492 1364
rect 5564 1356 5572 1364
rect 5532 1336 5540 1344
rect 5628 1336 5636 1344
rect 5436 1316 5444 1324
rect 5452 1316 5460 1324
rect 5580 1316 5588 1324
rect 5404 1236 5412 1244
rect 5372 1216 5380 1224
rect 5340 1176 5348 1184
rect 5356 1176 5364 1184
rect 5244 1096 5252 1104
rect 5292 1076 5300 1084
rect 5251 1006 5259 1014
rect 5261 1006 5269 1014
rect 5271 1006 5279 1014
rect 5281 1006 5289 1014
rect 5291 1006 5299 1014
rect 5301 1006 5309 1014
rect 5244 976 5252 984
rect 5340 836 5348 844
rect 5228 756 5236 764
rect 5308 716 5316 724
rect 5340 796 5348 804
rect 5356 756 5364 764
rect 5324 696 5332 704
rect 5212 656 5220 664
rect 5116 636 5124 644
rect 5164 616 5172 624
rect 5116 556 5124 564
rect 5148 556 5156 564
rect 5084 516 5092 524
rect 5052 476 5060 484
rect 5020 336 5028 344
rect 5052 336 5060 344
rect 5004 316 5012 324
rect 5148 536 5156 544
rect 5164 536 5172 544
rect 5180 516 5188 524
rect 5212 596 5220 604
rect 5251 606 5259 614
rect 5261 606 5269 614
rect 5271 606 5279 614
rect 5281 606 5289 614
rect 5291 606 5299 614
rect 5301 606 5309 614
rect 5228 576 5236 584
rect 5308 576 5316 584
rect 5436 1196 5444 1204
rect 5580 1276 5588 1284
rect 5612 1256 5620 1264
rect 5612 1196 5620 1204
rect 5468 1116 5476 1124
rect 5628 1136 5636 1144
rect 5500 1096 5508 1104
rect 5420 1076 5428 1084
rect 5420 1056 5428 1064
rect 5452 996 5460 1004
rect 5436 936 5444 944
rect 5596 1016 5604 1024
rect 5516 996 5524 1004
rect 5612 976 5620 984
rect 5468 916 5476 924
rect 5436 896 5444 904
rect 5452 856 5460 864
rect 5500 776 5508 784
rect 5628 916 5636 924
rect 5612 896 5620 904
rect 5564 736 5572 744
rect 5788 2016 5796 2024
rect 5820 2636 5828 2644
rect 5884 2616 5892 2624
rect 5900 2616 5908 2624
rect 5836 2556 5844 2564
rect 5948 2656 5956 2664
rect 5980 2636 5988 2644
rect 6252 2736 6260 2744
rect 6348 2716 6356 2724
rect 6236 2696 6244 2704
rect 6332 2696 6340 2704
rect 6396 2916 6404 2924
rect 6620 3316 6628 3324
rect 6588 3296 6596 3304
rect 6572 3096 6580 3104
rect 6476 3076 6484 3084
rect 6572 3076 6580 3084
rect 6460 3036 6468 3044
rect 6460 2936 6468 2944
rect 6524 2976 6532 2984
rect 6492 2956 6500 2964
rect 6508 2916 6516 2924
rect 6572 2956 6580 2964
rect 6572 2936 6580 2944
rect 6556 2896 6564 2904
rect 6636 3216 6644 3224
rect 6700 3416 6708 3424
rect 6716 3376 6724 3384
rect 6748 3376 6756 3384
rect 6620 3176 6628 3184
rect 6636 3176 6644 3184
rect 6684 3176 6692 3184
rect 6652 3116 6660 3124
rect 6604 3076 6612 3084
rect 6620 3076 6628 3084
rect 6620 3016 6628 3024
rect 6652 3016 6660 3024
rect 6684 3016 6692 3024
rect 6604 2956 6612 2964
rect 6636 2956 6644 2964
rect 6604 2936 6612 2944
rect 6588 2876 6596 2884
rect 6476 2836 6484 2844
rect 6572 2836 6580 2844
rect 6428 2776 6436 2784
rect 6076 2656 6084 2664
rect 6172 2656 6180 2664
rect 6380 2656 6388 2664
rect 6012 2616 6020 2624
rect 6044 2616 6052 2624
rect 5948 2536 5956 2544
rect 6028 2536 6036 2544
rect 5932 2516 5940 2524
rect 6028 2496 6036 2504
rect 5980 2336 5988 2344
rect 5900 2316 5908 2324
rect 5932 2316 5940 2324
rect 5820 2296 5828 2304
rect 5916 2276 5924 2284
rect 5852 2256 5860 2264
rect 5948 2256 5956 2264
rect 5996 2256 6004 2264
rect 5820 2236 5828 2244
rect 5868 2216 5876 2224
rect 5996 2236 6004 2244
rect 5964 2196 5972 2204
rect 6028 2236 6036 2244
rect 6012 2176 6020 2184
rect 6012 2156 6020 2164
rect 5852 2136 5860 2144
rect 5900 2136 5908 2144
rect 5836 2036 5844 2044
rect 5804 1936 5812 1944
rect 5740 1916 5748 1924
rect 6108 2576 6116 2584
rect 6156 2576 6164 2584
rect 6076 2556 6084 2564
rect 6156 2556 6164 2564
rect 6124 2536 6132 2544
rect 6220 2636 6228 2644
rect 6284 2636 6292 2644
rect 6204 2616 6212 2624
rect 6156 2516 6164 2524
rect 6236 2516 6244 2524
rect 6252 2516 6260 2524
rect 6268 2516 6276 2524
rect 6284 2496 6292 2504
rect 6428 2716 6436 2724
rect 6412 2696 6420 2704
rect 6444 2696 6452 2704
rect 6428 2676 6436 2684
rect 6412 2616 6420 2624
rect 6380 2536 6388 2544
rect 6460 2616 6468 2624
rect 6540 2816 6548 2824
rect 6684 2976 6692 2984
rect 6684 2956 6692 2964
rect 6956 3496 6964 3504
rect 6956 3476 6964 3484
rect 6876 3416 6884 3424
rect 6908 3356 6916 3364
rect 6940 3356 6948 3364
rect 6940 3336 6948 3344
rect 6764 3236 6772 3244
rect 6940 3216 6948 3224
rect 6755 3206 6763 3214
rect 6765 3206 6773 3214
rect 6775 3206 6783 3214
rect 6785 3206 6793 3214
rect 6795 3206 6803 3214
rect 6805 3206 6813 3214
rect 6908 3196 6916 3204
rect 6716 3056 6724 3064
rect 6716 3036 6724 3044
rect 6732 3036 6740 3044
rect 6860 3136 6868 3144
rect 7100 3936 7108 3944
rect 7164 3916 7172 3924
rect 7180 3916 7188 3924
rect 7100 3896 7108 3904
rect 7148 3896 7156 3904
rect 7052 3736 7060 3744
rect 7036 3716 7044 3724
rect 7324 5056 7332 5064
rect 7404 5056 7412 5064
rect 7388 5016 7396 5024
rect 7340 4976 7348 4984
rect 7244 4736 7252 4744
rect 7276 4736 7284 4744
rect 7260 4696 7268 4704
rect 7276 4676 7284 4684
rect 7388 4876 7396 4884
rect 7356 4716 7364 4724
rect 7372 4676 7380 4684
rect 7324 4656 7332 4664
rect 7340 4656 7348 4664
rect 7244 4576 7252 4584
rect 7372 4576 7380 4584
rect 7308 4556 7316 4564
rect 7356 4556 7364 4564
rect 7260 4536 7268 4544
rect 7308 4536 7316 4544
rect 7308 4516 7316 4524
rect 7292 4336 7300 4344
rect 7228 4316 7236 4324
rect 7276 4316 7284 4324
rect 7340 4296 7348 4304
rect 7228 4276 7236 4284
rect 7260 4276 7268 4284
rect 7292 4276 7300 4284
rect 7372 4276 7380 4284
rect 7212 4116 7220 4124
rect 7276 4196 7284 4204
rect 7340 4196 7348 4204
rect 7340 4176 7348 4184
rect 7372 4176 7380 4184
rect 7244 4156 7252 4164
rect 7308 4156 7316 4164
rect 7292 4116 7300 4124
rect 7228 4036 7236 4044
rect 7164 3876 7172 3884
rect 7196 3876 7204 3884
rect 7212 3876 7220 3884
rect 7196 3776 7204 3784
rect 7212 3676 7220 3684
rect 7100 3636 7108 3644
rect 7148 3636 7156 3644
rect 7020 3576 7028 3584
rect 7180 3576 7188 3584
rect 7068 3496 7076 3504
rect 7068 3476 7076 3484
rect 6924 3176 6932 3184
rect 6956 3176 6964 3184
rect 6972 3176 6980 3184
rect 6748 3016 6756 3024
rect 6828 3036 6836 3044
rect 6796 2976 6804 2984
rect 6844 2976 6852 2984
rect 6700 2936 6708 2944
rect 6620 2896 6628 2904
rect 6508 2776 6516 2784
rect 6604 2776 6612 2784
rect 6492 2656 6500 2664
rect 6460 2576 6468 2584
rect 6476 2576 6484 2584
rect 6332 2516 6340 2524
rect 6348 2456 6356 2464
rect 6124 2436 6132 2444
rect 6060 2316 6068 2324
rect 6108 2256 6116 2264
rect 6092 2196 6100 2204
rect 6076 2136 6084 2144
rect 5900 2116 5908 2124
rect 5964 2116 5972 2124
rect 6044 2116 6052 2124
rect 5884 2056 5892 2064
rect 5852 1956 5860 1964
rect 6076 2096 6084 2104
rect 6108 2076 6116 2084
rect 6060 2016 6068 2024
rect 5996 1956 6004 1964
rect 6060 1956 6068 1964
rect 5884 1936 5892 1944
rect 6044 1936 6052 1944
rect 5740 1896 5748 1904
rect 5804 1896 5812 1904
rect 5836 1896 5844 1904
rect 5932 1896 5940 1904
rect 5964 1896 5972 1904
rect 5724 1716 5732 1724
rect 5756 1876 5764 1884
rect 5772 1856 5780 1864
rect 6092 1896 6100 1904
rect 5916 1876 5924 1884
rect 5852 1816 5860 1824
rect 5804 1736 5812 1744
rect 6172 2356 6180 2364
rect 6252 2356 6260 2364
rect 6156 2336 6164 2344
rect 6460 2516 6468 2524
rect 6492 2516 6500 2524
rect 6444 2436 6452 2444
rect 6588 2736 6596 2744
rect 6604 2716 6612 2724
rect 6588 2656 6596 2664
rect 6540 2616 6548 2624
rect 6524 2596 6532 2604
rect 6572 2576 6580 2584
rect 6572 2536 6580 2544
rect 6828 2936 6836 2944
rect 6748 2916 6756 2924
rect 6716 2876 6724 2884
rect 6684 2816 6692 2824
rect 6636 2796 6644 2804
rect 6700 2776 6708 2784
rect 6636 2736 6644 2744
rect 6700 2696 6708 2704
rect 6755 2806 6763 2814
rect 6765 2806 6773 2814
rect 6775 2806 6783 2814
rect 6785 2806 6793 2814
rect 6795 2806 6803 2814
rect 6805 2806 6813 2814
rect 6780 2696 6788 2704
rect 6732 2676 6740 2684
rect 6652 2636 6660 2644
rect 6684 2576 6692 2584
rect 6620 2536 6628 2544
rect 6556 2476 6564 2484
rect 6604 2476 6612 2484
rect 6508 2416 6516 2424
rect 6540 2396 6548 2404
rect 6364 2336 6372 2344
rect 6252 2316 6260 2324
rect 6348 2316 6356 2324
rect 6460 2316 6468 2324
rect 6188 2296 6196 2304
rect 6476 2296 6484 2304
rect 6540 2296 6548 2304
rect 6284 2276 6292 2284
rect 6428 2276 6436 2284
rect 6476 2276 6484 2284
rect 6508 2276 6516 2284
rect 6236 2236 6244 2244
rect 6156 2216 6164 2224
rect 6236 2216 6244 2224
rect 6252 2216 6260 2224
rect 6332 2256 6340 2264
rect 6444 2256 6452 2264
rect 6412 2236 6420 2244
rect 6380 2216 6388 2224
rect 6188 2156 6196 2164
rect 6236 2156 6244 2164
rect 6316 2156 6324 2164
rect 6220 2056 6228 2064
rect 6396 2196 6404 2204
rect 6428 2156 6436 2164
rect 6460 2156 6468 2164
rect 6524 2156 6532 2164
rect 6268 2116 6276 2124
rect 6316 2116 6324 2124
rect 6252 2056 6260 2064
rect 6380 2096 6388 2104
rect 6332 2056 6340 2064
rect 6396 2016 6404 2024
rect 6476 2136 6484 2144
rect 6476 2116 6484 2124
rect 6620 2376 6628 2384
rect 6572 2356 6580 2364
rect 6812 2656 6820 2664
rect 6860 2876 6868 2884
rect 6844 2856 6852 2864
rect 6940 3136 6948 3144
rect 6972 3136 6980 3144
rect 7132 3476 7140 3484
rect 7164 3476 7172 3484
rect 7052 3336 7060 3344
rect 7052 3316 7060 3324
rect 7164 3416 7172 3424
rect 7244 3936 7252 3944
rect 7260 3916 7268 3924
rect 7276 3876 7284 3884
rect 7260 3796 7268 3804
rect 7356 4136 7364 4144
rect 7372 4116 7380 4124
rect 7340 3876 7348 3884
rect 7516 5056 7524 5064
rect 7500 5016 7508 5024
rect 7452 4996 7460 5004
rect 7484 4956 7492 4964
rect 7532 4956 7540 4964
rect 7500 4936 7508 4944
rect 7532 4936 7540 4944
rect 7516 4916 7524 4924
rect 7436 4876 7444 4884
rect 7420 4856 7428 4864
rect 7420 4716 7428 4724
rect 7404 4696 7412 4704
rect 7404 4656 7412 4664
rect 7436 4676 7444 4684
rect 7500 4896 7508 4904
rect 7468 4796 7476 4804
rect 7468 4696 7476 4704
rect 7452 4656 7460 4664
rect 7420 4636 7428 4644
rect 7420 4596 7428 4604
rect 7404 4536 7412 4544
rect 7404 4296 7412 4304
rect 7404 4276 7412 4284
rect 7484 4596 7492 4604
rect 7484 4536 7492 4544
rect 7452 4516 7460 4524
rect 7548 4896 7556 4904
rect 7516 4756 7524 4764
rect 7516 4716 7524 4724
rect 7436 4316 7444 4324
rect 7468 4496 7476 4504
rect 7436 4276 7444 4284
rect 7436 4256 7444 4264
rect 7468 4256 7476 4264
rect 7404 4156 7412 4164
rect 7388 4076 7396 4084
rect 7420 4136 7428 4144
rect 7404 4036 7412 4044
rect 7388 3916 7396 3924
rect 7404 3896 7412 3904
rect 7532 4516 7540 4524
rect 7532 4496 7540 4504
rect 7500 4296 7508 4304
rect 7452 4156 7460 4164
rect 7452 4116 7460 4124
rect 7452 4096 7460 4104
rect 7452 3916 7460 3924
rect 7356 3856 7364 3864
rect 7372 3856 7380 3864
rect 7436 3856 7444 3864
rect 7308 3836 7316 3844
rect 7372 3836 7380 3844
rect 7340 3796 7348 3804
rect 7308 3776 7316 3784
rect 7404 3756 7412 3764
rect 7388 3736 7396 3744
rect 7436 3736 7444 3744
rect 7452 3736 7460 3744
rect 7420 3696 7428 3704
rect 7452 3696 7460 3704
rect 7420 3676 7428 3684
rect 7388 3656 7396 3664
rect 7404 3656 7412 3664
rect 7356 3636 7364 3644
rect 7340 3576 7348 3584
rect 7276 3536 7284 3544
rect 7308 3536 7316 3544
rect 7260 3516 7268 3524
rect 7212 3496 7220 3504
rect 7116 3336 7124 3344
rect 7148 3336 7156 3344
rect 7132 3316 7140 3324
rect 7164 3316 7172 3324
rect 7244 3476 7252 3484
rect 7260 3356 7268 3364
rect 7244 3336 7252 3344
rect 7260 3336 7268 3344
rect 7308 3516 7316 3524
rect 7324 3516 7332 3524
rect 7292 3496 7300 3504
rect 7308 3476 7316 3484
rect 7308 3456 7316 3464
rect 7292 3376 7300 3384
rect 7308 3376 7316 3384
rect 7244 3316 7252 3324
rect 7036 3296 7044 3304
rect 7116 3276 7124 3284
rect 7084 3256 7092 3264
rect 7084 3136 7092 3144
rect 7004 3116 7012 3124
rect 6988 3096 6996 3104
rect 6972 3076 6980 3084
rect 6924 3016 6932 3024
rect 6908 2976 6916 2984
rect 6908 2936 6916 2944
rect 6892 2876 6900 2884
rect 6876 2756 6884 2764
rect 6876 2676 6884 2684
rect 6860 2656 6868 2664
rect 6844 2636 6852 2644
rect 6668 2536 6676 2544
rect 6780 2536 6788 2544
rect 6700 2516 6708 2524
rect 6748 2516 6756 2524
rect 6780 2516 6788 2524
rect 6716 2496 6724 2504
rect 6828 2476 6836 2484
rect 6828 2416 6836 2424
rect 6755 2406 6763 2414
rect 6765 2406 6773 2414
rect 6775 2406 6783 2414
rect 6785 2406 6793 2414
rect 6795 2406 6803 2414
rect 6805 2406 6813 2414
rect 6876 2556 6884 2564
rect 6796 2336 6804 2344
rect 6860 2336 6868 2344
rect 6636 2316 6644 2324
rect 6668 2296 6676 2304
rect 6572 2216 6580 2224
rect 6732 2316 6740 2324
rect 6828 2316 6836 2324
rect 6636 2256 6644 2264
rect 6684 2236 6692 2244
rect 6636 2216 6644 2224
rect 6700 2216 6708 2224
rect 6700 2196 6708 2204
rect 6588 2176 6596 2184
rect 6636 2176 6644 2184
rect 6572 2136 6580 2144
rect 6428 2096 6436 2104
rect 6524 2096 6532 2104
rect 6620 2096 6628 2104
rect 6572 2076 6580 2084
rect 6428 2056 6436 2064
rect 6620 2036 6628 2044
rect 6460 1976 6468 1984
rect 6508 1916 6516 1924
rect 6540 1916 6548 1924
rect 6188 1896 6196 1904
rect 6236 1896 6244 1904
rect 6300 1896 6308 1904
rect 6364 1896 6372 1904
rect 6412 1896 6420 1904
rect 6476 1896 6484 1904
rect 6524 1896 6532 1904
rect 6588 1896 6596 1904
rect 6156 1876 6164 1884
rect 6124 1856 6132 1864
rect 6012 1796 6020 1804
rect 6124 1796 6132 1804
rect 5916 1776 5924 1784
rect 5900 1756 5908 1764
rect 6108 1776 6116 1784
rect 6060 1756 6068 1764
rect 6140 1756 6148 1764
rect 5740 1636 5748 1644
rect 5708 1596 5716 1604
rect 5660 1416 5668 1424
rect 5740 1476 5748 1484
rect 5708 1456 5716 1464
rect 5820 1716 5828 1724
rect 5836 1716 5844 1724
rect 5836 1676 5844 1684
rect 5772 1636 5780 1644
rect 5836 1496 5844 1504
rect 5772 1456 5780 1464
rect 5820 1456 5828 1464
rect 5788 1416 5796 1424
rect 5756 1356 5764 1364
rect 5772 1336 5780 1344
rect 5740 1256 5748 1264
rect 5772 1136 5780 1144
rect 5836 1136 5844 1144
rect 5788 1116 5796 1124
rect 5900 1736 5908 1744
rect 5884 1596 5892 1604
rect 6220 1876 6228 1884
rect 6348 1876 6356 1884
rect 6412 1876 6420 1884
rect 6492 1876 6500 1884
rect 6508 1876 6516 1884
rect 6220 1856 6228 1864
rect 6332 1856 6340 1864
rect 6172 1736 6180 1744
rect 6252 1736 6260 1744
rect 6092 1716 6100 1724
rect 6140 1716 6148 1724
rect 6220 1716 6228 1724
rect 6364 1796 6372 1804
rect 6460 1776 6468 1784
rect 6332 1716 6340 1724
rect 5932 1696 5940 1704
rect 6204 1696 6212 1704
rect 6300 1696 6308 1704
rect 5932 1676 5940 1684
rect 5916 1496 5924 1504
rect 6028 1676 6036 1684
rect 5980 1636 5988 1644
rect 6188 1576 6196 1584
rect 5948 1516 5956 1524
rect 5996 1516 6004 1524
rect 6092 1516 6100 1524
rect 6140 1516 6148 1524
rect 6012 1496 6020 1504
rect 6044 1496 6052 1504
rect 5980 1476 5988 1484
rect 5964 1436 5972 1444
rect 5948 1416 5956 1424
rect 5996 1416 6004 1424
rect 6028 1416 6036 1424
rect 5900 1376 5908 1384
rect 6012 1356 6020 1364
rect 5932 1336 5940 1344
rect 5868 1316 5876 1324
rect 5996 1316 6004 1324
rect 5884 1296 5892 1304
rect 5884 1156 5892 1164
rect 5868 1116 5876 1124
rect 5788 1076 5796 1084
rect 5740 1016 5748 1024
rect 5836 1056 5844 1064
rect 5724 896 5732 904
rect 6076 1476 6084 1484
rect 6124 1476 6132 1484
rect 6172 1476 6180 1484
rect 6060 1396 6068 1404
rect 6284 1556 6292 1564
rect 6332 1556 6340 1564
rect 6236 1536 6244 1544
rect 6332 1536 6340 1544
rect 6540 1856 6548 1864
rect 6604 1856 6612 1864
rect 6412 1676 6420 1684
rect 6364 1516 6372 1524
rect 6220 1476 6228 1484
rect 6236 1476 6244 1484
rect 6300 1476 6308 1484
rect 6332 1496 6340 1504
rect 6364 1496 6372 1504
rect 6396 1496 6404 1504
rect 6588 1776 6596 1784
rect 6716 2176 6724 2184
rect 6652 2156 6660 2164
rect 6700 2156 6708 2164
rect 6668 2096 6676 2104
rect 6684 2096 6692 2104
rect 6652 2076 6660 2084
rect 6716 2076 6724 2084
rect 6716 1996 6724 2004
rect 6684 1936 6692 1944
rect 6700 1916 6708 1924
rect 6844 2296 6852 2304
rect 6780 2276 6788 2284
rect 6988 2956 6996 2964
rect 6972 2836 6980 2844
rect 6940 2656 6948 2664
rect 6988 2656 6996 2664
rect 6940 2616 6948 2624
rect 6956 2576 6964 2584
rect 6908 2516 6916 2524
rect 6924 2516 6932 2524
rect 6972 2516 6980 2524
rect 7020 3096 7028 3104
rect 7052 3096 7060 3104
rect 7068 3096 7076 3104
rect 7036 2976 7044 2984
rect 7052 2976 7060 2984
rect 7036 2936 7044 2944
rect 7100 2976 7108 2984
rect 7084 2956 7092 2964
rect 7100 2956 7108 2964
rect 7132 3096 7140 3104
rect 7132 3076 7140 3084
rect 7164 3076 7172 3084
rect 7148 2996 7156 3004
rect 7132 2956 7140 2964
rect 7100 2936 7108 2944
rect 7116 2936 7124 2944
rect 7020 2916 7028 2924
rect 7116 2896 7124 2904
rect 7068 2756 7076 2764
rect 7100 2736 7108 2744
rect 7324 3356 7332 3364
rect 7372 3496 7380 3504
rect 7436 3516 7444 3524
rect 7404 3496 7412 3504
rect 7420 3496 7428 3504
rect 7452 3496 7460 3504
rect 7516 4256 7524 4264
rect 7500 4156 7508 4164
rect 7516 4156 7524 4164
rect 7500 4136 7508 4144
rect 7484 4096 7492 4104
rect 7484 4076 7492 4084
rect 7516 4076 7524 4084
rect 7548 4156 7556 4164
rect 7548 4096 7556 4104
rect 7548 4076 7556 4084
rect 7500 3856 7508 3864
rect 7500 3716 7508 3724
rect 7500 3696 7508 3704
rect 7484 3656 7492 3664
rect 7532 3856 7540 3864
rect 7532 3696 7540 3704
rect 7516 3616 7524 3624
rect 7500 3576 7508 3584
rect 7500 3556 7508 3564
rect 7516 3556 7524 3564
rect 7404 3476 7412 3484
rect 7388 3456 7396 3464
rect 7452 3456 7460 3464
rect 7436 3436 7444 3444
rect 7372 3416 7380 3424
rect 7388 3396 7396 3404
rect 7356 3376 7364 3384
rect 7388 3376 7396 3384
rect 7500 3436 7508 3444
rect 7324 3336 7332 3344
rect 7340 3316 7348 3324
rect 7308 3256 7316 3264
rect 7340 3256 7348 3264
rect 7276 3156 7284 3164
rect 7212 3116 7220 3124
rect 7468 3356 7476 3364
rect 7404 3336 7412 3344
rect 7436 3336 7444 3344
rect 7388 3316 7396 3324
rect 7420 3296 7428 3304
rect 7372 3276 7380 3284
rect 7388 3116 7396 3124
rect 7436 3116 7444 3124
rect 7356 3096 7364 3104
rect 7196 3076 7204 3084
rect 7244 3076 7252 3084
rect 7356 3076 7364 3084
rect 7388 3076 7396 3084
rect 7228 3056 7236 3064
rect 7180 2996 7188 3004
rect 7164 2956 7172 2964
rect 7228 3016 7236 3024
rect 7340 2976 7348 2984
rect 7164 2936 7172 2944
rect 7228 2936 7236 2944
rect 7196 2916 7204 2924
rect 7228 2916 7236 2924
rect 7132 2876 7140 2884
rect 7132 2756 7140 2764
rect 7148 2716 7156 2724
rect 7036 2696 7044 2704
rect 7116 2696 7124 2704
rect 7148 2676 7156 2684
rect 7212 2736 7220 2744
rect 7180 2696 7188 2704
rect 7020 2636 7028 2644
rect 7036 2636 7044 2644
rect 7084 2636 7092 2644
rect 7052 2536 7060 2544
rect 7100 2616 7108 2624
rect 7004 2496 7012 2504
rect 6908 2456 6916 2464
rect 6924 2456 6932 2464
rect 7116 2456 7124 2464
rect 7052 2436 7060 2444
rect 7116 2416 7124 2424
rect 6940 2376 6948 2384
rect 7084 2336 7092 2344
rect 7132 2336 7140 2344
rect 6972 2316 6980 2324
rect 7132 2316 7140 2324
rect 7116 2296 7124 2304
rect 7132 2296 7140 2304
rect 7164 2636 7172 2644
rect 7212 2596 7220 2604
rect 7196 2576 7204 2584
rect 7196 2536 7204 2544
rect 7180 2476 7188 2484
rect 7164 2376 7172 2384
rect 7196 2316 7204 2324
rect 6940 2276 6948 2284
rect 6892 2256 6900 2264
rect 6892 2216 6900 2224
rect 6876 2176 6884 2184
rect 6892 2176 6900 2184
rect 6764 2136 6772 2144
rect 6860 2136 6868 2144
rect 6748 2096 6756 2104
rect 6876 2096 6884 2104
rect 6755 2006 6763 2014
rect 6765 2006 6773 2014
rect 6775 2006 6783 2014
rect 6785 2006 6793 2014
rect 6795 2006 6803 2014
rect 6805 2006 6813 2014
rect 6732 1896 6740 1904
rect 7004 2216 7012 2224
rect 6972 2176 6980 2184
rect 6988 2176 6996 2184
rect 6956 2156 6964 2164
rect 6988 2156 6996 2164
rect 6988 2136 6996 2144
rect 6940 2096 6948 2104
rect 7084 2256 7092 2264
rect 7036 2196 7044 2204
rect 7084 2216 7092 2224
rect 7100 2196 7108 2204
rect 7020 2116 7028 2124
rect 7004 2096 7012 2104
rect 6924 1976 6932 1984
rect 6956 1976 6964 1984
rect 6924 1956 6932 1964
rect 6828 1896 6836 1904
rect 6684 1856 6692 1864
rect 6476 1696 6484 1704
rect 6444 1676 6452 1684
rect 6508 1696 6516 1704
rect 6556 1696 6564 1704
rect 6444 1516 6452 1524
rect 6460 1516 6468 1524
rect 6444 1496 6452 1504
rect 6396 1476 6404 1484
rect 6428 1476 6436 1484
rect 6316 1456 6324 1464
rect 6428 1456 6436 1464
rect 6268 1436 6276 1444
rect 6236 1416 6244 1424
rect 6460 1436 6468 1444
rect 6444 1396 6452 1404
rect 6108 1376 6116 1384
rect 6124 1356 6132 1364
rect 6140 1356 6148 1364
rect 6204 1356 6212 1364
rect 6284 1356 6292 1364
rect 6332 1356 6340 1364
rect 6444 1356 6452 1364
rect 6060 1336 6068 1344
rect 6108 1336 6116 1344
rect 6092 1316 6100 1324
rect 6156 1316 6164 1324
rect 6188 1316 6196 1324
rect 6220 1316 6228 1324
rect 6252 1316 6260 1324
rect 6156 1176 6164 1184
rect 6044 1116 6052 1124
rect 6412 1336 6420 1344
rect 6316 1316 6324 1324
rect 6348 1316 6356 1324
rect 6332 1296 6340 1304
rect 6572 1496 6580 1504
rect 6524 1476 6532 1484
rect 6492 1456 6500 1464
rect 6524 1456 6532 1464
rect 6508 1316 6516 1324
rect 6732 1776 6740 1784
rect 6684 1756 6692 1764
rect 6892 1856 6900 1864
rect 6860 1796 6868 1804
rect 6892 1796 6900 1804
rect 6828 1756 6836 1764
rect 6860 1736 6868 1744
rect 6828 1716 6836 1724
rect 6860 1716 6868 1724
rect 6988 1776 6996 1784
rect 6940 1756 6948 1764
rect 6972 1756 6980 1764
rect 6860 1696 6868 1704
rect 6924 1696 6932 1704
rect 6620 1676 6628 1684
rect 6652 1676 6660 1684
rect 6748 1676 6756 1684
rect 6700 1656 6708 1664
rect 6636 1636 6644 1644
rect 6748 1636 6756 1644
rect 6755 1606 6763 1614
rect 6765 1606 6773 1614
rect 6775 1606 6783 1614
rect 6785 1606 6793 1614
rect 6795 1606 6803 1614
rect 6805 1606 6813 1614
rect 6732 1516 6740 1524
rect 7004 1716 7012 1724
rect 7068 2156 7076 2164
rect 7180 2296 7188 2304
rect 7180 2276 7188 2284
rect 7148 2176 7156 2184
rect 7196 2256 7204 2264
rect 7212 2236 7220 2244
rect 7276 2776 7284 2784
rect 7244 2756 7252 2764
rect 7260 2596 7268 2604
rect 7244 2576 7252 2584
rect 7260 2556 7268 2564
rect 7260 2536 7268 2544
rect 7292 2756 7300 2764
rect 7372 2996 7380 3004
rect 7372 2976 7380 2984
rect 7356 2796 7364 2804
rect 7420 3056 7428 3064
rect 7468 3316 7476 3324
rect 7532 3436 7540 3444
rect 7516 3356 7524 3364
rect 7532 3316 7540 3324
rect 7484 3176 7492 3184
rect 7516 3076 7524 3084
rect 7452 2976 7460 2984
rect 7388 2896 7396 2904
rect 7468 2876 7476 2884
rect 7372 2776 7380 2784
rect 7452 2756 7460 2764
rect 7324 2736 7332 2744
rect 7388 2736 7396 2744
rect 7372 2716 7380 2724
rect 7292 2696 7300 2704
rect 7308 2696 7316 2704
rect 7324 2676 7332 2684
rect 7420 2696 7428 2704
rect 7404 2676 7412 2684
rect 7436 2676 7444 2684
rect 7484 2856 7492 2864
rect 7516 2876 7524 2884
rect 7468 2716 7476 2724
rect 7500 2756 7508 2764
rect 7484 2676 7492 2684
rect 7340 2656 7348 2664
rect 7388 2656 7396 2664
rect 7308 2636 7316 2644
rect 7356 2636 7364 2644
rect 7468 2636 7476 2644
rect 7468 2616 7476 2624
rect 7340 2596 7348 2604
rect 7308 2576 7316 2584
rect 7356 2556 7364 2564
rect 7292 2536 7300 2544
rect 7452 2536 7460 2544
rect 7388 2516 7396 2524
rect 7452 2516 7460 2524
rect 7340 2376 7348 2384
rect 7436 2356 7444 2364
rect 7276 2316 7284 2324
rect 7244 2256 7252 2264
rect 7260 2256 7268 2264
rect 7132 2116 7140 2124
rect 7180 2116 7188 2124
rect 7116 2096 7124 2104
rect 7244 2156 7252 2164
rect 7228 2096 7236 2104
rect 7100 2076 7108 2084
rect 7180 2076 7188 2084
rect 7212 2076 7220 2084
rect 7052 1916 7060 1924
rect 7084 1896 7092 1904
rect 7052 1876 7060 1884
rect 7196 1896 7204 1904
rect 7212 1876 7220 1884
rect 7244 1876 7252 1884
rect 7068 1836 7076 1844
rect 7116 1836 7124 1844
rect 7148 1836 7156 1844
rect 7180 1836 7188 1844
rect 7116 1816 7124 1824
rect 7100 1756 7108 1764
rect 7036 1696 7044 1704
rect 6940 1676 6948 1684
rect 7004 1676 7012 1684
rect 6908 1536 6916 1544
rect 7004 1536 7012 1544
rect 6972 1516 6980 1524
rect 6988 1516 6996 1524
rect 6700 1496 6708 1504
rect 6860 1496 6868 1504
rect 6940 1496 6948 1504
rect 6636 1476 6644 1484
rect 6636 1456 6644 1464
rect 6668 1456 6676 1464
rect 6732 1476 6740 1484
rect 6908 1476 6916 1484
rect 6684 1416 6692 1424
rect 7084 1716 7092 1724
rect 7068 1676 7076 1684
rect 7132 1656 7140 1664
rect 7052 1516 7060 1524
rect 7132 1516 7140 1524
rect 7020 1496 7028 1504
rect 6988 1476 6996 1484
rect 7116 1476 7124 1484
rect 6956 1456 6964 1464
rect 7020 1456 7028 1464
rect 7116 1456 7124 1464
rect 6924 1416 6932 1424
rect 7100 1436 7108 1444
rect 7052 1416 7060 1424
rect 7052 1396 7060 1404
rect 6604 1356 6612 1364
rect 6652 1356 6660 1364
rect 6684 1356 6692 1364
rect 6876 1356 6884 1364
rect 7036 1356 7044 1364
rect 6588 1336 6596 1344
rect 6524 1296 6532 1304
rect 6556 1296 6564 1304
rect 6588 1296 6596 1304
rect 6428 1276 6436 1284
rect 6476 1276 6484 1284
rect 6588 1256 6596 1264
rect 6636 1296 6644 1304
rect 6668 1296 6676 1304
rect 6908 1256 6916 1264
rect 6755 1206 6763 1214
rect 6765 1206 6773 1214
rect 6775 1206 6783 1214
rect 6785 1206 6793 1214
rect 6795 1206 6803 1214
rect 6805 1206 6813 1214
rect 6796 1176 6804 1184
rect 6332 1136 6340 1144
rect 6476 1136 6484 1144
rect 6604 1136 6612 1144
rect 6652 1136 6660 1144
rect 6716 1136 6724 1144
rect 6252 1116 6260 1124
rect 6284 1116 6292 1124
rect 6348 1116 6356 1124
rect 6508 1116 6516 1124
rect 6012 1096 6020 1104
rect 6124 1096 6132 1104
rect 6204 1096 6212 1104
rect 6268 1096 6276 1104
rect 6364 1096 6372 1104
rect 6460 1096 6468 1104
rect 5932 1076 5940 1084
rect 5996 1076 6004 1084
rect 6108 1076 6116 1084
rect 5916 996 5924 1004
rect 5948 976 5956 984
rect 5884 956 5892 964
rect 6140 1036 6148 1044
rect 6268 1076 6276 1084
rect 6460 1076 6468 1084
rect 6188 1056 6196 1064
rect 6220 1056 6228 1064
rect 6172 1036 6180 1044
rect 6252 1036 6260 1044
rect 6156 976 6164 984
rect 6156 956 6164 964
rect 6332 1056 6340 1064
rect 6300 1036 6308 1044
rect 5836 936 5844 944
rect 5900 936 5908 944
rect 5964 936 5972 944
rect 6028 936 6036 944
rect 6156 936 6164 944
rect 5772 916 5780 924
rect 5804 916 5812 924
rect 6316 936 6324 944
rect 6380 1036 6388 1044
rect 6428 1036 6436 1044
rect 6668 1096 6676 1104
rect 6652 1076 6660 1084
rect 6636 1056 6644 1064
rect 6700 1076 6708 1084
rect 6572 1036 6580 1044
rect 6540 1016 6548 1024
rect 6572 1016 6580 1024
rect 6508 996 6516 1004
rect 7068 1336 7076 1344
rect 7004 1316 7012 1324
rect 7052 1276 7060 1284
rect 6972 1256 6980 1264
rect 6956 1176 6964 1184
rect 6892 1116 6900 1124
rect 6908 1116 6916 1124
rect 6972 1116 6980 1124
rect 6748 1096 6756 1104
rect 6732 1056 6740 1064
rect 6812 1056 6820 1064
rect 6844 1056 6852 1064
rect 6732 1036 6740 1044
rect 6604 976 6612 984
rect 6380 956 6388 964
rect 6444 956 6452 964
rect 6364 936 6372 944
rect 6396 940 6404 944
rect 6396 936 6404 940
rect 5948 916 5956 924
rect 6012 916 6020 924
rect 6108 916 6116 924
rect 6540 916 6548 924
rect 5820 876 5828 884
rect 5756 856 5764 864
rect 5644 716 5652 724
rect 5660 716 5668 724
rect 5452 696 5460 704
rect 5388 676 5396 684
rect 5436 676 5444 684
rect 5324 536 5332 544
rect 5356 536 5364 544
rect 5196 496 5204 504
rect 5100 436 5108 444
rect 5932 896 5940 904
rect 6060 896 6068 904
rect 6044 876 6052 884
rect 5932 836 5940 844
rect 6060 796 6068 804
rect 5964 716 5972 724
rect 6012 716 6020 724
rect 5484 676 5492 684
rect 5532 676 5540 684
rect 5548 676 5556 684
rect 5788 676 5796 684
rect 5420 556 5428 564
rect 5388 516 5396 524
rect 5340 496 5348 504
rect 5404 496 5412 504
rect 5676 636 5684 644
rect 5708 636 5716 644
rect 5724 636 5732 644
rect 5788 656 5796 664
rect 5852 656 5860 664
rect 5644 616 5652 624
rect 5564 576 5572 584
rect 5596 556 5604 564
rect 5516 536 5524 544
rect 5500 516 5508 524
rect 5532 516 5540 524
rect 5468 496 5476 504
rect 5500 496 5508 504
rect 5420 476 5428 484
rect 5388 456 5396 464
rect 5308 416 5316 424
rect 5164 396 5172 404
rect 5100 356 5108 364
rect 5132 356 5140 364
rect 5068 276 5076 284
rect 4972 256 4980 264
rect 4796 136 4804 144
rect 5004 236 5012 244
rect 4988 156 4996 164
rect 4780 116 4788 124
rect 4828 116 4836 124
rect 4844 116 4852 124
rect 4876 116 4884 124
rect 4940 116 4948 124
rect 4796 96 4804 104
rect 4812 96 4820 104
rect 4860 96 4868 104
rect 5084 216 5092 224
rect 5148 276 5156 284
rect 5196 356 5204 364
rect 5260 336 5268 344
rect 5356 316 5364 324
rect 5212 276 5220 284
rect 5116 256 5124 264
rect 5132 256 5140 264
rect 5164 256 5172 264
rect 5100 196 5108 204
rect 5068 176 5076 184
rect 5052 136 5060 144
rect 5180 216 5188 224
rect 5212 216 5220 224
rect 5196 196 5204 204
rect 5100 156 5108 164
rect 5196 156 5204 164
rect 5084 136 5092 144
rect 5340 296 5348 304
rect 5244 276 5252 284
rect 5260 276 5268 284
rect 5292 276 5300 284
rect 5340 276 5348 284
rect 5324 236 5332 244
rect 5251 206 5259 214
rect 5261 206 5269 214
rect 5271 206 5279 214
rect 5281 206 5289 214
rect 5291 206 5299 214
rect 5301 206 5309 214
rect 5468 436 5476 444
rect 5420 336 5428 344
rect 5612 516 5620 524
rect 5660 516 5668 524
rect 5580 496 5588 504
rect 5628 496 5636 504
rect 5644 496 5652 504
rect 5772 636 5780 644
rect 5852 636 5860 644
rect 5932 696 5940 704
rect 6028 696 6036 704
rect 5996 656 6004 664
rect 5900 636 5908 644
rect 5980 636 5988 644
rect 5868 616 5876 624
rect 5900 616 5908 624
rect 6028 576 6036 584
rect 5740 536 5748 544
rect 5868 536 5876 544
rect 5980 536 5988 544
rect 5548 476 5556 484
rect 5612 476 5620 484
rect 5516 396 5524 404
rect 5644 416 5652 424
rect 5404 316 5412 324
rect 5468 316 5476 324
rect 5388 296 5396 304
rect 5500 296 5508 304
rect 5484 276 5492 284
rect 5548 276 5556 284
rect 5596 256 5604 264
rect 5436 236 5444 244
rect 5484 236 5492 244
rect 5596 236 5604 244
rect 5356 216 5364 224
rect 5404 216 5412 224
rect 5324 196 5332 204
rect 5228 176 5236 184
rect 5420 196 5428 204
rect 5132 96 5140 104
rect 5196 96 5204 104
rect 5212 96 5220 104
rect 5484 156 5492 164
rect 5644 296 5652 304
rect 5740 496 5748 504
rect 5708 436 5716 444
rect 5708 396 5716 404
rect 5692 356 5700 364
rect 5692 316 5700 324
rect 5676 276 5684 284
rect 5644 236 5652 244
rect 5660 176 5668 184
rect 5692 176 5700 184
rect 5804 456 5812 464
rect 6140 876 6148 884
rect 6508 896 6516 904
rect 6332 816 6340 824
rect 6732 956 6740 964
rect 6668 936 6676 944
rect 6588 916 6596 924
rect 6652 916 6660 924
rect 6556 896 6564 904
rect 6540 856 6548 864
rect 6332 776 6340 784
rect 6508 756 6516 764
rect 6476 736 6484 744
rect 6348 716 6356 724
rect 6412 716 6420 724
rect 6188 696 6196 704
rect 6236 696 6244 704
rect 6316 696 6324 704
rect 6364 696 6372 704
rect 6412 696 6420 704
rect 6444 696 6452 704
rect 6092 676 6100 684
rect 6172 676 6180 684
rect 6284 676 6292 684
rect 6460 676 6468 684
rect 6124 656 6132 664
rect 6220 656 6228 664
rect 6348 656 6356 664
rect 6396 656 6404 664
rect 6092 596 6100 604
rect 6268 596 6276 604
rect 6076 536 6084 544
rect 6044 496 6052 504
rect 5948 376 5956 384
rect 5868 316 5876 324
rect 5916 316 5924 324
rect 5756 296 5764 304
rect 5836 296 5844 304
rect 5724 276 5732 284
rect 5740 276 5748 284
rect 5788 276 5796 284
rect 5820 276 5828 284
rect 5916 276 5924 284
rect 5932 276 5940 284
rect 5756 176 5764 184
rect 5884 256 5892 264
rect 5852 196 5860 204
rect 5788 156 5796 164
rect 5884 156 5892 164
rect 5804 136 5812 144
rect 5628 116 5636 124
rect 5516 96 5524 104
rect 5964 316 5972 324
rect 6028 316 6036 324
rect 5980 296 5988 304
rect 6060 296 6068 304
rect 6124 576 6132 584
rect 6108 536 6116 544
rect 6188 536 6196 544
rect 6268 536 6276 544
rect 6172 516 6180 524
rect 6204 516 6212 524
rect 6220 516 6228 524
rect 6156 496 6164 504
rect 6140 476 6148 484
rect 6108 456 6116 464
rect 6140 456 6148 464
rect 6252 476 6260 484
rect 6252 356 6260 364
rect 6332 636 6340 644
rect 6300 616 6308 624
rect 6316 556 6324 564
rect 6556 776 6564 784
rect 6588 776 6596 784
rect 6572 696 6580 704
rect 6572 676 6580 684
rect 6540 656 6548 664
rect 6412 576 6420 584
rect 6476 576 6484 584
rect 6380 556 6388 564
rect 6460 556 6468 564
rect 6412 536 6420 544
rect 6556 556 6564 564
rect 6572 556 6580 564
rect 6524 536 6532 544
rect 6396 516 6404 524
rect 6412 516 6420 524
rect 6364 496 6372 504
rect 6396 356 6404 364
rect 6348 316 6356 324
rect 6284 296 6292 304
rect 6444 336 6452 344
rect 6556 336 6564 344
rect 6412 316 6420 324
rect 6476 316 6484 324
rect 6524 316 6532 324
rect 6604 696 6612 704
rect 6636 696 6644 704
rect 6620 676 6628 684
rect 6876 1036 6884 1044
rect 6860 936 6868 944
rect 6828 916 6836 924
rect 6732 896 6740 904
rect 6716 716 6724 724
rect 6924 1056 6932 1064
rect 6940 1056 6948 1064
rect 6908 940 6916 944
rect 6908 936 6916 940
rect 6940 936 6948 944
rect 6956 896 6964 904
rect 6892 876 6900 884
rect 7084 1116 7092 1124
rect 7244 1796 7252 1804
rect 7260 1736 7268 1744
rect 7196 1716 7204 1724
rect 7324 2276 7332 2284
rect 7420 2276 7428 2284
rect 7292 2256 7300 2264
rect 7356 2236 7364 2244
rect 7324 2216 7332 2224
rect 7308 2136 7316 2144
rect 7308 1916 7316 1924
rect 7292 1896 7300 1904
rect 7308 1896 7316 1904
rect 7308 1736 7316 1744
rect 7164 1676 7172 1684
rect 7180 1656 7188 1664
rect 7164 1516 7172 1524
rect 7276 1696 7284 1704
rect 7292 1676 7300 1684
rect 7308 1676 7316 1684
rect 7260 1636 7268 1644
rect 7340 2176 7348 2184
rect 7388 2176 7396 2184
rect 7372 2116 7380 2124
rect 7388 2096 7396 2104
rect 7468 2476 7476 2484
rect 7468 2316 7476 2324
rect 7452 2236 7460 2244
rect 7484 2276 7492 2284
rect 7484 2256 7492 2264
rect 7532 2856 7540 2864
rect 7532 2836 7540 2844
rect 7532 2696 7540 2704
rect 7516 2656 7524 2664
rect 7532 2476 7540 2484
rect 7564 3916 7572 3924
rect 7564 3896 7572 3904
rect 7564 3716 7572 3724
rect 7564 3696 7572 3704
rect 7548 2396 7556 2404
rect 7516 2336 7524 2344
rect 7516 2296 7524 2304
rect 7548 2256 7556 2264
rect 7548 2236 7556 2244
rect 7500 2176 7508 2184
rect 7532 2156 7540 2164
rect 7436 2136 7444 2144
rect 7436 2116 7444 2124
rect 7404 1936 7412 1944
rect 7340 1916 7348 1924
rect 7388 1916 7396 1924
rect 7340 1876 7348 1884
rect 7420 1796 7428 1804
rect 7372 1776 7380 1784
rect 7356 1736 7364 1744
rect 7388 1736 7396 1744
rect 7468 2096 7476 2104
rect 7452 1916 7460 1924
rect 7484 1916 7492 1924
rect 7516 1896 7524 1904
rect 7500 1876 7508 1884
rect 7500 1856 7508 1864
rect 7452 1776 7460 1784
rect 7340 1676 7348 1684
rect 7388 1656 7396 1664
rect 7276 1616 7284 1624
rect 7324 1616 7332 1624
rect 7212 1536 7220 1544
rect 7132 1356 7140 1364
rect 7148 1356 7156 1364
rect 7164 1336 7172 1344
rect 7116 1296 7124 1304
rect 7148 1316 7156 1324
rect 7180 1316 7188 1324
rect 7244 1436 7252 1444
rect 7228 1356 7236 1364
rect 7164 1296 7172 1304
rect 7196 1296 7204 1304
rect 7132 1176 7140 1184
rect 7068 1036 7076 1044
rect 7004 996 7012 1004
rect 7004 956 7012 964
rect 6988 936 6996 944
rect 6988 916 6996 924
rect 6972 856 6980 864
rect 6972 836 6980 844
rect 6755 806 6763 814
rect 6765 806 6773 814
rect 6775 806 6783 814
rect 6785 806 6793 814
rect 6795 806 6803 814
rect 6805 806 6813 814
rect 6876 736 6884 744
rect 6908 736 6916 744
rect 6924 716 6932 724
rect 6748 696 6756 704
rect 6828 696 6836 704
rect 6700 676 6708 684
rect 6620 656 6628 664
rect 6620 596 6628 604
rect 6652 596 6660 604
rect 6956 696 6964 704
rect 6956 676 6964 684
rect 6924 656 6932 664
rect 6940 596 6948 604
rect 6700 576 6708 584
rect 6700 556 6708 564
rect 6812 556 6820 564
rect 6876 556 6884 564
rect 6508 296 6516 304
rect 5964 276 5972 284
rect 6012 276 6020 284
rect 6076 276 6084 284
rect 6172 276 6180 284
rect 6220 276 6228 284
rect 6268 276 6276 284
rect 6508 276 6516 284
rect 6124 256 6132 264
rect 6204 256 6212 264
rect 6252 256 6260 264
rect 6028 236 6036 244
rect 5932 116 5940 124
rect 5980 116 5988 124
rect 6044 116 6052 124
rect 6156 136 6164 144
rect 6140 116 6148 124
rect 6236 216 6244 224
rect 6220 136 6228 144
rect 6268 136 6276 144
rect 6316 136 6324 144
rect 6380 136 6388 144
rect 6204 116 6212 124
rect 6284 116 6292 124
rect 6316 116 6324 124
rect 6476 236 6484 244
rect 6636 516 6644 524
rect 7068 936 7076 944
rect 7036 916 7044 924
rect 7052 896 7060 904
rect 7036 856 7044 864
rect 7004 716 7012 724
rect 6988 576 6996 584
rect 6668 536 6676 544
rect 6940 536 6948 544
rect 6668 516 6676 524
rect 6780 516 6788 524
rect 6892 516 6900 524
rect 6755 406 6763 414
rect 6765 406 6773 414
rect 6775 406 6783 414
rect 6785 406 6793 414
rect 6795 406 6803 414
rect 6805 406 6813 414
rect 6668 356 6676 364
rect 6716 316 6724 324
rect 6876 316 6884 324
rect 6636 296 6644 304
rect 6684 276 6692 284
rect 6844 276 6852 284
rect 6636 256 6644 264
rect 6828 256 6836 264
rect 6860 256 6868 264
rect 6588 236 6596 244
rect 6620 236 6628 244
rect 6572 136 6580 144
rect 6668 236 6676 244
rect 6716 236 6724 244
rect 6636 136 6644 144
rect 6684 136 6692 144
rect 6748 216 6756 224
rect 6844 136 6852 144
rect 6924 436 6932 444
rect 6940 316 6948 324
rect 6924 256 6932 264
rect 6908 236 6916 244
rect 6940 236 6948 244
rect 6892 196 6900 204
rect 5964 96 5972 104
rect 6188 96 6196 104
rect 6332 96 6340 104
rect 6668 96 6676 104
rect 6700 96 6708 104
rect 7020 676 7028 684
rect 7052 676 7060 684
rect 7100 1056 7108 1064
rect 7116 1036 7124 1044
rect 7132 896 7140 904
rect 7100 876 7108 884
rect 7132 876 7140 884
rect 7180 1276 7188 1284
rect 7228 1276 7236 1284
rect 7388 1576 7396 1584
rect 7292 1496 7300 1504
rect 7292 1476 7300 1484
rect 7308 1456 7316 1464
rect 7340 1456 7348 1464
rect 7292 1356 7300 1364
rect 7276 1336 7284 1344
rect 7324 1436 7332 1444
rect 7356 1376 7364 1384
rect 7404 1376 7412 1384
rect 7324 1356 7332 1364
rect 7340 1356 7348 1364
rect 7436 1356 7444 1364
rect 7484 1716 7492 1724
rect 7484 1696 7492 1704
rect 7532 1876 7540 1884
rect 7548 1856 7556 1864
rect 7548 1796 7556 1804
rect 7516 1776 7524 1784
rect 7516 1756 7524 1764
rect 7548 1756 7556 1764
rect 7500 1676 7508 1684
rect 7468 1516 7476 1524
rect 7468 1456 7476 1464
rect 7516 1496 7524 1504
rect 7500 1476 7508 1484
rect 7500 1456 7508 1464
rect 7324 1336 7332 1344
rect 7452 1336 7460 1344
rect 7308 1316 7316 1324
rect 7292 1296 7300 1304
rect 7260 1276 7268 1284
rect 7180 1096 7188 1104
rect 7228 1056 7236 1064
rect 7244 996 7252 1004
rect 7196 976 7204 984
rect 7180 936 7188 944
rect 7196 936 7204 944
rect 7292 1056 7300 1064
rect 7308 996 7316 1004
rect 7292 956 7300 964
rect 7260 916 7268 924
rect 7196 856 7204 864
rect 7116 656 7124 664
rect 7068 556 7076 564
rect 7052 536 7060 544
rect 7100 536 7108 544
rect 7164 676 7172 684
rect 7164 516 7172 524
rect 7132 436 7140 444
rect 7180 496 7188 504
rect 7308 736 7316 744
rect 7212 716 7220 724
rect 7276 676 7284 684
rect 7340 1316 7348 1324
rect 7388 1316 7396 1324
rect 7452 1316 7460 1324
rect 7500 1316 7508 1324
rect 7484 1276 7492 1284
rect 7468 1256 7476 1264
rect 7372 1096 7380 1104
rect 7404 1096 7412 1104
rect 7468 1096 7476 1104
rect 7484 1096 7492 1104
rect 7516 1076 7524 1084
rect 7468 1056 7476 1064
rect 7500 1056 7508 1064
rect 7372 1036 7380 1044
rect 7356 956 7364 964
rect 7516 1016 7524 1024
rect 7564 1496 7572 1504
rect 7564 1296 7572 1304
rect 7564 1256 7572 1264
rect 7532 996 7540 1004
rect 7340 936 7348 944
rect 7340 916 7348 924
rect 7340 716 7348 724
rect 7484 956 7492 964
rect 7532 936 7540 944
rect 7420 916 7428 924
rect 7532 916 7540 924
rect 7404 776 7412 784
rect 7500 776 7508 784
rect 7388 736 7396 744
rect 7388 696 7396 704
rect 7436 696 7444 704
rect 7356 676 7364 684
rect 7420 676 7428 684
rect 7324 636 7332 644
rect 7228 616 7236 624
rect 7212 536 7220 544
rect 7548 776 7556 784
rect 7452 636 7460 644
rect 7292 556 7300 564
rect 7356 556 7364 564
rect 7420 556 7428 564
rect 7324 516 7332 524
rect 7228 496 7236 504
rect 7292 496 7300 504
rect 6988 276 6996 284
rect 6972 256 6980 264
rect 7004 256 7012 264
rect 6972 196 6980 204
rect 7148 316 7156 324
rect 7020 216 7028 224
rect 7372 436 7380 444
rect 7228 316 7236 324
rect 7292 316 7300 324
rect 7372 316 7380 324
rect 7212 296 7220 304
rect 7196 236 7204 244
rect 7148 196 7156 204
rect 6924 156 6932 164
rect 7004 156 7012 164
rect 7036 156 7044 164
rect 7052 156 7060 164
rect 7148 156 7156 164
rect 6956 136 6964 144
rect 7052 136 7060 144
rect 7100 136 7108 144
rect 7212 156 7220 164
rect 7260 296 7268 304
rect 7308 296 7316 304
rect 7356 296 7364 304
rect 7404 296 7412 304
rect 7340 256 7348 264
rect 7244 156 7252 164
rect 7308 156 7316 164
rect 7500 576 7508 584
rect 7484 556 7492 564
rect 7500 536 7508 544
rect 7468 336 7476 344
rect 7484 316 7492 324
rect 7436 276 7444 284
rect 7484 276 7492 284
rect 7420 256 7428 264
rect 7388 236 7396 244
rect 7388 156 7396 164
rect 7516 296 7524 304
rect 7564 336 7572 344
rect 7532 276 7540 284
rect 7532 256 7540 264
rect 7276 136 7284 144
rect 7516 136 7524 144
rect 7004 116 7012 124
rect 7116 116 7124 124
rect 7468 116 7476 124
rect 7532 116 7540 124
rect 7276 96 7284 104
rect 7308 96 7316 104
rect 4460 76 4468 84
rect 4492 76 4500 84
rect 4508 76 4516 84
rect 4572 76 4580 84
rect 4588 76 4596 84
rect 4684 76 4692 84
rect 5052 76 5060 84
rect 5420 76 5428 84
rect 4428 56 4436 64
rect 4476 56 4484 64
rect 3747 6 3755 14
rect 3757 6 3765 14
rect 3767 6 3775 14
rect 3777 6 3785 14
rect 3787 6 3795 14
rect 3797 6 3805 14
rect 5676 16 5684 24
rect 6755 6 6763 14
rect 6765 6 6773 14
rect 6775 6 6783 14
rect 6785 6 6793 14
rect 6795 6 6803 14
rect 6805 6 6813 14
<< metal3 >>
rect 3860 5217 3884 5223
rect 4756 5217 4764 5223
rect 738 5214 798 5216
rect 738 5206 739 5214
rect 748 5206 749 5214
rect 787 5206 788 5214
rect 797 5206 798 5214
rect 738 5204 798 5206
rect 3746 5214 3806 5216
rect 3746 5206 3747 5214
rect 3756 5206 3757 5214
rect 3795 5206 3796 5214
rect 3805 5206 3806 5214
rect 3746 5204 3806 5206
rect 6754 5214 6814 5216
rect 6754 5206 6755 5214
rect 6764 5206 6765 5214
rect 6803 5206 6804 5214
rect 6813 5206 6814 5214
rect 6754 5204 6814 5206
rect 4212 5157 5907 5163
rect 5901 5144 5907 5157
rect 6036 5157 6156 5163
rect 4452 5137 4636 5143
rect 4644 5137 4684 5143
rect 4932 5137 4956 5143
rect 5444 5137 5532 5143
rect 5556 5137 5724 5143
rect 5908 5137 6732 5143
rect 388 5117 476 5123
rect 1028 5117 1100 5123
rect 2740 5117 2892 5123
rect 3428 5117 3580 5123
rect 4740 5117 4780 5123
rect 4804 5117 4828 5123
rect 4884 5117 4972 5123
rect 4980 5117 5036 5123
rect 5044 5117 5068 5123
rect 5156 5117 5180 5123
rect 5524 5117 5612 5123
rect 6020 5117 6076 5123
rect 6084 5117 6188 5123
rect 6196 5117 6220 5123
rect 6308 5117 6332 5123
rect 7060 5117 7180 5123
rect 212 5097 844 5103
rect 852 5097 1036 5103
rect 1268 5097 1292 5103
rect 1524 5097 1740 5103
rect 1748 5097 1804 5103
rect 1844 5097 1964 5103
rect 2116 5097 2236 5103
rect 2420 5097 2492 5103
rect 2516 5097 2604 5103
rect 2612 5097 2764 5103
rect 2868 5097 3036 5103
rect 3060 5097 3212 5103
rect 3284 5097 3532 5103
rect 3716 5097 3948 5103
rect 3988 5097 4076 5103
rect 4500 5097 4604 5103
rect 4612 5097 5340 5103
rect 5348 5097 5404 5103
rect 5412 5097 5468 5103
rect 6068 5097 6092 5103
rect 6612 5097 6828 5103
rect 6884 5097 6940 5103
rect 7140 5097 7164 5103
rect 7316 5097 7356 5103
rect 132 5077 444 5083
rect 452 5077 684 5083
rect 692 5077 1068 5083
rect 1508 5077 1660 5083
rect 1780 5077 1836 5083
rect 1892 5077 2012 5083
rect 2020 5077 2172 5083
rect 2180 5077 2252 5083
rect 2484 5077 2572 5083
rect 2644 5077 3084 5083
rect 3364 5077 3436 5083
rect 3460 5077 3660 5083
rect 4260 5077 4556 5083
rect 4756 5077 4796 5083
rect 4820 5077 4876 5083
rect 5012 5077 5116 5083
rect 5124 5077 5180 5083
rect 5188 5077 5228 5083
rect 5364 5077 5532 5083
rect 5540 5077 5580 5083
rect 5732 5077 5772 5083
rect 5924 5077 6060 5083
rect 6084 5077 6124 5083
rect 6276 5077 6332 5083
rect 6964 5077 7036 5083
rect 7092 5077 7276 5083
rect 7284 5077 7308 5083
rect 7316 5077 7324 5083
rect 228 5057 268 5063
rect 276 5057 316 5063
rect 324 5057 396 5063
rect 900 5057 972 5063
rect 980 5057 1468 5063
rect 1476 5057 1516 5063
rect 1684 5057 2060 5063
rect 2356 5057 2540 5063
rect 3396 5057 3468 5063
rect 4100 5057 4316 5063
rect 4660 5057 4700 5063
rect 4708 5057 4716 5063
rect 4772 5057 4812 5063
rect 4836 5057 4924 5063
rect 5076 5057 5148 5063
rect 5204 5057 5212 5063
rect 5396 5057 5452 5063
rect 5732 5057 5852 5063
rect 5860 5057 5916 5063
rect 5972 5057 6092 5063
rect 6228 5057 6300 5063
rect 6340 5057 6380 5063
rect 6388 5057 6476 5063
rect 6484 5057 6588 5063
rect 6596 5057 6668 5063
rect 6676 5057 6716 5063
rect 6852 5057 7004 5063
rect 7012 5057 7084 5063
rect 7236 5057 7324 5063
rect 7348 5057 7404 5063
rect 7524 5057 7532 5063
rect 84 5037 236 5043
rect 356 5037 604 5043
rect 756 5037 908 5043
rect 1108 5037 1420 5043
rect 1444 5037 1548 5043
rect 1588 5037 1772 5043
rect 1780 5037 1852 5043
rect 2148 5037 2412 5043
rect 2484 5037 2716 5043
rect 3156 5037 3244 5043
rect 3252 5037 3340 5043
rect 4564 5037 4588 5043
rect 4596 5037 6700 5043
rect 6868 5037 7244 5043
rect 196 5017 300 5023
rect 1060 5017 1260 5023
rect 1284 5017 2140 5023
rect 2452 5017 2700 5023
rect 2724 5017 2972 5023
rect 5652 5017 5740 5023
rect 5748 5017 6028 5023
rect 6292 5017 6364 5023
rect 6372 5017 6412 5023
rect 6420 5017 6460 5023
rect 6468 5017 6492 5023
rect 7028 5017 7132 5023
rect 7204 5017 7244 5023
rect 7252 5017 7388 5023
rect 7396 5017 7500 5023
rect 2242 5014 2302 5016
rect 2242 5006 2243 5014
rect 2252 5006 2253 5014
rect 2291 5006 2292 5014
rect 2301 5006 2302 5014
rect 2242 5004 2302 5006
rect 5250 5014 5310 5016
rect 5250 5006 5251 5014
rect 5260 5006 5261 5014
rect 5299 5006 5300 5014
rect 5309 5006 5310 5014
rect 5250 5004 5310 5006
rect 932 4997 1228 5003
rect 1716 4997 1884 5003
rect 2500 4997 3548 5003
rect 3556 4997 3596 5003
rect 3604 4997 3676 5003
rect 3684 4997 3724 5003
rect 4964 4997 4988 5003
rect 5924 4997 5980 5003
rect 6100 4997 6188 5003
rect 7316 4997 7452 5003
rect 420 4977 1011 4983
rect 1005 4964 1011 4977
rect 1172 4977 1612 4983
rect 1620 4977 1788 4983
rect 1796 4977 2044 4983
rect 2573 4977 2780 4983
rect 2573 4964 2579 4977
rect 2900 4977 2924 4983
rect 2932 4977 3004 4983
rect 3124 4977 3148 4983
rect 3348 4977 3420 4983
rect 3428 4977 3756 4983
rect 4180 4977 4492 4983
rect 4900 4977 4972 4983
rect 5012 4977 5372 4983
rect 5876 4977 6108 4983
rect 6116 4977 6188 4983
rect 6356 4977 6428 4983
rect 6452 4977 6636 4983
rect 7204 4977 7340 4983
rect 84 4957 236 4963
rect 1012 4957 1532 4963
rect 1668 4957 1724 4963
rect 2388 4957 2460 4963
rect 2468 4957 2572 4963
rect 2772 4957 3036 4963
rect 3044 4957 3084 4963
rect 3092 4957 3356 4963
rect 3796 4957 3900 4963
rect 3972 4957 4236 4963
rect 4868 4957 5020 4963
rect 5028 4957 5164 4963
rect 5572 4957 5612 4963
rect 6372 4957 6396 4963
rect 6564 4957 6620 4963
rect 6900 4957 6940 4963
rect 6948 4957 7004 4963
rect 7012 4957 7100 4963
rect 7236 4957 7484 4963
rect 7540 4957 7564 4963
rect 196 4937 268 4943
rect 276 4937 380 4943
rect 388 4937 476 4943
rect 628 4937 716 4943
rect 724 4937 876 4943
rect 884 4937 940 4943
rect 1124 4937 1180 4943
rect 1220 4937 1404 4943
rect 1412 4937 1532 4943
rect 1732 4937 2492 4943
rect 2500 4937 2764 4943
rect 2788 4937 2940 4943
rect 3204 4937 3292 4943
rect 3300 4937 3516 4943
rect 3524 4937 3628 4943
rect 3732 4937 4060 4943
rect 4148 4937 4300 4943
rect 4308 4937 4348 4943
rect 4356 4937 4396 4943
rect 4404 4937 4588 4943
rect 4804 4937 5196 4943
rect 5236 4937 5340 4943
rect 5348 4937 5628 4943
rect 5780 4937 5804 4943
rect 5812 4937 5836 4943
rect 5844 4937 5852 4943
rect 5956 4937 6076 4943
rect 6292 4937 6412 4943
rect 6420 4937 6492 4943
rect 6500 4937 6636 4943
rect 6644 4937 6684 4943
rect 7012 4937 7052 4943
rect 7060 4937 7116 4943
rect 7508 4937 7532 4943
rect 228 4917 300 4923
rect 324 4917 428 4923
rect 772 4917 924 4923
rect 1028 4917 1075 4923
rect 1069 4904 1075 4917
rect 1140 4917 1292 4923
rect 1492 4917 1580 4923
rect 1668 4917 1820 4923
rect 2052 4917 2108 4923
rect 2116 4917 2124 4923
rect 2132 4917 2156 4923
rect 2356 4917 2364 4923
rect 2452 4917 2524 4923
rect 2628 4917 2668 4923
rect 2900 4917 2972 4923
rect 3236 4917 3500 4923
rect 3588 4917 3740 4923
rect 3956 4917 4028 4923
rect 4036 4917 4076 4923
rect 4084 4917 4172 4923
rect 5060 4917 5388 4923
rect 5604 4917 5660 4923
rect 5668 4917 5708 4923
rect 5716 4917 5804 4923
rect 6148 4917 6204 4923
rect 6324 4917 6364 4923
rect 6468 4917 6604 4923
rect 6612 4917 6652 4923
rect 6708 4917 6908 4923
rect 6916 4917 6956 4923
rect 7076 4917 7148 4923
rect 7476 4917 7516 4923
rect 580 4897 812 4903
rect 1076 4897 1148 4903
rect 1348 4897 1516 4903
rect 1764 4897 1948 4903
rect 1956 4897 1980 4903
rect 1988 4897 2076 4903
rect 3844 4897 3916 4903
rect 3924 4897 3996 4903
rect 4116 4897 4428 4903
rect 4884 4897 5148 4903
rect 5156 4897 5612 4903
rect 5636 4897 5740 4903
rect 6244 4897 6428 4903
rect 6596 4897 6860 4903
rect 6868 4897 7020 4903
rect 7028 4897 7068 4903
rect 7508 4897 7548 4903
rect 756 4877 828 4883
rect 1940 4877 1964 4883
rect 1972 4877 2348 4883
rect 2596 4877 3132 4883
rect 3140 4877 3228 4883
rect 3236 4877 3404 4883
rect 3636 4877 3980 4883
rect 4052 4877 4620 4883
rect 5076 4877 5484 4883
rect 5492 4877 5564 4883
rect 7396 4877 7436 4883
rect 308 4857 1628 4863
rect 2228 4857 3932 4863
rect 4004 4857 4124 4863
rect 4916 4857 5884 4863
rect 6669 4857 7420 4863
rect 6669 4844 6675 4857
rect 660 4837 684 4843
rect 692 4837 892 4843
rect 3316 4837 3452 4843
rect 3572 4837 6060 4843
rect 500 4817 556 4823
rect 564 4817 700 4823
rect 868 4817 1020 4823
rect 1204 4817 3724 4823
rect 5220 4817 5500 4823
rect 5524 4817 5676 4823
rect 5812 4817 5996 4823
rect 738 4814 798 4816
rect 738 4806 739 4814
rect 748 4806 749 4814
rect 787 4806 788 4814
rect 797 4806 798 4814
rect 738 4804 798 4806
rect 3746 4814 3806 4816
rect 3746 4806 3747 4814
rect 3756 4806 3757 4814
rect 3795 4806 3796 4814
rect 3805 4806 3806 4814
rect 3746 4804 3806 4806
rect 6754 4814 6814 4816
rect 6754 4806 6755 4814
rect 6764 4806 6765 4814
rect 6803 4806 6804 4814
rect 6813 4806 6814 4814
rect 6754 4804 6814 4806
rect 612 4797 684 4803
rect 1588 4797 1676 4803
rect 2564 4797 2620 4803
rect 2660 4797 2700 4803
rect 2916 4797 3020 4803
rect 3028 4797 3612 4803
rect 3620 4797 3628 4803
rect 4372 4797 4588 4803
rect 4596 4797 4972 4803
rect 5316 4797 5548 4803
rect 5684 4797 5692 4803
rect 6964 4797 7468 4803
rect 708 4777 1340 4783
rect 1348 4777 1596 4783
rect 1604 4777 1804 4783
rect 1812 4777 1948 4783
rect 1956 4777 2060 4783
rect 2100 4777 2236 4783
rect 2589 4777 3507 4783
rect 116 4757 204 4763
rect 500 4757 1212 4763
rect 2589 4763 2595 4777
rect 1556 4757 2595 4763
rect 2612 4757 2956 4763
rect 3501 4763 3507 4777
rect 3524 4777 3644 4783
rect 3652 4777 3836 4783
rect 4196 4777 4252 4783
rect 4260 4777 4364 4783
rect 4756 4777 4988 4783
rect 4996 4777 6076 4783
rect 6084 4777 7100 4783
rect 3501 4757 3708 4763
rect 3725 4757 3948 4763
rect 356 4737 412 4743
rect 420 4737 572 4743
rect 580 4737 860 4743
rect 916 4737 1116 4743
rect 1572 4737 1868 4743
rect 1908 4737 2188 4743
rect 2580 4737 2684 4743
rect 3172 4737 3292 4743
rect 3309 4737 3580 4743
rect 468 4717 700 4723
rect 820 4717 860 4723
rect 868 4717 1308 4723
rect 1316 4717 1356 4723
rect 1524 4717 1708 4723
rect 3309 4723 3315 4737
rect 3725 4743 3731 4757
rect 3956 4757 4092 4763
rect 4132 4757 4204 4763
rect 4980 4757 5052 4763
rect 5204 4757 5996 4763
rect 7188 4757 7196 4763
rect 7284 4757 7516 4763
rect 3700 4737 3731 4743
rect 3828 4737 4067 4743
rect 1844 4717 3315 4723
rect 3332 4717 3356 4723
rect 3396 4717 3452 4723
rect 3508 4717 3948 4723
rect 4061 4723 4067 4737
rect 4084 4737 4588 4743
rect 4596 4737 6035 4743
rect 6029 4724 6035 4737
rect 6388 4737 6604 4743
rect 6612 4737 6956 4743
rect 7108 4737 7212 4743
rect 7252 4737 7276 4743
rect 4061 4717 4108 4723
rect 4164 4717 4252 4723
rect 4756 4717 4796 4723
rect 5044 4717 5420 4723
rect 5428 4717 5724 4723
rect 5732 4717 5804 4723
rect 5812 4717 5980 4723
rect 6036 4717 6259 4723
rect 372 4697 460 4703
rect 564 4697 604 4703
rect 644 4697 716 4703
rect 740 4697 844 4703
rect 900 4697 1004 4703
rect 1156 4697 1164 4703
rect 1364 4697 1452 4703
rect 1572 4697 1644 4703
rect 1828 4697 1916 4703
rect 1972 4697 2044 4703
rect 2068 4697 2172 4703
rect 2180 4697 3404 4703
rect 3412 4697 3436 4703
rect 3732 4697 3868 4703
rect 3876 4697 4092 4703
rect 4100 4697 4172 4703
rect 4212 4697 4444 4703
rect 4740 4697 4780 4703
rect 5005 4697 5148 4703
rect 5005 4684 5011 4697
rect 5172 4697 5228 4703
rect 5508 4697 5532 4703
rect 5556 4697 5628 4703
rect 5636 4697 5756 4703
rect 5780 4697 5836 4703
rect 6116 4697 6220 4703
rect 6253 4703 6259 4717
rect 6500 4717 6556 4723
rect 6676 4717 6732 4723
rect 6852 4717 6924 4723
rect 7140 4717 7196 4723
rect 7204 4717 7356 4723
rect 7412 4717 7420 4723
rect 7444 4717 7516 4723
rect 6253 4697 6508 4703
rect 6516 4697 6556 4703
rect 6660 4697 6716 4703
rect 6740 4697 6876 4703
rect 6964 4697 7052 4703
rect 7156 4697 7260 4703
rect 7412 4697 7468 4703
rect 132 4677 268 4683
rect 452 4677 524 4683
rect 628 4677 668 4683
rect 916 4677 1372 4683
rect 1476 4677 1644 4683
rect 1780 4677 1932 4683
rect 1972 4677 1996 4683
rect 2036 4677 2156 4683
rect 2228 4677 2284 4683
rect 2292 4677 2716 4683
rect 3124 4677 3164 4683
rect 3476 4677 3548 4683
rect 3556 4677 3596 4683
rect 3604 4677 3676 4683
rect 3780 4677 3980 4683
rect 3988 4677 4220 4683
rect 4916 4677 4972 4683
rect 4980 4677 5004 4683
rect 5108 4677 5212 4683
rect 5396 4677 5660 4683
rect 5668 4677 5788 4683
rect 5796 4677 5900 4683
rect 6068 4677 6284 4683
rect 6548 4677 6620 4683
rect 6628 4677 7020 4683
rect 7028 4677 7180 4683
rect 7188 4677 7276 4683
rect 7380 4677 7436 4683
rect 196 4657 572 4663
rect 836 4657 924 4663
rect 948 4657 972 4663
rect 1060 4657 1132 4663
rect 1581 4657 1660 4663
rect 1581 4644 1587 4657
rect 1668 4657 1788 4663
rect 1860 4657 1916 4663
rect 1924 4657 1980 4663
rect 1988 4657 2108 4663
rect 2516 4657 2556 4663
rect 2596 4657 2684 4663
rect 2708 4657 2860 4663
rect 3156 4657 3196 4663
rect 3332 4657 3372 4663
rect 3604 4657 3660 4663
rect 3892 4657 4972 4663
rect 4980 4657 5036 4663
rect 5140 4657 5244 4663
rect 5444 4657 5740 4663
rect 6020 4657 6380 4663
rect 6708 4657 6892 4663
rect 6900 4657 7068 4663
rect 7076 4657 7212 4663
rect 7220 4657 7324 4663
rect 7332 4657 7340 4663
rect 7348 4657 7404 4663
rect 7460 4657 7500 4663
rect 340 4637 396 4643
rect 436 4637 556 4643
rect 708 4637 908 4643
rect 932 4637 1084 4643
rect 1124 4637 1164 4643
rect 1396 4637 1580 4643
rect 1620 4637 2892 4643
rect 2900 4637 2940 4643
rect 2948 4637 3500 4643
rect 3508 4637 3580 4643
rect 4068 4637 4588 4643
rect 4596 4637 4620 4643
rect 4628 4637 4908 4643
rect 4916 4637 5196 4643
rect 5204 4637 5228 4643
rect 6196 4637 6236 4643
rect 6916 4637 6956 4643
rect 6964 4637 7116 4643
rect 7172 4637 7420 4643
rect 964 4617 1548 4623
rect 1652 4617 1772 4623
rect 1908 4617 2012 4623
rect 2068 4617 2140 4623
rect 2516 4617 2604 4623
rect 2644 4617 3260 4623
rect 3268 4617 3340 4623
rect 3348 4617 3388 4623
rect 3412 4617 3468 4623
rect 4660 4617 4716 4623
rect 4724 4617 4796 4623
rect 4964 4617 5212 4623
rect 5620 4617 5932 4623
rect 6772 4617 6924 4623
rect 2242 4614 2302 4616
rect 2242 4606 2243 4614
rect 2252 4606 2253 4614
rect 2291 4606 2292 4614
rect 2301 4606 2302 4614
rect 2242 4604 2302 4606
rect 5250 4614 5310 4616
rect 5250 4606 5251 4614
rect 5260 4606 5261 4614
rect 5299 4606 5300 4614
rect 5309 4606 5310 4614
rect 5250 4604 5310 4606
rect 564 4597 988 4603
rect 1012 4597 1148 4603
rect 1332 4597 1468 4603
rect 1476 4597 1548 4603
rect 2404 4597 2540 4603
rect 2628 4597 3452 4603
rect 4852 4597 5132 4603
rect 5396 4597 5564 4603
rect 5780 4597 5948 4603
rect 7220 4597 7308 4603
rect 7428 4597 7484 4603
rect 164 4577 236 4583
rect 244 4577 1356 4583
rect 1396 4577 1436 4583
rect 1444 4577 1564 4583
rect 1748 4577 1820 4583
rect 1876 4577 1980 4583
rect 2132 4577 2316 4583
rect 2580 4577 2668 4583
rect 3220 4577 3532 4583
rect 3540 4577 3612 4583
rect 4676 4577 4764 4583
rect 4772 4577 4780 4583
rect 4804 4577 5036 4583
rect 5172 4577 5196 4583
rect 5220 4577 5372 4583
rect 5428 4577 5708 4583
rect 5860 4577 6028 4583
rect 6068 4577 6236 4583
rect 6276 4577 6396 4583
rect 6436 4577 6492 4583
rect 7076 4577 7180 4583
rect 7252 4577 7372 4583
rect 20 4557 188 4563
rect 564 4557 668 4563
rect 996 4557 1228 4563
rect 1556 4557 1612 4563
rect 1716 4557 1772 4563
rect 1812 4557 2060 4563
rect 2164 4557 2268 4563
rect 2276 4557 2508 4563
rect 2516 4557 2524 4563
rect 2564 4557 2604 4563
rect 2612 4557 2668 4563
rect 2724 4557 3868 4563
rect 4196 4557 4284 4563
rect 4324 4557 4396 4563
rect 4404 4557 4540 4563
rect 4548 4557 4556 4563
rect 4772 4557 4828 4563
rect 5012 4557 6124 4563
rect 6141 4557 6284 4563
rect 228 4537 300 4543
rect 340 4537 380 4543
rect 388 4537 396 4543
rect 468 4537 604 4543
rect 804 4537 860 4543
rect 1124 4537 1196 4543
rect 1204 4537 1244 4543
rect 1412 4537 1484 4543
rect 1492 4537 1500 4543
rect 1508 4537 1676 4543
rect 1684 4537 1932 4543
rect 2004 4537 2044 4543
rect 2052 4537 2124 4543
rect 2420 4537 2732 4543
rect 3060 4537 3084 4543
rect 3364 4537 3436 4543
rect 3684 4537 3980 4543
rect 3988 4537 4028 4543
rect 4164 4537 4220 4543
rect 4228 4537 4300 4543
rect 4644 4537 4876 4543
rect 5028 4537 5116 4543
rect 5156 4537 5244 4543
rect 5492 4537 5516 4543
rect 5524 4537 5612 4543
rect 5620 4537 5804 4543
rect 6141 4543 6147 4557
rect 6372 4557 6476 4563
rect 7156 4557 7212 4563
rect 7316 4557 7356 4563
rect 6004 4537 6147 4543
rect 6340 4537 6396 4543
rect 6404 4537 6476 4543
rect 6548 4537 6620 4543
rect 6708 4537 6908 4543
rect 7012 4537 7052 4543
rect 7060 4537 7196 4543
rect 7220 4537 7260 4543
rect 7268 4537 7308 4543
rect 7412 4537 7484 4543
rect 52 4517 92 4523
rect 100 4517 236 4523
rect 244 4517 268 4523
rect 276 4517 284 4523
rect 420 4517 508 4523
rect 548 4517 588 4523
rect 644 4517 860 4523
rect 1028 4517 1116 4523
rect 1140 4517 1148 4523
rect 1172 4517 1244 4523
rect 1252 4517 1308 4523
rect 1364 4517 1500 4523
rect 1540 4517 1612 4523
rect 1652 4517 1740 4523
rect 1780 4517 1804 4523
rect 1901 4517 1964 4523
rect 1901 4504 1907 4517
rect 2020 4517 2076 4523
rect 2212 4517 2428 4523
rect 2516 4517 2540 4523
rect 2692 4517 2764 4523
rect 2852 4517 3228 4523
rect 3412 4517 3436 4523
rect 3572 4517 3724 4523
rect 3940 4517 4092 4523
rect 4276 4517 4412 4523
rect 4580 4517 4588 4523
rect 4820 4517 5004 4523
rect 5012 4517 5036 4523
rect 5188 4517 5260 4523
rect 5412 4517 5516 4523
rect 5524 4517 5676 4523
rect 5908 4517 6060 4523
rect 6084 4517 6092 4523
rect 6164 4517 6188 4523
rect 6388 4517 6444 4523
rect 6477 4517 6572 4523
rect 388 4497 508 4503
rect 516 4497 524 4503
rect 532 4497 1052 4503
rect 1060 4497 1212 4503
rect 1284 4497 1420 4503
rect 1476 4497 1708 4503
rect 1716 4497 1900 4503
rect 1940 4497 2028 4503
rect 2116 4497 2396 4503
rect 2532 4497 2540 4503
rect 2548 4497 2572 4503
rect 2724 4497 2780 4503
rect 2788 4497 2796 4503
rect 2804 4497 2924 4503
rect 3060 4497 3116 4503
rect 3188 4497 3292 4503
rect 3396 4497 3420 4503
rect 4036 4497 4060 4503
rect 4788 4497 4940 4503
rect 4948 4497 5020 4503
rect 5108 4497 5420 4503
rect 5428 4497 5660 4503
rect 5972 4497 6172 4503
rect 6292 4497 6332 4503
rect 6477 4503 6483 4517
rect 6756 4517 6828 4523
rect 6932 4517 6956 4523
rect 7140 4517 7308 4523
rect 7460 4517 7532 4523
rect 6452 4497 6483 4503
rect 6500 4497 6556 4503
rect 6596 4497 6668 4503
rect 6804 4497 6924 4503
rect 6980 4497 7036 4503
rect 7092 4497 7148 4503
rect 7476 4497 7532 4503
rect 708 4477 828 4483
rect 1076 4477 1164 4483
rect 2180 4477 2188 4483
rect 2196 4477 2236 4483
rect 2516 4477 4140 4483
rect 4388 4477 4748 4483
rect 4756 4477 4844 4483
rect 4852 4477 5340 4483
rect 5348 4477 5388 4483
rect 5476 4477 5548 4483
rect 5556 4477 5580 4483
rect 5588 4477 5644 4483
rect 5652 4477 5868 4483
rect 6020 4477 6076 4483
rect 6100 4477 6204 4483
rect 6468 4477 6572 4483
rect 6660 4477 6796 4483
rect 6804 4477 6908 4483
rect 6948 4477 6988 4483
rect 356 4457 396 4463
rect 701 4463 707 4476
rect 452 4457 707 4463
rect 1300 4457 1548 4463
rect 1556 4457 2156 4463
rect 2164 4457 2252 4463
rect 2340 4457 2700 4463
rect 2708 4457 2828 4463
rect 2932 4457 3260 4463
rect 3268 4457 3340 4463
rect 3348 4457 3644 4463
rect 3860 4457 4076 4463
rect 4244 4457 4620 4463
rect 4628 4457 5436 4463
rect 6228 4457 6380 4463
rect 6532 4457 6636 4463
rect 6644 4457 6988 4463
rect 964 4437 1196 4443
rect 1204 4437 1388 4443
rect 1860 4437 2508 4443
rect 2525 4437 3116 4443
rect 2525 4424 2531 4437
rect 3140 4437 3372 4443
rect 3492 4437 3580 4443
rect 3725 4437 3868 4443
rect 852 4417 1804 4423
rect 2100 4417 2332 4423
rect 2516 4417 2524 4423
rect 2612 4417 2620 4423
rect 2660 4417 2988 4423
rect 3204 4417 3260 4423
rect 3725 4423 3731 4437
rect 4564 4437 4940 4443
rect 4948 4437 6220 4443
rect 6228 4437 7020 4443
rect 3332 4417 3731 4423
rect 4436 4417 4700 4423
rect 5684 4417 5884 4423
rect 6500 4417 6540 4423
rect 6596 4417 6684 4423
rect 738 4414 798 4416
rect 738 4406 739 4414
rect 748 4406 749 4414
rect 787 4406 788 4414
rect 797 4406 798 4414
rect 738 4404 798 4406
rect 3746 4414 3806 4416
rect 3746 4406 3747 4414
rect 3756 4406 3757 4414
rect 3795 4406 3796 4414
rect 3805 4406 3806 4414
rect 3746 4404 3806 4406
rect 6754 4414 6814 4416
rect 6754 4406 6755 4414
rect 6764 4406 6765 4414
rect 6803 4406 6804 4414
rect 6813 4406 6814 4414
rect 6754 4404 6814 4406
rect 1028 4397 1660 4403
rect 1748 4397 3731 4403
rect 564 4377 1756 4383
rect 3725 4383 3731 4397
rect 4052 4397 4956 4403
rect 5364 4397 5772 4403
rect 5780 4397 5916 4403
rect 2813 4377 3715 4383
rect 3725 4377 4012 4383
rect 468 4357 812 4363
rect 916 4357 1068 4363
rect 2813 4363 2819 4377
rect 1652 4357 2819 4363
rect 2836 4357 3148 4363
rect 3156 4357 3196 4363
rect 3412 4357 3468 4363
rect 3709 4363 3715 4377
rect 4884 4377 4924 4383
rect 5412 4377 5452 4383
rect 5572 4377 5612 4383
rect 5732 4377 5964 4383
rect 6644 4377 6828 4383
rect 6836 4377 6876 4383
rect 3709 4357 4204 4363
rect 4756 4357 4812 4363
rect 5444 4357 5772 4363
rect 5844 4357 5948 4363
rect 6436 4357 6844 4363
rect 404 4337 636 4343
rect 692 4337 732 4343
rect 868 4337 908 4343
rect 1188 4337 1324 4343
rect 1460 4337 1484 4343
rect 1524 4337 1612 4343
rect 2404 4337 2460 4343
rect 2772 4337 3084 4343
rect 3188 4337 3724 4343
rect 4836 4337 4908 4343
rect 4980 4337 5084 4343
rect 5172 4337 5868 4343
rect 6036 4337 6156 4343
rect 6468 4337 7052 4343
rect 7156 4337 7292 4343
rect 436 4317 860 4323
rect 1268 4317 1516 4323
rect 1524 4317 2684 4323
rect 3188 4317 3228 4323
rect 3236 4317 3500 4323
rect 3508 4317 3612 4323
rect 3716 4317 3820 4323
rect 4180 4317 4444 4323
rect 4692 4317 5452 4323
rect 5556 4317 5724 4323
rect 5828 4317 5852 4323
rect 6036 4317 6060 4323
rect 6068 4317 6140 4323
rect 6276 4317 6316 4323
rect 6356 4317 6604 4323
rect 6612 4317 6700 4323
rect 6772 4317 6844 4323
rect 6852 4317 6924 4323
rect 7028 4317 7180 4323
rect 7236 4317 7276 4323
rect 7380 4317 7436 4323
rect 228 4297 300 4303
rect 388 4297 428 4303
rect 788 4297 1020 4303
rect 1380 4297 1868 4303
rect 1876 4297 2060 4303
rect 2100 4297 2172 4303
rect 2356 4297 2428 4303
rect 2516 4297 2556 4303
rect 2756 4297 2812 4303
rect 2820 4297 2844 4303
rect 2884 4297 3011 4303
rect 84 4277 236 4283
rect 372 4277 524 4283
rect 772 4277 876 4283
rect 1172 4277 1196 4283
rect 1220 4277 1260 4283
rect 1268 4277 1276 4283
rect 1460 4277 1532 4283
rect 1588 4277 1628 4283
rect 2052 4277 2364 4283
rect 2420 4277 2460 4283
rect 2484 4277 2572 4283
rect 2644 4277 2668 4283
rect 2804 4277 2844 4283
rect 2900 4277 2956 4283
rect 3005 4283 3011 4297
rect 3028 4297 3804 4303
rect 4036 4297 4284 4303
rect 4292 4297 4300 4303
rect 4308 4297 4332 4303
rect 4372 4297 4428 4303
rect 4612 4297 4652 4303
rect 4788 4297 4860 4303
rect 4900 4297 5100 4303
rect 5108 4297 5148 4303
rect 5172 4297 6284 4303
rect 6532 4297 6556 4303
rect 6852 4297 6860 4303
rect 6996 4297 7084 4303
rect 7348 4297 7404 4303
rect 7453 4297 7500 4303
rect 3005 4277 3036 4283
rect 3396 4277 3420 4283
rect 3476 4277 3564 4283
rect 3629 4277 3676 4283
rect 196 4257 268 4263
rect 276 4257 380 4263
rect 420 4257 428 4263
rect 436 4257 668 4263
rect 804 4257 828 4263
rect 980 4257 1052 4263
rect 1076 4257 1324 4263
rect 1396 4257 1500 4263
rect 1508 4257 1548 4263
rect 1940 4257 2076 4263
rect 2100 4257 2348 4263
rect 2436 4257 2460 4263
rect 2484 4257 2524 4263
rect 2596 4257 2732 4263
rect 2820 4257 3004 4263
rect 3156 4257 3196 4263
rect 3421 4263 3427 4276
rect 3421 4257 3516 4263
rect 3629 4263 3635 4277
rect 4372 4277 4460 4283
rect 4468 4277 4604 4283
rect 4612 4277 4636 4283
rect 4756 4277 4780 4283
rect 5028 4277 5084 4283
rect 5140 4277 5212 4283
rect 5252 4277 6012 4283
rect 6036 4277 6172 4283
rect 6212 4277 6348 4283
rect 6452 4277 6508 4283
rect 6724 4277 6860 4283
rect 6916 4277 7091 4283
rect 7085 4264 7091 4277
rect 7172 4277 7228 4283
rect 7236 4277 7260 4283
rect 7268 4277 7292 4283
rect 7300 4277 7372 4283
rect 7412 4277 7436 4283
rect 3556 4257 3635 4263
rect 3652 4257 3724 4263
rect 4308 4257 4524 4263
rect 4532 4257 4572 4263
rect 4580 4257 4700 4263
rect 5156 4257 5356 4263
rect 5636 4257 5676 4263
rect 5940 4257 5996 4263
rect 6196 4257 6252 4263
rect 6420 4257 6556 4263
rect 6564 4257 6668 4263
rect 6676 4257 6812 4263
rect 6868 4257 7052 4263
rect 7092 4257 7132 4263
rect 7453 4263 7459 4297
rect 7444 4257 7459 4263
rect 7476 4257 7516 4263
rect 356 4237 572 4243
rect 868 4237 908 4243
rect 916 4237 1356 4243
rect 1364 4237 1532 4243
rect 1572 4237 1980 4243
rect 1988 4237 2188 4243
rect 2548 4237 3052 4243
rect 3492 4237 3596 4243
rect 4068 4237 4108 4243
rect 4308 4237 4364 4243
rect 5076 4237 5436 4243
rect 6020 4237 6236 4243
rect 6484 4237 6540 4243
rect 6548 4237 6604 4243
rect 6836 4237 6892 4243
rect 340 4217 476 4223
rect 532 4217 540 4223
rect 628 4217 828 4223
rect 836 4217 876 4223
rect 1060 4217 1100 4223
rect 1172 4217 1292 4223
rect 1300 4217 1596 4223
rect 1604 4217 1692 4223
rect 1700 4217 1788 4223
rect 1892 4217 1996 4223
rect 2004 4217 2140 4223
rect 2500 4217 3107 4223
rect 2242 4214 2302 4216
rect 2242 4206 2243 4214
rect 2252 4206 2253 4214
rect 2291 4206 2292 4214
rect 2301 4206 2302 4214
rect 2242 4204 2302 4206
rect 500 4197 588 4203
rect 596 4197 908 4203
rect 916 4197 956 4203
rect 964 4197 1628 4203
rect 1684 4197 1788 4203
rect 2020 4197 2108 4203
rect 2580 4197 2796 4203
rect 2804 4197 2828 4203
rect 2836 4197 3084 4203
rect 3101 4203 3107 4217
rect 3124 4217 4316 4223
rect 4548 4217 5100 4223
rect 5428 4217 6012 4223
rect 6020 4217 6156 4223
rect 6356 4217 6492 4223
rect 5250 4214 5310 4216
rect 5250 4206 5251 4214
rect 5260 4206 5261 4214
rect 5299 4206 5300 4214
rect 5309 4206 5310 4214
rect 5250 4204 5310 4206
rect 3101 4197 3404 4203
rect 3908 4197 3948 4203
rect 3956 4197 4092 4203
rect 4516 4197 4556 4203
rect 4564 4197 4988 4203
rect 4996 4197 5164 4203
rect 5812 4197 6124 4203
rect 6196 4197 6252 4203
rect 6260 4197 6508 4203
rect 6548 4197 6572 4203
rect 6580 4197 6620 4203
rect 6836 4197 7116 4203
rect 7124 4197 7180 4203
rect 7188 4197 7276 4203
rect 7284 4197 7340 4203
rect 356 4177 492 4183
rect 500 4177 652 4183
rect 660 4177 684 4183
rect 804 4177 876 4183
rect 1604 4177 1836 4183
rect 2100 4177 2124 4183
rect 2132 4177 2236 4183
rect 2452 4177 2476 4183
rect 2484 4177 2588 4183
rect 3588 4177 3772 4183
rect 3972 4177 3996 4183
rect 4388 4177 4748 4183
rect 4980 4177 5036 4183
rect 5236 4177 5260 4183
rect 5300 4177 5324 4183
rect 5700 4177 5788 4183
rect 5844 4177 6076 4183
rect 6116 4177 6124 4183
rect 6228 4177 6252 4183
rect 6356 4177 6700 4183
rect 6868 4177 7020 4183
rect 7348 4177 7372 4183
rect 7421 4177 7500 4183
rect 196 4157 268 4163
rect 276 4157 332 4163
rect 372 4157 604 4163
rect 612 4157 652 4163
rect 804 4157 892 4163
rect 1620 4157 1660 4163
rect 1828 4157 1900 4163
rect 2196 4157 2220 4163
rect 2548 4157 2572 4163
rect 2580 4157 3020 4163
rect 3092 4157 3276 4163
rect 3284 4157 3484 4163
rect 4020 4157 4044 4163
rect 4084 4157 4140 4163
rect 4356 4157 4476 4163
rect 4836 4157 4972 4163
rect 4980 4157 5228 4163
rect 5236 4157 5340 4163
rect 5380 4157 5484 4163
rect 5492 4157 5548 4163
rect 5556 4157 5644 4163
rect 5716 4157 5804 4163
rect 6260 4157 6380 4163
rect 6948 4157 7004 4163
rect 7252 4157 7308 4163
rect 7421 4163 7427 4177
rect 7412 4157 7427 4163
rect 7444 4157 7452 4163
rect 7460 4157 7500 4163
rect 7524 4157 7548 4163
rect 228 4137 307 4143
rect 301 4124 307 4137
rect 820 4137 924 4143
rect 948 4137 1004 4143
rect 1300 4137 1404 4143
rect 1540 4137 1580 4143
rect 1684 4137 1756 4143
rect 1812 4137 1948 4143
rect 2756 4137 2908 4143
rect 3332 4137 3612 4143
rect 3924 4137 3996 4143
rect 4004 4137 4044 4143
rect 4196 4137 4284 4143
rect 4292 4137 4380 4143
rect 4388 4137 4412 4143
rect 4436 4137 5036 4143
rect 5108 4137 5308 4143
rect 5341 4143 5347 4156
rect 5341 4137 5500 4143
rect 5540 4137 5612 4143
rect 5668 4137 5740 4143
rect 5748 4137 5820 4143
rect 5828 4137 5852 4143
rect 6148 4137 6284 4143
rect 6308 4137 6332 4143
rect 6724 4137 7356 4143
rect 7364 4137 7420 4143
rect 7428 4137 7500 4143
rect 84 4117 236 4123
rect 308 4117 332 4123
rect 580 4117 620 4123
rect 884 4117 956 4123
rect 964 4117 1004 4123
rect 1204 4117 1292 4123
rect 1476 4117 1740 4123
rect 1940 4117 2028 4123
rect 2036 4117 2092 4123
rect 2132 4117 2348 4123
rect 2404 4117 2780 4123
rect 3028 4117 3244 4123
rect 3300 4117 3340 4123
rect 3556 4117 3644 4123
rect 3700 4117 3836 4123
rect 3844 4117 3852 4123
rect 4132 4117 4172 4123
rect 4180 4117 4332 4123
rect 4564 4117 4732 4123
rect 5060 4117 5116 4123
rect 5316 4117 5388 4123
rect 5652 4117 5692 4123
rect 5716 4117 5756 4123
rect 5764 4117 5820 4123
rect 6132 4117 6140 4123
rect 6436 4117 6892 4123
rect 7220 4117 7292 4123
rect 7380 4117 7452 4123
rect 484 4097 572 4103
rect 692 4097 764 4103
rect 852 4097 924 4103
rect 996 4097 1196 4103
rect 1204 4097 1740 4103
rect 1748 4097 2460 4103
rect 2516 4097 2556 4103
rect 2964 4097 3036 4103
rect 3508 4097 3548 4103
rect 3892 4097 3964 4103
rect 3972 4097 4140 4103
rect 4148 4097 4268 4103
rect 4276 4097 4300 4103
rect 5428 4097 5532 4103
rect 5636 4097 5708 4103
rect 5748 4097 6188 4103
rect 6196 4097 6284 4103
rect 6292 4097 6396 4103
rect 6820 4097 6860 4103
rect 6868 4097 6924 4103
rect 6996 4097 7052 4103
rect 7460 4097 7484 4103
rect 7492 4097 7548 4103
rect 212 4077 812 4083
rect 932 4077 1452 4083
rect 1684 4077 1708 4083
rect 1732 4077 1836 4083
rect 1860 4077 2140 4083
rect 2436 4077 2508 4083
rect 2564 4077 2700 4083
rect 4084 4077 4236 4083
rect 4244 4077 5004 4083
rect 5076 4077 5180 4083
rect 5188 4077 5212 4083
rect 5460 4077 6732 4083
rect 7396 4077 7484 4083
rect 7524 4077 7548 4083
rect 676 4057 1036 4063
rect 1044 4057 1180 4063
rect 1396 4057 1436 4063
rect 1492 4057 4028 4063
rect 5069 4063 5075 4076
rect 4868 4057 5075 4063
rect 5508 4057 5804 4063
rect 564 4037 716 4043
rect 724 4037 1260 4043
rect 1444 4037 2163 4043
rect 1380 4017 1532 4023
rect 2157 4023 2163 4037
rect 2180 4037 2572 4043
rect 2580 4037 3292 4043
rect 3396 4037 3404 4043
rect 3725 4037 3900 4043
rect 3725 4023 3731 4037
rect 5492 4037 6012 4043
rect 6020 4037 6028 4043
rect 7140 4037 7228 4043
rect 7412 4037 7500 4043
rect 1540 4017 1987 4023
rect 2157 4017 3731 4023
rect 738 4014 798 4016
rect 738 4006 739 4014
rect 748 4006 749 4014
rect 787 4006 788 4014
rect 797 4006 798 4014
rect 738 4004 798 4006
rect 1284 3997 1484 4003
rect 1492 3997 1852 4003
rect 1876 3997 1964 4003
rect 1981 4003 1987 4017
rect 5076 4017 5580 4023
rect 5588 4017 5868 4023
rect 5876 4017 6028 4023
rect 3746 4014 3806 4016
rect 3746 4006 3747 4014
rect 3756 4006 3757 4014
rect 3795 4006 3796 4014
rect 3805 4006 3806 4014
rect 3746 4004 3806 4006
rect 6754 4014 6814 4016
rect 6754 4006 6755 4014
rect 6764 4006 6765 4014
rect 6803 4006 6804 4014
rect 6813 4006 6814 4014
rect 6754 4004 6814 4006
rect 1981 3997 2044 4003
rect 2052 3997 3132 4003
rect 4276 3997 4396 4003
rect 4669 3997 5692 4003
rect 4669 3984 4675 3997
rect 5700 3997 5740 4003
rect 5908 3997 6316 4003
rect 868 3977 956 3983
rect 1332 3977 1516 3983
rect 1636 3977 1788 3983
rect 2148 3977 2332 3983
rect 2356 3977 2812 3983
rect 2820 3977 2988 3983
rect 3060 3977 3196 3983
rect 4132 3977 4668 3983
rect 4916 3977 4972 3983
rect 5012 3977 5036 3983
rect 5204 3977 5388 3983
rect 5396 3977 5644 3983
rect 6244 3977 6684 3983
rect 6692 3977 6748 3983
rect 1156 3957 1420 3963
rect 1428 3957 2396 3963
rect 2676 3957 3036 3963
rect 3860 3957 4012 3963
rect 4020 3957 4204 3963
rect 4212 3957 4236 3963
rect 4244 3957 4284 3963
rect 4292 3957 4364 3963
rect 4468 3957 4492 3963
rect 4628 3957 4652 3963
rect 6237 3963 6243 3976
rect 4948 3957 6243 3963
rect 276 3937 1116 3943
rect 1300 3937 1356 3943
rect 1524 3937 1548 3943
rect 1588 3937 1612 3943
rect 1620 3937 1772 3943
rect 2228 3937 2396 3943
rect 2612 3937 2668 3943
rect 2676 3937 2940 3943
rect 2948 3937 2972 3943
rect 3188 3937 3244 3943
rect 3764 3937 4124 3943
rect 4148 3937 4172 3943
rect 4180 3937 4476 3943
rect 4484 3937 4652 3943
rect 4740 3937 5020 3943
rect 5124 3937 5212 3943
rect 5348 3937 5820 3943
rect 5828 3937 5884 3943
rect 5924 3937 5996 3943
rect 6164 3937 6284 3943
rect 6308 3937 6652 3943
rect 7108 3937 7244 3943
rect 7412 3937 7436 3943
rect 84 3917 252 3923
rect 340 3917 364 3923
rect 548 3917 636 3923
rect 1060 3917 1148 3923
rect 1268 3917 1420 3923
rect 1549 3917 2060 3923
rect 1549 3904 1555 3917
rect 2372 3917 2508 3923
rect 2628 3917 2716 3923
rect 2724 3917 2780 3923
rect 3044 3917 3244 3923
rect 4212 3917 4396 3923
rect 4420 3917 4428 3923
rect 4452 3917 4828 3923
rect 4836 3917 4876 3923
rect 4884 3917 4924 3923
rect 4932 3917 5436 3923
rect 5444 3917 5484 3923
rect 5796 3917 6348 3923
rect 6356 3917 6444 3923
rect 6916 3917 7004 3923
rect 7044 3917 7164 3923
rect 7188 3917 7260 3923
rect 7396 3917 7452 3923
rect 7549 3917 7564 3923
rect 244 3897 284 3903
rect 292 3897 412 3903
rect 420 3897 524 3903
rect 532 3897 620 3903
rect 980 3897 1292 3903
rect 1300 3897 1324 3903
rect 1364 3897 1548 3903
rect 1812 3897 1820 3903
rect 1908 3897 1996 3903
rect 2468 3897 2508 3903
rect 2516 3897 2636 3903
rect 2660 3897 2684 3903
rect 2756 3897 2844 3903
rect 2916 3897 3116 3903
rect 3316 3897 3356 3903
rect 3444 3897 3516 3903
rect 3572 3897 3628 3903
rect 4196 3897 4444 3903
rect 4484 3897 4620 3903
rect 4701 3897 4979 3903
rect 4701 3884 4707 3897
rect 132 3877 332 3883
rect 340 3877 588 3883
rect 916 3877 1036 3883
rect 1060 3877 1484 3883
rect 1524 3877 1644 3883
rect 1828 3877 1932 3883
rect 1940 3877 2012 3883
rect 2164 3877 2700 3883
rect 2932 3877 2988 3883
rect 2996 3877 3148 3883
rect 3220 3877 3324 3883
rect 3332 3877 3388 3883
rect 3540 3877 3820 3883
rect 3844 3877 4092 3883
rect 3917 3864 3923 3877
rect 4100 3877 4156 3883
rect 4356 3877 4540 3883
rect 4644 3877 4700 3883
rect 4868 3877 4876 3883
rect 4916 3877 4956 3883
rect 4973 3883 4979 3897
rect 4996 3897 5004 3903
rect 5044 3897 5084 3903
rect 5364 3897 5500 3903
rect 5780 3897 6140 3903
rect 6148 3897 6268 3903
rect 6500 3897 6716 3903
rect 6900 3897 6940 3903
rect 7028 3897 7100 3903
rect 7108 3897 7148 3903
rect 4973 3877 5100 3883
rect 5108 3877 5228 3883
rect 5636 3877 5708 3883
rect 5940 3877 5980 3883
rect 5988 3877 6124 3883
rect 6244 3877 6371 3883
rect 228 3857 508 3863
rect 516 3857 1116 3863
rect 1124 3857 1468 3863
rect 1476 3857 1644 3863
rect 1700 3857 2188 3863
rect 2196 3857 2252 3863
rect 2260 3857 2364 3863
rect 2564 3857 2764 3863
rect 2772 3857 2780 3863
rect 3044 3857 3308 3863
rect 3572 3857 3868 3863
rect 4404 3857 4572 3863
rect 4580 3857 4844 3863
rect 4852 3857 5068 3863
rect 5188 3857 5404 3863
rect 5428 3857 5548 3863
rect 5556 3857 5692 3863
rect 5732 3857 5772 3863
rect 5844 3857 6252 3863
rect 6365 3863 6371 3877
rect 6388 3877 6412 3883
rect 6516 3877 6668 3883
rect 6868 3877 6908 3883
rect 6916 3877 6924 3883
rect 6932 3877 6956 3883
rect 7172 3877 7196 3883
rect 7220 3877 7276 3883
rect 7316 3877 7340 3883
rect 6365 3857 6380 3863
rect 6500 3857 6556 3863
rect 6564 3857 6684 3863
rect 6980 3857 7356 3863
rect 7380 3857 7436 3863
rect 7444 3857 7500 3863
rect 7549 3863 7555 3917
rect 7572 3897 7603 3903
rect 7540 3857 7555 3863
rect 564 3837 844 3843
rect 1140 3837 1356 3843
rect 2132 3837 2540 3843
rect 2548 3837 2844 3843
rect 3332 3837 3452 3843
rect 3908 3837 5052 3843
rect 5300 3837 5324 3843
rect 5476 3837 5500 3843
rect 5620 3837 5916 3843
rect 5956 3837 6172 3843
rect 6212 3837 6380 3843
rect 7316 3837 7372 3843
rect 868 3817 876 3823
rect 884 3817 1692 3823
rect 1892 3817 2140 3823
rect 2340 3817 2780 3823
rect 2788 3817 3020 3823
rect 3268 3817 3308 3823
rect 4100 3817 4940 3823
rect 5940 3817 6236 3823
rect 6260 3817 6492 3823
rect 2242 3814 2302 3816
rect 2242 3806 2243 3814
rect 2252 3806 2253 3814
rect 2291 3806 2292 3814
rect 2301 3806 2302 3814
rect 2242 3804 2302 3806
rect 5250 3814 5310 3816
rect 5250 3806 5251 3814
rect 5260 3806 5261 3814
rect 5299 3806 5300 3814
rect 5309 3806 5310 3814
rect 5250 3804 5310 3806
rect 324 3797 1132 3803
rect 1236 3797 1340 3803
rect 2724 3797 2812 3803
rect 2820 3797 3324 3803
rect 5325 3797 6412 3803
rect 532 3777 716 3783
rect 724 3777 876 3783
rect 884 3777 924 3783
rect 1236 3777 1420 3783
rect 1428 3777 1852 3783
rect 1860 3777 1948 3783
rect 2164 3777 2252 3783
rect 2452 3777 2636 3783
rect 2644 3777 2748 3783
rect 2884 3777 3132 3783
rect 3140 3777 3212 3783
rect 3220 3777 3340 3783
rect 3508 3777 3612 3783
rect 4468 3777 4636 3783
rect 5325 3783 5331 3797
rect 6420 3797 6572 3803
rect 6580 3797 6668 3803
rect 7268 3797 7340 3803
rect 5044 3777 5331 3783
rect 5524 3777 5580 3783
rect 5972 3777 5996 3783
rect 6020 3777 6604 3783
rect 7204 3777 7308 3783
rect 212 3757 796 3763
rect 948 3757 988 3763
rect 1012 3757 1052 3763
rect 1956 3757 1964 3763
rect 1972 3757 1980 3763
rect 2004 3757 2076 3763
rect 2084 3757 2220 3763
rect 2356 3757 2380 3763
rect 2948 3757 3596 3763
rect 3604 3757 3628 3763
rect 3636 3757 3660 3763
rect 4132 3757 4156 3763
rect 4180 3757 4284 3763
rect 4356 3757 4444 3763
rect 4612 3757 4668 3763
rect 5108 3757 5148 3763
rect 5236 3757 5260 3763
rect 5540 3757 5564 3763
rect 5668 3757 5740 3763
rect 5956 3757 6188 3763
rect 6260 3757 6412 3763
rect 6756 3757 6844 3763
rect 6852 3757 6876 3763
rect 6884 3757 6988 3763
rect 7380 3757 7404 3763
rect 244 3737 268 3743
rect 276 3737 284 3743
rect 308 3737 428 3743
rect 804 3737 1020 3743
rect 1140 3737 1404 3743
rect 1412 3737 1484 3743
rect 1812 3737 1836 3743
rect 1844 3737 2028 3743
rect 2148 3737 2188 3743
rect 2260 3737 2476 3743
rect 2484 3737 2972 3743
rect 3220 3737 3260 3743
rect 3284 3737 3308 3743
rect 3860 3737 3932 3743
rect 4148 3737 4268 3743
rect 4452 3737 4540 3743
rect 4548 3737 4556 3743
rect 4564 3737 4796 3743
rect 4804 3737 5036 3743
rect 5220 3737 5388 3743
rect 5396 3737 5596 3743
rect 5604 3737 5724 3743
rect 5732 3737 5772 3743
rect 6036 3737 6076 3743
rect 6084 3737 6156 3743
rect 6164 3737 6220 3743
rect 6484 3737 6556 3743
rect 6612 3737 6700 3743
rect 6740 3737 6924 3743
rect 6932 3737 7004 3743
rect 7060 3737 7388 3743
rect 7396 3737 7436 3743
rect 7460 3737 7523 3743
rect 84 3717 252 3723
rect 500 3717 588 3723
rect 612 3717 908 3723
rect 1044 3717 1180 3723
rect 1204 3717 1292 3723
rect 1892 3717 1916 3723
rect 2004 3717 2044 3723
rect 2372 3717 2412 3723
rect 2420 3717 2620 3723
rect 2740 3717 2892 3723
rect 2916 3717 3004 3723
rect 3172 3717 3180 3723
rect 3204 3717 3324 3723
rect 3412 3717 3500 3723
rect 3540 3717 3548 3723
rect 3556 3717 3580 3723
rect 4068 3717 4332 3723
rect 4340 3717 4380 3723
rect 4772 3717 4844 3723
rect 5028 3717 5084 3723
rect 5140 3717 5212 3723
rect 5524 3717 5612 3723
rect 5700 3717 5868 3723
rect 5876 3717 5980 3723
rect 6036 3717 6268 3723
rect 6276 3717 6332 3723
rect 6404 3717 6508 3723
rect 6580 3717 6668 3723
rect 6692 3717 6764 3723
rect 6980 3717 7036 3723
rect 7380 3717 7500 3723
rect 244 3697 332 3703
rect 436 3697 492 3703
rect 516 3697 956 3703
rect 1140 3697 1196 3703
rect 1476 3697 1612 3703
rect 1652 3697 1836 3703
rect 1844 3697 1932 3703
rect 2404 3697 2508 3703
rect 2852 3697 2924 3703
rect 3156 3697 3292 3703
rect 3588 3697 3724 3703
rect 4868 3697 5068 3703
rect 5076 3697 5132 3703
rect 5428 3697 5436 3703
rect 5652 3697 6012 3703
rect 6164 3697 6188 3703
rect 6212 3697 6364 3703
rect 6372 3697 6444 3703
rect 6948 3697 7404 3703
rect 7428 3697 7452 3703
rect 7517 3703 7523 3737
rect 7572 3717 7603 3723
rect 7508 3697 7523 3703
rect 7540 3697 7564 3703
rect 500 3677 556 3683
rect 852 3677 924 3683
rect 948 3677 1724 3683
rect 1748 3677 2140 3683
rect 2436 3677 3532 3683
rect 3924 3677 4892 3683
rect 4900 3677 5116 3683
rect 6941 3683 6947 3696
rect 5124 3677 6947 3683
rect 7220 3677 7420 3683
rect 7444 3677 7603 3683
rect 1108 3657 2380 3663
rect 2388 3657 2572 3663
rect 3508 3657 3708 3663
rect 4148 3657 4396 3663
rect 4404 3657 4476 3663
rect 5620 3657 5820 3663
rect 6324 3657 6524 3663
rect 7220 3657 7388 3663
rect 308 3637 348 3643
rect 388 3637 940 3643
rect 1396 3637 2172 3643
rect 3188 3637 3388 3643
rect 3732 3637 4860 3643
rect 5060 3637 6572 3643
rect 6580 3637 6636 3643
rect 6676 3637 7100 3643
rect 7156 3637 7356 3643
rect 7485 3643 7491 3656
rect 7444 3637 7491 3643
rect 884 3617 940 3623
rect 948 3617 988 3623
rect 996 3617 1068 3623
rect 1076 3617 1260 3623
rect 1268 3617 1363 3623
rect 738 3614 798 3616
rect 738 3606 739 3614
rect 748 3606 749 3614
rect 787 3606 788 3614
rect 797 3606 798 3614
rect 738 3604 798 3606
rect 1357 3603 1363 3617
rect 1476 3617 1500 3623
rect 1652 3617 3580 3623
rect 3956 3617 4012 3623
rect 4020 3617 4044 3623
rect 6148 3617 6492 3623
rect 6500 3617 6556 3623
rect 6964 3617 6972 3623
rect 7348 3617 7516 3623
rect 3746 3614 3806 3616
rect 3746 3606 3747 3614
rect 3756 3606 3757 3614
rect 3795 3606 3796 3614
rect 3805 3606 3806 3614
rect 3746 3604 3806 3606
rect 6754 3614 6814 3616
rect 6754 3606 6755 3614
rect 6764 3606 6765 3614
rect 6803 3606 6804 3614
rect 6813 3606 6814 3614
rect 6754 3604 6814 3606
rect 1357 3597 1772 3603
rect 1780 3597 1996 3603
rect 2036 3597 2348 3603
rect 2628 3597 3292 3603
rect 3300 3597 3340 3603
rect 3348 3597 3436 3603
rect 4244 3597 4828 3603
rect 5508 3597 6572 3603
rect 948 3577 1644 3583
rect 1668 3577 1740 3583
rect 1828 3577 2028 3583
rect 2052 3577 2876 3583
rect 2884 3577 2956 3583
rect 2964 3577 3356 3583
rect 3364 3577 3372 3583
rect 4452 3577 4588 3583
rect 6212 3577 6476 3583
rect 6596 3577 6860 3583
rect 7028 3577 7180 3583
rect 7284 3577 7340 3583
rect 7508 3577 7523 3583
rect 7517 3564 7523 3577
rect 804 3557 1340 3563
rect 1588 3557 1660 3563
rect 1684 3557 1900 3563
rect 1917 3557 2092 3563
rect 644 3537 812 3543
rect 820 3537 844 3543
rect 852 3537 1084 3543
rect 1092 3537 1452 3543
rect 1917 3543 1923 3557
rect 2669 3557 2908 3563
rect 2669 3544 2675 3557
rect 2916 3557 3052 3563
rect 4708 3557 4716 3563
rect 5044 3557 5244 3563
rect 6020 3557 6124 3563
rect 6260 3557 6316 3563
rect 6404 3557 7084 3563
rect 7092 3557 7500 3563
rect 1732 3537 1923 3543
rect 1988 3537 2012 3543
rect 2372 3537 2428 3543
rect 2436 3537 2444 3543
rect 2484 3537 2668 3543
rect 2804 3537 2988 3543
rect 3108 3537 3404 3543
rect 4100 3537 4364 3543
rect 4420 3537 4444 3543
rect 4660 3537 4748 3543
rect 4804 3537 4860 3543
rect 5044 3537 5100 3543
rect 5684 3537 5724 3543
rect 5748 3537 5756 3543
rect 5956 3537 6172 3543
rect 6180 3537 6268 3543
rect 6468 3537 6540 3543
rect 6580 3537 6892 3543
rect 6932 3537 6956 3543
rect 7284 3537 7308 3543
rect 340 3517 483 3523
rect 477 3504 483 3517
rect 868 3517 883 3523
rect 372 3497 412 3503
rect 420 3497 460 3503
rect 484 3497 620 3503
rect 660 3497 700 3503
rect 756 3497 860 3503
rect 877 3503 883 3517
rect 900 3517 1388 3523
rect 1732 3517 1948 3523
rect 2020 3517 2092 3523
rect 2164 3517 2380 3523
rect 2692 3517 2748 3523
rect 2868 3517 3084 3523
rect 3092 3517 3196 3523
rect 3204 3517 3212 3523
rect 3332 3517 3436 3523
rect 3636 3517 3692 3523
rect 3940 3517 3948 3523
rect 3956 3517 4012 3523
rect 4148 3517 4300 3523
rect 4372 3517 4380 3523
rect 4468 3517 4908 3523
rect 5044 3517 5068 3523
rect 5140 3517 5228 3523
rect 5492 3517 5756 3523
rect 5828 3517 5996 3523
rect 6084 3517 6156 3523
rect 6420 3517 6572 3523
rect 6852 3517 6860 3523
rect 7268 3517 7308 3523
rect 7332 3517 7436 3523
rect 877 3497 908 3503
rect 932 3497 1052 3503
rect 1124 3497 1308 3503
rect 1364 3497 1436 3503
rect 1460 3497 1628 3503
rect 1636 3497 1676 3503
rect 1700 3497 1756 3503
rect 1764 3497 1836 3503
rect 1860 3497 2124 3503
rect 2180 3497 2220 3503
rect 2452 3497 2540 3503
rect 2740 3497 2860 3503
rect 2980 3497 3100 3503
rect 3108 3497 3500 3503
rect 3620 3497 3868 3503
rect 3876 3497 4060 3503
rect 4276 3497 4444 3503
rect 4612 3497 4620 3503
rect 4628 3497 4716 3503
rect 4820 3497 4828 3503
rect 4948 3497 5404 3503
rect 5460 3497 5516 3503
rect 5620 3497 5788 3503
rect 5796 3497 5948 3503
rect 5988 3497 6444 3503
rect 6484 3497 6524 3503
rect 6900 3497 6956 3503
rect 7076 3497 7107 3503
rect -35 3477 12 3483
rect 132 3477 172 3483
rect 180 3477 316 3483
rect 564 3477 1100 3483
rect 1108 3477 1180 3483
rect 1188 3477 1500 3483
rect 1556 3477 1708 3483
rect 1876 3477 1932 3483
rect 2196 3477 2364 3483
rect 2708 3477 2764 3483
rect 2804 3477 2860 3483
rect 2964 3477 3020 3483
rect 3044 3477 3084 3483
rect 3172 3477 3180 3483
rect 3220 3477 3276 3483
rect 3380 3477 3564 3483
rect 3908 3477 3964 3483
rect 4308 3477 4476 3483
rect 4532 3477 4588 3483
rect 4717 3483 4723 3496
rect 4717 3477 5548 3483
rect 5940 3477 5980 3483
rect 5988 3477 6028 3483
rect 6052 3477 6108 3483
rect 6164 3477 6412 3483
rect 6692 3477 6828 3483
rect 6964 3477 7068 3483
rect 7101 3483 7107 3497
rect 7220 3497 7292 3503
rect 7380 3497 7404 3503
rect 7428 3497 7452 3503
rect 7101 3477 7132 3483
rect 7172 3477 7244 3483
rect 7316 3477 7404 3483
rect 340 3457 380 3463
rect 452 3457 524 3463
rect 820 3457 988 3463
rect 1044 3457 1116 3463
rect 1252 3457 1356 3463
rect 1540 3457 2012 3463
rect 2196 3457 2332 3463
rect 2644 3457 2748 3463
rect 2820 3457 2924 3463
rect 2948 3457 3084 3463
rect 3268 3457 3372 3463
rect 3412 3457 3660 3463
rect 4292 3457 4364 3463
rect 4484 3457 4796 3463
rect 4836 3457 4892 3463
rect 4916 3457 5004 3463
rect 5044 3457 5116 3463
rect 5172 3457 5228 3463
rect 5348 3457 5356 3463
rect 5364 3457 5420 3463
rect 5773 3463 5779 3476
rect 5716 3457 6620 3463
rect 6628 3457 7308 3463
rect 7396 3457 7452 3463
rect 20 3437 1740 3443
rect 1876 3437 1996 3443
rect 2148 3437 2252 3443
rect 2356 3437 2844 3443
rect 2852 3437 2860 3443
rect 2868 3437 3100 3443
rect 3108 3437 3228 3443
rect 3236 3437 3260 3443
rect 4212 3437 4412 3443
rect 4692 3437 4716 3443
rect 5005 3443 5011 3456
rect 5005 3437 5052 3443
rect 5060 3437 5100 3443
rect 5156 3437 5180 3443
rect 6388 3437 6428 3443
rect 6452 3437 6652 3443
rect 6660 3437 7203 3443
rect 660 3417 1900 3423
rect 1924 3417 2060 3423
rect 2141 3423 2147 3436
rect 2068 3417 2147 3423
rect 2388 3417 2748 3423
rect 2756 3417 3180 3423
rect 3380 3417 3484 3423
rect 4052 3417 4460 3423
rect 4660 3417 5180 3423
rect 5428 3417 5820 3423
rect 5828 3417 5964 3423
rect 6308 3417 6412 3423
rect 6420 3417 6524 3423
rect 6564 3417 6700 3423
rect 6884 3417 7164 3423
rect 7197 3423 7203 3437
rect 7220 3437 7436 3443
rect 7508 3437 7532 3443
rect 7197 3417 7372 3423
rect 2242 3414 2302 3416
rect 2242 3406 2243 3414
rect 2252 3406 2253 3414
rect 2291 3406 2292 3414
rect 2301 3406 2302 3414
rect 2242 3404 2302 3406
rect 5250 3414 5310 3416
rect 5250 3406 5251 3414
rect 5260 3406 5261 3414
rect 5299 3406 5300 3414
rect 5309 3406 5310 3414
rect 5250 3404 5310 3406
rect 532 3397 860 3403
rect 1028 3397 1052 3403
rect 1396 3397 1884 3403
rect 1892 3397 2227 3403
rect 692 3377 764 3383
rect 772 3377 940 3383
rect 948 3377 1036 3383
rect 1252 3377 1436 3383
rect 1444 3377 1532 3383
rect 1572 3377 2188 3383
rect 2221 3383 2227 3397
rect 2692 3397 2732 3403
rect 3220 3397 3612 3403
rect 4356 3397 5052 3403
rect 5140 3397 5164 3403
rect 6244 3397 6316 3403
rect 6404 3397 7388 3403
rect 2221 3377 2396 3383
rect 2740 3377 2892 3383
rect 2900 3377 3244 3383
rect 3252 3377 3468 3383
rect 4068 3377 4108 3383
rect 4532 3377 4556 3383
rect 4740 3377 4780 3383
rect 4820 3377 4844 3383
rect 4900 3377 4963 3383
rect 196 3357 332 3363
rect 468 3357 1516 3363
rect 1524 3357 1676 3363
rect 1684 3357 1708 3363
rect 1716 3357 1724 3363
rect 1764 3357 1948 3363
rect 1972 3357 2348 3363
rect 2388 3357 3116 3363
rect 3156 3357 3212 3363
rect 3316 3357 3596 3363
rect 4132 3357 4172 3363
rect 4276 3357 4460 3363
rect 4564 3357 4812 3363
rect 4957 3363 4963 3377
rect 5172 3377 5212 3383
rect 5348 3377 5612 3383
rect 5812 3377 5868 3383
rect 6100 3377 6220 3383
rect 6276 3377 6460 3383
rect 6468 3377 6588 3383
rect 6612 3377 6716 3383
rect 6756 3377 7292 3383
rect 7316 3377 7356 3383
rect 7396 3377 7436 3383
rect 4957 3357 5276 3363
rect 5300 3357 5356 3363
rect 5380 3357 5404 3363
rect 5508 3357 5836 3363
rect 6260 3357 6476 3363
rect 6484 3357 6652 3363
rect 6916 3357 6940 3363
rect 6996 3357 7260 3363
rect 7332 3357 7340 3363
rect 7476 3357 7516 3363
rect 420 3337 524 3343
rect 932 3337 956 3343
rect 964 3337 972 3343
rect 980 3337 1356 3343
rect 1364 3337 1852 3343
rect 1924 3337 2220 3343
rect 2228 3337 2492 3343
rect 2500 3337 2828 3343
rect 3140 3337 3324 3343
rect 3492 3337 3532 3343
rect 3700 3337 3788 3343
rect 3892 3337 3932 3343
rect 4116 3337 4204 3343
rect 4452 3337 4540 3343
rect 4612 3337 4668 3343
rect 4724 3337 4732 3343
rect 4788 3337 4876 3343
rect 4941 3343 4947 3356
rect 4941 3337 4988 3343
rect 5012 3337 5132 3343
rect 5140 3337 5404 3343
rect 5412 3337 5596 3343
rect 5620 3337 5628 3343
rect 5636 3337 5708 3343
rect 5716 3337 5788 3343
rect 5860 3337 5948 3343
rect 5956 3337 6076 3343
rect 6084 3337 6252 3343
rect 6388 3337 6508 3343
rect 6548 3337 6572 3343
rect 6948 3337 7052 3343
rect 7124 3337 7148 3343
rect 7188 3337 7244 3343
rect 7252 3337 7260 3343
rect 7332 3337 7404 3343
rect 7412 3337 7436 3343
rect 132 3317 156 3323
rect 164 3317 236 3323
rect 580 3317 1052 3323
rect 1076 3317 1116 3323
rect 1124 3317 1164 3323
rect 1172 3317 1212 3323
rect 1428 3317 1436 3323
rect 1988 3317 2028 3323
rect 2052 3317 2156 3323
rect 2356 3317 2572 3323
rect 2804 3317 2860 3323
rect 3012 3317 3404 3323
rect 3412 3317 3516 3323
rect 3588 3317 3628 3323
rect 3636 3317 3820 3323
rect 3828 3317 3948 3323
rect 4116 3317 4188 3323
rect 4260 3317 4364 3323
rect 4436 3317 4444 3323
rect 4468 3317 4604 3323
rect 4628 3317 4684 3323
rect 4724 3317 4748 3323
rect 4820 3317 4924 3323
rect 4964 3317 5084 3323
rect 5092 3317 5452 3323
rect 5588 3317 5660 3323
rect 5668 3317 5740 3323
rect 5748 3317 6012 3323
rect 6084 3317 6124 3323
rect 6532 3317 6620 3323
rect 7060 3317 7132 3323
rect 7172 3317 7244 3323
rect 7284 3317 7340 3323
rect 7348 3317 7388 3323
rect 7476 3317 7500 3323
rect 7508 3317 7532 3323
rect 724 3297 876 3303
rect 916 3297 972 3303
rect 1204 3297 1308 3303
rect 1460 3297 1788 3303
rect 1796 3297 1852 3303
rect 1908 3297 2380 3303
rect 2612 3297 2620 3303
rect 2740 3297 2796 3303
rect 3204 3297 3244 3303
rect 3364 3297 3404 3303
rect 3428 3297 3500 3303
rect 3668 3297 3996 3303
rect 4228 3297 4252 3303
rect 4420 3297 4940 3303
rect 5012 3297 5036 3303
rect 5140 3297 5164 3303
rect 5476 3297 5548 3303
rect 5572 3297 5660 3303
rect 5732 3297 6300 3303
rect 6356 3297 6444 3303
rect 6532 3297 6588 3303
rect 6708 3297 7036 3303
rect 7252 3297 7420 3303
rect 708 3277 892 3283
rect 1156 3277 1404 3283
rect 1412 3277 2220 3283
rect 2612 3277 3932 3283
rect 4292 3277 4460 3283
rect 4500 3277 4732 3283
rect 4836 3277 4860 3283
rect 5204 3277 5692 3283
rect 5732 3277 5772 3283
rect 6068 3277 6108 3283
rect 7124 3277 7372 3283
rect 660 3257 1427 3263
rect 692 3237 1148 3243
rect 1421 3243 1427 3257
rect 1492 3257 1628 3263
rect 1748 3257 2044 3263
rect 2644 3257 2700 3263
rect 2708 3257 3020 3263
rect 3028 3257 3228 3263
rect 3236 3257 3340 3263
rect 3652 3257 4812 3263
rect 5076 3257 5788 3263
rect 5844 3257 7084 3263
rect 7316 3257 7340 3263
rect 1421 3237 1564 3243
rect 1732 3237 3884 3243
rect 3908 3237 5484 3243
rect 5940 3237 6764 3243
rect 1204 3217 1468 3223
rect 1476 3217 1612 3223
rect 1892 3217 1996 3223
rect 2068 3217 3068 3223
rect 3284 3217 3660 3223
rect 4660 3217 5580 3223
rect 5604 3217 6332 3223
rect 6564 3217 6636 3223
rect 6932 3217 6940 3223
rect 738 3214 798 3216
rect 738 3206 739 3214
rect 748 3206 749 3214
rect 787 3206 788 3214
rect 797 3206 798 3214
rect 738 3204 798 3206
rect 3746 3214 3806 3216
rect 3746 3206 3747 3214
rect 3756 3206 3757 3214
rect 3795 3206 3796 3214
rect 3805 3206 3806 3214
rect 3746 3204 3806 3206
rect 6754 3214 6814 3216
rect 6754 3206 6755 3214
rect 6764 3206 6765 3214
rect 6803 3206 6804 3214
rect 6813 3206 6814 3214
rect 6754 3204 6814 3206
rect 1284 3197 1324 3203
rect 1812 3197 1820 3203
rect 1828 3197 2028 3203
rect 2036 3197 2316 3203
rect 2372 3197 2636 3203
rect 2660 3197 2668 3203
rect 2772 3197 2940 3203
rect 3044 3197 3340 3203
rect 3380 3197 3580 3203
rect 4084 3197 4268 3203
rect 4580 3197 4620 3203
rect 4756 3197 5516 3203
rect 5764 3197 5868 3203
rect 6420 3197 6739 3203
rect 964 3177 1068 3183
rect 1844 3177 1868 3183
rect 2116 3177 2636 3183
rect 2660 3177 2924 3183
rect 2932 3177 2972 3183
rect 3060 3177 3388 3183
rect 3396 3177 3564 3183
rect 3700 3177 3756 3183
rect 4084 3177 4220 3183
rect 4749 3183 4755 3196
rect 4228 3177 4755 3183
rect 5204 3177 5708 3183
rect 5748 3177 5756 3183
rect 5780 3177 6060 3183
rect 6340 3177 6620 3183
rect 6644 3177 6684 3183
rect 6733 3183 6739 3197
rect 6916 3197 6988 3203
rect 6733 3177 6924 3183
rect 6980 3177 7020 3183
rect 7492 3177 7500 3183
rect 180 3157 1660 3163
rect 2212 3157 2380 3163
rect 2788 3157 3196 3163
rect 3220 3157 3420 3163
rect 3444 3157 4316 3163
rect 4404 3157 4604 3163
rect 4628 3157 5036 3163
rect 5220 3157 6220 3163
rect 6237 3157 6364 3163
rect 612 3137 636 3143
rect 676 3137 700 3143
rect 717 3137 1116 3143
rect 436 3117 572 3123
rect 717 3123 723 3137
rect 1124 3137 1420 3143
rect 1428 3137 1923 3143
rect 628 3117 723 3123
rect 948 3117 1196 3123
rect 1252 3117 1292 3123
rect 1300 3117 1388 3123
rect 1396 3117 1596 3123
rect 1917 3123 1923 3137
rect 2052 3137 2076 3143
rect 2084 3137 2499 3143
rect 1917 3117 2108 3123
rect 2180 3117 2236 3123
rect 2452 3117 2476 3123
rect 2493 3123 2499 3137
rect 2548 3137 2572 3143
rect 2580 3137 2652 3143
rect 2756 3137 2892 3143
rect 2964 3137 3100 3143
rect 3508 3137 3676 3143
rect 4276 3137 4300 3143
rect 4532 3137 4556 3143
rect 4724 3137 4764 3143
rect 5108 3137 5212 3143
rect 5380 3137 5420 3143
rect 5501 3137 5964 3143
rect 5501 3124 5507 3137
rect 6237 3143 6243 3157
rect 6388 3157 7276 3163
rect 5988 3137 6243 3143
rect 6324 3137 6396 3143
rect 6436 3137 6460 3143
rect 6484 3137 6860 3143
rect 6948 3137 6972 3143
rect 2493 3117 2668 3123
rect 2772 3117 2988 3123
rect 3076 3117 3132 3123
rect 3140 3117 3148 3123
rect 3252 3117 3324 3123
rect 3508 3117 3548 3123
rect 3988 3117 4108 3123
rect 4244 3117 4348 3123
rect 4532 3117 4588 3123
rect 4692 3117 4748 3123
rect 4916 3117 5036 3123
rect 5044 3117 5484 3123
rect 5492 3117 5500 3123
rect 5652 3117 5820 3123
rect 5908 3117 6060 3123
rect 6228 3117 6268 3123
rect 6317 3117 6652 3123
rect 6317 3104 6323 3117
rect 6660 3117 7004 3123
rect 7012 3117 7212 3123
rect 7396 3117 7436 3123
rect 52 3097 92 3103
rect 164 3097 172 3103
rect 180 3097 204 3103
rect 260 3097 348 3103
rect 356 3097 556 3103
rect 564 3097 684 3103
rect 724 3097 748 3103
rect 868 3097 1452 3103
rect 1940 3097 1948 3103
rect 2004 3097 2252 3103
rect 2724 3097 2780 3103
rect 2948 3097 3100 3103
rect 3108 3097 3356 3103
rect 3396 3097 3500 3103
rect 3556 3097 3628 3103
rect 3636 3097 3820 3103
rect 3956 3097 4044 3103
rect 4180 3097 4236 3103
rect 4292 3097 4396 3103
rect 4452 3097 4748 3103
rect 5028 3097 5212 3103
rect 5684 3097 5692 3103
rect 5700 3097 5772 3103
rect 6020 3097 6316 3103
rect 6452 3097 6540 3103
rect 6580 3097 6988 3103
rect 6996 3097 7020 3103
rect 7060 3097 7068 3103
rect 7076 3097 7132 3103
rect 7364 3097 7404 3103
rect 564 3077 636 3083
rect 644 3077 1356 3083
rect 1364 3077 2732 3083
rect 2740 3077 2796 3083
rect 2804 3077 3148 3083
rect 3156 3077 3180 3083
rect 3549 3083 3555 3096
rect 3460 3077 3555 3083
rect 4004 3077 4012 3083
rect 4212 3077 4252 3083
rect 4324 3077 4364 3083
rect 5076 3077 5084 3083
rect 5428 3077 5900 3083
rect 6004 3077 6108 3083
rect 6132 3077 6220 3083
rect 6308 3077 6316 3083
rect 6484 3077 6572 3083
rect 6628 3077 6924 3083
rect 6932 3077 6972 3083
rect 7140 3077 7164 3083
rect 7204 3077 7244 3083
rect 7364 3077 7388 3083
rect 7476 3077 7516 3083
rect 852 3057 908 3063
rect 916 3057 988 3063
rect 1012 3057 1068 3063
rect 1076 3057 1132 3063
rect 1140 3057 1308 3063
rect 1652 3057 1676 3063
rect 1972 3057 2172 3063
rect 2196 3057 2508 3063
rect 2516 3057 2796 3063
rect 3268 3057 3308 3063
rect 3316 3057 3612 3063
rect 3620 3057 3740 3063
rect 4052 3057 4316 3063
rect 4404 3057 4444 3063
rect 4468 3057 4492 3063
rect 4532 3057 4972 3063
rect 5140 3057 5164 3063
rect 5188 3057 5260 3063
rect 5620 3057 6076 3063
rect 6084 3057 6364 3063
rect 6372 3057 6716 3063
rect 6724 3057 6892 3063
rect 6900 3057 7180 3063
rect 7236 3057 7420 3063
rect 372 3037 476 3043
rect 548 3037 668 3043
rect 676 3037 796 3043
rect 1396 3037 1756 3043
rect 1764 3037 1875 3043
rect 1316 3017 1404 3023
rect 1869 3023 1875 3037
rect 1892 3037 2060 3043
rect 2148 3037 2540 3043
rect 2548 3037 2652 3043
rect 2660 3037 3052 3043
rect 3252 3037 3468 3043
rect 3636 3037 4380 3043
rect 4420 3037 4492 3043
rect 4644 3037 4739 3043
rect 1869 3017 1932 3023
rect 2068 3017 2156 3023
rect 2644 3017 3315 3023
rect 2242 3014 2302 3016
rect 2242 3006 2243 3014
rect 2252 3006 2253 3014
rect 2291 3006 2292 3014
rect 2301 3006 2302 3014
rect 2242 3004 2302 3006
rect 804 2997 1004 3003
rect 1300 2997 1724 3003
rect 1748 2997 1868 3003
rect 2068 2997 2092 3003
rect 2644 2997 2668 3003
rect 3092 2997 3116 3003
rect 3124 2997 3164 3003
rect 3309 3003 3315 3017
rect 3332 3017 3836 3023
rect 4436 3017 4716 3023
rect 4733 3023 4739 3037
rect 4756 3037 4876 3043
rect 5108 3037 5148 3043
rect 5172 3037 5331 3043
rect 4733 3017 5196 3023
rect 5325 3023 5331 3037
rect 5364 3037 5507 3043
rect 5325 3017 5356 3023
rect 5444 3017 5484 3023
rect 5501 3023 5507 3037
rect 5556 3037 5628 3043
rect 5652 3037 5980 3043
rect 6004 3037 6460 3043
rect 6708 3037 6716 3043
rect 6740 3037 6828 3043
rect 5501 3017 6476 3023
rect 6628 3017 6636 3023
rect 6660 3017 6684 3023
rect 6756 3017 6924 3023
rect 7124 3017 7228 3023
rect 5250 3014 5310 3016
rect 5250 3006 5251 3014
rect 5260 3006 5261 3014
rect 5299 3006 5300 3014
rect 5309 3006 5310 3014
rect 5250 3004 5310 3006
rect 3309 2997 3468 3003
rect 3668 2997 3884 3003
rect 4260 2997 4972 3003
rect 5325 2997 5660 3003
rect 20 2977 428 2983
rect 676 2977 1068 2983
rect 1076 2977 1388 2983
rect 1780 2977 2092 2983
rect 2388 2977 2700 2983
rect 2852 2977 2892 2983
rect 2900 2977 2972 2983
rect 3348 2977 3628 2983
rect 3700 2977 3740 2983
rect 4596 2977 4844 2983
rect 5325 2983 5331 2997
rect 5860 2997 5923 3003
rect 4884 2977 5331 2983
rect 5540 2977 5564 2983
rect 5636 2977 5900 2983
rect 5917 2983 5923 2997
rect 6308 2997 7123 3003
rect 5917 2977 6515 2983
rect 244 2957 252 2963
rect 308 2957 348 2963
rect 596 2957 620 2963
rect 836 2957 860 2963
rect 932 2957 972 2963
rect 1508 2957 1548 2963
rect 1556 2957 1580 2963
rect 1684 2957 1740 2963
rect 1780 2957 1788 2963
rect 1940 2957 2124 2963
rect 2164 2957 2540 2963
rect 2612 2957 2668 2963
rect 2804 2957 2844 2963
rect 2868 2957 2940 2963
rect 3236 2957 3276 2963
rect 3332 2957 3372 2963
rect 3476 2957 3708 2963
rect 4116 2957 4940 2963
rect 5060 2957 5100 2963
rect 5124 2957 5196 2963
rect 5220 2957 5276 2963
rect 5348 2957 5372 2963
rect 5396 2957 5452 2963
rect 5556 2957 5580 2963
rect 5684 2957 5708 2963
rect 5844 2957 5932 2963
rect 5956 2957 6028 2963
rect 6164 2957 6284 2963
rect 6420 2957 6492 2963
rect 6509 2963 6515 2977
rect 6532 2977 6684 2983
rect 6804 2977 6844 2983
rect 6852 2977 6908 2983
rect 6916 2977 7036 2983
rect 7044 2977 7052 2983
rect 7060 2977 7100 2983
rect 7117 2983 7123 2997
rect 7156 2997 7180 3003
rect 7188 2997 7372 3003
rect 7117 2977 7340 2983
rect 7380 2977 7452 2983
rect 6509 2957 6572 2963
rect 6612 2957 6636 2963
rect 6692 2957 6956 2963
rect 6996 2957 7084 2963
rect 7108 2957 7116 2963
rect 7140 2957 7164 2963
rect 100 2937 284 2943
rect 436 2937 524 2943
rect 868 2937 972 2943
rect 1236 2937 1340 2943
rect 1364 2937 1388 2943
rect 1428 2937 1516 2943
rect 1716 2937 1788 2943
rect 1796 2937 1900 2943
rect 1908 2937 1980 2943
rect 2004 2937 2060 2943
rect 2132 2937 2460 2943
rect 2468 2937 2492 2943
rect 2660 2937 2684 2943
rect 2708 2937 2860 2943
rect 3220 2937 3340 2943
rect 3524 2937 3628 2943
rect 3668 2937 3692 2943
rect 4132 2937 4204 2943
rect 4276 2937 4332 2943
rect 4420 2937 4428 2943
rect 4436 2937 4700 2943
rect 4708 2937 4988 2943
rect 4996 2937 5356 2943
rect 5364 2937 5404 2943
rect 5412 2937 5548 2943
rect 5604 2937 5708 2943
rect 5924 2937 5980 2943
rect 6020 2937 6172 2943
rect 6196 2937 6284 2943
rect 6468 2937 6572 2943
rect 6708 2937 6828 2943
rect 6868 2937 6908 2943
rect 7044 2937 7100 2943
rect 7124 2937 7164 2943
rect 7236 2937 7372 2943
rect 228 2917 236 2923
rect 244 2917 268 2923
rect 276 2917 300 2923
rect 356 2917 380 2923
rect 388 2917 476 2923
rect 644 2917 716 2923
rect 916 2917 1036 2923
rect 1124 2917 1260 2923
rect 1540 2917 1676 2923
rect 1780 2917 1948 2923
rect 1972 2917 2348 2923
rect 2436 2917 2476 2923
rect 2580 2917 2732 2923
rect 2932 2917 3068 2923
rect 3268 2917 3548 2923
rect 3604 2917 3676 2923
rect 3812 2917 3916 2923
rect 3988 2917 4060 2923
rect 4196 2917 4252 2923
rect 4260 2917 4620 2923
rect 4756 2917 5084 2923
rect 5108 2917 5372 2923
rect 5396 2917 5420 2923
rect 5469 2917 5500 2923
rect 452 2897 956 2903
rect 980 2897 988 2903
rect 1412 2897 1804 2903
rect 1860 2897 1980 2903
rect 1988 2897 2620 2903
rect 2724 2897 2796 2903
rect 2836 2897 2908 2903
rect 3092 2897 3212 2903
rect 3316 2897 4092 2903
rect 4452 2897 4476 2903
rect 4500 2897 4796 2903
rect 4932 2897 4940 2903
rect 5012 2897 5132 2903
rect 5469 2903 5475 2917
rect 5524 2917 5548 2923
rect 5604 2917 5804 2923
rect 5908 2917 5996 2923
rect 6404 2917 6412 2923
rect 6516 2917 6748 2923
rect 7028 2917 7196 2923
rect 7236 2917 7244 2923
rect 5188 2897 5475 2903
rect 5492 2897 5516 2903
rect 5540 2897 6300 2903
rect 6564 2897 6572 2903
rect 6628 2897 6636 2903
rect 7124 2897 7388 2903
rect 308 2877 1468 2883
rect 1476 2877 2076 2883
rect 2084 2877 2124 2883
rect 2276 2877 2556 2883
rect 2708 2877 2764 2883
rect 3332 2877 3532 2883
rect 3572 2877 3756 2883
rect 4196 2877 4284 2883
rect 4580 2877 4780 2883
rect 4788 2877 4908 2883
rect 4948 2877 6204 2883
rect 6596 2877 6716 2883
rect 6868 2877 6892 2883
rect 6900 2877 7132 2883
rect 7476 2877 7516 2883
rect 116 2857 204 2863
rect 212 2857 300 2863
rect 548 2857 892 2863
rect 900 2857 956 2863
rect 964 2857 1212 2863
rect 1220 2857 1452 2863
rect 1460 2857 1500 2863
rect 1892 2857 1964 2863
rect 2004 2857 2172 2863
rect 2228 2857 2364 2863
rect 2772 2857 3420 2863
rect 3508 2857 3692 2863
rect 3716 2857 4076 2863
rect 4164 2857 4572 2863
rect 4644 2857 4700 2863
rect 4756 2857 5027 2863
rect 468 2837 876 2843
rect 900 2837 1244 2843
rect 1316 2837 1468 2843
rect 1572 2837 1724 2843
rect 1844 2837 2028 2843
rect 2068 2837 2172 2843
rect 2596 2837 3004 2843
rect 3204 2837 3372 2843
rect 3380 2837 3468 2843
rect 3508 2837 3596 2843
rect 3725 2837 3836 2843
rect 852 2817 1340 2823
rect 1364 2817 1420 2823
rect 1668 2817 1964 2823
rect 3725 2823 3731 2837
rect 4228 2837 4828 2843
rect 4868 2837 5004 2843
rect 5021 2843 5027 2857
rect 5044 2857 6844 2863
rect 6852 2857 7484 2863
rect 7492 2857 7532 2863
rect 5021 2837 5059 2843
rect 3236 2817 3731 2823
rect 4292 2817 5036 2823
rect 5053 2823 5059 2837
rect 5076 2837 5756 2843
rect 5764 2837 6476 2843
rect 6580 2837 6604 2843
rect 6612 2837 6972 2843
rect 7092 2837 7340 2843
rect 7508 2837 7532 2843
rect 5053 2817 5148 2823
rect 5204 2817 5420 2823
rect 5444 2817 5836 2823
rect 5860 2817 5932 2823
rect 6324 2817 6540 2823
rect 6676 2817 6684 2823
rect 738 2814 798 2816
rect 738 2806 739 2814
rect 748 2806 749 2814
rect 787 2806 788 2814
rect 797 2806 798 2814
rect 738 2804 798 2806
rect 3746 2814 3806 2816
rect 3746 2806 3747 2814
rect 3756 2806 3757 2814
rect 3795 2806 3796 2814
rect 3805 2806 3806 2814
rect 3746 2804 3806 2806
rect 6754 2814 6814 2816
rect 6754 2806 6755 2814
rect 6764 2806 6765 2814
rect 6803 2806 6804 2814
rect 6813 2806 6814 2814
rect 6754 2804 6814 2806
rect 852 2797 972 2803
rect 1060 2797 1292 2803
rect 1300 2797 1692 2803
rect 1700 2797 1884 2803
rect 1892 2797 2204 2803
rect 2932 2797 2940 2803
rect 3556 2797 3731 2803
rect 564 2777 1116 2783
rect 1364 2777 1484 2783
rect 1540 2777 1747 2783
rect 420 2757 851 2763
rect 468 2737 572 2743
rect 845 2743 851 2757
rect 868 2757 1052 2763
rect 1348 2757 1628 2763
rect 1741 2763 1747 2777
rect 1764 2777 1868 2783
rect 2532 2777 2572 2783
rect 2644 2777 2828 2783
rect 2852 2777 3132 2783
rect 3140 2777 3244 2783
rect 3412 2777 3708 2783
rect 3725 2783 3731 2797
rect 3892 2797 5100 2803
rect 5124 2797 6636 2803
rect 7156 2797 7356 2803
rect 3725 2777 3996 2783
rect 4356 2777 4652 2783
rect 4788 2777 4796 2783
rect 4836 2777 4956 2783
rect 4980 2777 5244 2783
rect 5252 2777 5404 2783
rect 5588 2777 5980 2783
rect 6436 2777 6508 2783
rect 6612 2777 6700 2783
rect 7284 2777 7372 2783
rect 1741 2757 2156 2763
rect 2900 2757 3036 2763
rect 3044 2757 3228 2763
rect 3636 2757 3900 2763
rect 3988 2757 4332 2763
rect 4436 2757 4492 2763
rect 4628 2757 5116 2763
rect 5188 2757 5356 2763
rect 5380 2757 5436 2763
rect 5492 2757 5532 2763
rect 5540 2757 5580 2763
rect 5812 2757 5868 2763
rect 6212 2757 6876 2763
rect 6884 2757 7068 2763
rect 7140 2757 7244 2763
rect 7252 2757 7292 2763
rect 7300 2757 7452 2763
rect 845 2737 1340 2743
rect 1444 2737 1452 2743
rect 1716 2737 1788 2743
rect 1924 2737 2012 2743
rect 2068 2737 2300 2743
rect 3028 2737 3116 2743
rect 3124 2737 3148 2743
rect 3156 2737 3340 2743
rect 3364 2737 3436 2743
rect 3661 2737 4124 2743
rect 3661 2724 3667 2737
rect 4324 2737 5100 2743
rect 5108 2737 5596 2743
rect 5604 2737 6060 2743
rect 6180 2737 6252 2743
rect 6260 2737 6588 2743
rect 6644 2737 6739 2743
rect 372 2717 396 2723
rect 516 2717 844 2723
rect 868 2717 876 2723
rect 1028 2717 1068 2723
rect 1284 2717 1292 2723
rect 1524 2717 1564 2723
rect 1572 2717 1948 2723
rect 1956 2717 2076 2723
rect 2084 2717 2716 2723
rect 3380 2717 3420 2723
rect 3444 2717 3452 2723
rect 3492 2717 3564 2723
rect 3572 2717 3660 2723
rect 3764 2717 3900 2723
rect 4020 2717 4060 2723
rect 4068 2717 4140 2723
rect 4148 2717 4316 2723
rect 4340 2717 4588 2723
rect 4644 2717 4700 2723
rect 4772 2717 4956 2723
rect 5028 2717 5068 2723
rect 5236 2717 5388 2723
rect 5428 2717 5436 2723
rect 5444 2717 5644 2723
rect 5764 2717 6044 2723
rect 6356 2717 6428 2723
rect 6580 2717 6604 2723
rect 6733 2723 6739 2737
rect 7108 2737 7180 2743
rect 7188 2737 7212 2743
rect 7220 2737 7324 2743
rect 7332 2737 7388 2743
rect 6733 2717 7148 2723
rect 7156 2717 7372 2723
rect 7476 2717 7571 2723
rect 324 2697 364 2703
rect 436 2697 524 2703
rect 548 2697 588 2703
rect 628 2697 652 2703
rect 1044 2697 1084 2703
rect 1156 2697 1196 2703
rect 1220 2697 1404 2703
rect 1604 2697 1660 2703
rect 1844 2697 2140 2703
rect 2228 2697 2540 2703
rect 2676 2697 2684 2703
rect 2788 2697 2844 2703
rect 2964 2697 3436 2703
rect 3476 2697 3516 2703
rect 3524 2697 3612 2703
rect 3700 2697 4012 2703
rect 4100 2697 4348 2703
rect 4404 2697 4460 2703
rect 4548 2697 4668 2703
rect 4676 2697 4748 2703
rect 4772 2697 4844 2703
rect 4868 2697 4908 2703
rect 4948 2697 5036 2703
rect 5108 2697 5132 2703
rect 5204 2697 5724 2703
rect 5732 2697 5756 2703
rect 5796 2697 5852 2703
rect 6004 2697 6124 2703
rect 6244 2697 6332 2703
rect 6452 2697 6700 2703
rect 6788 2697 6892 2703
rect 7044 2697 7116 2703
rect 7284 2697 7292 2703
rect 7316 2697 7420 2703
rect 7540 2697 7555 2703
rect 132 2677 620 2683
rect 900 2677 940 2683
rect 1012 2677 1132 2683
rect 1140 2677 1180 2683
rect 1188 2677 1244 2683
rect 1252 2677 1372 2683
rect 1380 2677 1436 2683
rect 1444 2677 1644 2683
rect 1652 2677 1708 2683
rect 1748 2677 1820 2683
rect 1860 2677 1900 2683
rect 1940 2677 2108 2683
rect 2132 2677 2412 2683
rect 2516 2677 2803 2683
rect 20 2657 204 2663
rect 212 2657 428 2663
rect 484 2657 572 2663
rect 916 2657 1043 2663
rect 452 2637 524 2643
rect 612 2637 620 2643
rect 724 2637 780 2643
rect 948 2637 1020 2643
rect 1037 2643 1043 2657
rect 1172 2657 1196 2663
rect 1364 2657 1388 2663
rect 1396 2657 1676 2663
rect 1684 2657 2044 2663
rect 2052 2657 2428 2663
rect 2436 2657 2748 2663
rect 2797 2663 2803 2677
rect 2820 2677 3052 2683
rect 3124 2677 3260 2683
rect 3284 2677 3372 2683
rect 3412 2677 4236 2683
rect 4349 2683 4355 2696
rect 4349 2677 4396 2683
rect 4461 2683 4467 2696
rect 4461 2677 5212 2683
rect 5220 2677 6156 2683
rect 6164 2677 6428 2683
rect 6436 2677 6732 2683
rect 7037 2683 7043 2696
rect 6884 2677 7043 2683
rect 7181 2683 7187 2696
rect 7156 2677 7187 2683
rect 7252 2677 7324 2683
rect 7412 2677 7436 2683
rect 7444 2677 7468 2683
rect 7492 2677 7532 2683
rect 2797 2657 2876 2663
rect 2932 2657 2988 2663
rect 3060 2657 3868 2663
rect 3908 2657 4060 2663
rect 4372 2657 5052 2663
rect 5060 2657 5084 2663
rect 5092 2657 5452 2663
rect 5460 2657 5500 2663
rect 5796 2657 5948 2663
rect 5956 2657 6076 2663
rect 6084 2657 6172 2663
rect 6388 2657 6492 2663
rect 6596 2657 6812 2663
rect 6820 2657 6860 2663
rect 6900 2657 6940 2663
rect 6996 2657 7340 2663
rect 7396 2657 7516 2663
rect 1037 2637 1484 2643
rect 1492 2637 1516 2643
rect 1524 2637 1676 2643
rect 1684 2637 1900 2643
rect 2052 2637 2060 2643
rect 2692 2637 2812 2643
rect 2980 2637 3068 2643
rect 3476 2637 4044 2643
rect 4388 2637 4636 2643
rect 4644 2637 5564 2643
rect 5588 2637 5644 2643
rect 5684 2637 5724 2643
rect 5828 2637 5980 2643
rect 5988 2637 6220 2643
rect 6228 2637 6284 2643
rect 6589 2643 6595 2656
rect 6292 2637 6595 2643
rect 6644 2637 6652 2643
rect 6852 2637 7020 2643
rect 7044 2637 7084 2643
rect 7092 2637 7164 2643
rect 7172 2637 7308 2643
rect 7364 2637 7468 2643
rect 7549 2643 7555 2697
rect 7540 2637 7555 2643
rect 372 2617 588 2623
rect 596 2617 636 2623
rect 644 2617 972 2623
rect 980 2617 1020 2623
rect 1172 2617 1260 2623
rect 1364 2617 1420 2623
rect 1444 2617 1532 2623
rect 1556 2617 1660 2623
rect 1668 2617 1859 2623
rect 20 2597 364 2603
rect 788 2597 956 2603
rect 1124 2597 1356 2603
rect 1428 2597 1500 2603
rect 1780 2597 1836 2603
rect 1853 2603 1859 2617
rect 2020 2617 2076 2623
rect 2660 2617 2668 2623
rect 3364 2617 3372 2623
rect 3444 2617 4131 2623
rect 2242 2614 2302 2616
rect 2242 2606 2243 2614
rect 2252 2606 2253 2614
rect 2291 2606 2292 2614
rect 2301 2606 2302 2614
rect 2242 2604 2302 2606
rect 1853 2597 2060 2603
rect 2580 2597 2924 2603
rect 3117 2597 3212 2603
rect 3117 2584 3123 2597
rect 3268 2597 3388 2603
rect 3604 2597 3692 2603
rect 4036 2597 4108 2603
rect 4125 2603 4131 2617
rect 4324 2617 4428 2623
rect 4580 2617 4716 2623
rect 4756 2617 5180 2623
rect 5364 2617 5548 2623
rect 5588 2617 5884 2623
rect 5908 2617 6012 2623
rect 6052 2617 6204 2623
rect 6420 2617 6460 2623
rect 6548 2617 6940 2623
rect 7357 2623 7363 2636
rect 7108 2617 7363 2623
rect 7565 2623 7571 2717
rect 7476 2617 7571 2623
rect 5250 2614 5310 2616
rect 5250 2606 5251 2614
rect 5260 2606 5261 2614
rect 5299 2606 5300 2614
rect 5309 2606 5310 2614
rect 5250 2604 5310 2606
rect 4125 2597 4732 2603
rect 4756 2597 4892 2603
rect 4916 2597 5228 2603
rect 5364 2597 5388 2603
rect 5412 2597 5436 2603
rect 5572 2597 6524 2603
rect 6532 2597 7212 2603
rect 7220 2597 7260 2603
rect 7348 2597 7404 2603
rect 148 2577 220 2583
rect 244 2577 300 2583
rect 404 2577 556 2583
rect 1060 2577 1068 2583
rect 1268 2577 1356 2583
rect 1364 2577 1452 2583
rect 1668 2577 1852 2583
rect 1860 2577 1916 2583
rect 2180 2577 3004 2583
rect 3428 2577 3452 2583
rect 3629 2577 3884 2583
rect 308 2557 332 2563
rect 372 2557 476 2563
rect 557 2563 563 2576
rect 557 2557 1372 2563
rect 1380 2557 1404 2563
rect 1428 2557 1580 2563
rect 1684 2557 1932 2563
rect 1972 2557 2204 2563
rect 2340 2557 2652 2563
rect 2804 2557 2972 2563
rect 2980 2557 2988 2563
rect 3053 2557 3356 2563
rect 3053 2544 3059 2557
rect 3629 2563 3635 2577
rect 3956 2577 3996 2583
rect 4100 2577 4172 2583
rect 4196 2577 4684 2583
rect 4708 2577 4780 2583
rect 4884 2577 4940 2583
rect 5044 2577 5187 2583
rect 3460 2557 3635 2563
rect 3732 2557 3820 2563
rect 4068 2557 4220 2563
rect 4372 2557 5068 2563
rect 5124 2557 5164 2563
rect 5181 2563 5187 2577
rect 5236 2577 5612 2583
rect 5636 2577 5740 2583
rect 5764 2577 6108 2583
rect 6164 2577 6460 2583
rect 6580 2577 6684 2583
rect 6964 2577 7196 2583
rect 7252 2577 7308 2583
rect 7316 2577 7372 2583
rect 5181 2557 5372 2563
rect 5380 2557 5468 2563
rect 5533 2557 5660 2563
rect 180 2537 492 2543
rect 500 2537 764 2543
rect 820 2537 988 2543
rect 1348 2537 1484 2543
rect 1508 2537 1516 2543
rect 1652 2537 1724 2543
rect 1828 2537 1852 2543
rect 2148 2537 2684 2543
rect 2692 2537 2700 2543
rect 2772 2537 2860 2543
rect 3012 2537 3052 2543
rect 3284 2537 3500 2543
rect 3508 2537 3580 2543
rect 3604 2537 3660 2543
rect 3668 2537 3740 2543
rect 4020 2537 5132 2543
rect 5533 2543 5539 2557
rect 5844 2557 6076 2563
rect 6084 2557 6156 2563
rect 6260 2557 6876 2563
rect 7188 2557 7260 2563
rect 7268 2557 7340 2563
rect 7364 2557 7564 2563
rect 5348 2537 5539 2543
rect 5556 2537 5676 2543
rect 5956 2537 6028 2543
rect 6036 2537 6124 2543
rect 6132 2537 6380 2543
rect 6420 2537 6476 2543
rect 6484 2537 6572 2543
rect 6628 2537 6668 2543
rect 6788 2537 6988 2543
rect 7060 2537 7196 2543
rect 7204 2537 7244 2543
rect 7268 2537 7292 2543
rect 7444 2537 7452 2543
rect 148 2517 236 2523
rect 292 2517 332 2523
rect 356 2517 428 2523
rect 1108 2517 1132 2523
rect 1460 2517 1532 2523
rect 1572 2517 1852 2523
rect 1860 2517 2124 2523
rect 2132 2517 2588 2523
rect 2724 2517 2764 2523
rect 2772 2517 3180 2523
rect 3188 2517 3228 2523
rect 3508 2517 3596 2523
rect 3684 2517 3948 2523
rect 4004 2517 4108 2523
rect 4132 2517 4252 2523
rect 4692 2517 4828 2523
rect 4836 2517 4860 2523
rect 5092 2517 5132 2523
rect 5204 2517 5292 2523
rect 5396 2517 5436 2523
rect 5556 2517 5676 2523
rect 5684 2517 5932 2523
rect 6164 2517 6236 2523
rect 6276 2517 6332 2523
rect 6468 2517 6492 2523
rect 6708 2517 6748 2523
rect 6788 2517 6908 2523
rect 6932 2517 6956 2523
rect 6980 2517 7388 2523
rect 7460 2517 7532 2523
rect 468 2497 1068 2503
rect 1124 2497 1228 2503
rect 1876 2497 1948 2503
rect 1956 2497 2012 2503
rect 2020 2497 2092 2503
rect 2100 2497 2140 2503
rect 2148 2497 2300 2503
rect 2324 2497 2380 2503
rect 2500 2497 2508 2503
rect 2708 2497 2956 2503
rect 3012 2497 3068 2503
rect 3348 2497 3468 2503
rect 3604 2497 3676 2503
rect 4308 2497 4508 2503
rect 4884 2497 4908 2503
rect 5124 2497 5212 2503
rect 5396 2497 5484 2503
rect 5492 2497 5516 2503
rect 6036 2497 6284 2503
rect 6724 2497 7004 2503
rect 7012 2497 7052 2503
rect 1108 2477 1132 2483
rect 1508 2477 1564 2483
rect 1796 2477 1868 2483
rect 1924 2477 3484 2483
rect 3588 2477 3708 2483
rect 4372 2477 4940 2483
rect 5245 2477 5612 2483
rect 324 2457 2156 2463
rect 2164 2457 2492 2463
rect 2500 2457 2700 2463
rect 3236 2457 3372 2463
rect 3444 2457 3788 2463
rect 4436 2457 4524 2463
rect 5245 2463 5251 2477
rect 6548 2477 6556 2483
rect 6612 2477 6828 2483
rect 6909 2477 7180 2483
rect 6909 2464 6915 2477
rect 7476 2477 7532 2483
rect 4692 2457 5251 2463
rect 5364 2457 5436 2463
rect 5588 2457 6060 2463
rect 6356 2457 6908 2463
rect 6932 2457 7116 2463
rect 7156 2457 7180 2463
rect 244 2437 332 2443
rect 340 2437 412 2443
rect 948 2437 1772 2443
rect 1933 2437 2620 2443
rect 516 2417 588 2423
rect 1933 2423 1939 2437
rect 3396 2437 3692 2443
rect 4212 2437 4604 2443
rect 4628 2437 5036 2443
rect 5428 2437 6124 2443
rect 6132 2437 6444 2443
rect 6452 2437 6668 2443
rect 6685 2437 7052 2443
rect 1492 2417 1939 2423
rect 1956 2417 1964 2423
rect 2004 2417 2524 2423
rect 3316 2417 3596 2423
rect 4164 2417 4396 2423
rect 4509 2417 4716 2423
rect 738 2414 798 2416
rect 738 2406 739 2414
rect 748 2406 749 2414
rect 787 2406 788 2414
rect 797 2406 798 2414
rect 738 2404 798 2406
rect 3746 2414 3806 2416
rect 3746 2406 3747 2414
rect 3756 2406 3757 2414
rect 3795 2406 3796 2414
rect 3805 2406 3806 2414
rect 3746 2404 3806 2406
rect 372 2397 396 2403
rect 1428 2397 1548 2403
rect 1636 2397 1795 2403
rect 260 2377 1100 2383
rect 1476 2377 1564 2383
rect 1716 2377 1772 2383
rect 1789 2383 1795 2397
rect 1812 2397 1964 2403
rect 2196 2397 3228 2403
rect 3588 2397 3628 2403
rect 3828 2397 4108 2403
rect 4509 2403 4515 2417
rect 4724 2417 4812 2423
rect 4820 2417 4844 2423
rect 4852 2417 4924 2423
rect 5204 2417 5420 2423
rect 5460 2417 5772 2423
rect 6685 2423 6691 2437
rect 6516 2417 6691 2423
rect 6836 2417 7116 2423
rect 6754 2414 6814 2416
rect 6754 2406 6755 2414
rect 6764 2406 6765 2414
rect 6803 2406 6804 2414
rect 6813 2406 6814 2414
rect 6754 2404 6814 2406
rect 4116 2397 4515 2403
rect 4532 2397 4588 2403
rect 4964 2397 5116 2403
rect 5172 2397 5388 2403
rect 5460 2397 6540 2403
rect 7540 2397 7548 2403
rect 1789 2377 1996 2383
rect 2404 2377 2460 2383
rect 2468 2377 2508 2383
rect 2516 2377 2732 2383
rect 3124 2377 3180 2383
rect 3220 2377 3260 2383
rect 3284 2377 3468 2383
rect 3524 2377 4092 2383
rect 4292 2377 4588 2383
rect 4596 2377 4764 2383
rect 4996 2377 5171 2383
rect 276 2357 572 2363
rect 580 2357 604 2363
rect 612 2357 812 2363
rect 820 2357 1308 2363
rect 1316 2357 2604 2363
rect 2644 2357 3404 2363
rect 3636 2357 3676 2363
rect 3684 2357 3724 2363
rect 3732 2357 3884 2363
rect 3892 2357 4060 2363
rect 4596 2357 4652 2363
rect 5012 2357 5148 2363
rect 5165 2363 5171 2377
rect 5284 2377 5404 2383
rect 5428 2377 5612 2383
rect 6628 2377 6940 2383
rect 7172 2377 7340 2383
rect 5165 2357 5516 2363
rect 5540 2357 5644 2363
rect 6180 2357 6252 2363
rect 6580 2357 7436 2363
rect 996 2337 1196 2343
rect 1300 2337 1372 2343
rect 1380 2337 1555 2343
rect 500 2317 620 2323
rect 836 2317 876 2323
rect 1076 2317 1171 2323
rect 52 2297 156 2303
rect 180 2297 204 2303
rect 228 2297 252 2303
rect 276 2297 828 2303
rect 868 2297 924 2303
rect 1165 2303 1171 2317
rect 1188 2317 1324 2323
rect 1396 2317 1484 2323
rect 1549 2323 1555 2337
rect 1572 2337 2124 2343
rect 2196 2337 2860 2343
rect 2932 2337 3324 2343
rect 3533 2337 3948 2343
rect 1549 2317 1628 2323
rect 1636 2317 1660 2323
rect 1748 2317 1964 2323
rect 2020 2317 2172 2323
rect 2388 2317 2428 2323
rect 2436 2317 2476 2323
rect 2484 2317 2796 2323
rect 2804 2317 3004 2323
rect 3428 2317 3436 2323
rect 3533 2323 3539 2337
rect 4100 2337 4332 2343
rect 4340 2337 4444 2343
rect 4452 2337 4492 2343
rect 4788 2337 5004 2343
rect 5204 2337 5356 2343
rect 5412 2337 5539 2343
rect 5533 2324 5539 2337
rect 5988 2337 6156 2343
rect 6164 2337 6364 2343
rect 6804 2337 6860 2343
rect 7092 2337 7132 2343
rect 7284 2337 7516 2343
rect 3460 2317 3539 2323
rect 3556 2317 3628 2323
rect 3844 2317 4140 2323
rect 4276 2317 4284 2323
rect 4532 2317 4572 2323
rect 4804 2317 4876 2323
rect 4948 2317 5132 2323
rect 5140 2317 5196 2323
rect 5236 2317 5340 2323
rect 5428 2317 5500 2323
rect 5684 2317 5708 2323
rect 5908 2317 5932 2323
rect 6068 2317 6252 2323
rect 6356 2317 6460 2323
rect 6644 2317 6732 2323
rect 6836 2317 6972 2323
rect 6980 2317 7116 2323
rect 7140 2317 7196 2323
rect 7284 2317 7468 2323
rect 1165 2297 1324 2303
rect 1332 2297 1756 2303
rect 1780 2297 1852 2303
rect 2164 2297 2252 2303
rect 2260 2297 2844 2303
rect 3300 2297 3372 2303
rect 3380 2297 3420 2303
rect 3508 2297 3548 2303
rect 4084 2297 4124 2303
rect 4132 2297 5820 2303
rect 5828 2297 6188 2303
rect 6196 2297 6476 2303
rect 6484 2297 6540 2303
rect 6676 2297 6844 2303
rect 7092 2297 7116 2303
rect 7140 2297 7180 2303
rect 7508 2297 7516 2303
rect 7549 2297 7603 2303
rect 196 2277 236 2283
rect 244 2277 332 2283
rect 868 2277 1340 2283
rect 1412 2277 1692 2283
rect 1716 2277 1804 2283
rect 1828 2277 1884 2283
rect 1908 2277 2380 2283
rect 2468 2277 2620 2283
rect 2676 2277 2700 2283
rect 2708 2277 2908 2283
rect 3252 2277 3276 2283
rect 3300 2277 3308 2283
rect 3364 2277 3468 2283
rect 3476 2277 3628 2283
rect 3636 2277 3788 2283
rect 3892 2277 3980 2283
rect 4164 2277 4348 2283
rect 4356 2277 4476 2283
rect 4484 2277 4604 2283
rect 4756 2277 4796 2283
rect 4980 2277 5020 2283
rect 5092 2277 5244 2283
rect 5380 2277 5388 2283
rect 5444 2277 5875 2283
rect 436 2257 540 2263
rect 548 2257 572 2263
rect 1300 2257 1372 2263
rect 1428 2257 1740 2263
rect 1972 2257 2076 2263
rect 2084 2257 2268 2263
rect 2276 2257 2444 2263
rect 2516 2257 2620 2263
rect 3284 2257 3324 2263
rect 3556 2257 3692 2263
rect 3716 2257 4156 2263
rect 4244 2257 4348 2263
rect 4532 2257 4652 2263
rect 4900 2257 4988 2263
rect 4996 2257 5436 2263
rect 5668 2257 5708 2263
rect 5716 2257 5772 2263
rect 5780 2257 5852 2263
rect 5869 2263 5875 2277
rect 5924 2277 6284 2283
rect 6292 2277 6428 2283
rect 6436 2277 6476 2283
rect 6484 2277 6508 2283
rect 6516 2277 6780 2283
rect 6948 2277 7180 2283
rect 7188 2277 7324 2283
rect 7332 2277 7420 2283
rect 7549 2283 7555 2297
rect 7492 2277 7555 2283
rect 5869 2257 5948 2263
rect 6004 2257 6108 2263
rect 6116 2257 6332 2263
rect 6452 2257 6636 2263
rect 6900 2257 6924 2263
rect 7204 2257 7244 2263
rect 7268 2257 7292 2263
rect 7476 2257 7484 2263
rect 7492 2257 7548 2263
rect 1492 2237 1724 2243
rect 1748 2237 1932 2243
rect 2100 2237 2204 2243
rect 2212 2237 2492 2243
rect 2548 2237 3532 2243
rect 3588 2237 3644 2243
rect 3876 2237 3884 2243
rect 4356 2237 4540 2243
rect 4580 2237 4620 2243
rect 4637 2237 4972 2243
rect 692 2217 732 2223
rect 740 2217 1484 2223
rect 1572 2217 1708 2223
rect 1844 2217 2220 2223
rect 2580 2217 2652 2223
rect 2836 2217 3660 2223
rect 4637 2223 4643 2237
rect 5012 2237 5052 2243
rect 5060 2237 5404 2243
rect 5604 2237 5676 2243
rect 5732 2237 5820 2243
rect 5828 2237 5996 2243
rect 6004 2237 6028 2243
rect 6244 2237 6412 2243
rect 6692 2237 7011 2243
rect 3732 2217 4643 2223
rect 5005 2223 5011 2236
rect 7005 2224 7011 2237
rect 7220 2237 7356 2243
rect 7460 2237 7548 2243
rect 4772 2217 5011 2223
rect 5348 2217 5452 2223
rect 5556 2217 5868 2223
rect 6164 2217 6188 2223
rect 6228 2217 6236 2223
rect 6260 2217 6380 2223
rect 6388 2217 6572 2223
rect 6644 2217 6700 2223
rect 6708 2217 6892 2223
rect 7012 2217 7084 2223
rect 7220 2217 7324 2223
rect 2242 2214 2302 2216
rect 2242 2206 2243 2214
rect 2252 2206 2253 2214
rect 2291 2206 2292 2214
rect 2301 2206 2302 2214
rect 2242 2204 2302 2206
rect 5250 2214 5310 2216
rect 5250 2206 5251 2214
rect 5260 2206 5261 2214
rect 5299 2206 5300 2214
rect 5309 2206 5310 2214
rect 5250 2204 5310 2206
rect 564 2197 1100 2203
rect 1108 2197 1404 2203
rect 1540 2197 1612 2203
rect 1636 2197 1836 2203
rect 1844 2197 1900 2203
rect 1988 2197 2188 2203
rect 2388 2197 2716 2203
rect 2852 2197 2892 2203
rect 3220 2197 4060 2203
rect 4420 2197 4956 2203
rect 4980 2197 5196 2203
rect 5325 2197 5756 2203
rect 1108 2177 1388 2183
rect 1476 2177 1484 2183
rect 1604 2177 1724 2183
rect 1748 2177 3532 2183
rect 3572 2177 3932 2183
rect 4052 2177 4188 2183
rect 5325 2183 5331 2197
rect 6100 2197 6396 2203
rect 6708 2197 7036 2203
rect 7044 2197 7100 2203
rect 4196 2177 5331 2183
rect 5396 2177 5427 2183
rect 20 2157 44 2163
rect 164 2157 204 2163
rect 324 2157 444 2163
rect 452 2157 476 2163
rect 1204 2157 1404 2163
rect 1444 2157 1708 2163
rect 2388 2157 2556 2163
rect 2596 2157 2748 2163
rect 2916 2157 2988 2163
rect 3044 2157 3084 2163
rect 3156 2157 3340 2163
rect 3412 2157 3612 2163
rect 3668 2157 3708 2163
rect 4276 2157 4492 2163
rect 4516 2157 4739 2163
rect 52 2137 92 2143
rect 100 2137 172 2143
rect 253 2137 284 2143
rect 253 2124 259 2137
rect 388 2137 668 2143
rect 676 2137 812 2143
rect 1076 2137 1132 2143
rect 1140 2137 1180 2143
rect 1236 2137 1532 2143
rect 1700 2137 1900 2143
rect 2116 2137 2332 2143
rect 2388 2137 2636 2143
rect 2644 2137 2668 2143
rect 2708 2137 2764 2143
rect 2964 2137 2988 2143
rect 2996 2137 3068 2143
rect 3076 2137 3116 2143
rect 3268 2137 3468 2143
rect 3540 2137 3660 2143
rect 3924 2137 4012 2143
rect 4116 2137 4300 2143
rect 4580 2137 4604 2143
rect 4733 2143 4739 2157
rect 4756 2157 4844 2163
rect 4868 2157 4892 2163
rect 5028 2157 5148 2163
rect 5300 2157 5404 2163
rect 5421 2163 5427 2177
rect 5492 2177 5596 2183
rect 5620 2177 5660 2183
rect 5764 2177 6012 2183
rect 6020 2177 6588 2183
rect 6596 2177 6636 2183
rect 6724 2177 6876 2183
rect 6900 2177 6972 2183
rect 6996 2177 7148 2183
rect 7348 2177 7388 2183
rect 5421 2157 5628 2163
rect 5901 2157 6012 2163
rect 5901 2144 5907 2157
rect 6196 2157 6236 2163
rect 6324 2157 6428 2163
rect 6468 2157 6524 2163
rect 6532 2157 6652 2163
rect 6660 2157 6700 2163
rect 6964 2157 6988 2163
rect 7076 2157 7244 2163
rect 7252 2157 7532 2163
rect 4733 2137 5276 2143
rect 5396 2137 5452 2143
rect 5860 2137 5900 2143
rect 6084 2137 6476 2143
rect 6580 2137 6636 2143
rect 6772 2137 6860 2143
rect 6996 2137 7308 2143
rect 7316 2137 7436 2143
rect 84 2117 124 2123
rect 196 2117 252 2123
rect 276 2117 332 2123
rect 340 2117 524 2123
rect 548 2117 652 2123
rect 660 2117 684 2123
rect 932 2117 988 2123
rect 1172 2117 1260 2123
rect 1364 2117 1740 2123
rect 1764 2117 1980 2123
rect 2020 2117 2124 2123
rect 2548 2117 2588 2123
rect 2701 2123 2707 2136
rect 2605 2117 2707 2123
rect 84 2097 348 2103
rect 356 2097 396 2103
rect 564 2097 972 2103
rect 1396 2097 1500 2103
rect 1700 2097 1724 2103
rect 1748 2097 1804 2103
rect 2605 2103 2611 2117
rect 2788 2117 2796 2123
rect 3060 2117 3276 2123
rect 3316 2117 3436 2123
rect 3636 2117 3644 2123
rect 3764 2117 4140 2123
rect 4580 2117 4652 2123
rect 4708 2117 4780 2123
rect 4788 2117 4860 2123
rect 4868 2117 4908 2123
rect 4916 2117 4988 2123
rect 4996 2117 5132 2123
rect 5188 2117 5212 2123
rect 5348 2117 5500 2123
rect 5620 2117 5660 2123
rect 5716 2117 5788 2123
rect 5844 2117 5900 2123
rect 5972 2117 6044 2123
rect 6276 2117 6284 2123
rect 6484 2117 7020 2123
rect 7124 2117 7132 2123
rect 7156 2117 7180 2123
rect 7380 2117 7436 2123
rect 1892 2097 2611 2103
rect 2708 2097 3036 2103
rect 3108 2097 3212 2103
rect 3572 2097 3596 2103
rect 3780 2097 4332 2103
rect 4468 2097 4508 2103
rect 4612 2097 4812 2103
rect 5060 2097 5116 2103
rect 5140 2097 5148 2103
rect 5156 2097 5196 2103
rect 5284 2097 6076 2103
rect 6388 2097 6428 2103
rect 6484 2097 6524 2103
rect 6628 2097 6668 2103
rect 6692 2097 6748 2103
rect 6884 2097 6940 2103
rect 7012 2097 7052 2103
rect 7124 2097 7228 2103
rect 7396 2097 7468 2103
rect 116 2077 476 2083
rect 484 2077 540 2083
rect 580 2077 588 2083
rect 612 2077 652 2083
rect 660 2077 732 2083
rect 916 2077 1715 2083
rect 884 2057 924 2063
rect 964 2057 1036 2063
rect 1044 2057 1548 2063
rect 1709 2063 1715 2077
rect 1885 2083 1891 2096
rect 1732 2077 1891 2083
rect 1940 2077 2012 2083
rect 2532 2077 3356 2083
rect 3572 2077 3820 2083
rect 3860 2077 4476 2083
rect 4484 2077 4492 2083
rect 4500 2077 4691 2083
rect 1709 2057 1740 2063
rect 1757 2057 1852 2063
rect 740 2037 972 2043
rect 980 2037 1324 2043
rect 1460 2037 1516 2043
rect 1757 2043 1763 2057
rect 1860 2057 2172 2063
rect 2180 2057 2508 2063
rect 2612 2057 2940 2063
rect 3316 2057 4236 2063
rect 4308 2057 4428 2063
rect 4436 2057 4604 2063
rect 4685 2063 4691 2077
rect 4724 2077 5004 2083
rect 5012 2077 5100 2083
rect 5108 2077 6108 2083
rect 6196 2077 6572 2083
rect 6660 2077 6716 2083
rect 7108 2077 7116 2083
rect 7188 2077 7212 2083
rect 4685 2057 4844 2063
rect 5044 2057 5340 2063
rect 5357 2057 5884 2063
rect 5357 2044 5363 2057
rect 5972 2057 6220 2063
rect 6228 2057 6252 2063
rect 6260 2057 6332 2063
rect 6340 2057 6428 2063
rect 1524 2037 1763 2043
rect 1828 2037 2028 2043
rect 2868 2037 3164 2043
rect 3396 2037 3468 2043
rect 3604 2037 3676 2043
rect 3700 2037 3836 2043
rect 3844 2037 3868 2043
rect 4244 2037 5356 2043
rect 5476 2037 5836 2043
rect 6628 2037 6892 2043
rect 1380 2017 1539 2023
rect 738 2014 798 2016
rect 738 2006 739 2014
rect 748 2006 749 2014
rect 787 2006 788 2014
rect 797 2006 798 2014
rect 738 2004 798 2006
rect 1012 1997 1516 2003
rect 1533 2003 1539 2017
rect 1588 2017 2524 2023
rect 2548 2017 2956 2023
rect 3844 2017 4700 2023
rect 5012 2017 5036 2023
rect 5108 2017 5148 2023
rect 5236 2017 5788 2023
rect 6068 2017 6396 2023
rect 3746 2014 3806 2016
rect 3746 2006 3747 2014
rect 3756 2006 3757 2014
rect 3795 2006 3796 2014
rect 3805 2006 3806 2014
rect 3746 2004 3806 2006
rect 6754 2014 6814 2016
rect 6754 2006 6755 2014
rect 6764 2006 6765 2014
rect 6803 2006 6804 2014
rect 6813 2006 6814 2014
rect 6754 2004 6814 2006
rect 1533 1997 1580 2003
rect 1613 1997 1628 2003
rect 1613 1983 1619 1997
rect 1940 1997 2028 2003
rect 2772 1997 2988 2003
rect 3012 1997 3580 2003
rect 3828 1997 4204 2003
rect 4564 1997 4684 2003
rect 4788 1997 6716 2003
rect 420 1977 1619 1983
rect 1844 1977 2028 1983
rect 2036 1977 2812 1983
rect 2820 1977 3068 1983
rect 3085 1977 3404 1983
rect 500 1957 524 1963
rect 660 1957 1260 1963
rect 1284 1957 1468 1963
rect 1476 1957 1660 1963
rect 1972 1957 2083 1963
rect 20 1937 300 1943
rect 308 1937 1484 1943
rect 2077 1943 2083 1957
rect 3085 1963 3091 1977
rect 3428 1977 3436 1983
rect 3604 1977 3708 1983
rect 3748 1977 3964 1983
rect 4292 1977 4956 1983
rect 4964 1977 6460 1983
rect 6468 1977 6924 1983
rect 6932 1977 6956 1983
rect 2388 1957 3091 1963
rect 3348 1957 3836 1963
rect 4084 1957 5388 1963
rect 5396 1957 5852 1963
rect 5860 1957 5996 1963
rect 6004 1957 6060 1963
rect 7028 1957 7564 1963
rect 2077 1937 2828 1943
rect 2868 1937 3347 1943
rect 228 1917 268 1923
rect 276 1917 556 1923
rect 980 1917 1052 1923
rect 1140 1917 1292 1923
rect 1316 1917 1388 1923
rect 1460 1917 1564 1923
rect 1572 1917 1580 1923
rect 1652 1917 1868 1923
rect 1924 1917 2060 1923
rect 2100 1917 2300 1923
rect 2356 1917 2867 1923
rect 148 1897 236 1903
rect 516 1897 803 1903
rect 180 1877 332 1883
rect 340 1877 620 1883
rect 628 1877 780 1883
rect 797 1883 803 1897
rect 836 1897 988 1903
rect 1268 1897 1340 1903
rect 1428 1897 1468 1903
rect 1588 1897 1804 1903
rect 1876 1897 1900 1903
rect 1908 1897 1964 1903
rect 2500 1897 2540 1903
rect 2596 1897 2620 1903
rect 2804 1897 2844 1903
rect 2861 1903 2867 1917
rect 3076 1917 3324 1923
rect 3341 1923 3347 1937
rect 3364 1937 3468 1943
rect 3684 1937 3820 1943
rect 3956 1937 5804 1943
rect 5892 1937 6044 1943
rect 6692 1937 7404 1943
rect 3341 1917 3644 1923
rect 3684 1917 3724 1923
rect 4148 1917 4284 1923
rect 4420 1917 4460 1923
rect 4500 1917 4627 1923
rect 2861 1897 3244 1903
rect 3300 1897 3388 1903
rect 3396 1897 3452 1903
rect 3460 1897 3516 1903
rect 3524 1897 3580 1903
rect 3588 1897 3644 1903
rect 3652 1897 3708 1903
rect 4148 1897 4364 1903
rect 4452 1897 4556 1903
rect 4596 1897 4604 1903
rect 4621 1903 4627 1917
rect 4644 1917 4668 1923
rect 4916 1917 5068 1923
rect 5076 1917 5340 1923
rect 5348 1917 5484 1923
rect 5524 1917 5532 1923
rect 5540 1917 5740 1923
rect 6516 1917 6540 1923
rect 6708 1917 7052 1923
rect 7316 1917 7340 1923
rect 7396 1917 7452 1923
rect 7460 1917 7484 1923
rect 4621 1897 4844 1903
rect 4980 1897 5004 1903
rect 5060 1897 5468 1903
rect 5700 1897 5740 1903
rect 5748 1897 5804 1903
rect 5844 1897 5932 1903
rect 5972 1897 6092 1903
rect 6196 1897 6236 1903
rect 6308 1897 6364 1903
rect 6420 1897 6476 1903
rect 6484 1897 6524 1903
rect 6532 1897 6588 1903
rect 6740 1897 6828 1903
rect 7092 1897 7196 1903
rect 7204 1897 7276 1903
rect 7284 1897 7292 1903
rect 7316 1897 7516 1903
rect 797 1877 1068 1883
rect 1124 1877 1372 1883
rect 1501 1877 1596 1883
rect 212 1857 371 1863
rect 365 1844 371 1857
rect 532 1857 668 1863
rect 948 1857 988 1863
rect 996 1857 1020 1863
rect 1108 1857 1180 1863
rect 1501 1863 1507 1877
rect 1604 1877 1676 1883
rect 1716 1877 1820 1883
rect 1876 1877 1932 1883
rect 1972 1877 2204 1883
rect 2228 1877 2428 1883
rect 2436 1877 2460 1883
rect 2468 1877 2748 1883
rect 2804 1877 2876 1883
rect 2900 1877 2972 1883
rect 3236 1877 3260 1883
rect 3316 1877 3404 1883
rect 3444 1877 3500 1883
rect 3508 1877 3564 1883
rect 3572 1877 3628 1883
rect 3636 1877 3692 1883
rect 3716 1877 4332 1883
rect 4436 1877 4908 1883
rect 4948 1877 4995 1883
rect 1188 1857 1507 1863
rect 1524 1857 1932 1863
rect 2004 1857 2188 1863
rect 2196 1857 2268 1863
rect 2532 1857 2588 1863
rect 2612 1857 2620 1863
rect 2740 1857 3004 1863
rect 3428 1857 3532 1863
rect 3668 1857 3948 1863
rect 4244 1857 4300 1863
rect 4404 1857 4412 1863
rect 4420 1857 4844 1863
rect 4900 1857 4972 1863
rect 4989 1863 4995 1877
rect 5012 1877 5116 1883
rect 5380 1877 5516 1883
rect 5764 1877 5916 1883
rect 6228 1877 6348 1883
rect 6420 1877 6492 1883
rect 6516 1877 6988 1883
rect 6996 1877 7052 1883
rect 7220 1877 7244 1883
rect 7348 1877 7500 1883
rect 4989 1857 5436 1863
rect 5684 1857 5772 1863
rect 6132 1857 6220 1863
rect 6228 1857 6332 1863
rect 6548 1857 6604 1863
rect 6612 1857 6684 1863
rect 6900 1857 6956 1863
rect 7508 1857 7548 1863
rect 180 1837 316 1843
rect 372 1837 956 1843
rect 964 1837 1212 1843
rect 1252 1837 1356 1843
rect 1492 1837 2412 1843
rect 2596 1837 2812 1843
rect 3012 1837 3484 1843
rect 3508 1837 3740 1843
rect 3892 1837 4252 1843
rect 4340 1837 4508 1843
rect 4532 1837 4572 1843
rect 4756 1837 4812 1843
rect 4852 1837 5036 1843
rect 5044 1837 5052 1843
rect 5172 1837 5612 1843
rect 7076 1837 7116 1843
rect 7156 1837 7180 1843
rect 852 1817 908 1823
rect 980 1817 1036 1823
rect 1204 1817 1388 1823
rect 1684 1817 1804 1823
rect 1812 1817 2060 1823
rect 2164 1817 2188 1823
rect 2340 1817 3548 1823
rect 3588 1817 3708 1823
rect 3748 1817 4028 1823
rect 4084 1817 4156 1823
rect 4324 1817 4492 1823
rect 4564 1817 4620 1823
rect 4708 1817 4988 1823
rect 5108 1817 5212 1823
rect 5396 1817 5596 1823
rect 5844 1817 5852 1823
rect 2242 1814 2302 1816
rect 2242 1806 2243 1814
rect 2252 1806 2253 1814
rect 2291 1806 2292 1814
rect 2301 1806 2302 1814
rect 2242 1804 2302 1806
rect 20 1797 300 1803
rect 308 1797 572 1803
rect 596 1797 1356 1803
rect 1428 1797 1548 1803
rect 1572 1797 1644 1803
rect 1924 1797 2220 1803
rect 2564 1797 2860 1803
rect 3268 1797 3308 1803
rect 3316 1797 3372 1803
rect 3380 1797 3436 1803
rect 3668 1797 3692 1803
rect 3700 1797 3964 1803
rect 3972 1797 4076 1803
rect 4260 1797 4460 1803
rect 4493 1803 4499 1816
rect 5250 1814 5310 1816
rect 5250 1806 5251 1814
rect 5260 1806 5261 1814
rect 5299 1806 5300 1814
rect 5309 1806 5310 1814
rect 5250 1804 5310 1806
rect 4493 1797 4636 1803
rect 4932 1797 5212 1803
rect 5332 1797 5404 1803
rect 5476 1797 5628 1803
rect 6020 1797 6124 1803
rect 6372 1797 6412 1803
rect 6420 1797 6860 1803
rect 6868 1797 6892 1803
rect 7252 1797 7420 1803
rect 7428 1797 7548 1803
rect 580 1777 652 1783
rect 660 1777 1692 1783
rect 1700 1777 1900 1783
rect 1908 1777 2556 1783
rect 2708 1777 2764 1783
rect 2788 1777 3324 1783
rect 3341 1777 3500 1783
rect 484 1757 588 1763
rect 852 1757 988 1763
rect 1012 1757 1228 1763
rect 1396 1757 1468 1763
rect 1492 1757 1580 1763
rect 1636 1757 1692 1763
rect 1860 1757 1932 1763
rect 1988 1757 2044 1763
rect 2052 1757 2460 1763
rect 2468 1757 2764 1763
rect 2788 1757 3228 1763
rect 3341 1763 3347 1777
rect 3604 1777 3900 1783
rect 4052 1777 4140 1783
rect 4148 1777 4556 1783
rect 4804 1777 4876 1783
rect 4932 1777 5372 1783
rect 5444 1777 5548 1783
rect 5588 1777 5916 1783
rect 6116 1777 6460 1783
rect 6596 1777 6604 1783
rect 6740 1777 6988 1783
rect 7380 1777 7452 1783
rect 7524 1777 7532 1783
rect 3252 1757 3347 1763
rect 3380 1757 3468 1763
rect 3572 1757 3644 1763
rect 3652 1757 3724 1763
rect 3732 1757 3868 1763
rect 3876 1757 3932 1763
rect 4100 1757 4172 1763
rect 4180 1757 4428 1763
rect 4436 1757 4492 1763
rect 4500 1757 4540 1763
rect 4884 1757 4956 1763
rect 5236 1757 5324 1763
rect 5364 1757 5420 1763
rect 5460 1757 5676 1763
rect 5684 1757 5900 1763
rect 6068 1757 6140 1763
rect 6692 1757 6828 1763
rect 6948 1757 6972 1763
rect 7108 1757 7116 1763
rect 7252 1757 7516 1763
rect 7524 1757 7548 1763
rect 148 1737 236 1743
rect 692 1737 1004 1743
rect 1076 1737 1260 1743
rect 1300 1737 1324 1743
rect 1332 1737 1452 1743
rect 1508 1737 1516 1743
rect 1524 1737 1644 1743
rect 1716 1737 2060 1743
rect 2100 1737 2172 1743
rect 2196 1737 2348 1743
rect 2580 1737 2620 1743
rect 2628 1737 3468 1743
rect 3476 1737 3820 1743
rect 4068 1737 4188 1743
rect 4196 1737 4396 1743
rect 4484 1737 4572 1743
rect 4804 1737 5116 1743
rect 5124 1737 5452 1743
rect 5812 1737 5900 1743
rect 6180 1737 6252 1743
rect 6260 1737 6860 1743
rect 7268 1737 7308 1743
rect 7364 1737 7388 1743
rect 116 1717 220 1723
rect 228 1717 268 1723
rect 276 1717 332 1723
rect 388 1717 428 1723
rect 548 1717 700 1723
rect 900 1717 972 1723
rect 1076 1717 1612 1723
rect 1796 1717 1836 1723
rect 2052 1717 2108 1723
rect 2132 1717 2188 1723
rect 2404 1717 2572 1723
rect 2852 1717 2860 1723
rect 3124 1717 3292 1723
rect 3620 1717 3836 1723
rect 3860 1717 4236 1723
rect 4276 1717 4284 1723
rect 4292 1717 4668 1723
rect 4676 1717 4844 1723
rect 4884 1717 5020 1723
rect 5156 1717 5436 1723
rect 5508 1717 5564 1723
rect 5652 1717 5676 1723
rect 5732 1717 5820 1723
rect 5844 1717 6092 1723
rect 6148 1717 6220 1723
rect 6340 1717 6828 1723
rect 6868 1717 7004 1723
rect 7092 1717 7196 1723
rect 7492 1717 7500 1723
rect 228 1697 508 1703
rect 516 1697 556 1703
rect 916 1697 1004 1703
rect 1044 1697 1116 1703
rect 1124 1697 1132 1703
rect 1348 1697 1548 1703
rect 1620 1697 1964 1703
rect 2036 1697 2108 1703
rect 2164 1697 2204 1703
rect 2228 1697 2348 1703
rect 2436 1697 2732 1703
rect 2756 1697 2860 1703
rect 2868 1697 3020 1703
rect 3028 1697 3084 1703
rect 3284 1697 3308 1703
rect 3540 1697 3660 1703
rect 3828 1697 3900 1703
rect 3988 1697 4012 1703
rect 4292 1697 4684 1703
rect 4852 1697 5164 1703
rect 5412 1697 5436 1703
rect 5460 1697 5532 1703
rect 5540 1697 5596 1703
rect 5604 1697 5676 1703
rect 5684 1697 5932 1703
rect 6212 1697 6300 1703
rect 6484 1697 6508 1703
rect 6564 1697 6860 1703
rect 7044 1697 7052 1703
rect 7220 1697 7276 1703
rect 7444 1697 7484 1703
rect 756 1677 892 1683
rect 900 1677 1068 1683
rect 1092 1677 1148 1683
rect 1236 1677 1244 1683
rect 1252 1677 1404 1683
rect 1412 1677 1532 1683
rect 1540 1677 1804 1683
rect 1821 1677 1868 1683
rect 964 1657 1052 1663
rect 1108 1657 1148 1663
rect 1364 1657 1404 1663
rect 1476 1657 1724 1663
rect 1821 1663 1827 1677
rect 1940 1677 2060 1683
rect 2084 1677 2364 1683
rect 2388 1677 2412 1683
rect 2484 1677 3052 1683
rect 3076 1677 3212 1683
rect 3284 1677 3308 1683
rect 3524 1677 3596 1683
rect 3668 1677 4028 1683
rect 4036 1677 4140 1683
rect 4148 1677 4259 1683
rect 1780 1657 1827 1663
rect 1844 1657 2268 1663
rect 2308 1657 2828 1663
rect 3556 1657 4236 1663
rect 4253 1663 4259 1677
rect 4484 1677 4652 1683
rect 4980 1677 5132 1683
rect 5396 1677 5484 1683
rect 5524 1677 5836 1683
rect 5940 1677 6028 1683
rect 6420 1677 6444 1683
rect 6628 1677 6652 1683
rect 6756 1677 6940 1683
rect 7012 1677 7068 1683
rect 7172 1677 7292 1683
rect 7316 1677 7340 1683
rect 4253 1657 4396 1663
rect 4404 1657 4588 1663
rect 4996 1657 5196 1663
rect 5252 1657 6700 1663
rect 7140 1657 7180 1663
rect 7188 1657 7388 1663
rect 516 1637 860 1643
rect 1028 1637 1356 1643
rect 1364 1637 1644 1643
rect 1764 1637 2332 1643
rect 2356 1637 3308 1643
rect 3732 1637 4124 1643
rect 4132 1637 4236 1643
rect 4244 1637 4444 1643
rect 4468 1637 4732 1643
rect 4852 1637 5692 1643
rect 5700 1637 5740 1643
rect 5780 1637 5980 1643
rect 6644 1637 6748 1643
rect 7268 1637 7276 1643
rect 1076 1617 1212 1623
rect 1220 1617 1500 1623
rect 1508 1617 1772 1623
rect 1780 1617 1964 1623
rect 2068 1617 2252 1623
rect 2692 1617 2764 1623
rect 2804 1617 3132 1623
rect 3236 1617 3708 1623
rect 4228 1617 4300 1623
rect 4340 1617 5500 1623
rect 5524 1617 5548 1623
rect 7284 1617 7324 1623
rect 738 1614 798 1616
rect 738 1606 739 1614
rect 748 1606 749 1614
rect 787 1606 788 1614
rect 797 1606 798 1614
rect 738 1604 798 1606
rect 3746 1614 3806 1616
rect 3746 1606 3747 1614
rect 3756 1606 3757 1614
rect 3795 1606 3796 1614
rect 3805 1606 3806 1614
rect 3746 1604 3806 1606
rect 6754 1614 6814 1616
rect 6754 1606 6755 1614
rect 6764 1606 6765 1614
rect 6803 1606 6804 1614
rect 6813 1606 6814 1614
rect 6754 1604 6814 1606
rect 1188 1597 1820 1603
rect 1844 1597 1932 1603
rect 2020 1597 2163 1603
rect 564 1577 1132 1583
rect 1316 1577 1516 1583
rect 1748 1577 1868 1583
rect 1924 1577 1948 1583
rect 1988 1577 2028 1583
rect 2100 1577 2140 1583
rect 2157 1583 2163 1597
rect 2276 1597 2700 1603
rect 2740 1597 2988 1603
rect 3012 1597 3212 1603
rect 3476 1597 3596 1603
rect 3821 1597 5228 1603
rect 2157 1577 2252 1583
rect 2292 1577 2412 1583
rect 2564 1577 2732 1583
rect 2772 1577 2860 1583
rect 2884 1577 2924 1583
rect 3028 1577 3052 1583
rect 3821 1583 3827 1597
rect 5492 1597 5596 1603
rect 5604 1597 5708 1603
rect 5716 1597 5884 1603
rect 3636 1577 3827 1583
rect 3837 1577 4044 1583
rect 1012 1557 1116 1563
rect 1133 1563 1139 1576
rect 1133 1557 1388 1563
rect 1396 1557 1532 1563
rect 1588 1557 1996 1563
rect 2084 1557 2508 1563
rect 2740 1557 3020 1563
rect 3572 1557 3603 1563
rect 420 1537 636 1543
rect 644 1537 1283 1543
rect 1277 1524 1283 1537
rect 1316 1537 1980 1543
rect 2004 1537 2060 1543
rect 2068 1537 2204 1543
rect 2212 1537 2236 1543
rect 2244 1537 2380 1543
rect 2388 1537 2444 1543
rect 2532 1537 2556 1543
rect 2692 1537 2956 1543
rect 3044 1537 3132 1543
rect 3597 1543 3603 1557
rect 3837 1563 3843 1577
rect 4116 1577 4348 1583
rect 4356 1577 4652 1583
rect 4660 1577 4892 1583
rect 4900 1577 5100 1583
rect 5124 1577 5180 1583
rect 5268 1577 5388 1583
rect 5412 1577 6188 1583
rect 6292 1577 7388 1583
rect 3812 1557 3843 1563
rect 3876 1557 3884 1563
rect 3956 1557 5644 1563
rect 6292 1557 6332 1563
rect 3597 1537 4243 1543
rect 525 1517 604 1523
rect 525 1504 531 1517
rect 1012 1517 1043 1523
rect 1037 1504 1043 1517
rect 1124 1517 1260 1523
rect 1284 1517 1372 1523
rect 1524 1517 2172 1523
rect 2196 1517 2396 1523
rect 2404 1517 2540 1523
rect 2548 1517 2620 1523
rect 2628 1517 2700 1523
rect 2708 1517 2748 1523
rect 2836 1517 2940 1523
rect 3044 1517 3084 1523
rect 3124 1517 3244 1523
rect 3380 1517 3596 1523
rect 3684 1517 3724 1523
rect 3764 1517 4108 1523
rect 4116 1517 4220 1523
rect 4237 1523 4243 1537
rect 4260 1537 4284 1543
rect 4301 1537 4460 1543
rect 4301 1523 4307 1537
rect 4516 1537 4572 1543
rect 4628 1537 4684 1543
rect 4756 1537 6236 1543
rect 6340 1537 6908 1543
rect 7012 1537 7212 1543
rect 4237 1517 4307 1523
rect 4356 1517 4380 1523
rect 4404 1517 4796 1523
rect 4804 1517 4940 1523
rect 4948 1517 5004 1523
rect 5044 1517 5068 1523
rect 5108 1517 5148 1523
rect 5156 1517 5228 1523
rect 5380 1517 5500 1523
rect 5572 1517 5612 1523
rect 5956 1517 5996 1523
rect 6100 1517 6140 1523
rect 6372 1517 6444 1523
rect 6468 1517 6732 1523
rect 6749 1517 6972 1523
rect 52 1497 108 1503
rect 148 1497 220 1503
rect 452 1497 492 1503
rect 500 1497 524 1503
rect 548 1497 652 1503
rect 820 1497 1020 1503
rect 1044 1497 1132 1503
rect 1156 1497 1340 1503
rect 1348 1497 1436 1503
rect 1524 1497 1644 1503
rect 1764 1497 1788 1503
rect 1892 1497 2012 1503
rect 2052 1497 2220 1503
rect 2228 1497 2380 1503
rect 2388 1497 2444 1503
rect 2532 1497 2860 1503
rect 2964 1497 3084 1503
rect 3092 1497 3212 1503
rect 3677 1503 3683 1516
rect 3252 1497 3683 1503
rect 3716 1497 3884 1503
rect 4116 1497 4172 1503
rect 4180 1497 4188 1503
rect 4276 1497 4364 1503
rect 4516 1497 4524 1503
rect 4532 1497 4876 1503
rect 4884 1497 5356 1503
rect 5364 1497 5532 1503
rect 5540 1497 5548 1503
rect 5844 1497 5916 1503
rect 5924 1497 6012 1503
rect 6020 1497 6044 1503
rect 6061 1497 6332 1503
rect 340 1477 668 1483
rect 676 1477 716 1483
rect 1092 1477 1180 1483
rect 1188 1477 1452 1483
rect 1460 1477 1564 1483
rect 1924 1477 2284 1483
rect 2308 1477 2348 1483
rect 2516 1477 2764 1483
rect 2957 1483 2963 1496
rect 2852 1477 2963 1483
rect 3348 1477 3644 1483
rect 3652 1477 3699 1483
rect 3693 1464 3699 1477
rect 3732 1477 3868 1483
rect 3876 1477 4012 1483
rect 4020 1477 4092 1483
rect 4212 1477 4236 1483
rect 4260 1477 4396 1483
rect 4484 1477 4924 1483
rect 4932 1477 5052 1483
rect 5060 1477 5324 1483
rect 5332 1477 5500 1483
rect 5556 1477 5740 1483
rect 6061 1483 6067 1497
rect 6372 1497 6396 1503
rect 6452 1497 6572 1503
rect 6749 1503 6755 1517
rect 6996 1517 7052 1523
rect 7140 1517 7164 1523
rect 7380 1517 7468 1523
rect 6708 1497 6755 1503
rect 6868 1497 6940 1503
rect 7028 1497 7292 1503
rect 7524 1497 7532 1503
rect 7572 1497 7603 1503
rect 5988 1477 6067 1483
rect 6084 1477 6124 1483
rect 6180 1477 6220 1483
rect 6244 1477 6300 1483
rect 6404 1477 6428 1483
rect 6436 1477 6524 1483
rect 6532 1477 6636 1483
rect 6740 1477 6908 1483
rect 6916 1477 6988 1483
rect 7124 1477 7292 1483
rect 7348 1477 7500 1483
rect 308 1457 572 1463
rect 877 1457 1212 1463
rect 877 1443 883 1457
rect 1492 1457 1548 1463
rect 1604 1457 1756 1463
rect 1796 1457 1868 1463
rect 1940 1457 1948 1463
rect 2004 1457 2156 1463
rect 2180 1457 2236 1463
rect 2260 1457 2380 1463
rect 2644 1457 2684 1463
rect 2708 1457 2828 1463
rect 2948 1457 3068 1463
rect 3284 1457 3580 1463
rect 3652 1457 3660 1463
rect 3700 1457 3740 1463
rect 4036 1457 4172 1463
rect 4180 1457 4236 1463
rect 4308 1457 4380 1463
rect 5428 1457 5708 1463
rect 5780 1457 5820 1463
rect 6324 1457 6428 1463
rect 6500 1457 6524 1463
rect 6644 1457 6668 1463
rect 6964 1457 7020 1463
rect 7316 1457 7340 1463
rect 7476 1457 7500 1463
rect 388 1437 883 1443
rect 1044 1437 1068 1443
rect 1092 1437 1100 1443
rect 1556 1437 1660 1443
rect 2036 1437 2156 1443
rect 2180 1437 2300 1443
rect 2324 1437 3548 1443
rect 3636 1437 3820 1443
rect 3828 1437 4108 1443
rect 4116 1437 4364 1443
rect 4381 1437 5388 1443
rect 132 1417 428 1423
rect 436 1417 988 1423
rect 996 1417 1324 1423
rect 1332 1417 1628 1423
rect 1636 1417 1996 1423
rect 2404 1417 2716 1423
rect 3028 1417 3180 1423
rect 3188 1417 3756 1423
rect 4381 1423 4387 1437
rect 5428 1437 5964 1443
rect 6276 1437 6460 1443
rect 6964 1437 6988 1443
rect 7060 1437 7100 1443
rect 7252 1437 7324 1443
rect 3780 1417 4387 1423
rect 4452 1417 4684 1423
rect 4692 1417 4780 1423
rect 4788 1417 4908 1423
rect 4916 1417 5100 1423
rect 5668 1417 5788 1423
rect 5796 1417 5948 1423
rect 5956 1417 5996 1423
rect 6004 1417 6028 1423
rect 6244 1417 6684 1423
rect 6932 1417 7052 1423
rect 2242 1414 2302 1416
rect 2242 1406 2243 1414
rect 2252 1406 2253 1414
rect 2291 1406 2292 1414
rect 2301 1406 2302 1414
rect 2242 1404 2302 1406
rect 5250 1414 5310 1416
rect 5250 1406 5251 1414
rect 5260 1406 5261 1414
rect 5299 1406 5300 1414
rect 5309 1406 5310 1414
rect 5250 1404 5310 1406
rect 532 1397 579 1403
rect 573 1384 579 1397
rect 756 1397 1020 1403
rect 1028 1397 1148 1403
rect 1236 1397 1340 1403
rect 1348 1397 1580 1403
rect 1604 1397 1724 1403
rect 1940 1397 2220 1403
rect 2452 1397 3276 1403
rect 4180 1397 4316 1403
rect 4548 1397 4764 1403
rect 4788 1397 4876 1403
rect 4884 1397 5164 1403
rect 6068 1397 6444 1403
rect 6932 1397 6956 1403
rect 7060 1397 7180 1403
rect 196 1377 380 1383
rect 580 1377 659 1383
rect 653 1364 659 1377
rect 916 1377 1068 1383
rect 1108 1377 1260 1383
rect 1268 1377 1420 1383
rect 1460 1377 1532 1383
rect 1588 1377 1692 1383
rect 1764 1377 2028 1383
rect 2068 1377 2124 1383
rect 2148 1377 2188 1383
rect 2596 1377 2700 1383
rect 2756 1377 2844 1383
rect 2884 1377 2956 1383
rect 3220 1377 3308 1383
rect 3348 1377 3548 1383
rect 3604 1377 3772 1383
rect 3796 1377 4284 1383
rect 4548 1377 4716 1383
rect 4740 1377 4972 1383
rect 5188 1377 5388 1383
rect 5908 1377 6108 1383
rect 7364 1377 7404 1383
rect 20 1357 611 1363
rect 605 1344 611 1357
rect 660 1357 748 1363
rect 1252 1357 1324 1363
rect 1524 1357 1564 1363
rect 1588 1357 1708 1363
rect 1748 1357 1788 1363
rect 1972 1357 2540 1363
rect 2564 1357 3372 1363
rect 3396 1357 3404 1363
rect 3828 1357 3916 1363
rect 4228 1357 4364 1363
rect 4452 1357 4492 1363
rect 4500 1357 4588 1363
rect 4708 1357 4844 1363
rect 4964 1357 4988 1363
rect 5124 1357 5196 1363
rect 5492 1357 5564 1363
rect 5764 1357 5939 1363
rect 5933 1344 5939 1357
rect 6020 1357 6124 1363
rect 6148 1357 6204 1363
rect 6292 1357 6332 1363
rect 6452 1357 6604 1363
rect 6660 1357 6684 1363
rect 6884 1357 7036 1363
rect 7044 1357 7132 1363
rect 7156 1357 7180 1363
rect 7236 1357 7292 1363
rect 7300 1357 7324 1363
rect 7348 1357 7436 1363
rect 292 1337 412 1343
rect 612 1337 684 1343
rect 708 1337 892 1343
rect 916 1337 1052 1343
rect 1060 1337 1100 1343
rect 1140 1337 1148 1343
rect 1156 1337 1356 1343
rect 1684 1337 1756 1343
rect 1812 1337 1948 1343
rect 1972 1337 1980 1343
rect 2004 1337 2044 1343
rect 2196 1337 2332 1343
rect 2372 1337 2412 1343
rect 2484 1337 2668 1343
rect 2692 1337 2892 1343
rect 2900 1337 2924 1343
rect 3076 1337 3292 1343
rect 3300 1337 3356 1343
rect 3364 1337 3420 1343
rect 3428 1337 3484 1343
rect 3748 1337 4124 1343
rect 4132 1337 4188 1343
rect 4340 1337 4492 1343
rect 4580 1337 4636 1343
rect 4836 1337 4860 1343
rect 4996 1337 5020 1343
rect 5037 1337 5532 1343
rect 5037 1324 5043 1337
rect 5540 1337 5628 1343
rect 5636 1337 5772 1343
rect 5940 1337 6060 1343
rect 6116 1337 6412 1343
rect 6420 1337 6588 1343
rect 7076 1337 7164 1343
rect 7172 1337 7276 1343
rect 7332 1337 7452 1343
rect 180 1317 252 1323
rect 516 1317 1836 1323
rect 2004 1317 2012 1323
rect 2036 1317 2300 1323
rect 2340 1317 2556 1323
rect 2628 1317 2732 1323
rect 2820 1317 3212 1323
rect 3316 1317 3372 1323
rect 3380 1317 3436 1323
rect 3444 1317 3468 1323
rect 3492 1317 3532 1323
rect 3556 1317 3580 1323
rect 3780 1317 3916 1323
rect 3956 1317 4179 1323
rect 4173 1304 4179 1317
rect 4228 1317 4236 1323
rect 4244 1317 4332 1323
rect 4468 1317 4604 1323
rect 4740 1317 4828 1323
rect 4836 1317 5020 1323
rect 5172 1317 5308 1323
rect 5412 1317 5436 1323
rect 5460 1317 5580 1323
rect 5876 1317 5964 1323
rect 6004 1317 6092 1323
rect 6100 1317 6156 1323
rect 6196 1317 6220 1323
rect 6324 1317 6348 1323
rect 6356 1317 6508 1323
rect 7012 1317 7148 1323
rect 7156 1317 7180 1323
rect 7316 1317 7340 1323
rect 7396 1317 7452 1323
rect 7460 1317 7500 1323
rect 724 1297 1244 1303
rect 1268 1297 1292 1303
rect 1364 1297 1452 1303
rect 1524 1297 1564 1303
rect 1668 1297 1676 1303
rect 1700 1297 1756 1303
rect 1764 1297 1820 1303
rect 2164 1297 2316 1303
rect 2356 1297 2460 1303
rect 2468 1297 2524 1303
rect 2564 1297 2796 1303
rect 2820 1297 2844 1303
rect 3028 1297 3500 1303
rect 3540 1297 3596 1303
rect 3684 1297 4044 1303
rect 4132 1297 4156 1303
rect 4180 1297 4332 1303
rect 4372 1297 4652 1303
rect 4660 1297 4723 1303
rect 644 1277 1164 1283
rect 1204 1277 1276 1283
rect 1412 1277 1644 1283
rect 1700 1277 1804 1283
rect 2036 1277 2492 1283
rect 2516 1277 2540 1283
rect 2701 1277 3004 1283
rect 1188 1257 1292 1263
rect 1332 1257 1795 1263
rect 372 1237 1187 1243
rect 1181 1223 1187 1237
rect 1204 1237 1612 1243
rect 1789 1243 1795 1257
rect 1812 1257 1852 1263
rect 1908 1257 2044 1263
rect 2701 1263 2707 1277
rect 3028 1277 3052 1283
rect 3124 1277 3196 1283
rect 3220 1277 3372 1283
rect 3412 1277 3788 1283
rect 4212 1277 4435 1283
rect 2228 1257 2707 1263
rect 2724 1257 3132 1263
rect 3140 1257 3244 1263
rect 3284 1257 3308 1263
rect 3332 1257 3948 1263
rect 3972 1257 4412 1263
rect 4429 1263 4435 1277
rect 4468 1277 4700 1283
rect 4717 1283 4723 1297
rect 4948 1297 5116 1303
rect 5156 1297 5884 1303
rect 6340 1297 6524 1303
rect 6532 1297 6556 1303
rect 6596 1297 6636 1303
rect 6676 1297 7116 1303
rect 7172 1297 7180 1303
rect 7204 1297 7292 1303
rect 7572 1297 7603 1303
rect 4717 1277 5356 1283
rect 6436 1277 6476 1283
rect 6580 1277 6636 1283
rect 7060 1277 7084 1283
rect 7188 1277 7228 1283
rect 7268 1277 7484 1283
rect 4429 1257 5612 1263
rect 6596 1257 6908 1263
rect 6916 1257 6972 1263
rect 7476 1257 7564 1263
rect 1789 1237 1900 1243
rect 1972 1237 2172 1243
rect 2196 1237 2428 1243
rect 2516 1237 2796 1243
rect 2900 1237 3676 1243
rect 3700 1237 3827 1243
rect 1181 1217 1308 1223
rect 1348 1217 1532 1223
rect 1540 1217 1676 1223
rect 1684 1217 1852 1223
rect 1860 1217 2092 1223
rect 2100 1217 2604 1223
rect 2660 1217 3372 1223
rect 3821 1223 3827 1237
rect 4084 1237 4268 1243
rect 4308 1237 4332 1243
rect 4340 1237 4428 1243
rect 4612 1237 5404 1243
rect 3821 1217 4780 1223
rect 5012 1217 5052 1223
rect 5076 1217 5212 1223
rect 5380 1217 5420 1223
rect 738 1214 798 1216
rect 738 1206 739 1214
rect 748 1206 749 1214
rect 787 1206 788 1214
rect 797 1206 798 1214
rect 738 1204 798 1206
rect 3746 1214 3806 1216
rect 3746 1206 3747 1214
rect 3756 1206 3757 1214
rect 3795 1206 3796 1214
rect 3805 1206 3806 1214
rect 3746 1204 3806 1206
rect 6754 1214 6814 1216
rect 6754 1206 6755 1214
rect 6764 1206 6765 1214
rect 6803 1206 6804 1214
rect 6813 1206 6814 1214
rect 6754 1204 6814 1206
rect 1117 1197 2108 1203
rect 1117 1183 1123 1197
rect 2180 1197 2348 1203
rect 2580 1197 2620 1203
rect 2980 1197 3724 1203
rect 4324 1197 5436 1203
rect 5620 1197 6540 1203
rect 388 1177 1123 1183
rect 1172 1177 1212 1183
rect 1556 1177 2092 1183
rect 2132 1177 2188 1183
rect 2276 1177 2508 1183
rect 2532 1177 2732 1183
rect 2749 1177 2892 1183
rect 468 1157 2188 1163
rect 2749 1163 2755 1177
rect 2932 1177 2972 1183
rect 3204 1177 3276 1183
rect 3316 1177 3916 1183
rect 4164 1177 4204 1183
rect 4212 1177 4732 1183
rect 5076 1177 5340 1183
rect 5364 1177 6156 1183
rect 6804 1177 6956 1183
rect 6964 1177 7132 1183
rect 2308 1157 2755 1163
rect 2772 1157 3372 1163
rect 3956 1157 4060 1163
rect 4228 1157 4268 1163
rect 4276 1157 5884 1163
rect 788 1137 2003 1143
rect 644 1117 700 1123
rect 1012 1117 1052 1123
rect 1060 1117 1084 1123
rect 1108 1117 1203 1123
rect 637 1103 643 1116
rect -35 1097 643 1103
rect 692 1097 876 1103
rect 980 1097 1011 1103
rect 868 1077 988 1083
rect 1005 1083 1011 1097
rect 1108 1097 1116 1103
rect 1197 1103 1203 1117
rect 1220 1117 1228 1123
rect 1524 1117 1644 1123
rect 1652 1117 1724 1123
rect 1812 1117 1964 1123
rect 1997 1123 2003 1137
rect 2020 1137 2076 1143
rect 2084 1137 2140 1143
rect 2148 1137 2204 1143
rect 2212 1137 2364 1143
rect 2372 1137 2444 1143
rect 2452 1137 2508 1143
rect 2740 1137 2940 1143
rect 3284 1137 3308 1143
rect 3876 1137 4348 1143
rect 4356 1137 5004 1143
rect 5028 1137 5196 1143
rect 5220 1137 5628 1143
rect 5780 1137 5836 1143
rect 6340 1137 6476 1143
rect 6484 1137 6604 1143
rect 6660 1137 6716 1143
rect 1997 1117 2476 1123
rect 2740 1117 2764 1123
rect 2836 1117 3020 1123
rect 3044 1117 3180 1123
rect 3284 1117 3420 1123
rect 3508 1117 3628 1123
rect 3732 1117 3964 1123
rect 4004 1117 4252 1123
rect 4276 1117 4364 1123
rect 4420 1117 4684 1123
rect 4820 1117 4876 1123
rect 5044 1117 5196 1123
rect 5204 1117 5468 1123
rect 5476 1117 5612 1123
rect 5796 1117 5836 1123
rect 5876 1117 6044 1123
rect 6260 1117 6284 1123
rect 6292 1117 6348 1123
rect 6516 1117 6892 1123
rect 6916 1117 6972 1123
rect 1197 1097 1548 1103
rect 1556 1097 1596 1103
rect 1972 1097 2140 1103
rect 2164 1097 2236 1103
rect 2420 1097 2476 1103
rect 2548 1097 2636 1103
rect 2644 1097 2684 1103
rect 2772 1097 2796 1103
rect 2900 1097 3836 1103
rect 3892 1097 4060 1103
rect 4068 1097 4140 1103
rect 4308 1097 4396 1103
rect 4404 1097 4828 1103
rect 4836 1097 4844 1103
rect 5140 1097 5235 1103
rect 1005 1077 1100 1083
rect 1108 1077 1164 1083
rect 1444 1077 1516 1083
rect 1652 1077 1980 1083
rect 2004 1077 2060 1083
rect 2068 1077 2124 1083
rect 2132 1077 2188 1083
rect 2196 1077 2364 1083
rect 2372 1077 2428 1083
rect 2436 1077 2492 1083
rect 2516 1077 2604 1083
rect 2756 1077 2780 1083
rect 2788 1077 2828 1083
rect 2852 1077 2892 1083
rect 3092 1077 3132 1083
rect 3172 1077 3196 1083
rect 3284 1077 3308 1083
rect 3396 1077 3539 1083
rect 596 1057 2764 1063
rect 2916 1057 3244 1063
rect 3309 1063 3315 1076
rect 3309 1057 3404 1063
rect 3412 1057 3420 1063
rect 3428 1057 3468 1063
rect 3476 1057 3484 1063
rect 3492 1057 3516 1063
rect 3533 1063 3539 1077
rect 3556 1077 3564 1083
rect 3668 1077 3708 1083
rect 3716 1077 3820 1083
rect 3940 1077 3980 1083
rect 4132 1077 4316 1083
rect 4388 1077 4412 1083
rect 4436 1077 4460 1083
rect 4516 1077 4652 1083
rect 4852 1077 4924 1083
rect 4932 1077 5084 1083
rect 5229 1083 5235 1097
rect 5252 1097 5500 1103
rect 6020 1097 6124 1103
rect 6212 1097 6220 1103
rect 6228 1097 6268 1103
rect 6372 1097 6460 1103
rect 6676 1097 6748 1103
rect 7188 1097 7372 1103
rect 7380 1097 7404 1103
rect 7444 1097 7468 1103
rect 7492 1097 7564 1103
rect 5229 1077 5292 1083
rect 5428 1077 5788 1083
rect 5940 1077 5996 1083
rect 6004 1077 6108 1083
rect 6260 1077 6268 1083
rect 6468 1077 6652 1083
rect 7316 1077 7516 1083
rect 3533 1057 3724 1063
rect 3821 1063 3827 1076
rect 3821 1057 3884 1063
rect 3892 1057 3916 1063
rect 3924 1057 3948 1063
rect 4148 1057 4332 1063
rect 4628 1057 4860 1063
rect 4868 1057 5212 1063
rect 5293 1063 5299 1076
rect 5293 1057 5420 1063
rect 5844 1057 6188 1063
rect 6228 1057 6332 1063
rect 6644 1057 6732 1063
rect 6820 1057 6844 1063
rect 6852 1057 6924 1063
rect 6932 1057 6940 1063
rect 6948 1057 7100 1063
rect 7236 1057 7292 1063
rect 7300 1057 7468 1063
rect 7476 1057 7500 1063
rect 164 1037 204 1043
rect 212 1037 316 1043
rect 1412 1037 2844 1043
rect 2884 1037 2956 1043
rect 2980 1037 3052 1043
rect 3124 1037 3196 1043
rect 3252 1037 3324 1043
rect 3380 1037 3388 1043
rect 3540 1037 5964 1043
rect 6148 1037 6172 1043
rect 6180 1037 6252 1043
rect 6260 1037 6300 1043
rect 6308 1037 6380 1043
rect 6436 1037 6572 1043
rect 6580 1037 6700 1043
rect 6740 1037 6876 1043
rect 7076 1037 7116 1043
rect 7124 1037 7372 1043
rect 20 1017 460 1023
rect 820 1017 860 1023
rect 1220 1017 1964 1023
rect 2068 1017 2092 1023
rect 2148 1017 2156 1023
rect 2596 1017 2812 1023
rect 2868 1017 3020 1023
rect 3076 1017 3148 1023
rect 3156 1017 3164 1023
rect 3236 1017 3900 1023
rect 3972 1017 4220 1023
rect 4756 1017 4924 1023
rect 4932 1017 5148 1023
rect 5588 1017 5596 1023
rect 6548 1017 6572 1023
rect 7092 1017 7516 1023
rect 2242 1014 2302 1016
rect 2242 1006 2243 1014
rect 2252 1006 2253 1014
rect 2291 1006 2292 1014
rect 2301 1006 2302 1014
rect 2242 1004 2302 1006
rect 5250 1014 5310 1016
rect 5250 1006 5251 1014
rect 5260 1006 5261 1014
rect 5299 1006 5300 1014
rect 5309 1006 5310 1014
rect 5250 1004 5310 1006
rect -35 997 268 1003
rect 916 997 1116 1003
rect 1124 997 1244 1003
rect 1364 997 1452 1003
rect 1524 997 1708 1003
rect 2084 997 2172 1003
rect 2404 997 2556 1003
rect 2628 997 2684 1003
rect 2692 997 3356 1003
rect 3380 997 3859 1003
rect 388 977 444 983
rect 884 977 940 983
rect 964 977 1388 983
rect 1588 977 1667 983
rect -35 957 12 963
rect 292 957 396 963
rect 420 957 476 963
rect 516 957 620 963
rect 628 957 652 963
rect 1204 957 1260 963
rect 1428 957 1612 963
rect 1661 963 1667 977
rect 1684 977 2476 983
rect 2516 977 2540 983
rect 2557 977 2588 983
rect 1661 957 1836 963
rect 2004 957 2099 963
rect 228 937 252 943
rect 308 937 428 943
rect 436 937 604 943
rect 612 937 1148 943
rect 1188 937 1228 943
rect 1236 937 1292 943
rect 1316 937 1372 943
rect 1476 937 1859 943
rect -35 903 -29 923
rect 276 917 348 923
rect 388 917 428 923
rect 484 917 604 923
rect 756 917 812 923
rect 1092 917 1180 923
rect 1252 917 1324 923
rect 1444 917 1484 923
rect 1492 917 1644 923
rect 1853 923 1859 937
rect 1876 937 1964 943
rect 1972 937 2060 943
rect 2093 943 2099 957
rect 2228 957 2252 963
rect 2260 957 2380 963
rect 2388 957 2460 963
rect 2557 963 2563 977
rect 2628 977 2652 983
rect 2685 977 2876 983
rect 2548 957 2563 963
rect 2685 963 2691 977
rect 3060 977 3084 983
rect 3108 977 3228 983
rect 3316 977 3324 983
rect 3508 977 3836 983
rect 3853 983 3859 997
rect 3876 997 4716 1003
rect 5460 997 5516 1003
rect 5524 997 5916 1003
rect 6516 997 7004 1003
rect 7252 997 7308 1003
rect 3853 977 4140 983
rect 4340 977 4652 983
rect 4804 977 5244 983
rect 5620 977 5948 983
rect 6164 977 6604 983
rect 6708 977 7196 983
rect 2580 957 2691 963
rect 2708 957 2748 963
rect 2772 957 3004 963
rect 3012 957 3340 963
rect 3572 957 3580 963
rect 3604 957 3644 963
rect 3652 957 3708 963
rect 3716 957 3740 963
rect 3764 957 4316 963
rect 4372 957 4403 963
rect 2093 937 2764 943
rect 2788 937 2812 943
rect 2820 937 2844 943
rect 2884 937 3052 943
rect 3076 937 3164 943
rect 3213 937 3276 943
rect 1853 917 2012 923
rect 2036 917 2076 923
rect 2084 917 2188 923
rect 2356 917 2412 923
rect 2420 917 2556 923
rect 2596 917 2636 923
rect 2676 917 2716 923
rect 2868 917 2908 923
rect 2964 917 3116 923
rect 3213 923 3219 937
rect 3341 943 3347 956
rect 3341 937 3612 943
rect 3620 937 3628 943
rect 3636 937 3996 943
rect 4036 937 4108 943
rect 4116 937 4156 943
rect 4164 937 4172 943
rect 4180 937 4252 943
rect 4308 937 4332 943
rect 4397 943 4403 957
rect 4420 957 4428 963
rect 4788 957 4835 963
rect 4397 937 4444 943
rect 4468 937 4508 943
rect 4708 937 4780 943
rect 4829 943 4835 957
rect 4852 957 4860 963
rect 4868 957 5116 963
rect 5892 957 6092 963
rect 6388 957 6444 963
rect 6740 957 7004 963
rect 7300 957 7356 963
rect 7364 957 7484 963
rect 4829 937 5084 943
rect 5156 937 5436 943
rect 5844 937 5900 943
rect 5908 937 5964 943
rect 6036 937 6156 943
rect 6164 937 6316 943
rect 6324 937 6364 943
rect 6372 937 6396 943
rect 6676 937 6860 943
rect 6868 937 6908 943
rect 6916 937 6940 943
rect 6996 937 7068 943
rect 7076 937 7180 943
rect 7204 937 7244 943
rect 7348 937 7532 943
rect 3156 917 3219 923
rect 3236 917 3596 923
rect 3700 917 3971 923
rect -35 897 396 903
rect 1188 897 1196 903
rect 1204 897 1212 903
rect 1332 897 1372 903
rect 1380 897 1580 903
rect 1588 897 1724 903
rect 1940 897 1964 903
rect 2068 897 2364 903
rect 2372 897 2572 903
rect 2948 897 3004 903
rect 3060 897 3244 903
rect 3268 897 3500 903
rect 3524 897 3692 903
rect 3732 897 3852 903
rect 3892 897 3948 903
rect 3965 903 3971 917
rect 4100 917 4851 923
rect 3965 897 4108 903
rect 4148 897 4620 903
rect 4692 897 4700 903
rect 4845 903 4851 917
rect 4868 917 4940 923
rect 5124 917 5180 923
rect 5476 917 5628 923
rect 5636 917 5772 923
rect 5812 917 5948 923
rect 6020 917 6108 923
rect 6548 917 6588 923
rect 6660 917 6828 923
rect 6996 917 7036 923
rect 7268 917 7340 923
rect 7348 917 7420 923
rect 7428 917 7532 923
rect 4845 897 5436 903
rect 5620 897 5724 903
rect 5940 897 6060 903
rect 6516 897 6556 903
rect 6564 897 6732 903
rect 6964 897 7052 903
rect 7060 897 7132 903
rect 196 877 268 883
rect 276 877 348 883
rect 356 877 540 883
rect 1236 877 1468 883
rect 1492 877 1516 883
rect 1540 877 1580 883
rect 1604 877 3084 883
rect 3124 877 3180 883
rect 3268 877 3292 883
rect 3364 877 3564 883
rect 3949 883 3955 896
rect 3780 877 3891 883
rect 3949 877 4691 883
rect 3885 864 3891 877
rect 468 857 2588 863
rect 2836 857 3660 863
rect 3748 857 3868 863
rect 3988 857 4060 863
rect 4292 857 4332 863
rect 4404 857 4476 863
rect 4685 863 4691 877
rect 4708 877 4812 883
rect 5828 877 6044 883
rect 6100 877 6140 883
rect 6148 877 6892 883
rect 6900 877 7100 883
rect 7140 877 7276 883
rect 4685 857 5452 863
rect 5764 857 5772 863
rect 6548 857 6972 863
rect 7044 857 7196 863
rect 1508 837 1612 843
rect 1620 837 2860 843
rect 2964 837 2988 843
rect 3236 837 3308 843
rect 3588 837 5340 843
rect 5684 837 5932 843
rect 6964 837 6972 843
rect 244 817 316 823
rect 324 817 412 823
rect 1268 817 1900 823
rect 1940 817 2092 823
rect 2100 817 2828 823
rect 2836 817 3340 823
rect 3556 817 3708 823
rect 3860 817 3948 823
rect 4260 817 4316 823
rect 4324 817 4652 823
rect 4660 817 4732 823
rect 4900 817 6332 823
rect 738 814 798 816
rect 738 806 739 814
rect 748 806 749 814
rect 787 806 788 814
rect 797 806 798 814
rect 738 804 798 806
rect 3746 814 3806 816
rect 3746 806 3747 814
rect 3756 806 3757 814
rect 3795 806 3796 814
rect 3805 806 3806 814
rect 3746 804 3806 806
rect 6754 814 6814 816
rect 6754 806 6755 814
rect 6764 806 6765 814
rect 6803 806 6804 814
rect 6813 806 6814 814
rect 6754 804 6814 806
rect 404 797 412 803
rect 1556 797 1932 803
rect 2020 797 2268 803
rect 2388 797 2476 803
rect 2500 797 2524 803
rect 2612 797 2892 803
rect 3108 797 3724 803
rect 3972 797 4348 803
rect 4436 797 4668 803
rect 4836 797 4908 803
rect 5348 797 6060 803
rect 6068 797 6700 803
rect 20 777 44 783
rect 52 777 156 783
rect 1124 777 1324 783
rect 1668 777 1820 783
rect 1908 777 2332 783
rect 2372 777 2396 783
rect 2436 777 2595 783
rect 1309 757 1628 763
rect 1309 744 1315 757
rect 2084 757 2508 763
rect 2589 763 2595 777
rect 2644 777 3228 783
rect 3252 777 3372 783
rect 3620 777 4092 783
rect 4404 777 4636 783
rect 4644 777 4764 783
rect 4788 777 4844 783
rect 5012 777 5500 783
rect 6340 777 6556 783
rect 6564 777 6588 783
rect 7412 777 7500 783
rect 7508 777 7548 783
rect 2589 757 3724 763
rect 3748 757 4236 763
rect 4372 757 4492 763
rect 4612 757 5020 763
rect 5236 757 5356 763
rect 868 737 1164 743
rect 1172 737 1308 743
rect 1652 737 2028 743
rect 2068 737 2124 743
rect 2132 737 2204 743
rect 2212 737 2348 743
rect 2500 737 2908 743
rect 2916 737 3404 743
rect 3412 737 3580 743
rect 3588 737 3836 743
rect 3892 737 3948 743
rect 4020 737 4108 743
rect 4116 737 4204 743
rect 4212 737 4444 743
rect 4724 737 4819 743
rect 436 717 684 723
rect 692 717 828 723
rect 1060 717 1276 723
rect 1284 717 1548 723
rect 1844 717 2092 723
rect 2996 717 3020 723
rect 3204 717 3292 723
rect 3332 717 3388 723
rect 3396 717 3420 723
rect 3476 717 3516 723
rect 3684 717 3916 723
rect 4004 717 4220 723
rect 4372 717 4380 723
rect 4628 717 4796 723
rect 4813 723 4819 737
rect 4868 737 4924 743
rect 5572 737 6220 743
rect 6228 737 6476 743
rect 6884 737 6908 743
rect 7316 737 7388 743
rect 7396 737 7436 743
rect 4813 717 4988 723
rect 5028 717 5100 723
rect 5172 717 5196 723
rect 5316 717 5644 723
rect 5652 717 5660 723
rect 5972 717 6012 723
rect 6356 717 6412 723
rect 6724 717 6924 723
rect 6996 717 7004 723
rect 7220 717 7340 723
rect 148 697 252 703
rect 372 697 412 703
rect 900 697 924 703
rect 1172 697 1740 703
rect 1828 697 1852 703
rect 2052 697 2108 703
rect 2116 697 2204 703
rect 2212 697 2332 703
rect 2404 697 2444 703
rect 2468 697 2508 703
rect 2580 697 2604 703
rect 2756 697 2876 703
rect 2900 697 2940 703
rect 2957 697 3020 703
rect 228 677 348 683
rect 356 677 396 683
rect 1300 677 1340 683
rect 1396 677 1516 683
rect 1588 677 1692 683
rect 1924 677 1948 683
rect 1956 677 2572 683
rect 2957 683 2963 697
rect 3060 697 3100 703
rect 3124 697 3228 703
rect 3245 697 3404 703
rect 2948 677 2963 683
rect 3028 677 3084 683
rect 3245 683 3251 697
rect 3412 697 3564 703
rect 3572 697 4060 703
rect 4276 697 4316 703
rect 4420 697 4604 703
rect 4644 697 4716 703
rect 4724 697 4828 703
rect 5332 697 5452 703
rect 5940 697 6028 703
rect 6164 697 6188 703
rect 6228 697 6236 703
rect 6324 697 6364 703
rect 6420 697 6444 703
rect 6580 697 6604 703
rect 6644 697 6748 703
rect 6756 697 6828 703
rect 6836 697 6956 703
rect 7396 697 7436 703
rect 3092 677 3251 683
rect 3300 677 3372 683
rect 3476 677 3564 683
rect 3876 677 3932 683
rect 3972 677 4028 683
rect 4637 683 4643 696
rect 4292 677 4643 683
rect 4660 677 4956 683
rect 4964 677 5036 683
rect 5108 677 5164 683
rect 5396 677 5436 683
rect 5444 677 5484 683
rect 5492 677 5532 683
rect 5556 677 5788 683
rect 6100 677 6172 683
rect 6180 677 6284 683
rect 6468 677 6572 683
rect 6628 677 6700 683
rect 6964 677 7020 683
rect 7060 677 7164 683
rect 7284 677 7356 683
rect 7364 677 7420 683
rect 260 657 316 663
rect 676 657 1164 663
rect 1412 657 1516 663
rect 1524 657 1660 663
rect 1716 657 1996 663
rect 2020 657 2220 663
rect 2228 657 2620 663
rect 2868 657 3004 663
rect 3012 657 3036 663
rect 3044 657 3260 663
rect 3268 657 3340 663
rect 3428 657 3612 663
rect 3684 657 3708 663
rect 3716 657 3964 663
rect 4068 657 4364 663
rect 4372 657 4396 663
rect 4404 657 4476 663
rect 4484 657 4812 663
rect 4820 657 4844 663
rect 4852 657 4924 663
rect 5220 657 5699 663
rect 212 637 268 643
rect 308 637 476 643
rect 516 637 732 643
rect 1156 637 2396 643
rect 2468 637 2572 643
rect 3076 637 3132 643
rect 3140 637 3164 643
rect 3220 637 3388 643
rect 3812 637 3916 643
rect 4340 637 4380 643
rect 4692 637 4732 643
rect 4772 637 5004 643
rect 5012 637 5116 643
rect 5124 637 5676 643
rect 5693 643 5699 657
rect 5780 657 5788 663
rect 5860 657 5996 663
rect 6132 657 6220 663
rect 6228 657 6348 663
rect 6356 657 6396 663
rect 6548 657 6620 663
rect 6932 657 7116 663
rect 5693 637 5708 643
rect 5732 637 5772 643
rect 5860 637 5900 643
rect 5908 637 5980 643
rect 5988 637 6332 643
rect 7332 637 7452 643
rect 740 617 940 623
rect 948 617 1244 623
rect 1684 617 1820 623
rect 1860 617 1900 623
rect 1924 617 2012 623
rect 2148 617 2188 623
rect 2324 617 2524 623
rect 2532 617 2556 623
rect 2884 617 3084 623
rect 3108 617 3292 623
rect 3316 617 3852 623
rect 3885 617 4124 623
rect 2242 614 2302 616
rect 2242 606 2243 614
rect 2252 606 2253 614
rect 2291 606 2292 614
rect 2301 606 2302 614
rect 2242 604 2302 606
rect 84 597 236 603
rect 292 597 332 603
rect 388 597 460 603
rect 916 597 1116 603
rect 1364 597 1676 603
rect 1892 597 2220 603
rect 3076 597 3148 603
rect 3885 603 3891 617
rect 4196 617 4492 623
rect 4900 617 5036 623
rect 5060 617 5164 623
rect 5652 617 5868 623
rect 5876 617 5900 623
rect 5972 617 6300 623
rect 6308 617 7228 623
rect 5250 614 5310 616
rect 5250 606 5251 614
rect 5260 606 5261 614
rect 5299 606 5300 614
rect 5309 606 5310 614
rect 5250 604 5310 606
rect 3412 597 3891 603
rect 3908 597 4044 603
rect 4228 597 5212 603
rect 6100 597 6268 603
rect 6276 597 6620 603
rect 6660 597 6940 603
rect 196 577 300 583
rect 404 577 588 583
rect 596 577 652 583
rect 916 577 1212 583
rect 1396 577 1500 583
rect 1508 577 1596 583
rect 1828 577 2188 583
rect 3188 577 3196 583
rect 3204 577 3244 583
rect 3284 577 3484 583
rect 3492 577 3539 583
rect 708 557 764 563
rect 772 557 892 563
rect 900 557 956 563
rect 964 557 1196 563
rect 1444 557 1532 563
rect 1652 557 1692 563
rect 1780 557 1868 563
rect 2004 557 2076 563
rect 2180 557 2364 563
rect 2372 557 2460 563
rect 2564 557 2572 563
rect 2580 557 2700 563
rect 2708 557 2828 563
rect 3060 557 3116 563
rect 3156 557 3292 563
rect 3533 563 3539 577
rect 4221 583 4227 596
rect 3556 577 4227 583
rect 4237 577 4684 583
rect 3533 557 3708 563
rect 3732 557 3820 563
rect 4237 563 4243 577
rect 5236 577 5308 583
rect 5325 577 5564 583
rect 3956 557 4243 563
rect 4676 557 5068 563
rect 5076 557 5116 563
rect 5325 563 5331 577
rect 6036 577 6124 583
rect 6420 577 6476 583
rect 6708 577 6988 583
rect 7380 577 7500 583
rect 5156 557 5331 563
rect 5428 557 5596 563
rect 6189 557 6316 563
rect 6189 544 6195 557
rect 6388 557 6460 563
rect 6468 557 6556 563
rect 6580 557 6636 563
rect 6708 557 6812 563
rect 6884 557 7068 563
rect 7300 557 7356 563
rect 7364 557 7420 563
rect 7428 557 7484 563
rect 132 537 220 543
rect 228 537 460 543
rect 820 537 860 543
rect 868 537 924 543
rect 1204 537 1404 543
rect 1524 537 1564 543
rect 1572 537 1612 543
rect 1652 537 1676 543
rect 1684 537 1708 543
rect 1844 537 1980 543
rect 1988 537 1996 543
rect 2004 537 2188 543
rect 2308 537 2691 543
rect 532 517 588 523
rect 596 517 620 523
rect 628 517 1052 523
rect 1060 517 1068 523
rect 1284 517 1404 523
rect 1428 517 1644 523
rect 1716 517 1788 523
rect 1796 517 1820 523
rect 2084 517 2156 523
rect 2372 517 2476 523
rect 2685 523 2691 537
rect 2708 537 2764 543
rect 2996 537 3228 543
rect 3236 537 3532 543
rect 3540 537 3756 543
rect 3764 537 3900 543
rect 3908 537 4364 543
rect 4372 537 4396 543
rect 4404 537 4684 543
rect 4692 537 4732 543
rect 4740 537 4972 543
rect 4996 537 5020 543
rect 5028 537 5148 543
rect 5172 537 5324 543
rect 5524 537 5612 543
rect 5748 537 5868 543
rect 5988 537 6076 543
rect 6084 537 6108 543
rect 6116 537 6188 543
rect 6276 537 6412 543
rect 6532 537 6668 543
rect 6948 537 7052 543
rect 7108 537 7212 543
rect 2685 517 2716 523
rect 2900 517 3276 523
rect 3364 517 3484 523
rect 3716 517 3852 523
rect 3860 517 4252 523
rect 4260 517 4316 523
rect 4324 517 4348 523
rect 4356 517 4684 523
rect 4692 517 4940 523
rect 4948 517 5084 523
rect 5188 517 5363 523
rect 436 497 588 503
rect 692 497 796 503
rect 964 497 1020 503
rect 1037 497 1628 503
rect 372 477 716 483
rect 1037 483 1043 497
rect 2020 497 2316 503
rect 3044 497 3068 503
rect 3188 497 3436 503
rect 3444 497 3548 503
rect 3604 497 3980 503
rect 4084 497 4204 503
rect 4484 497 4540 503
rect 4820 497 4876 503
rect 5204 497 5340 503
rect 5357 503 5363 517
rect 5508 517 5532 523
rect 5620 517 5660 523
rect 6180 517 6204 523
rect 6228 517 6396 523
rect 6420 517 6636 523
rect 6676 517 6780 523
rect 6900 517 7164 523
rect 7252 517 7324 523
rect 5357 497 5404 503
rect 5476 497 5500 503
rect 5588 497 5628 503
rect 5652 497 5740 503
rect 6052 497 6156 503
rect 6164 497 6364 503
rect 6893 503 6899 516
rect 6372 497 6899 503
rect 7188 497 7228 503
rect 7236 497 7292 503
rect 836 477 1043 483
rect 1540 477 1836 483
rect 2804 477 3212 483
rect 3284 477 3436 483
rect 3476 477 3532 483
rect 3540 477 3628 483
rect 3636 477 4108 483
rect 4116 477 4172 483
rect 4436 477 4492 483
rect 4900 477 5052 483
rect 5428 477 5548 483
rect 5556 477 5612 483
rect 6148 477 6252 483
rect 660 457 1347 463
rect 1341 443 1347 457
rect 1396 457 1804 463
rect 1892 457 2652 463
rect 3380 457 4092 463
rect 4100 457 4300 463
rect 4308 457 4476 463
rect 4948 457 5388 463
rect 5428 457 5804 463
rect 6116 457 6140 463
rect 1341 437 1932 443
rect 1972 437 2188 443
rect 2228 437 3404 443
rect 3508 437 3612 443
rect 3620 437 3708 443
rect 3764 437 3916 443
rect 4036 437 4108 443
rect 4132 437 4268 443
rect 4340 437 4940 443
rect 5108 437 5468 443
rect 5716 437 6924 443
rect 6932 437 7132 443
rect 7140 437 7372 443
rect 452 417 556 423
rect 1140 417 1324 423
rect 1332 417 1884 423
rect 2052 417 2156 423
rect 2180 417 2380 423
rect 2740 417 2908 423
rect 4084 417 4300 423
rect 4852 417 4876 423
rect 4884 417 5308 423
rect 5316 417 5644 423
rect 738 414 798 416
rect 738 406 739 414
rect 748 406 749 414
rect 787 406 788 414
rect 797 406 798 414
rect 738 404 798 406
rect 3746 414 3806 416
rect 3746 406 3747 414
rect 3756 406 3757 414
rect 3795 406 3796 414
rect 3805 406 3806 414
rect 3746 404 3806 406
rect 6754 414 6814 416
rect 6754 406 6755 414
rect 6764 406 6765 414
rect 6803 406 6804 414
rect 6813 406 6814 414
rect 6754 404 6814 406
rect 1172 397 1196 403
rect 1476 397 1516 403
rect 1604 397 1644 403
rect 1652 397 2140 403
rect 2196 397 2204 403
rect 2212 397 2396 403
rect 2404 397 2876 403
rect 2884 397 3244 403
rect 4932 397 5164 403
rect 5524 397 5708 403
rect 468 377 1036 383
rect 1044 377 1964 383
rect 2084 377 2492 383
rect 3172 377 3340 383
rect 3348 377 3884 383
rect 4420 377 4572 383
rect 4580 377 4620 383
rect 4628 377 4668 383
rect 4676 377 5948 383
rect 116 357 188 363
rect 196 357 1708 363
rect 1748 357 1964 363
rect 1972 357 2739 363
rect 2733 344 2739 357
rect 3124 357 3324 363
rect 3876 357 3932 363
rect 3940 357 4172 363
rect 4180 357 4332 363
rect 4804 357 4812 363
rect 4916 357 5100 363
rect 5140 357 5196 363
rect 5684 357 5692 363
rect 6260 357 6396 363
rect 6404 357 6668 363
rect 1012 337 1084 343
rect 1092 337 1484 343
rect 1492 337 1612 343
rect 1620 337 1724 343
rect 2036 337 2147 343
rect 2141 324 2147 337
rect 2468 337 2620 343
rect 2628 337 2700 343
rect 2740 337 2764 343
rect 2772 337 3052 343
rect 3076 337 3116 343
rect 3220 337 3852 343
rect 3892 337 3996 343
rect 4516 337 4636 343
rect 4708 337 5020 343
rect 5060 337 5260 343
rect 5268 337 5420 343
rect 6452 337 6556 343
rect 7476 337 7564 343
rect 196 317 588 323
rect 596 317 620 323
rect 676 317 716 323
rect 724 317 908 323
rect 964 317 1740 323
rect 1812 317 1868 323
rect 1876 317 2076 323
rect 2148 317 2300 323
rect 2372 317 2428 323
rect 2660 317 2707 323
rect 2701 304 2707 317
rect 2820 317 2828 323
rect 2996 317 3116 323
rect 3124 317 3139 323
rect 564 297 636 303
rect 644 297 812 303
rect 884 297 1004 303
rect 1172 297 1196 303
rect 1572 297 1708 303
rect 1780 297 1948 303
rect 2068 297 2108 303
rect 2164 297 2508 303
rect 2516 297 2604 303
rect 2612 297 2684 303
rect 2708 297 2780 303
rect 2964 297 3116 303
rect 3133 303 3139 317
rect 3908 317 3980 323
rect 3988 317 4428 323
rect 4484 317 4652 323
rect 4660 317 4732 323
rect 4756 317 4796 323
rect 4804 317 5004 323
rect 5012 317 5356 323
rect 5412 317 5468 323
rect 5620 317 5692 323
rect 5876 317 5916 323
rect 5972 317 6028 323
rect 6356 317 6412 323
rect 6484 317 6524 323
rect 6724 317 6876 323
rect 6884 317 6940 323
rect 7156 317 7228 323
rect 7236 317 7292 323
rect 7380 317 7484 323
rect 3133 297 3388 303
rect 3396 297 3532 303
rect 3556 297 3660 303
rect 3860 297 3900 303
rect 3924 297 3932 303
rect 3972 297 4092 303
rect 4404 297 4492 303
rect 4500 297 4540 303
rect 4644 297 4700 303
rect 4756 297 4828 303
rect 4916 297 5340 303
rect 5396 297 5500 303
rect 5652 297 5756 303
rect 5764 297 5836 303
rect 5917 303 5923 316
rect 5917 297 5980 303
rect 5988 297 6060 303
rect 6292 297 6508 303
rect 6548 297 6636 303
rect 6644 297 7212 303
rect 7268 297 7308 303
rect 7364 297 7404 303
rect 7412 297 7516 303
rect 276 277 540 283
rect 548 277 668 283
rect 676 277 684 283
rect 692 277 700 283
rect 932 277 1020 283
rect 1268 277 1580 283
rect 1652 277 1804 283
rect 1860 277 1932 283
rect 2196 277 2236 283
rect 2244 277 2444 283
rect 2452 277 2860 283
rect 2980 277 3068 283
rect 3124 277 3164 283
rect 3268 277 3356 283
rect 3396 277 3468 283
rect 3508 277 3548 283
rect 3556 277 3724 283
rect 3844 277 4140 283
rect 4148 277 4220 283
rect 4260 277 4380 283
rect 4820 277 4924 283
rect 4932 277 5068 283
rect 5156 277 5187 283
rect 596 257 684 263
rect 820 257 892 263
rect 1172 257 1548 263
rect 2420 257 2524 263
rect 2548 257 2572 263
rect 2596 257 2636 263
rect 2692 257 2732 263
rect 2740 257 2828 263
rect 2948 257 2988 263
rect 3060 257 3180 263
rect 3364 257 3580 263
rect 3588 257 3644 263
rect 3732 257 3884 263
rect 4388 257 4540 263
rect 4564 257 4700 263
rect 4708 257 4924 263
rect 4980 257 5116 263
rect 5140 257 5164 263
rect 5181 263 5187 277
rect 5220 277 5244 283
rect 5268 277 5292 283
rect 5348 277 5484 283
rect 5492 277 5548 283
rect 5684 277 5724 283
rect 5748 277 5788 283
rect 5828 277 5916 283
rect 5940 277 5964 283
rect 6020 277 6076 283
rect 6180 277 6220 283
rect 6228 277 6268 283
rect 6516 277 6684 283
rect 6852 277 6988 283
rect 7156 277 7436 283
rect 7492 277 7532 283
rect 5181 257 5596 263
rect 5892 257 6124 263
rect 6132 257 6204 263
rect 6212 257 6252 263
rect 6644 257 6828 263
rect 6868 257 6924 263
rect 6932 257 6972 263
rect 7012 257 7340 263
rect 7428 257 7532 263
rect 228 237 380 243
rect 868 237 972 243
rect 1156 237 1164 243
rect 1236 237 1516 243
rect 1652 237 2364 243
rect 2372 237 2460 243
rect 2468 237 2588 243
rect 3620 237 3692 243
rect 4132 237 4188 243
rect 4196 237 4444 243
rect 4596 237 4668 243
rect 4676 237 5004 243
rect 5012 237 5324 243
rect 5444 237 5484 243
rect 5604 237 5644 243
rect 5652 237 6028 243
rect 6484 237 6588 243
rect 6596 237 6620 243
rect 6628 237 6668 243
rect 6676 237 6716 243
rect 6916 237 6940 243
rect 7204 237 7388 243
rect 148 217 252 223
rect 996 217 1196 223
rect 1284 217 1436 223
rect 2884 217 3036 223
rect 3044 217 3372 223
rect 4276 217 4460 223
rect 4500 217 5084 223
rect 5188 217 5212 223
rect 5364 217 5404 223
rect 5412 217 6236 223
rect 6756 217 7020 223
rect 2242 214 2302 216
rect 2242 206 2243 214
rect 2252 206 2253 214
rect 2291 206 2292 214
rect 2301 206 2302 214
rect 2242 204 2302 206
rect 5250 214 5310 216
rect 5250 206 5251 214
rect 5260 206 5261 214
rect 5299 206 5300 214
rect 5309 206 5310 214
rect 5250 204 5310 206
rect 1220 197 1484 203
rect 1636 197 2044 203
rect 2628 197 2812 203
rect 2836 197 2956 203
rect 2964 197 3228 203
rect 3236 197 3484 203
rect 4196 197 4236 203
rect 5108 197 5196 203
rect 5332 197 5420 203
rect 5428 197 5852 203
rect 6900 197 6972 203
rect 6980 197 7148 203
rect 68 177 124 183
rect 132 177 556 183
rect 1476 177 1516 183
rect 1892 177 2140 183
rect 2148 177 2428 183
rect 2468 177 2508 183
rect 2564 177 2732 183
rect 2756 177 2892 183
rect 2932 177 3420 183
rect 3428 177 3676 183
rect 4740 177 5068 183
rect 5076 177 5228 183
rect 5364 177 5660 183
rect 5700 177 5756 183
rect 1140 157 1196 163
rect 1396 157 1468 163
rect 1540 157 1596 163
rect 1604 157 1660 163
rect 2068 157 2172 163
rect 2180 157 2300 163
rect 2404 157 2796 163
rect 2804 157 2860 163
rect 3108 157 3132 163
rect 3956 157 4044 163
rect 4180 157 4364 163
rect 4388 157 4396 163
rect 4452 157 4668 163
rect 4996 157 5100 163
rect 5204 157 5484 163
rect 5796 157 5884 163
rect 6932 157 7004 163
rect 7044 157 7052 163
rect 7060 157 7148 163
rect 7156 157 7212 163
rect 7220 157 7244 163
rect 7316 157 7388 163
rect 36 137 156 143
rect 164 137 236 143
rect 308 137 492 143
rect 500 137 796 143
rect 804 137 988 143
rect 1012 137 1052 143
rect 1060 137 1100 143
rect 1108 137 1180 143
rect 1188 137 1228 143
rect 1444 137 1772 143
rect 2084 137 2140 143
rect 2148 137 2284 143
rect 2500 137 2627 143
rect 20 117 76 123
rect 356 117 844 123
rect 1476 117 1692 123
rect 1700 117 1852 123
rect 1860 117 2572 123
rect 2621 123 2627 137
rect 2644 137 2668 143
rect 2724 137 2844 143
rect 2852 137 2892 143
rect 3172 137 3260 143
rect 3396 137 3420 143
rect 4004 137 4060 143
rect 4356 137 4364 143
rect 4484 137 4524 143
rect 4548 137 4668 143
rect 4676 137 4732 143
rect 4804 137 5011 143
rect 2621 117 2652 123
rect 2692 117 3324 123
rect 3332 117 4076 123
rect 4292 117 4364 123
rect 4372 117 4780 123
rect 4820 117 4828 123
rect 4852 117 4876 123
rect 5005 123 5011 137
rect 5060 137 5084 143
rect 5396 137 5804 143
rect 6164 137 6220 143
rect 6228 137 6268 143
rect 6324 137 6380 143
rect 6580 137 6636 143
rect 6692 137 6844 143
rect 6964 137 7052 143
rect 7108 137 7276 143
rect 7476 137 7516 143
rect 5005 117 5628 123
rect 5940 117 5980 123
rect 6052 117 6140 123
rect 6173 117 6204 123
rect 84 97 188 103
rect 772 97 1068 103
rect 1076 97 1276 103
rect 1508 97 2140 103
rect 2148 97 2220 103
rect 2340 97 2700 103
rect 2708 97 2732 103
rect 4077 103 4083 116
rect 4077 97 4796 103
rect 4820 97 4860 103
rect 5140 97 5196 103
rect 5220 97 5516 103
rect 6173 103 6179 117
rect 6292 117 6316 123
rect 7012 117 7116 123
rect 7348 117 7468 123
rect 5972 97 6179 103
rect 6196 97 6332 103
rect 6676 97 6700 103
rect 7284 97 7308 103
rect 1044 77 1372 83
rect 1700 77 1756 83
rect 1972 77 2092 83
rect 2260 77 2316 83
rect 4356 77 4412 83
rect 4468 77 4492 83
rect 4516 77 4572 83
rect 4596 77 4684 83
rect 4692 77 5052 83
rect 5060 77 5420 83
rect 260 57 1228 63
rect 4436 57 4476 63
rect 852 37 940 43
rect 1172 37 1196 43
rect 1268 37 1340 43
rect 692 17 716 23
rect 836 17 860 23
rect 996 17 1404 23
rect 1572 17 1596 23
rect 738 14 798 16
rect 738 6 739 14
rect 748 6 749 14
rect 787 6 788 14
rect 797 6 798 14
rect 738 4 798 6
rect 3746 14 3806 16
rect 3746 6 3747 14
rect 3756 6 3757 14
rect 3795 6 3796 14
rect 3805 6 3806 14
rect 3746 4 3806 6
rect 6754 14 6814 16
rect 6754 6 6755 14
rect 6764 6 6765 14
rect 6803 6 6804 14
rect 6813 6 6814 14
rect 6754 4 6814 6
<< m4contact >>
rect 4748 5216 4756 5224
rect 740 5206 747 5214
rect 747 5206 748 5214
rect 752 5206 757 5214
rect 757 5206 759 5214
rect 759 5206 760 5214
rect 764 5206 767 5214
rect 767 5206 769 5214
rect 769 5206 772 5214
rect 776 5206 777 5214
rect 777 5206 779 5214
rect 779 5206 784 5214
rect 788 5206 789 5214
rect 789 5206 796 5214
rect 3748 5206 3755 5214
rect 3755 5206 3756 5214
rect 3760 5206 3765 5214
rect 3765 5206 3767 5214
rect 3767 5206 3768 5214
rect 3772 5206 3775 5214
rect 3775 5206 3777 5214
rect 3777 5206 3780 5214
rect 3784 5206 3785 5214
rect 3785 5206 3787 5214
rect 3787 5206 3792 5214
rect 3796 5206 3797 5214
rect 3797 5206 3804 5214
rect 6756 5206 6763 5214
rect 6763 5206 6764 5214
rect 6768 5206 6773 5214
rect 6773 5206 6775 5214
rect 6775 5206 6776 5214
rect 6780 5206 6783 5214
rect 6783 5206 6785 5214
rect 6785 5206 6788 5214
rect 6792 5206 6793 5214
rect 6793 5206 6795 5214
rect 6795 5206 6800 5214
rect 6804 5206 6805 5214
rect 6805 5206 6812 5214
rect 4684 5136 4692 5144
rect 1260 5096 1268 5104
rect 3980 5096 3988 5104
rect 5004 5076 5012 5084
rect 1676 5056 1684 5064
rect 4716 5056 4724 5064
rect 5196 5056 5204 5064
rect 7340 5056 7348 5064
rect 7532 5056 7540 5064
rect 6860 5036 6868 5044
rect 1260 5016 1268 5024
rect 6284 5016 6292 5024
rect 2244 5006 2251 5014
rect 2251 5006 2252 5014
rect 2256 5006 2261 5014
rect 2261 5006 2263 5014
rect 2263 5006 2264 5014
rect 2268 5006 2271 5014
rect 2271 5006 2273 5014
rect 2273 5006 2276 5014
rect 2280 5006 2281 5014
rect 2281 5006 2283 5014
rect 2283 5006 2288 5014
rect 2292 5006 2293 5014
rect 2293 5006 2300 5014
rect 5252 5006 5259 5014
rect 5259 5006 5260 5014
rect 5264 5006 5269 5014
rect 5269 5006 5271 5014
rect 5271 5006 5272 5014
rect 5276 5006 5279 5014
rect 5279 5006 5281 5014
rect 5281 5006 5284 5014
rect 5288 5006 5289 5014
rect 5289 5006 5291 5014
rect 5291 5006 5296 5014
rect 5300 5006 5301 5014
rect 5301 5006 5308 5014
rect 7308 4996 7316 5004
rect 2924 4976 2932 4984
rect 7564 4956 7572 4964
rect 5740 4936 5748 4944
rect 5836 4936 5844 4944
rect 2348 4916 2356 4924
rect 7468 4916 7476 4924
rect 5612 4896 5620 4904
rect 1932 4876 1940 4884
rect 2348 4876 2356 4884
rect 3980 4876 3988 4884
rect 4908 4856 4916 4864
rect 6668 4836 6676 4844
rect 5516 4816 5524 4824
rect 5804 4816 5812 4824
rect 6316 4816 6324 4824
rect 740 4806 747 4814
rect 747 4806 748 4814
rect 752 4806 757 4814
rect 757 4806 759 4814
rect 759 4806 760 4814
rect 764 4806 767 4814
rect 767 4806 769 4814
rect 769 4806 772 4814
rect 776 4806 777 4814
rect 777 4806 779 4814
rect 779 4806 784 4814
rect 788 4806 789 4814
rect 789 4806 796 4814
rect 3748 4806 3755 4814
rect 3755 4806 3756 4814
rect 3760 4806 3765 4814
rect 3765 4806 3767 4814
rect 3767 4806 3768 4814
rect 3772 4806 3775 4814
rect 3775 4806 3777 4814
rect 3777 4806 3780 4814
rect 3784 4806 3785 4814
rect 3785 4806 3787 4814
rect 3787 4806 3792 4814
rect 3796 4806 3797 4814
rect 3797 4806 3804 4814
rect 6756 4806 6763 4814
rect 6763 4806 6764 4814
rect 6768 4806 6773 4814
rect 6773 4806 6775 4814
rect 6775 4806 6776 4814
rect 6780 4806 6783 4814
rect 6783 4806 6785 4814
rect 6785 4806 6788 4814
rect 6792 4806 6793 4814
rect 6793 4806 6795 4814
rect 6795 4806 6800 4814
rect 6804 4806 6805 4814
rect 6805 4806 6812 4814
rect 1004 4796 1012 4804
rect 1580 4796 1588 4804
rect 3628 4796 3636 4804
rect 5676 4796 5684 4804
rect 6956 4796 6964 4804
rect 1548 4756 1556 4764
rect 4364 4776 4372 4784
rect 3948 4756 3956 4764
rect 4748 4756 4756 4764
rect 7180 4756 7188 4764
rect 7276 4756 7284 4764
rect 4588 4736 4596 4744
rect 4108 4716 4116 4724
rect 4748 4716 4756 4724
rect 1164 4696 1172 4704
rect 2060 4696 2068 4704
rect 3404 4696 3412 4704
rect 4204 4696 4212 4704
rect 4780 4696 4788 4704
rect 5164 4696 5172 4704
rect 7404 4716 7412 4724
rect 7436 4716 7444 4724
rect 1644 4676 1652 4684
rect 3116 4676 3124 4684
rect 5004 4676 5012 4684
rect 6284 4676 6292 4684
rect 940 4656 948 4664
rect 7500 4656 7508 4664
rect 332 4636 340 4644
rect 556 4636 564 4644
rect 908 4636 916 4644
rect 1612 4636 1620 4644
rect 5196 4636 5204 4644
rect 1548 4616 1556 4624
rect 4716 4616 4724 4624
rect 2244 4606 2251 4614
rect 2251 4606 2252 4614
rect 2256 4606 2261 4614
rect 2261 4606 2263 4614
rect 2263 4606 2264 4614
rect 2268 4606 2271 4614
rect 2271 4606 2273 4614
rect 2273 4606 2276 4614
rect 2280 4606 2281 4614
rect 2281 4606 2283 4614
rect 2283 4606 2288 4614
rect 2292 4606 2293 4614
rect 2293 4606 2300 4614
rect 5252 4606 5259 4614
rect 5259 4606 5260 4614
rect 5264 4606 5269 4614
rect 5269 4606 5271 4614
rect 5271 4606 5272 4614
rect 5276 4606 5279 4614
rect 5279 4606 5281 4614
rect 5281 4606 5284 4614
rect 5288 4606 5289 4614
rect 5289 4606 5291 4614
rect 5291 4606 5296 4614
rect 5300 4606 5301 4614
rect 5301 4606 5308 4614
rect 556 4596 564 4604
rect 1004 4596 1012 4604
rect 7212 4596 7220 4604
rect 7308 4596 7316 4604
rect 236 4576 244 4584
rect 2572 4576 2580 4584
rect 6060 4576 6068 4584
rect 7180 4576 7188 4584
rect 1804 4556 1812 4564
rect 2508 4556 2516 4564
rect 5004 4556 5012 4564
rect 1196 4536 1204 4544
rect 1932 4536 1940 4544
rect 3084 4536 3092 4544
rect 6156 4536 6164 4544
rect 6700 4536 6708 4544
rect 268 4516 276 4524
rect 1132 4516 1140 4524
rect 1612 4516 1620 4524
rect 1644 4516 1652 4524
rect 1804 4516 1812 4524
rect 4588 4516 4596 4524
rect 6060 4516 6068 4524
rect 6092 4516 6100 4524
rect 2540 4496 2548 4504
rect 4780 4496 4788 4504
rect 2188 4476 2196 4484
rect 6092 4476 6100 4484
rect 3116 4436 3124 4444
rect 2508 4416 2516 4424
rect 2604 4416 2612 4424
rect 4428 4416 4436 4424
rect 5132 4416 5140 4424
rect 740 4406 747 4414
rect 747 4406 748 4414
rect 752 4406 757 4414
rect 757 4406 759 4414
rect 759 4406 760 4414
rect 764 4406 767 4414
rect 767 4406 769 4414
rect 769 4406 772 4414
rect 776 4406 777 4414
rect 777 4406 779 4414
rect 779 4406 784 4414
rect 788 4406 789 4414
rect 789 4406 796 4414
rect 3748 4406 3755 4414
rect 3755 4406 3756 4414
rect 3760 4406 3765 4414
rect 3765 4406 3767 4414
rect 3767 4406 3768 4414
rect 3772 4406 3775 4414
rect 3775 4406 3777 4414
rect 3777 4406 3780 4414
rect 3784 4406 3785 4414
rect 3785 4406 3787 4414
rect 3787 4406 3792 4414
rect 3796 4406 3797 4414
rect 3797 4406 3804 4414
rect 6756 4406 6763 4414
rect 6763 4406 6764 4414
rect 6768 4406 6773 4414
rect 6773 4406 6775 4414
rect 6775 4406 6776 4414
rect 6780 4406 6783 4414
rect 6783 4406 6785 4414
rect 6785 4406 6788 4414
rect 6792 4406 6793 4414
rect 6793 4406 6795 4414
rect 6795 4406 6800 4414
rect 6804 4406 6805 4414
rect 6805 4406 6812 4414
rect 2348 4376 2356 4384
rect 4876 4376 4884 4384
rect 5612 4376 5620 4384
rect 4748 4356 4756 4364
rect 4972 4336 4980 4344
rect 5868 4336 5876 4344
rect 6348 4336 6356 4344
rect 3180 4316 3188 4324
rect 4684 4316 4692 4324
rect 6316 4316 6324 4324
rect 7372 4316 7380 4324
rect 2060 4296 2068 4304
rect 2348 4296 2356 4304
rect 1260 4276 1268 4284
rect 2460 4276 2468 4284
rect 5100 4296 5108 4304
rect 5164 4296 5172 4304
rect 6860 4296 6868 4304
rect 1932 4256 1940 4264
rect 2092 4256 2100 4264
rect 2348 4256 2356 4264
rect 2476 4256 2484 4264
rect 4364 4276 4372 4284
rect 4460 4276 4468 4284
rect 6028 4276 6036 4284
rect 5932 4256 5940 4264
rect 6188 4256 6196 4264
rect 2540 4236 2548 4244
rect 524 4216 532 4224
rect 1164 4216 1172 4224
rect 1292 4216 1300 4224
rect 2244 4206 2251 4214
rect 2251 4206 2252 4214
rect 2256 4206 2261 4214
rect 2261 4206 2263 4214
rect 2263 4206 2264 4214
rect 2268 4206 2271 4214
rect 2271 4206 2273 4214
rect 2273 4206 2276 4214
rect 2280 4206 2281 4214
rect 2281 4206 2283 4214
rect 2283 4206 2288 4214
rect 2292 4206 2293 4214
rect 2293 4206 2300 4214
rect 908 4196 916 4204
rect 6156 4216 6164 4224
rect 5252 4206 5259 4214
rect 5259 4206 5260 4214
rect 5264 4206 5269 4214
rect 5269 4206 5271 4214
rect 5271 4206 5272 4214
rect 5276 4206 5279 4214
rect 5279 4206 5281 4214
rect 5281 4206 5284 4214
rect 5288 4206 5289 4214
rect 5289 4206 5291 4214
rect 5291 4206 5296 4214
rect 5300 4206 5301 4214
rect 5301 4206 5308 4214
rect 6252 4196 6260 4204
rect 1196 4176 1204 4184
rect 3020 4176 3028 4184
rect 3276 4176 3284 4184
rect 5036 4176 5044 4184
rect 6124 4176 6132 4184
rect 6220 4176 6228 4184
rect 6700 4176 6708 4184
rect 3084 4156 3092 4164
rect 4012 4156 4020 4164
rect 7500 4176 7508 4184
rect 7436 4156 7444 4164
rect 332 4116 340 4124
rect 1356 4116 1364 4124
rect 1388 4116 1396 4124
rect 2092 4116 2100 4124
rect 3692 4116 3700 4124
rect 5868 4116 5876 4124
rect 6124 4116 6132 4124
rect 1196 4096 1204 4104
rect 3148 4096 3156 4104
rect 3564 4096 3572 4104
rect 5164 4096 5172 4104
rect 1676 4076 1684 4084
rect 1708 4076 1716 4084
rect 1484 4056 1492 4064
rect 5804 4056 5812 4064
rect 2572 4036 2580 4044
rect 3404 4036 3412 4044
rect 7500 4036 7508 4044
rect 740 4006 747 4014
rect 747 4006 748 4014
rect 752 4006 757 4014
rect 757 4006 759 4014
rect 759 4006 760 4014
rect 764 4006 767 4014
rect 767 4006 769 4014
rect 769 4006 772 4014
rect 776 4006 777 4014
rect 777 4006 779 4014
rect 779 4006 784 4014
rect 788 4006 789 4014
rect 789 4006 796 4014
rect 6028 4016 6036 4024
rect 3748 4006 3755 4014
rect 3755 4006 3756 4014
rect 3760 4006 3765 4014
rect 3765 4006 3767 4014
rect 3767 4006 3768 4014
rect 3772 4006 3775 4014
rect 3775 4006 3777 4014
rect 3777 4006 3780 4014
rect 3784 4006 3785 4014
rect 3785 4006 3787 4014
rect 3787 4006 3792 4014
rect 3796 4006 3797 4014
rect 3797 4006 3804 4014
rect 6756 4006 6763 4014
rect 6763 4006 6764 4014
rect 6768 4006 6773 4014
rect 6773 4006 6775 4014
rect 6775 4006 6776 4014
rect 6780 4006 6783 4014
rect 6783 4006 6785 4014
rect 6785 4006 6788 4014
rect 6792 4006 6793 4014
rect 6793 4006 6795 4014
rect 6795 4006 6800 4014
rect 6804 4006 6805 4014
rect 6805 4006 6812 4014
rect 1324 3976 1332 3984
rect 2348 3976 2356 3984
rect 4972 3976 4980 3984
rect 3852 3956 3860 3964
rect 4492 3956 4500 3964
rect 268 3936 276 3944
rect 6156 3936 6164 3944
rect 7404 3936 7412 3944
rect 7436 3936 7444 3944
rect 364 3916 372 3924
rect 1420 3916 1428 3924
rect 4428 3916 4436 3924
rect 5484 3916 5492 3924
rect 908 3896 916 3904
rect 1292 3896 1300 3904
rect 1356 3896 1364 3904
rect 1804 3896 1812 3904
rect 2508 3896 2516 3904
rect 4460 3896 4468 3904
rect 1484 3876 1492 3884
rect 2924 3876 2932 3884
rect 4876 3876 4884 3884
rect 4908 3876 4916 3884
rect 5004 3896 5012 3904
rect 7404 3896 7412 3904
rect 5100 3876 5108 3884
rect 5932 3876 5940 3884
rect 1644 3856 1652 3864
rect 2188 3856 2196 3864
rect 2764 3856 2772 3864
rect 3916 3856 3924 3864
rect 7308 3876 7316 3884
rect 2540 3836 2548 3844
rect 5612 3836 5620 3844
rect 6380 3836 6388 3844
rect 876 3816 884 3824
rect 3308 3816 3316 3824
rect 2244 3806 2251 3814
rect 2251 3806 2252 3814
rect 2256 3806 2261 3814
rect 2261 3806 2263 3814
rect 2263 3806 2264 3814
rect 2268 3806 2271 3814
rect 2271 3806 2273 3814
rect 2273 3806 2276 3814
rect 2280 3806 2281 3814
rect 2281 3806 2283 3814
rect 2283 3806 2288 3814
rect 2292 3806 2293 3814
rect 2293 3806 2300 3814
rect 5252 3806 5259 3814
rect 5259 3806 5260 3814
rect 5264 3806 5269 3814
rect 5269 3806 5271 3814
rect 5271 3806 5272 3814
rect 5276 3806 5279 3814
rect 5279 3806 5281 3814
rect 5281 3806 5284 3814
rect 5288 3806 5289 3814
rect 5289 3806 5291 3814
rect 5291 3806 5296 3814
rect 5300 3806 5301 3814
rect 5301 3806 5308 3814
rect 1132 3796 1140 3804
rect 3564 3796 3572 3804
rect 364 3776 372 3784
rect 4364 3776 4372 3784
rect 4460 3776 4468 3784
rect 6412 3796 6420 3804
rect 5996 3776 6004 3784
rect 1964 3756 1972 3764
rect 3628 3756 3636 3764
rect 3660 3756 3668 3764
rect 4492 3756 4500 3764
rect 7372 3756 7380 3764
rect 268 3736 276 3744
rect 1132 3736 1140 3744
rect 1484 3736 1492 3744
rect 3276 3736 3284 3744
rect 3180 3716 3188 3724
rect 6668 3716 6676 3724
rect 7372 3716 7380 3724
rect 1644 3696 1652 3704
rect 1836 3696 1844 3704
rect 1932 3696 1940 3704
rect 5420 3696 5428 3704
rect 7404 3696 7412 3704
rect 556 3676 564 3684
rect 940 3676 948 3684
rect 1740 3676 1748 3684
rect 7436 3676 7444 3684
rect 2380 3656 2388 3664
rect 4140 3656 4148 3664
rect 7212 3656 7220 3664
rect 7404 3656 7412 3664
rect 940 3636 948 3644
rect 6572 3636 6580 3644
rect 7436 3636 7444 3644
rect 1260 3616 1268 3624
rect 740 3606 747 3614
rect 747 3606 748 3614
rect 752 3606 757 3614
rect 757 3606 759 3614
rect 759 3606 760 3614
rect 764 3606 767 3614
rect 767 3606 769 3614
rect 769 3606 772 3614
rect 776 3606 777 3614
rect 777 3606 779 3614
rect 779 3606 784 3614
rect 788 3606 789 3614
rect 789 3606 796 3614
rect 1644 3616 1652 3624
rect 4012 3616 4020 3624
rect 6956 3616 6964 3624
rect 7340 3616 7348 3624
rect 3748 3606 3755 3614
rect 3755 3606 3756 3614
rect 3760 3606 3765 3614
rect 3765 3606 3767 3614
rect 3767 3606 3768 3614
rect 3772 3606 3775 3614
rect 3775 3606 3777 3614
rect 3777 3606 3780 3614
rect 3784 3606 3785 3614
rect 3785 3606 3787 3614
rect 3787 3606 3792 3614
rect 3796 3606 3797 3614
rect 3797 3606 3804 3614
rect 6756 3606 6763 3614
rect 6763 3606 6764 3614
rect 6768 3606 6773 3614
rect 6773 3606 6775 3614
rect 6775 3606 6776 3614
rect 6780 3606 6783 3614
rect 6783 3606 6785 3614
rect 6785 3606 6788 3614
rect 6792 3606 6793 3614
rect 6793 3606 6795 3614
rect 6795 3606 6800 3614
rect 6804 3606 6805 3614
rect 6805 3606 6812 3614
rect 3436 3596 3444 3604
rect 1644 3576 1652 3584
rect 4588 3576 4596 3584
rect 7276 3576 7284 3584
rect 1580 3556 1588 3564
rect 4716 3556 4724 3564
rect 5036 3556 5044 3564
rect 7084 3556 7092 3564
rect 2092 3536 2100 3544
rect 5100 3536 5108 3544
rect 5676 3536 5684 3544
rect 5740 3536 5748 3544
rect 6540 3536 6548 3544
rect 172 3516 180 3524
rect 652 3496 660 3504
rect 1388 3516 1396 3524
rect 3084 3516 3092 3524
rect 3948 3516 3956 3524
rect 4364 3516 4372 3524
rect 4428 3516 4436 3524
rect 5132 3516 5140 3524
rect 5484 3516 5492 3524
rect 6860 3516 6868 3524
rect 1356 3496 1364 3504
rect 4620 3496 4628 3504
rect 4812 3496 4820 3504
rect 4940 3496 4948 3504
rect 5452 3496 5460 3504
rect 5516 3496 5524 3504
rect 6444 3496 6452 3504
rect 3180 3476 3188 3484
rect 5548 3476 5556 3484
rect 332 3456 340 3464
rect 2188 3456 2196 3464
rect 5164 3456 5172 3464
rect 5356 3456 5364 3464
rect 1740 3436 1748 3444
rect 2860 3436 2868 3444
rect 6444 3436 6452 3444
rect 1900 3416 1908 3424
rect 7212 3436 7220 3444
rect 2244 3406 2251 3414
rect 2251 3406 2252 3414
rect 2256 3406 2261 3414
rect 2261 3406 2263 3414
rect 2263 3406 2264 3414
rect 2268 3406 2271 3414
rect 2271 3406 2273 3414
rect 2273 3406 2276 3414
rect 2280 3406 2281 3414
rect 2281 3406 2283 3414
rect 2283 3406 2288 3414
rect 2292 3406 2293 3414
rect 2293 3406 2300 3414
rect 5252 3406 5259 3414
rect 5259 3406 5260 3414
rect 5264 3406 5269 3414
rect 5269 3406 5271 3414
rect 5271 3406 5272 3414
rect 5276 3406 5279 3414
rect 5279 3406 5281 3414
rect 5281 3406 5284 3414
rect 5288 3406 5289 3414
rect 5289 3406 5291 3414
rect 5291 3406 5296 3414
rect 5300 3406 5301 3414
rect 5301 3406 5308 3414
rect 524 3396 532 3404
rect 1388 3396 1396 3404
rect 2188 3376 2196 3384
rect 3212 3396 3220 3404
rect 5132 3396 5140 3404
rect 5164 3396 5172 3404
rect 5516 3396 5524 3404
rect 6316 3396 6324 3404
rect 2508 3376 2516 3384
rect 4524 3376 4532 3384
rect 4780 3376 4788 3384
rect 1708 3356 1716 3364
rect 3308 3356 3316 3364
rect 4492 3356 4500 3364
rect 4812 3356 4820 3364
rect 7436 3376 7444 3384
rect 5356 3356 5364 3364
rect 6988 3356 6996 3364
rect 7340 3356 7348 3364
rect 972 3336 980 3344
rect 3884 3336 3892 3344
rect 4716 3336 4724 3344
rect 5132 3336 5140 3344
rect 5612 3336 5620 3344
rect 6252 3336 6260 3344
rect 6380 3336 6388 3344
rect 6540 3336 6548 3344
rect 7180 3336 7188 3344
rect 7404 3336 7412 3344
rect 1420 3316 1428 3324
rect 3404 3316 3412 3324
rect 4428 3316 4436 3324
rect 4620 3316 4628 3324
rect 4748 3316 4756 3324
rect 7276 3316 7284 3324
rect 7500 3316 7508 3324
rect 1452 3296 1460 3304
rect 1900 3296 1908 3304
rect 2604 3296 2612 3304
rect 2860 3296 2868 3304
rect 4940 3296 4948 3304
rect 6348 3296 6356 3304
rect 6700 3296 6708 3304
rect 7244 3296 7252 3304
rect 4492 3276 4500 3284
rect 6060 3276 6068 3284
rect 6540 3276 6548 3284
rect 652 3256 660 3264
rect 1484 3256 1492 3264
rect 2700 3256 2708 3264
rect 3020 3256 3028 3264
rect 3884 3236 3892 3244
rect 5932 3236 5940 3244
rect 4652 3216 4660 3224
rect 6924 3216 6932 3224
rect 740 3206 747 3214
rect 747 3206 748 3214
rect 752 3206 757 3214
rect 757 3206 759 3214
rect 759 3206 760 3214
rect 764 3206 767 3214
rect 767 3206 769 3214
rect 769 3206 772 3214
rect 776 3206 777 3214
rect 777 3206 779 3214
rect 779 3206 784 3214
rect 788 3206 789 3214
rect 789 3206 796 3214
rect 3748 3206 3755 3214
rect 3755 3206 3756 3214
rect 3760 3206 3765 3214
rect 3765 3206 3767 3214
rect 3767 3206 3768 3214
rect 3772 3206 3775 3214
rect 3775 3206 3777 3214
rect 3777 3206 3780 3214
rect 3784 3206 3785 3214
rect 3785 3206 3787 3214
rect 3787 3206 3792 3214
rect 3796 3206 3797 3214
rect 3797 3206 3804 3214
rect 6756 3206 6763 3214
rect 6763 3206 6764 3214
rect 6768 3206 6773 3214
rect 6773 3206 6775 3214
rect 6775 3206 6776 3214
rect 6780 3206 6783 3214
rect 6783 3206 6785 3214
rect 6785 3206 6788 3214
rect 6792 3206 6793 3214
rect 6793 3206 6795 3214
rect 6795 3206 6800 3214
rect 6804 3206 6805 3214
rect 6805 3206 6812 3214
rect 1324 3196 1332 3204
rect 1804 3196 1812 3204
rect 2028 3196 2036 3204
rect 2636 3196 2644 3204
rect 2668 3196 2676 3204
rect 3340 3196 3348 3204
rect 4076 3196 4084 3204
rect 4748 3196 4756 3204
rect 5516 3196 5524 3204
rect 6412 3196 6420 3204
rect 1836 3176 1844 3184
rect 2924 3176 2932 3184
rect 5708 3176 5716 3184
rect 5740 3176 5748 3184
rect 5772 3176 5780 3184
rect 6988 3196 6996 3204
rect 6956 3176 6964 3184
rect 7020 3176 7028 3184
rect 7500 3176 7508 3184
rect 172 3156 180 3164
rect 5036 3156 5044 3164
rect 1388 3116 1396 3124
rect 2892 3136 2900 3144
rect 5100 3136 5108 3144
rect 5420 3136 5428 3144
rect 6316 3136 6324 3144
rect 6476 3136 6484 3144
rect 7084 3136 7092 3144
rect 3500 3116 3508 3124
rect 4524 3116 4532 3124
rect 5484 3116 5492 3124
rect 5644 3116 5652 3124
rect 6220 3116 6228 3124
rect 172 3096 180 3104
rect 204 3096 212 3104
rect 1452 3096 1460 3104
rect 1932 3096 1940 3104
rect 5676 3096 5684 3104
rect 7404 3096 7412 3104
rect 556 3076 564 3084
rect 1356 3076 1364 3084
rect 2796 3076 2804 3084
rect 3148 3076 3156 3084
rect 3372 3076 3380 3084
rect 4012 3076 4020 3084
rect 5068 3076 5076 3084
rect 5132 3076 5140 3084
rect 5996 3076 6004 3084
rect 6220 3076 6228 3084
rect 6316 3076 6324 3084
rect 6604 3076 6612 3084
rect 6924 3076 6932 3084
rect 7468 3076 7476 3084
rect 1068 3056 1076 3064
rect 1676 3056 1684 3064
rect 1964 3056 1972 3064
rect 4460 3056 4468 3064
rect 4524 3056 4532 3064
rect 4972 3056 4980 3064
rect 5612 3056 5620 3064
rect 6892 3056 6900 3064
rect 7180 3056 7188 3064
rect 3628 3036 3636 3044
rect 2244 3006 2251 3014
rect 2251 3006 2252 3014
rect 2256 3006 2261 3014
rect 2261 3006 2263 3014
rect 2263 3006 2264 3014
rect 2268 3006 2271 3014
rect 2271 3006 2273 3014
rect 2273 3006 2276 3014
rect 2280 3006 2281 3014
rect 2281 3006 2283 3014
rect 2283 3006 2288 3014
rect 2292 3006 2293 3014
rect 2293 3006 2300 3014
rect 2060 2996 2068 3004
rect 2092 2996 2100 3004
rect 4748 3036 4756 3044
rect 6700 3036 6708 3044
rect 6476 3016 6484 3024
rect 6636 3016 6644 3024
rect 7116 3016 7124 3024
rect 5252 3006 5259 3014
rect 5259 3006 5260 3014
rect 5264 3006 5269 3014
rect 5269 3006 5271 3014
rect 5271 3006 5272 3014
rect 5276 3006 5279 3014
rect 5279 3006 5281 3014
rect 5281 3006 5284 3014
rect 5288 3006 5289 3014
rect 5289 3006 5291 3014
rect 5291 3006 5296 3014
rect 5300 3006 5301 3014
rect 5301 3006 5308 3014
rect 3340 2976 3348 2984
rect 3628 2976 3636 2984
rect 5900 2976 5908 2984
rect 236 2956 244 2964
rect 588 2956 596 2964
rect 1772 2956 1780 2964
rect 1932 2956 1940 2964
rect 2860 2956 2868 2964
rect 3468 2956 3476 2964
rect 4108 2956 4116 2964
rect 5196 2956 5204 2964
rect 5548 2956 5556 2964
rect 6412 2956 6420 2964
rect 6956 2956 6964 2964
rect 7116 2956 7124 2964
rect 972 2936 980 2944
rect 3660 2936 3668 2944
rect 4428 2936 4436 2944
rect 6188 2936 6196 2944
rect 6572 2936 6580 2944
rect 6604 2936 6612 2944
rect 6860 2936 6868 2944
rect 7372 2936 7380 2944
rect 1356 2916 1364 2924
rect 4620 2916 4628 2924
rect 4748 2916 4756 2924
rect 972 2896 980 2904
rect 3084 2896 3092 2904
rect 4940 2896 4948 2904
rect 5516 2916 5524 2924
rect 5548 2916 5556 2924
rect 5580 2916 5588 2924
rect 5900 2916 5908 2924
rect 6412 2916 6420 2924
rect 7244 2916 7252 2924
rect 5484 2896 5492 2904
rect 6572 2896 6580 2904
rect 6636 2896 6644 2904
rect 1964 2856 1972 2864
rect 3468 2836 3476 2844
rect 3500 2836 3508 2844
rect 844 2816 852 2824
rect 5036 2856 5044 2864
rect 5036 2816 5044 2824
rect 5068 2836 5076 2844
rect 6604 2836 6612 2844
rect 7084 2836 7092 2844
rect 7340 2836 7348 2844
rect 7500 2836 7508 2844
rect 5164 2816 5172 2824
rect 5196 2816 5204 2824
rect 5932 2816 5940 2824
rect 6668 2816 6676 2824
rect 740 2806 747 2814
rect 747 2806 748 2814
rect 752 2806 757 2814
rect 757 2806 759 2814
rect 759 2806 760 2814
rect 764 2806 767 2814
rect 767 2806 769 2814
rect 769 2806 772 2814
rect 776 2806 777 2814
rect 777 2806 779 2814
rect 779 2806 784 2814
rect 788 2806 789 2814
rect 789 2806 796 2814
rect 3748 2806 3755 2814
rect 3755 2806 3756 2814
rect 3760 2806 3765 2814
rect 3765 2806 3767 2814
rect 3767 2806 3768 2814
rect 3772 2806 3775 2814
rect 3775 2806 3777 2814
rect 3777 2806 3780 2814
rect 3784 2806 3785 2814
rect 3785 2806 3787 2814
rect 3787 2806 3792 2814
rect 3796 2806 3797 2814
rect 3797 2806 3804 2814
rect 6756 2806 6763 2814
rect 6763 2806 6764 2814
rect 6768 2806 6773 2814
rect 6773 2806 6775 2814
rect 6775 2806 6776 2814
rect 6780 2806 6783 2814
rect 6783 2806 6785 2814
rect 6785 2806 6788 2814
rect 6792 2806 6793 2814
rect 6793 2806 6795 2814
rect 6795 2806 6800 2814
rect 6804 2806 6805 2814
rect 6805 2806 6812 2814
rect 2924 2796 2932 2804
rect 2572 2776 2580 2784
rect 2636 2776 2644 2784
rect 3884 2796 3892 2804
rect 7148 2796 7156 2804
rect 4780 2776 4788 2784
rect 4972 2776 4980 2784
rect 5452 2776 5460 2784
rect 5580 2776 5588 2784
rect 5356 2756 5364 2764
rect 7500 2756 7508 2764
rect 1452 2736 1460 2744
rect 396 2716 404 2724
rect 844 2716 852 2724
rect 876 2716 884 2724
rect 1292 2716 1300 2724
rect 1516 2716 1524 2724
rect 3436 2716 3444 2724
rect 4012 2716 4020 2724
rect 5420 2716 5428 2724
rect 5644 2716 5652 2724
rect 6572 2716 6580 2724
rect 7180 2736 7188 2744
rect 620 2696 628 2704
rect 1196 2696 1204 2704
rect 1772 2696 1780 2704
rect 1836 2696 1844 2704
rect 2668 2696 2676 2704
rect 3692 2696 3700 2704
rect 4396 2696 4404 2704
rect 4460 2696 4468 2704
rect 4748 2696 4756 2704
rect 5100 2696 5108 2704
rect 5196 2696 5204 2704
rect 6412 2696 6420 2704
rect 6892 2696 6900 2704
rect 7276 2696 7284 2704
rect 652 2656 660 2664
rect 620 2636 628 2644
rect 1356 2656 1364 2664
rect 6156 2676 6164 2684
rect 7244 2676 7252 2684
rect 7468 2676 7476 2684
rect 7532 2676 7540 2684
rect 6892 2656 6900 2664
rect 2060 2636 2068 2644
rect 3468 2636 3476 2644
rect 5580 2636 5588 2644
rect 6636 2636 6644 2644
rect 7532 2636 7540 2644
rect 1420 2616 1428 2624
rect 1356 2596 1364 2604
rect 1772 2596 1780 2604
rect 2668 2616 2676 2624
rect 3372 2616 3380 2624
rect 2244 2606 2251 2614
rect 2251 2606 2252 2614
rect 2256 2606 2261 2614
rect 2261 2606 2263 2614
rect 2263 2606 2264 2614
rect 2268 2606 2271 2614
rect 2271 2606 2273 2614
rect 2273 2606 2276 2614
rect 2280 2606 2281 2614
rect 2281 2606 2283 2614
rect 2283 2606 2288 2614
rect 2292 2606 2293 2614
rect 2293 2606 2300 2614
rect 3212 2596 3220 2604
rect 4716 2616 4724 2624
rect 5356 2616 5364 2624
rect 5252 2606 5259 2614
rect 5259 2606 5260 2614
rect 5264 2606 5269 2614
rect 5269 2606 5271 2614
rect 5271 2606 5272 2614
rect 5276 2606 5279 2614
rect 5279 2606 5281 2614
rect 5281 2606 5284 2614
rect 5288 2606 5289 2614
rect 5289 2606 5291 2614
rect 5291 2606 5296 2614
rect 5300 2606 5301 2614
rect 5301 2606 5308 2614
rect 4748 2596 4756 2604
rect 5388 2596 5396 2604
rect 7404 2596 7412 2604
rect 236 2576 244 2584
rect 1068 2576 1076 2584
rect 3116 2576 3124 2584
rect 332 2556 340 2564
rect 1420 2556 1428 2564
rect 1676 2556 1684 2564
rect 1932 2556 1940 2564
rect 3884 2576 3892 2584
rect 4364 2556 4372 2564
rect 5068 2556 5076 2564
rect 6476 2576 6484 2584
rect 7372 2576 7380 2584
rect 1516 2536 1524 2544
rect 2700 2536 2708 2544
rect 3052 2536 3060 2544
rect 3148 2536 3156 2544
rect 4012 2536 4020 2544
rect 5132 2536 5140 2544
rect 6252 2556 6260 2564
rect 7180 2556 7188 2564
rect 7340 2556 7348 2564
rect 7564 2556 7572 2564
rect 5676 2536 5684 2544
rect 6412 2536 6420 2544
rect 6476 2536 6484 2544
rect 6988 2536 6996 2544
rect 7244 2536 7252 2544
rect 7436 2536 7444 2544
rect 236 2516 244 2524
rect 1100 2516 1108 2524
rect 2124 2516 2132 2524
rect 3948 2516 3956 2524
rect 4108 2516 4116 2524
rect 4428 2516 4436 2524
rect 5388 2516 5396 2524
rect 5548 2516 5556 2524
rect 6252 2516 6260 2524
rect 6956 2516 6964 2524
rect 7532 2516 7540 2524
rect 1452 2496 1460 2504
rect 2508 2496 2516 2504
rect 2636 2496 2644 2504
rect 2700 2496 2708 2504
rect 3596 2496 3604 2504
rect 5484 2496 5492 2504
rect 5516 2496 5524 2504
rect 7052 2496 7060 2504
rect 2700 2456 2708 2464
rect 4428 2456 4436 2464
rect 4524 2456 4532 2464
rect 4684 2456 4692 2464
rect 5612 2476 5620 2484
rect 6540 2476 6548 2484
rect 5356 2456 5364 2464
rect 6060 2456 6068 2464
rect 7148 2456 7156 2464
rect 7180 2456 7188 2464
rect 332 2436 340 2444
rect 1772 2436 1780 2444
rect 588 2416 596 2424
rect 3692 2436 3700 2444
rect 4204 2436 4212 2444
rect 6668 2436 6676 2444
rect 1964 2416 1972 2424
rect 1996 2416 2004 2424
rect 740 2406 747 2414
rect 747 2406 748 2414
rect 752 2406 757 2414
rect 757 2406 759 2414
rect 759 2406 760 2414
rect 764 2406 767 2414
rect 767 2406 769 2414
rect 769 2406 772 2414
rect 776 2406 777 2414
rect 777 2406 779 2414
rect 779 2406 784 2414
rect 788 2406 789 2414
rect 789 2406 796 2414
rect 3748 2406 3755 2414
rect 3755 2406 3756 2414
rect 3760 2406 3765 2414
rect 3765 2406 3767 2414
rect 3767 2406 3768 2414
rect 3772 2406 3775 2414
rect 3775 2406 3777 2414
rect 3777 2406 3780 2414
rect 3784 2406 3785 2414
rect 3785 2406 3787 2414
rect 3787 2406 3792 2414
rect 3796 2406 3797 2414
rect 3797 2406 3804 2414
rect 396 2396 404 2404
rect 1804 2396 1812 2404
rect 3628 2396 3636 2404
rect 6756 2406 6763 2414
rect 6763 2406 6764 2414
rect 6768 2406 6773 2414
rect 6773 2406 6775 2414
rect 6775 2406 6776 2414
rect 6780 2406 6783 2414
rect 6783 2406 6785 2414
rect 6785 2406 6788 2414
rect 6792 2406 6793 2414
rect 6793 2406 6795 2414
rect 6795 2406 6800 2414
rect 6804 2406 6805 2414
rect 6805 2406 6812 2414
rect 4524 2396 4532 2404
rect 4588 2396 4596 2404
rect 7532 2396 7540 2404
rect 1996 2376 2004 2384
rect 2028 2376 2036 2384
rect 3276 2376 3284 2384
rect 3468 2376 3476 2384
rect 4588 2356 4596 2364
rect 4652 2356 4660 2364
rect 5004 2356 5012 2364
rect 5420 2376 5428 2384
rect 5612 2376 5620 2384
rect 876 2316 884 2324
rect 44 2296 52 2304
rect 172 2296 180 2304
rect 204 2296 212 2304
rect 268 2296 276 2304
rect 2860 2336 2868 2344
rect 3468 2336 3476 2344
rect 3436 2316 3444 2324
rect 5356 2336 5364 2344
rect 7276 2336 7284 2344
rect 4268 2316 4276 2324
rect 4876 2316 4884 2324
rect 5132 2316 5140 2324
rect 5196 2316 5204 2324
rect 7116 2316 7124 2324
rect 7084 2296 7092 2304
rect 7500 2296 7508 2304
rect 1804 2276 1812 2284
rect 1900 2276 1908 2284
rect 2380 2276 2388 2284
rect 3308 2276 3316 2284
rect 5388 2276 5396 2284
rect 1292 2256 1300 2264
rect 2508 2256 2516 2264
rect 6924 2256 6932 2264
rect 7084 2256 7092 2264
rect 7468 2256 7476 2264
rect 556 2236 564 2244
rect 3884 2236 3892 2244
rect 2572 2216 2580 2224
rect 3660 2216 3668 2224
rect 4972 2236 4980 2244
rect 5068 2216 5076 2224
rect 5452 2216 5460 2224
rect 6188 2216 6196 2224
rect 6220 2216 6228 2224
rect 7212 2216 7220 2224
rect 2244 2206 2251 2214
rect 2251 2206 2252 2214
rect 2256 2206 2261 2214
rect 2261 2206 2263 2214
rect 2263 2206 2264 2214
rect 2268 2206 2271 2214
rect 2271 2206 2273 2214
rect 2273 2206 2276 2214
rect 2280 2206 2281 2214
rect 2281 2206 2283 2214
rect 2283 2206 2288 2214
rect 2292 2206 2293 2214
rect 2293 2206 2300 2214
rect 5252 2206 5259 2214
rect 5259 2206 5260 2214
rect 5264 2206 5269 2214
rect 5269 2206 5271 2214
rect 5271 2206 5272 2214
rect 5276 2206 5279 2214
rect 5279 2206 5281 2214
rect 5281 2206 5284 2214
rect 5288 2206 5289 2214
rect 5289 2206 5291 2214
rect 5291 2206 5296 2214
rect 5300 2206 5301 2214
rect 5301 2206 5308 2214
rect 1100 2196 1108 2204
rect 1900 2196 1908 2204
rect 2380 2196 2388 2204
rect 3212 2196 3220 2204
rect 4972 2196 4980 2204
rect 1484 2176 1492 2184
rect 1740 2176 1748 2184
rect 3532 2176 3540 2184
rect 5964 2196 5972 2204
rect 5356 2176 5364 2184
rect 44 2156 52 2164
rect 1196 2156 1204 2164
rect 4076 2156 4084 2164
rect 2380 2136 2388 2144
rect 2636 2136 2644 2144
rect 2892 2136 2900 2144
rect 3148 2136 3156 2144
rect 3532 2136 3540 2144
rect 4524 2136 4532 2144
rect 4620 2136 4628 2144
rect 7500 2176 7508 2184
rect 6572 2136 6580 2144
rect 6636 2136 6644 2144
rect 1068 2116 1076 2124
rect 1356 2116 1364 2124
rect 1996 2116 2004 2124
rect 1388 2096 1396 2104
rect 2796 2116 2804 2124
rect 3052 2116 3060 2124
rect 3628 2116 3636 2124
rect 5612 2116 5620 2124
rect 5836 2116 5844 2124
rect 6284 2116 6292 2124
rect 6316 2116 6324 2124
rect 7116 2116 7124 2124
rect 7148 2116 7156 2124
rect 2668 2096 2676 2104
rect 2700 2096 2708 2104
rect 3596 2096 3604 2104
rect 4556 2096 4564 2104
rect 5132 2096 5140 2104
rect 5196 2096 5204 2104
rect 6476 2096 6484 2104
rect 7052 2096 7060 2104
rect 588 2076 596 2084
rect 3564 2076 3572 2084
rect 4492 2076 4500 2084
rect 1740 2056 1748 2064
rect 1516 2036 1524 2044
rect 2508 2056 2516 2064
rect 3308 2056 3316 2064
rect 4300 2056 4308 2064
rect 4428 2056 4436 2064
rect 6188 2076 6196 2084
rect 7116 2076 7124 2084
rect 5964 2056 5972 2064
rect 5356 2036 5364 2044
rect 6892 2036 6900 2044
rect 204 2016 212 2024
rect 740 2006 747 2014
rect 747 2006 748 2014
rect 752 2006 757 2014
rect 757 2006 759 2014
rect 759 2006 760 2014
rect 764 2006 767 2014
rect 767 2006 769 2014
rect 769 2006 772 2014
rect 776 2006 777 2014
rect 777 2006 779 2014
rect 779 2006 784 2014
rect 788 2006 789 2014
rect 789 2006 796 2014
rect 3404 2016 3412 2024
rect 5004 2016 5012 2024
rect 5100 2016 5108 2024
rect 3748 2006 3755 2014
rect 3755 2006 3756 2014
rect 3760 2006 3765 2014
rect 3765 2006 3767 2014
rect 3767 2006 3768 2014
rect 3772 2006 3775 2014
rect 3775 2006 3777 2014
rect 3777 2006 3780 2014
rect 3784 2006 3785 2014
rect 3785 2006 3787 2014
rect 3787 2006 3792 2014
rect 3796 2006 3797 2014
rect 3797 2006 3804 2014
rect 6756 2006 6763 2014
rect 6763 2006 6764 2014
rect 6768 2006 6773 2014
rect 6773 2006 6775 2014
rect 6775 2006 6776 2014
rect 6780 2006 6783 2014
rect 6783 2006 6785 2014
rect 6785 2006 6788 2014
rect 6792 2006 6793 2014
rect 6793 2006 6795 2014
rect 6795 2006 6800 2014
rect 6804 2006 6805 2014
rect 6805 2006 6812 2014
rect 1772 1996 1780 2004
rect 1932 1996 1940 2004
rect 2028 1996 2036 2004
rect 2764 1996 2772 2004
rect 1260 1956 1268 1964
rect 1964 1956 1972 1964
rect 3436 1976 3444 1984
rect 3596 1976 3604 1984
rect 4076 1956 4084 1964
rect 5388 1956 5396 1964
rect 6924 1956 6932 1964
rect 7020 1956 7028 1964
rect 7564 1956 7572 1964
rect 2860 1936 2868 1944
rect 268 1916 276 1924
rect 1308 1916 1316 1924
rect 1580 1916 1588 1924
rect 1644 1916 1652 1924
rect 2092 1916 2100 1924
rect 2348 1916 2356 1924
rect 1804 1896 1812 1904
rect 3468 1936 3476 1944
rect 3948 1936 3956 1944
rect 3244 1896 3252 1904
rect 4588 1896 4596 1904
rect 5484 1916 5492 1924
rect 5516 1916 5524 1924
rect 4844 1896 4852 1904
rect 7276 1896 7284 1904
rect 1068 1876 1076 1884
rect 1100 1856 1108 1864
rect 1868 1876 1876 1884
rect 3052 1876 3060 1884
rect 3308 1876 3316 1884
rect 4332 1876 4340 1884
rect 1932 1856 1940 1864
rect 2604 1856 2612 1864
rect 3180 1856 3188 1864
rect 3660 1856 3668 1864
rect 4396 1856 4404 1864
rect 5004 1876 5012 1884
rect 6156 1876 6164 1884
rect 6988 1876 6996 1884
rect 7212 1876 7220 1884
rect 7532 1876 7540 1884
rect 6956 1856 6964 1864
rect 172 1836 180 1844
rect 1356 1836 1364 1844
rect 1484 1836 1492 1844
rect 4300 1836 4308 1844
rect 4524 1836 4532 1844
rect 4844 1836 4852 1844
rect 5036 1836 5044 1844
rect 908 1816 916 1824
rect 4556 1816 4564 1824
rect 4620 1816 4628 1824
rect 5388 1816 5396 1824
rect 5836 1816 5844 1824
rect 7116 1816 7124 1824
rect 2244 1806 2251 1814
rect 2251 1806 2252 1814
rect 2256 1806 2261 1814
rect 2261 1806 2263 1814
rect 2263 1806 2264 1814
rect 2268 1806 2271 1814
rect 2271 1806 2273 1814
rect 2273 1806 2276 1814
rect 2280 1806 2281 1814
rect 2281 1806 2283 1814
rect 2283 1806 2288 1814
rect 2292 1806 2293 1814
rect 2293 1806 2300 1814
rect 4076 1796 4084 1804
rect 5252 1806 5259 1814
rect 5259 1806 5260 1814
rect 5264 1806 5269 1814
rect 5269 1806 5271 1814
rect 5271 1806 5272 1814
rect 5276 1806 5279 1814
rect 5279 1806 5281 1814
rect 5281 1806 5284 1814
rect 5288 1806 5289 1814
rect 5289 1806 5291 1814
rect 5291 1806 5296 1814
rect 5300 1806 5301 1814
rect 5301 1806 5308 1814
rect 6412 1796 6420 1804
rect 2764 1776 2772 1784
rect 1004 1756 1012 1764
rect 2780 1756 2788 1764
rect 3244 1756 3252 1764
rect 4140 1776 4148 1784
rect 4556 1776 4564 1784
rect 6604 1776 6612 1784
rect 7532 1776 7540 1784
rect 5452 1756 5460 1764
rect 5676 1756 5684 1764
rect 7116 1756 7124 1764
rect 7244 1756 7252 1764
rect 1292 1736 1300 1744
rect 1516 1736 1524 1744
rect 2444 1736 2452 1744
rect 2572 1736 2580 1744
rect 332 1716 340 1724
rect 1068 1716 1076 1724
rect 1836 1716 1844 1724
rect 2124 1716 2132 1724
rect 2764 1716 2772 1724
rect 2860 1716 2868 1724
rect 3404 1716 3412 1724
rect 4268 1716 4276 1724
rect 7500 1716 7508 1724
rect 1004 1696 1012 1704
rect 1132 1696 1140 1704
rect 2028 1696 2036 1704
rect 2348 1696 2356 1704
rect 3276 1696 3284 1704
rect 4012 1696 4020 1704
rect 4684 1696 4692 1704
rect 6924 1696 6932 1704
rect 7052 1696 7060 1704
rect 7212 1696 7220 1704
rect 7436 1696 7444 1704
rect 1356 1656 1364 1664
rect 1932 1676 1940 1684
rect 2060 1676 2068 1684
rect 3596 1676 3604 1684
rect 4268 1676 4276 1684
rect 7500 1676 7508 1684
rect 2348 1636 2356 1644
rect 3308 1636 3316 1644
rect 4460 1636 4468 1644
rect 4844 1636 4852 1644
rect 7276 1636 7284 1644
rect 1772 1616 1780 1624
rect 2060 1616 2068 1624
rect 4332 1616 4340 1624
rect 740 1606 747 1614
rect 747 1606 748 1614
rect 752 1606 757 1614
rect 757 1606 759 1614
rect 759 1606 760 1614
rect 764 1606 767 1614
rect 767 1606 769 1614
rect 769 1606 772 1614
rect 776 1606 777 1614
rect 777 1606 779 1614
rect 779 1606 784 1614
rect 788 1606 789 1614
rect 789 1606 796 1614
rect 3748 1606 3755 1614
rect 3755 1606 3756 1614
rect 3760 1606 3765 1614
rect 3765 1606 3767 1614
rect 3767 1606 3768 1614
rect 3772 1606 3775 1614
rect 3775 1606 3777 1614
rect 3777 1606 3780 1614
rect 3784 1606 3785 1614
rect 3785 1606 3787 1614
rect 3787 1606 3792 1614
rect 3796 1606 3797 1614
rect 3797 1606 3804 1614
rect 6756 1606 6763 1614
rect 6763 1606 6764 1614
rect 6768 1606 6773 1614
rect 6773 1606 6775 1614
rect 6775 1606 6776 1614
rect 6780 1606 6783 1614
rect 6783 1606 6785 1614
rect 6785 1606 6788 1614
rect 6792 1606 6793 1614
rect 6793 1606 6795 1614
rect 6795 1606 6800 1614
rect 6804 1606 6805 1614
rect 6805 1606 6812 1614
rect 556 1576 564 1584
rect 3212 1596 3220 1604
rect 3532 1576 3540 1584
rect 3628 1576 3636 1584
rect 5484 1596 5492 1604
rect 1388 1556 1396 1564
rect 1580 1556 1588 1564
rect 2732 1556 2740 1564
rect 5100 1576 5108 1584
rect 5388 1576 5396 1584
rect 6284 1576 6292 1584
rect 3884 1556 3892 1564
rect 1516 1516 1524 1524
rect 4460 1536 4468 1544
rect 4396 1516 4404 1524
rect 5004 1516 5012 1524
rect 5100 1516 5108 1524
rect 1644 1496 1652 1504
rect 1804 1496 1812 1504
rect 3244 1496 3252 1504
rect 4172 1496 4180 1504
rect 4364 1496 4372 1504
rect 4524 1496 4532 1504
rect 5548 1496 5556 1504
rect 332 1476 340 1484
rect 2348 1476 2356 1484
rect 3340 1476 3348 1484
rect 4204 1476 4212 1484
rect 4396 1476 4404 1484
rect 7372 1516 7380 1524
rect 7532 1496 7540 1504
rect 7340 1476 7348 1484
rect 1868 1456 1876 1464
rect 1932 1456 1940 1464
rect 1996 1456 2004 1464
rect 2156 1456 2164 1464
rect 3660 1456 3668 1464
rect 4236 1456 4244 1464
rect 7116 1456 7124 1464
rect 1100 1436 1108 1444
rect 1996 1416 2004 1424
rect 2764 1416 2772 1424
rect 3020 1416 3028 1424
rect 6956 1436 6964 1444
rect 6988 1436 6996 1444
rect 7052 1436 7060 1444
rect 2244 1406 2251 1414
rect 2251 1406 2252 1414
rect 2256 1406 2261 1414
rect 2261 1406 2263 1414
rect 2263 1406 2264 1414
rect 2268 1406 2271 1414
rect 2271 1406 2273 1414
rect 2273 1406 2276 1414
rect 2280 1406 2281 1414
rect 2281 1406 2283 1414
rect 2283 1406 2288 1414
rect 2292 1406 2293 1414
rect 2293 1406 2300 1414
rect 5252 1406 5259 1414
rect 5259 1406 5260 1414
rect 5264 1406 5269 1414
rect 5269 1406 5271 1414
rect 5271 1406 5272 1414
rect 5276 1406 5279 1414
rect 5279 1406 5281 1414
rect 5281 1406 5284 1414
rect 5288 1406 5289 1414
rect 5289 1406 5291 1414
rect 5291 1406 5296 1414
rect 5300 1406 5301 1414
rect 5301 1406 5308 1414
rect 1228 1396 1236 1404
rect 3276 1396 3284 1404
rect 4780 1396 4788 1404
rect 4876 1396 4884 1404
rect 5164 1396 5172 1404
rect 6924 1396 6932 1404
rect 6956 1396 6964 1404
rect 7180 1396 7188 1404
rect 1100 1376 1108 1384
rect 2028 1376 2036 1384
rect 3052 1376 3060 1384
rect 1580 1356 1588 1364
rect 3404 1356 3412 1364
rect 3628 1356 3636 1364
rect 4492 1356 4500 1364
rect 7180 1356 7188 1364
rect 908 1336 916 1344
rect 1132 1336 1140 1344
rect 1676 1336 1684 1344
rect 1964 1336 1972 1344
rect 2188 1336 2196 1344
rect 2412 1336 2420 1344
rect 4556 1336 4564 1344
rect 1836 1316 1844 1324
rect 1996 1316 2004 1324
rect 2028 1316 2036 1324
rect 3212 1316 3220 1324
rect 3948 1316 3956 1324
rect 4236 1316 4244 1324
rect 5036 1316 5044 1324
rect 5964 1316 5972 1324
rect 6252 1316 6260 1324
rect 1292 1296 1300 1304
rect 1676 1296 1684 1304
rect 4172 1296 4180 1304
rect 1900 1256 1908 1264
rect 3212 1276 3220 1284
rect 3276 1256 3284 1264
rect 3948 1256 3956 1264
rect 7180 1296 7188 1304
rect 5580 1276 5588 1284
rect 6572 1276 6580 1284
rect 6636 1276 6644 1284
rect 7084 1276 7092 1284
rect 5740 1256 5748 1264
rect 1964 1236 1972 1244
rect 2508 1236 2516 1244
rect 3692 1236 3700 1244
rect 2604 1216 2612 1224
rect 3372 1216 3380 1224
rect 4780 1216 4788 1224
rect 5068 1216 5076 1224
rect 5420 1216 5428 1224
rect 740 1206 747 1214
rect 747 1206 748 1214
rect 752 1206 757 1214
rect 757 1206 759 1214
rect 759 1206 760 1214
rect 764 1206 767 1214
rect 767 1206 769 1214
rect 769 1206 772 1214
rect 776 1206 777 1214
rect 777 1206 779 1214
rect 779 1206 784 1214
rect 788 1206 789 1214
rect 789 1206 796 1214
rect 3748 1206 3755 1214
rect 3755 1206 3756 1214
rect 3760 1206 3765 1214
rect 3765 1206 3767 1214
rect 3767 1206 3768 1214
rect 3772 1206 3775 1214
rect 3775 1206 3777 1214
rect 3777 1206 3780 1214
rect 3784 1206 3785 1214
rect 3785 1206 3787 1214
rect 3787 1206 3792 1214
rect 3796 1206 3797 1214
rect 3797 1206 3804 1214
rect 6756 1206 6763 1214
rect 6763 1206 6764 1214
rect 6768 1206 6773 1214
rect 6773 1206 6775 1214
rect 6775 1206 6776 1214
rect 6780 1206 6783 1214
rect 6783 1206 6785 1214
rect 6785 1206 6788 1214
rect 6792 1206 6793 1214
rect 6793 1206 6795 1214
rect 6795 1206 6800 1214
rect 6804 1206 6805 1214
rect 6805 1206 6812 1214
rect 3852 1196 3860 1204
rect 6540 1196 6548 1204
rect 1548 1176 1556 1184
rect 2092 1176 2100 1184
rect 2124 1176 2132 1184
rect 2508 1176 2516 1184
rect 2732 1176 2740 1184
rect 2188 1156 2196 1164
rect 3916 1176 3924 1184
rect 3948 1156 3956 1164
rect 4268 1156 4276 1164
rect 876 1096 884 1104
rect 1100 1096 1108 1104
rect 1228 1116 1236 1124
rect 1804 1116 1812 1124
rect 1964 1116 1972 1124
rect 3308 1136 3316 1144
rect 5004 1136 5012 1144
rect 3628 1116 3636 1124
rect 5196 1116 5204 1124
rect 5612 1116 5620 1124
rect 5836 1116 5844 1124
rect 7084 1116 7092 1124
rect 2476 1096 2484 1104
rect 2892 1096 2900 1104
rect 4844 1096 4852 1104
rect 3084 1076 3092 1084
rect 3564 1076 3572 1084
rect 3852 1076 3860 1084
rect 6220 1096 6228 1104
rect 7436 1096 7444 1104
rect 7564 1096 7572 1104
rect 6252 1076 6260 1084
rect 6700 1076 6708 1084
rect 7308 1076 7316 1084
rect 204 1036 212 1044
rect 3372 1036 3380 1044
rect 3532 1036 3540 1044
rect 5964 1036 5972 1044
rect 6700 1036 6708 1044
rect 12 1016 20 1024
rect 2124 1016 2132 1024
rect 2156 1016 2164 1024
rect 2412 1016 2420 1024
rect 2444 1016 2452 1024
rect 2860 1016 2868 1024
rect 3020 1016 3028 1024
rect 5580 1016 5588 1024
rect 5740 1016 5748 1024
rect 7084 1016 7092 1024
rect 2244 1006 2251 1014
rect 2251 1006 2252 1014
rect 2256 1006 2261 1014
rect 2261 1006 2263 1014
rect 2263 1006 2264 1014
rect 2268 1006 2271 1014
rect 2271 1006 2273 1014
rect 2273 1006 2276 1014
rect 2280 1006 2281 1014
rect 2281 1006 2283 1014
rect 2283 1006 2288 1014
rect 2292 1006 2293 1014
rect 2293 1006 2300 1014
rect 5252 1006 5259 1014
rect 5259 1006 5260 1014
rect 5264 1006 5269 1014
rect 5269 1006 5271 1014
rect 5271 1006 5272 1014
rect 5276 1006 5279 1014
rect 5279 1006 5281 1014
rect 5281 1006 5284 1014
rect 5288 1006 5289 1014
rect 5289 1006 5291 1014
rect 5291 1006 5296 1014
rect 5300 1006 5301 1014
rect 5301 1006 5308 1014
rect 396 996 404 1004
rect 876 976 884 984
rect 12 956 20 964
rect 1676 976 1684 984
rect 2476 976 2484 984
rect 1644 916 1652 924
rect 2060 936 2068 944
rect 3052 976 3060 984
rect 3308 976 3316 984
rect 3500 976 3508 984
rect 7532 996 7540 1004
rect 6700 976 6708 984
rect 3564 956 3572 964
rect 3052 936 3060 944
rect 4300 936 4308 944
rect 4428 956 4436 964
rect 4460 936 4468 944
rect 4844 956 4852 964
rect 6092 956 6100 964
rect 6156 956 6164 964
rect 7244 936 7252 944
rect 396 896 404 904
rect 1196 896 1204 904
rect 1580 896 1588 904
rect 1932 896 1940 904
rect 2060 896 2068 904
rect 3052 896 3060 904
rect 3244 896 3252 904
rect 3500 896 3508 904
rect 3692 896 3700 904
rect 3948 896 3956 904
rect 4076 916 4084 924
rect 4108 896 4116 904
rect 4620 896 4628 904
rect 4684 896 4692 904
rect 5612 896 5620 904
rect 1516 876 1524 884
rect 3084 876 3092 884
rect 3116 876 3124 884
rect 3884 856 3892 864
rect 4332 856 4340 864
rect 6092 876 6100 884
rect 7276 876 7284 884
rect 5772 856 5780 864
rect 3308 836 3316 844
rect 5676 836 5684 844
rect 6956 836 6964 844
rect 1900 816 1908 824
rect 1932 816 1940 824
rect 2828 816 2836 824
rect 3340 816 3348 824
rect 740 806 747 814
rect 747 806 748 814
rect 752 806 757 814
rect 757 806 759 814
rect 759 806 760 814
rect 764 806 767 814
rect 767 806 769 814
rect 769 806 772 814
rect 776 806 777 814
rect 777 806 779 814
rect 779 806 784 814
rect 788 806 789 814
rect 789 806 796 814
rect 3748 806 3755 814
rect 3755 806 3756 814
rect 3760 806 3765 814
rect 3765 806 3767 814
rect 3767 806 3768 814
rect 3772 806 3775 814
rect 3775 806 3777 814
rect 3777 806 3780 814
rect 3784 806 3785 814
rect 3785 806 3787 814
rect 3787 806 3792 814
rect 3796 806 3797 814
rect 3797 806 3804 814
rect 6756 806 6763 814
rect 6763 806 6764 814
rect 6768 806 6773 814
rect 6773 806 6775 814
rect 6775 806 6776 814
rect 6780 806 6783 814
rect 6783 806 6785 814
rect 6785 806 6788 814
rect 6792 806 6793 814
rect 6793 806 6795 814
rect 6795 806 6800 814
rect 6804 806 6805 814
rect 6805 806 6812 814
rect 396 796 404 804
rect 2380 796 2388 804
rect 2892 796 2900 804
rect 6700 796 6708 804
rect 44 776 52 784
rect 1900 776 1908 784
rect 3244 776 3252 784
rect 5004 776 5012 784
rect 6508 756 6516 764
rect 1644 736 1652 744
rect 3404 736 3412 744
rect 1548 716 1556 724
rect 1580 716 1588 724
rect 1836 716 1844 724
rect 3084 716 3092 724
rect 3628 716 3636 724
rect 3916 716 3924 724
rect 4364 716 4372 724
rect 4620 716 4628 724
rect 6220 736 6228 744
rect 7436 736 7444 744
rect 5164 716 5172 724
rect 6988 716 6996 724
rect 2572 676 2580 684
rect 3564 696 3572 704
rect 6156 696 6164 704
rect 6220 696 6228 704
rect 4396 656 4404 664
rect 4844 656 4852 664
rect 5772 656 5780 664
rect 1900 616 1908 624
rect 2188 616 2196 624
rect 3084 616 3092 624
rect 3308 616 3316 624
rect 2244 606 2251 614
rect 2251 606 2252 614
rect 2256 606 2261 614
rect 2261 606 2263 614
rect 2263 606 2264 614
rect 2268 606 2271 614
rect 2271 606 2273 614
rect 2273 606 2276 614
rect 2280 606 2281 614
rect 2281 606 2283 614
rect 2283 606 2288 614
rect 2292 606 2293 614
rect 2293 606 2300 614
rect 1676 596 1684 604
rect 3404 596 3412 604
rect 4492 616 4500 624
rect 5964 616 5972 624
rect 5252 606 5259 614
rect 5259 606 5260 614
rect 5264 606 5269 614
rect 5269 606 5271 614
rect 5271 606 5272 614
rect 5276 606 5279 614
rect 5279 606 5281 614
rect 5281 606 5284 614
rect 5288 606 5289 614
rect 5289 606 5291 614
rect 5291 606 5296 614
rect 5300 606 5301 614
rect 5301 606 5308 614
rect 588 576 596 584
rect 908 576 916 584
rect 3244 576 3252 584
rect 1932 556 1940 564
rect 2572 556 2580 564
rect 7372 576 7380 584
rect 6636 556 6644 564
rect 1996 536 2004 544
rect 1644 516 1652 524
rect 4364 536 4372 544
rect 4684 536 4692 544
rect 5356 536 5364 544
rect 5612 536 5620 544
rect 7500 536 7508 544
rect 4940 516 4948 524
rect 5388 516 5396 524
rect 7244 516 7252 524
rect 1836 476 1844 484
rect 1804 456 1812 464
rect 5420 456 5428 464
rect 1964 436 1972 444
rect 2188 436 2196 444
rect 3404 436 3412 444
rect 3916 436 3924 444
rect 4332 436 4340 444
rect 556 416 564 424
rect 4076 416 4084 424
rect 740 406 747 414
rect 747 406 748 414
rect 752 406 757 414
rect 757 406 759 414
rect 759 406 760 414
rect 764 406 767 414
rect 767 406 769 414
rect 769 406 772 414
rect 776 406 777 414
rect 777 406 779 414
rect 779 406 784 414
rect 788 406 789 414
rect 789 406 796 414
rect 3748 406 3755 414
rect 3755 406 3756 414
rect 3760 406 3765 414
rect 3765 406 3767 414
rect 3767 406 3768 414
rect 3772 406 3775 414
rect 3775 406 3777 414
rect 3777 406 3780 414
rect 3784 406 3785 414
rect 3785 406 3787 414
rect 3787 406 3792 414
rect 3796 406 3797 414
rect 3797 406 3804 414
rect 6756 406 6763 414
rect 6763 406 6764 414
rect 6768 406 6773 414
rect 6773 406 6775 414
rect 6775 406 6776 414
rect 6780 406 6783 414
rect 6783 406 6785 414
rect 6785 406 6788 414
rect 6792 406 6793 414
rect 6793 406 6795 414
rect 6795 406 6800 414
rect 6804 406 6805 414
rect 6805 406 6812 414
rect 1644 396 1652 404
rect 2188 396 2196 404
rect 1964 376 1972 384
rect 1740 356 1748 364
rect 3116 356 3124 364
rect 4812 356 4820 364
rect 5676 356 5684 364
rect 2732 336 2740 344
rect 3052 336 3060 344
rect 3852 336 3860 344
rect 3884 336 3892 344
rect 908 316 916 324
rect 1740 316 1748 324
rect 2828 316 2836 324
rect 1164 296 1172 304
rect 5612 316 5620 324
rect 3916 296 3924 304
rect 6540 296 6548 304
rect 2860 276 2868 284
rect 7148 276 7156 284
rect 1164 236 1172 244
rect 1228 236 1236 244
rect 4492 216 4500 224
rect 2244 206 2251 214
rect 2251 206 2252 214
rect 2256 206 2261 214
rect 2261 206 2263 214
rect 2263 206 2264 214
rect 2268 206 2271 214
rect 2271 206 2273 214
rect 2273 206 2276 214
rect 2280 206 2281 214
rect 2281 206 2283 214
rect 2283 206 2288 214
rect 2292 206 2293 214
rect 2293 206 2300 214
rect 5252 206 5259 214
rect 5259 206 5260 214
rect 5264 206 5269 214
rect 5269 206 5271 214
rect 5271 206 5272 214
rect 5276 206 5279 214
rect 5279 206 5281 214
rect 5281 206 5284 214
rect 5288 206 5289 214
rect 5289 206 5291 214
rect 5291 206 5296 214
rect 5300 206 5301 214
rect 5301 206 5308 214
rect 2732 176 2740 184
rect 5356 176 5364 184
rect 4396 156 4404 164
rect 4364 136 4372 144
rect 4812 116 4820 124
rect 4940 116 4948 124
rect 5388 136 5396 144
rect 7468 136 7476 144
rect 7340 116 7348 124
rect 7532 116 7540 124
rect 1228 56 1236 64
rect 1196 36 1204 44
rect 1644 36 1652 44
rect 5676 16 5684 24
rect 740 6 747 14
rect 747 6 748 14
rect 752 6 757 14
rect 757 6 759 14
rect 759 6 760 14
rect 764 6 767 14
rect 767 6 769 14
rect 769 6 772 14
rect 776 6 777 14
rect 777 6 779 14
rect 779 6 784 14
rect 788 6 789 14
rect 789 6 796 14
rect 3748 6 3755 14
rect 3755 6 3756 14
rect 3760 6 3765 14
rect 3765 6 3767 14
rect 3767 6 3768 14
rect 3772 6 3775 14
rect 3775 6 3777 14
rect 3777 6 3780 14
rect 3784 6 3785 14
rect 3785 6 3787 14
rect 3787 6 3792 14
rect 3796 6 3797 14
rect 3797 6 3804 14
rect 6756 6 6763 14
rect 6763 6 6764 14
rect 6768 6 6773 14
rect 6773 6 6775 14
rect 6775 6 6776 14
rect 6780 6 6783 14
rect 6783 6 6785 14
rect 6785 6 6788 14
rect 6792 6 6793 14
rect 6793 6 6795 14
rect 6795 6 6800 14
rect 6804 6 6805 14
rect 6805 6 6812 14
<< metal4 >>
rect 4746 5224 4758 5226
rect 4746 5216 4748 5224
rect 4756 5216 4758 5224
rect 736 5214 800 5216
rect 736 5206 740 5214
rect 748 5206 752 5214
rect 760 5206 764 5214
rect 772 5206 776 5214
rect 784 5206 788 5214
rect 796 5206 800 5214
rect 736 4814 800 5206
rect 1258 5104 1270 5106
rect 1258 5096 1260 5104
rect 1268 5096 1270 5104
rect 1258 5024 1270 5096
rect 1258 5016 1260 5024
rect 1268 5016 1270 5024
rect 1258 5014 1270 5016
rect 1674 5064 1686 5066
rect 1674 5056 1676 5064
rect 1684 5056 1686 5064
rect 736 4806 740 4814
rect 748 4806 752 4814
rect 760 4806 764 4814
rect 772 4806 776 4814
rect 784 4806 788 4814
rect 796 4806 800 4814
rect 330 4644 342 4646
rect 330 4636 332 4644
rect 340 4636 342 4644
rect 234 4584 246 4586
rect 234 4576 236 4584
rect 244 4576 246 4584
rect 170 3524 182 3526
rect 170 3516 172 3524
rect 180 3516 182 3524
rect 170 3164 182 3516
rect 170 3156 172 3164
rect 180 3156 182 3164
rect 170 3104 182 3156
rect 170 3096 172 3104
rect 180 3096 182 3104
rect 170 3094 182 3096
rect 202 3104 214 3106
rect 202 3096 204 3104
rect 212 3096 214 3104
rect 42 2304 54 2306
rect 42 2296 44 2304
rect 52 2296 54 2304
rect 42 2164 54 2296
rect 42 2156 44 2164
rect 52 2156 54 2164
rect 10 1024 22 1026
rect 10 1016 12 1024
rect 20 1016 22 1024
rect 10 964 22 1016
rect 10 956 12 964
rect 20 956 22 964
rect 10 954 22 956
rect 42 784 54 2156
rect 170 2304 182 2306
rect 170 2296 172 2304
rect 180 2296 182 2304
rect 170 1844 182 2296
rect 202 2304 214 3096
rect 234 2964 246 4576
rect 266 4524 278 4526
rect 266 4516 268 4524
rect 276 4516 278 4524
rect 266 3944 278 4516
rect 330 4124 342 4636
rect 554 4644 566 4646
rect 554 4636 556 4644
rect 564 4636 566 4644
rect 554 4604 566 4636
rect 554 4596 556 4604
rect 564 4596 566 4604
rect 330 4116 332 4124
rect 340 4116 342 4124
rect 330 4114 342 4116
rect 522 4224 534 4226
rect 522 4216 524 4224
rect 532 4216 534 4224
rect 266 3936 268 3944
rect 276 3936 278 3944
rect 266 3744 278 3936
rect 362 3924 374 3926
rect 362 3916 364 3924
rect 372 3916 374 3924
rect 362 3784 374 3916
rect 362 3776 364 3784
rect 372 3776 374 3784
rect 362 3774 374 3776
rect 266 3736 268 3744
rect 276 3736 278 3744
rect 266 3734 278 3736
rect 234 2956 236 2964
rect 244 2956 246 2964
rect 234 2954 246 2956
rect 330 3464 342 3466
rect 330 3456 332 3464
rect 340 3456 342 3464
rect 234 2584 246 2586
rect 234 2576 236 2584
rect 244 2576 246 2584
rect 234 2524 246 2576
rect 330 2564 342 3456
rect 522 3404 534 4216
rect 554 3684 566 4596
rect 554 3676 556 3684
rect 564 3676 566 3684
rect 554 3674 566 3676
rect 736 4414 800 4806
rect 1002 4804 1014 4806
rect 1002 4796 1004 4804
rect 1012 4796 1014 4804
rect 938 4664 950 4666
rect 938 4656 940 4664
rect 948 4656 950 4664
rect 938 4646 950 4656
rect 906 4644 950 4646
rect 906 4636 908 4644
rect 916 4636 950 4644
rect 906 4634 950 4636
rect 1002 4604 1014 4796
rect 1578 4804 1590 4806
rect 1578 4796 1580 4804
rect 1588 4796 1590 4804
rect 1546 4764 1558 4766
rect 1546 4756 1548 4764
rect 1556 4756 1558 4764
rect 1002 4596 1004 4604
rect 1012 4596 1014 4604
rect 1002 4594 1014 4596
rect 1162 4704 1174 4706
rect 1162 4696 1164 4704
rect 1172 4696 1174 4704
rect 736 4406 740 4414
rect 748 4406 752 4414
rect 760 4406 764 4414
rect 772 4406 776 4414
rect 784 4406 788 4414
rect 796 4406 800 4414
rect 736 4014 800 4406
rect 1130 4524 1142 4526
rect 1130 4516 1132 4524
rect 1140 4516 1142 4524
rect 736 4006 740 4014
rect 748 4006 752 4014
rect 760 4006 764 4014
rect 772 4006 776 4014
rect 784 4006 788 4014
rect 796 4006 800 4014
rect 736 3614 800 4006
rect 906 4204 918 4206
rect 906 4196 908 4204
rect 916 4196 918 4204
rect 906 3904 918 4196
rect 906 3896 908 3904
rect 916 3896 918 3904
rect 906 3894 918 3896
rect 736 3606 740 3614
rect 748 3606 752 3614
rect 760 3606 764 3614
rect 772 3606 776 3614
rect 784 3606 788 3614
rect 796 3606 800 3614
rect 522 3396 524 3404
rect 532 3396 534 3404
rect 522 3394 534 3396
rect 650 3504 662 3506
rect 650 3496 652 3504
rect 660 3496 662 3504
rect 650 3264 662 3496
rect 650 3256 652 3264
rect 660 3256 662 3264
rect 554 3084 566 3086
rect 554 3076 556 3084
rect 564 3076 566 3084
rect 330 2556 332 2564
rect 340 2556 342 2564
rect 330 2554 342 2556
rect 394 2724 406 2726
rect 394 2716 396 2724
rect 404 2716 406 2724
rect 234 2516 236 2524
rect 244 2516 246 2524
rect 234 2514 246 2516
rect 330 2444 342 2446
rect 330 2436 332 2444
rect 340 2436 342 2444
rect 202 2296 204 2304
rect 212 2296 214 2304
rect 202 2294 214 2296
rect 266 2304 278 2306
rect 266 2296 268 2304
rect 276 2296 278 2304
rect 170 1836 172 1844
rect 180 1836 182 1844
rect 170 1834 182 1836
rect 202 2024 214 2026
rect 202 2016 204 2024
rect 212 2016 214 2024
rect 202 1044 214 2016
rect 266 1924 278 2296
rect 266 1916 268 1924
rect 276 1916 278 1924
rect 266 1914 278 1916
rect 330 1724 342 2436
rect 394 2404 406 2716
rect 394 2396 396 2404
rect 404 2396 406 2404
rect 394 2394 406 2396
rect 554 2244 566 3076
rect 586 2964 598 2966
rect 586 2956 588 2964
rect 596 2956 598 2964
rect 586 2424 598 2956
rect 618 2704 630 2706
rect 618 2696 620 2704
rect 628 2696 630 2704
rect 618 2644 630 2696
rect 650 2664 662 3256
rect 650 2656 652 2664
rect 660 2656 662 2664
rect 650 2654 662 2656
rect 736 3214 800 3606
rect 736 3206 740 3214
rect 748 3206 752 3214
rect 760 3206 764 3214
rect 772 3206 776 3214
rect 784 3206 788 3214
rect 796 3206 800 3214
rect 736 2814 800 3206
rect 874 3824 886 3826
rect 874 3816 876 3824
rect 884 3816 886 3824
rect 736 2806 740 2814
rect 748 2806 752 2814
rect 760 2806 764 2814
rect 772 2806 776 2814
rect 784 2806 788 2814
rect 796 2806 800 2814
rect 618 2636 620 2644
rect 628 2636 630 2644
rect 618 2634 630 2636
rect 586 2416 588 2424
rect 596 2416 598 2424
rect 586 2414 598 2416
rect 736 2414 800 2806
rect 842 2824 854 2826
rect 842 2816 844 2824
rect 852 2816 854 2824
rect 842 2724 854 2816
rect 842 2716 844 2724
rect 852 2716 854 2724
rect 842 2714 854 2716
rect 874 2724 886 3816
rect 1130 3804 1142 4516
rect 1162 4224 1174 4696
rect 1546 4624 1558 4756
rect 1546 4616 1548 4624
rect 1556 4616 1558 4624
rect 1546 4614 1558 4616
rect 1162 4216 1164 4224
rect 1172 4216 1174 4224
rect 1162 4214 1174 4216
rect 1194 4544 1206 4546
rect 1194 4536 1196 4544
rect 1204 4536 1206 4544
rect 1194 4184 1206 4536
rect 1194 4176 1196 4184
rect 1204 4176 1206 4184
rect 1194 4174 1206 4176
rect 1258 4284 1270 4286
rect 1258 4276 1260 4284
rect 1268 4276 1270 4284
rect 1130 3796 1132 3804
rect 1140 3796 1142 3804
rect 1130 3744 1142 3796
rect 1130 3736 1132 3744
rect 1140 3736 1142 3744
rect 1130 3734 1142 3736
rect 1194 4104 1206 4106
rect 1194 4096 1196 4104
rect 1204 4096 1206 4104
rect 938 3684 950 3686
rect 938 3676 940 3684
rect 948 3676 950 3684
rect 938 3644 950 3676
rect 938 3636 940 3644
rect 948 3636 950 3644
rect 938 3634 950 3636
rect 970 3344 982 3346
rect 970 3336 972 3344
rect 980 3336 982 3344
rect 970 2944 982 3336
rect 970 2936 972 2944
rect 980 2936 982 2944
rect 970 2904 982 2936
rect 970 2896 972 2904
rect 980 2896 982 2904
rect 970 2894 982 2896
rect 1066 3064 1078 3066
rect 1066 3056 1068 3064
rect 1076 3056 1078 3064
rect 874 2716 876 2724
rect 884 2716 886 2724
rect 874 2714 886 2716
rect 1066 2584 1078 3056
rect 1066 2576 1068 2584
rect 1076 2576 1078 2584
rect 1066 2574 1078 2576
rect 1194 2704 1206 4096
rect 1258 3624 1270 4276
rect 1290 4224 1302 4226
rect 1290 4216 1292 4224
rect 1300 4216 1302 4224
rect 1290 3904 1302 4216
rect 1354 4124 1366 4126
rect 1354 4116 1356 4124
rect 1364 4116 1366 4124
rect 1290 3896 1292 3904
rect 1300 3896 1302 3904
rect 1290 3894 1302 3896
rect 1322 3984 1334 3986
rect 1322 3976 1324 3984
rect 1332 3976 1334 3984
rect 1258 3616 1260 3624
rect 1268 3616 1270 3624
rect 1258 3614 1270 3616
rect 1322 3204 1334 3976
rect 1322 3196 1324 3204
rect 1332 3196 1334 3204
rect 1322 3194 1334 3196
rect 1354 3904 1366 4116
rect 1354 3896 1356 3904
rect 1364 3896 1366 3904
rect 1354 3504 1366 3896
rect 1386 4124 1398 4126
rect 1386 4116 1388 4124
rect 1396 4116 1398 4124
rect 1386 3524 1398 4116
rect 1482 4064 1494 4066
rect 1482 4056 1484 4064
rect 1492 4056 1494 4064
rect 1386 3516 1388 3524
rect 1396 3516 1398 3524
rect 1386 3514 1398 3516
rect 1418 3924 1430 3926
rect 1418 3916 1420 3924
rect 1428 3916 1430 3924
rect 1354 3496 1356 3504
rect 1364 3496 1366 3504
rect 1354 3084 1366 3496
rect 1386 3404 1398 3406
rect 1386 3396 1388 3404
rect 1396 3396 1398 3404
rect 1386 3124 1398 3396
rect 1418 3324 1430 3916
rect 1482 3884 1494 4056
rect 1482 3876 1484 3884
rect 1492 3876 1494 3884
rect 1482 3874 1494 3876
rect 1418 3316 1420 3324
rect 1428 3316 1430 3324
rect 1418 3314 1430 3316
rect 1482 3744 1494 3746
rect 1482 3736 1484 3744
rect 1492 3736 1494 3744
rect 1386 3116 1388 3124
rect 1396 3116 1398 3124
rect 1386 3114 1398 3116
rect 1450 3304 1462 3306
rect 1450 3296 1452 3304
rect 1460 3296 1462 3304
rect 1450 3104 1462 3296
rect 1482 3264 1494 3736
rect 1578 3564 1590 4796
rect 1642 4684 1654 4686
rect 1642 4676 1644 4684
rect 1652 4676 1654 4684
rect 1610 4644 1622 4646
rect 1610 4636 1612 4644
rect 1620 4636 1622 4644
rect 1610 4524 1622 4636
rect 1610 4516 1612 4524
rect 1620 4516 1622 4524
rect 1610 4514 1622 4516
rect 1642 4524 1654 4676
rect 1642 4516 1644 4524
rect 1652 4516 1654 4524
rect 1642 4514 1654 4516
rect 1674 4084 1686 5056
rect 2240 5014 2304 5216
rect 2240 5006 2244 5014
rect 2252 5006 2256 5014
rect 2264 5006 2268 5014
rect 2276 5006 2280 5014
rect 2288 5006 2292 5014
rect 2300 5006 2304 5014
rect 1930 4884 1942 4886
rect 1930 4876 1932 4884
rect 1940 4876 1942 4884
rect 1802 4564 1814 4566
rect 1802 4556 1804 4564
rect 1812 4556 1814 4564
rect 1802 4524 1814 4556
rect 1930 4544 1942 4876
rect 1930 4536 1932 4544
rect 1940 4536 1942 4544
rect 1930 4534 1942 4536
rect 2058 4704 2070 4706
rect 2058 4696 2060 4704
rect 2068 4696 2070 4704
rect 1802 4516 1804 4524
rect 1812 4516 1814 4524
rect 1802 4514 1814 4516
rect 2058 4304 2070 4696
rect 2240 4614 2304 5006
rect 3744 5214 3808 5216
rect 3744 5206 3748 5214
rect 3756 5206 3760 5214
rect 3768 5206 3772 5214
rect 3780 5206 3784 5214
rect 3792 5206 3796 5214
rect 3804 5206 3808 5214
rect 2922 4984 2934 4986
rect 2922 4976 2924 4984
rect 2932 4976 2934 4984
rect 2240 4606 2244 4614
rect 2252 4606 2256 4614
rect 2264 4606 2268 4614
rect 2276 4606 2280 4614
rect 2288 4606 2292 4614
rect 2300 4606 2304 4614
rect 2058 4296 2060 4304
rect 2068 4296 2070 4304
rect 2058 4294 2070 4296
rect 2186 4484 2198 4486
rect 2186 4476 2188 4484
rect 2196 4476 2198 4484
rect 1930 4264 1942 4266
rect 1930 4256 1932 4264
rect 1940 4256 1942 4264
rect 1674 4076 1676 4084
rect 1684 4076 1686 4084
rect 1674 4074 1686 4076
rect 1706 4084 1718 4086
rect 1706 4076 1708 4084
rect 1716 4076 1718 4084
rect 1642 3864 1654 3866
rect 1642 3856 1644 3864
rect 1652 3856 1654 3864
rect 1642 3704 1654 3856
rect 1642 3696 1644 3704
rect 1652 3696 1654 3704
rect 1642 3694 1654 3696
rect 1642 3624 1654 3626
rect 1642 3616 1644 3624
rect 1652 3616 1654 3624
rect 1642 3584 1654 3616
rect 1642 3576 1644 3584
rect 1652 3576 1654 3584
rect 1642 3574 1654 3576
rect 1578 3556 1580 3564
rect 1588 3556 1590 3564
rect 1578 3554 1590 3556
rect 1706 3364 1718 4076
rect 1802 3904 1814 3906
rect 1802 3896 1804 3904
rect 1812 3896 1814 3904
rect 1738 3684 1750 3686
rect 1738 3676 1740 3684
rect 1748 3676 1750 3684
rect 1738 3444 1750 3676
rect 1738 3436 1740 3444
rect 1748 3436 1750 3444
rect 1738 3434 1750 3436
rect 1706 3356 1708 3364
rect 1716 3356 1718 3364
rect 1706 3354 1718 3356
rect 1482 3256 1484 3264
rect 1492 3256 1494 3264
rect 1482 3254 1494 3256
rect 1802 3204 1814 3896
rect 1802 3196 1804 3204
rect 1812 3196 1814 3204
rect 1802 3194 1814 3196
rect 1834 3704 1846 3706
rect 1834 3696 1836 3704
rect 1844 3696 1846 3704
rect 1834 3184 1846 3696
rect 1930 3704 1942 4256
rect 2090 4264 2102 4266
rect 2090 4256 2092 4264
rect 2100 4256 2102 4264
rect 2090 4124 2102 4256
rect 2090 4116 2092 4124
rect 2100 4116 2102 4124
rect 2090 4114 2102 4116
rect 2186 3864 2198 4476
rect 2186 3856 2188 3864
rect 2196 3856 2198 3864
rect 2186 3854 2198 3856
rect 2240 4214 2304 4606
rect 2346 4924 2358 4926
rect 2346 4916 2348 4924
rect 2356 4916 2358 4924
rect 2346 4884 2358 4916
rect 2346 4876 2348 4884
rect 2356 4876 2358 4884
rect 2346 4384 2358 4876
rect 2570 4584 2582 4586
rect 2570 4576 2572 4584
rect 2580 4576 2582 4584
rect 2506 4564 2518 4566
rect 2506 4556 2508 4564
rect 2516 4556 2518 4564
rect 2506 4424 2518 4556
rect 2506 4416 2508 4424
rect 2516 4416 2518 4424
rect 2506 4414 2518 4416
rect 2538 4504 2550 4506
rect 2538 4496 2540 4504
rect 2548 4496 2550 4504
rect 2346 4376 2348 4384
rect 2356 4376 2358 4384
rect 2346 4374 2358 4376
rect 2240 4206 2244 4214
rect 2252 4206 2256 4214
rect 2264 4206 2268 4214
rect 2276 4206 2280 4214
rect 2288 4206 2292 4214
rect 2300 4206 2304 4214
rect 2240 3814 2304 4206
rect 2346 4304 2358 4306
rect 2346 4296 2348 4304
rect 2356 4296 2358 4304
rect 2346 4264 2358 4296
rect 2458 4284 2486 4286
rect 2458 4276 2460 4284
rect 2468 4276 2486 4284
rect 2458 4274 2486 4276
rect 2346 4256 2348 4264
rect 2356 4256 2358 4264
rect 2346 3984 2358 4256
rect 2474 4264 2486 4274
rect 2474 4256 2476 4264
rect 2484 4256 2486 4264
rect 2474 4254 2486 4256
rect 2346 3976 2348 3984
rect 2356 3976 2358 3984
rect 2346 3974 2358 3976
rect 2538 4244 2550 4496
rect 2538 4236 2540 4244
rect 2548 4236 2550 4244
rect 2240 3806 2244 3814
rect 2252 3806 2256 3814
rect 2264 3806 2268 3814
rect 2276 3806 2280 3814
rect 2288 3806 2292 3814
rect 2300 3806 2304 3814
rect 1930 3696 1932 3704
rect 1940 3696 1942 3704
rect 1930 3694 1942 3696
rect 1962 3764 1974 3766
rect 1962 3756 1964 3764
rect 1972 3756 1974 3764
rect 1898 3424 1910 3426
rect 1898 3416 1900 3424
rect 1908 3416 1910 3424
rect 1898 3304 1910 3416
rect 1898 3296 1900 3304
rect 1908 3296 1910 3304
rect 1898 3294 1910 3296
rect 1834 3176 1836 3184
rect 1844 3176 1846 3184
rect 1834 3174 1846 3176
rect 1450 3096 1452 3104
rect 1460 3096 1462 3104
rect 1450 3094 1462 3096
rect 1930 3104 1942 3106
rect 1930 3096 1932 3104
rect 1940 3096 1942 3104
rect 1354 3076 1356 3084
rect 1364 3076 1366 3084
rect 1354 3074 1366 3076
rect 1674 3064 1686 3066
rect 1674 3056 1676 3064
rect 1684 3056 1686 3064
rect 1354 2924 1366 2926
rect 1354 2916 1356 2924
rect 1364 2916 1366 2924
rect 1194 2696 1196 2704
rect 1204 2696 1206 2704
rect 554 2236 556 2244
rect 564 2236 566 2244
rect 554 2234 566 2236
rect 736 2406 740 2414
rect 748 2406 752 2414
rect 760 2406 764 2414
rect 772 2406 776 2414
rect 784 2406 788 2414
rect 796 2406 800 2414
rect 330 1716 332 1724
rect 340 1716 342 1724
rect 330 1484 342 1716
rect 586 2084 598 2086
rect 586 2076 588 2084
rect 596 2076 598 2084
rect 330 1476 332 1484
rect 340 1476 342 1484
rect 330 1474 342 1476
rect 554 1584 566 1586
rect 554 1576 556 1584
rect 564 1576 566 1584
rect 202 1036 204 1044
rect 212 1036 214 1044
rect 202 1034 214 1036
rect 394 1004 406 1006
rect 394 996 396 1004
rect 404 996 406 1004
rect 394 904 406 996
rect 394 896 396 904
rect 404 896 406 904
rect 394 804 406 896
rect 394 796 396 804
rect 404 796 406 804
rect 394 794 406 796
rect 42 776 44 784
rect 52 776 54 784
rect 42 774 54 776
rect 554 424 566 1576
rect 586 584 598 2076
rect 586 576 588 584
rect 596 576 598 584
rect 586 574 598 576
rect 736 2014 800 2406
rect 1098 2524 1110 2526
rect 1098 2516 1100 2524
rect 1108 2516 1110 2524
rect 736 2006 740 2014
rect 748 2006 752 2014
rect 760 2006 764 2014
rect 772 2006 776 2014
rect 784 2006 788 2014
rect 796 2006 800 2014
rect 736 1614 800 2006
rect 736 1606 740 1614
rect 748 1606 752 1614
rect 760 1606 764 1614
rect 772 1606 776 1614
rect 784 1606 788 1614
rect 796 1606 800 1614
rect 736 1214 800 1606
rect 736 1206 740 1214
rect 748 1206 752 1214
rect 760 1206 764 1214
rect 772 1206 776 1214
rect 784 1206 788 1214
rect 796 1206 800 1214
rect 736 814 800 1206
rect 874 2324 886 2326
rect 874 2316 876 2324
rect 884 2316 886 2324
rect 874 1104 886 2316
rect 1098 2204 1110 2516
rect 1098 2196 1100 2204
rect 1108 2196 1110 2204
rect 1098 2194 1110 2196
rect 1194 2164 1206 2696
rect 1290 2724 1302 2726
rect 1290 2716 1292 2724
rect 1300 2716 1302 2724
rect 1290 2264 1302 2716
rect 1354 2664 1366 2916
rect 1354 2656 1356 2664
rect 1364 2656 1366 2664
rect 1354 2654 1366 2656
rect 1450 2744 1462 2746
rect 1450 2736 1452 2744
rect 1460 2736 1462 2744
rect 1418 2624 1430 2626
rect 1418 2616 1420 2624
rect 1428 2616 1430 2624
rect 1290 2256 1292 2264
rect 1300 2256 1302 2264
rect 1290 2254 1302 2256
rect 1354 2604 1366 2606
rect 1354 2596 1356 2604
rect 1364 2596 1366 2604
rect 1194 2156 1196 2164
rect 1204 2156 1206 2164
rect 1194 2154 1206 2156
rect 1066 2124 1078 2126
rect 1066 2116 1068 2124
rect 1076 2116 1078 2124
rect 1066 1884 1078 2116
rect 1354 2124 1366 2596
rect 1418 2564 1430 2616
rect 1418 2556 1420 2564
rect 1428 2556 1430 2564
rect 1418 2554 1430 2556
rect 1450 2504 1462 2736
rect 1514 2724 1526 2726
rect 1514 2716 1516 2724
rect 1524 2716 1526 2724
rect 1514 2544 1526 2716
rect 1674 2564 1686 3056
rect 1770 2964 1782 2966
rect 1770 2956 1772 2964
rect 1780 2956 1782 2964
rect 1770 2704 1782 2956
rect 1930 2964 1942 3096
rect 1962 3064 1974 3756
rect 2090 3544 2102 3546
rect 2090 3536 2092 3544
rect 2100 3536 2102 3544
rect 1962 3056 1964 3064
rect 1972 3056 1974 3064
rect 1962 3054 1974 3056
rect 2026 3204 2038 3206
rect 2026 3196 2028 3204
rect 2036 3196 2038 3204
rect 1930 2956 1932 2964
rect 1940 2956 1942 2964
rect 1930 2954 1942 2956
rect 1962 2864 1974 2866
rect 1962 2856 1964 2864
rect 1972 2856 1974 2864
rect 1770 2696 1772 2704
rect 1780 2696 1782 2704
rect 1770 2694 1782 2696
rect 1834 2704 1846 2706
rect 1834 2696 1836 2704
rect 1844 2696 1846 2704
rect 1674 2556 1676 2564
rect 1684 2556 1686 2564
rect 1674 2554 1686 2556
rect 1770 2604 1782 2606
rect 1770 2596 1772 2604
rect 1780 2596 1782 2604
rect 1514 2536 1516 2544
rect 1524 2536 1526 2544
rect 1514 2534 1526 2536
rect 1450 2496 1452 2504
rect 1460 2496 1462 2504
rect 1450 2494 1462 2496
rect 1770 2444 1782 2596
rect 1770 2436 1772 2444
rect 1780 2436 1782 2444
rect 1770 2434 1782 2436
rect 1802 2404 1814 2406
rect 1802 2396 1804 2404
rect 1812 2396 1814 2404
rect 1802 2284 1814 2396
rect 1802 2276 1804 2284
rect 1812 2276 1814 2284
rect 1802 2274 1814 2276
rect 1354 2116 1356 2124
rect 1364 2116 1366 2124
rect 1354 2114 1366 2116
rect 1482 2184 1494 2186
rect 1482 2176 1484 2184
rect 1492 2176 1494 2184
rect 1386 2104 1398 2106
rect 1386 2096 1388 2104
rect 1396 2096 1398 2104
rect 1258 1964 1270 1966
rect 1258 1956 1260 1964
rect 1268 1956 1270 1964
rect 1258 1926 1270 1956
rect 1258 1924 1318 1926
rect 1258 1916 1308 1924
rect 1316 1916 1318 1924
rect 1258 1914 1318 1916
rect 1066 1876 1068 1884
rect 1076 1876 1078 1884
rect 906 1824 918 1826
rect 906 1816 908 1824
rect 916 1816 918 1824
rect 906 1344 918 1816
rect 1002 1764 1014 1766
rect 1002 1756 1004 1764
rect 1012 1756 1014 1764
rect 1002 1704 1014 1756
rect 1066 1724 1078 1876
rect 1066 1716 1068 1724
rect 1076 1716 1078 1724
rect 1066 1714 1078 1716
rect 1098 1864 1110 1866
rect 1098 1856 1100 1864
rect 1108 1856 1110 1864
rect 1002 1696 1004 1704
rect 1012 1696 1014 1704
rect 1002 1694 1014 1696
rect 1098 1444 1110 1856
rect 1354 1844 1366 1846
rect 1354 1836 1356 1844
rect 1364 1836 1366 1844
rect 1290 1744 1302 1746
rect 1290 1736 1292 1744
rect 1300 1736 1302 1744
rect 1098 1436 1100 1444
rect 1108 1436 1110 1444
rect 1098 1434 1110 1436
rect 1130 1704 1142 1706
rect 1130 1696 1132 1704
rect 1140 1696 1142 1704
rect 906 1336 908 1344
rect 916 1336 918 1344
rect 906 1334 918 1336
rect 1098 1384 1110 1386
rect 1098 1376 1100 1384
rect 1108 1376 1110 1384
rect 874 1096 876 1104
rect 884 1096 886 1104
rect 874 984 886 1096
rect 1098 1104 1110 1376
rect 1130 1344 1142 1696
rect 1130 1336 1132 1344
rect 1140 1336 1142 1344
rect 1130 1334 1142 1336
rect 1226 1404 1238 1406
rect 1226 1396 1228 1404
rect 1236 1396 1238 1404
rect 1226 1124 1238 1396
rect 1290 1304 1302 1736
rect 1354 1664 1366 1836
rect 1354 1656 1356 1664
rect 1364 1656 1366 1664
rect 1354 1654 1366 1656
rect 1386 1564 1398 2096
rect 1482 1844 1494 2176
rect 1738 2184 1750 2186
rect 1738 2176 1740 2184
rect 1748 2176 1750 2184
rect 1738 2064 1750 2176
rect 1738 2056 1740 2064
rect 1748 2056 1750 2064
rect 1738 2054 1750 2056
rect 1482 1836 1484 1844
rect 1492 1836 1494 1844
rect 1482 1834 1494 1836
rect 1514 2044 1526 2046
rect 1514 2036 1516 2044
rect 1524 2036 1526 2044
rect 1514 1744 1526 2036
rect 1770 2004 1782 2006
rect 1770 1996 1772 2004
rect 1780 1996 1782 2004
rect 1514 1736 1516 1744
rect 1524 1736 1526 1744
rect 1514 1734 1526 1736
rect 1578 1924 1590 1926
rect 1578 1916 1580 1924
rect 1588 1916 1590 1924
rect 1386 1556 1388 1564
rect 1396 1556 1398 1564
rect 1386 1554 1398 1556
rect 1578 1564 1590 1916
rect 1578 1556 1580 1564
rect 1588 1556 1590 1564
rect 1290 1296 1292 1304
rect 1300 1296 1302 1304
rect 1290 1294 1302 1296
rect 1514 1524 1526 1526
rect 1514 1516 1516 1524
rect 1524 1516 1526 1524
rect 1226 1116 1228 1124
rect 1236 1116 1238 1124
rect 1226 1114 1238 1116
rect 1098 1096 1100 1104
rect 1108 1096 1110 1104
rect 1098 1094 1110 1096
rect 874 976 876 984
rect 884 976 886 984
rect 874 974 886 976
rect 736 806 740 814
rect 748 806 752 814
rect 760 806 764 814
rect 772 806 776 814
rect 784 806 788 814
rect 796 806 800 814
rect 554 416 556 424
rect 564 416 566 424
rect 554 414 566 416
rect 736 414 800 806
rect 1194 904 1206 906
rect 1194 896 1196 904
rect 1204 896 1206 904
rect 736 406 740 414
rect 748 406 752 414
rect 760 406 764 414
rect 772 406 776 414
rect 784 406 788 414
rect 796 406 800 414
rect 736 14 800 406
rect 906 584 918 586
rect 906 576 908 584
rect 916 576 918 584
rect 906 324 918 576
rect 906 316 908 324
rect 916 316 918 324
rect 906 314 918 316
rect 1162 304 1174 306
rect 1162 296 1164 304
rect 1172 296 1174 304
rect 1162 244 1174 296
rect 1162 236 1164 244
rect 1172 236 1174 244
rect 1162 234 1174 236
rect 1194 44 1206 896
rect 1514 884 1526 1516
rect 1578 1364 1590 1556
rect 1578 1356 1580 1364
rect 1588 1356 1590 1364
rect 1578 1354 1590 1356
rect 1642 1924 1654 1926
rect 1642 1916 1644 1924
rect 1652 1916 1654 1924
rect 1642 1504 1654 1916
rect 1770 1624 1782 1996
rect 1770 1616 1772 1624
rect 1780 1616 1782 1624
rect 1770 1614 1782 1616
rect 1802 1904 1814 1906
rect 1802 1896 1804 1904
rect 1812 1896 1814 1904
rect 1642 1496 1644 1504
rect 1652 1496 1654 1504
rect 1514 876 1516 884
rect 1524 876 1526 884
rect 1514 874 1526 876
rect 1546 1184 1558 1186
rect 1546 1176 1548 1184
rect 1556 1176 1558 1184
rect 1546 724 1558 1176
rect 1642 924 1654 1496
rect 1802 1504 1814 1896
rect 1802 1496 1804 1504
rect 1812 1496 1814 1504
rect 1802 1494 1814 1496
rect 1834 1724 1846 2696
rect 1930 2564 1942 2566
rect 1930 2556 1932 2564
rect 1940 2556 1942 2564
rect 1898 2284 1910 2286
rect 1898 2276 1900 2284
rect 1908 2276 1910 2284
rect 1898 2204 1910 2276
rect 1898 2196 1900 2204
rect 1908 2196 1910 2204
rect 1898 2194 1910 2196
rect 1930 2004 1942 2556
rect 1962 2424 1974 2856
rect 1962 2416 1964 2424
rect 1972 2416 1974 2424
rect 1962 2414 1974 2416
rect 1994 2424 2006 2426
rect 1994 2416 1996 2424
rect 2004 2416 2006 2424
rect 1994 2384 2006 2416
rect 1994 2376 1996 2384
rect 2004 2376 2006 2384
rect 1994 2374 2006 2376
rect 2026 2384 2038 3196
rect 2058 3004 2070 3006
rect 2058 2996 2060 3004
rect 2068 2996 2070 3004
rect 2058 2644 2070 2996
rect 2090 3004 2102 3536
rect 2186 3464 2198 3466
rect 2186 3456 2188 3464
rect 2196 3456 2198 3464
rect 2186 3384 2198 3456
rect 2186 3376 2188 3384
rect 2196 3376 2198 3384
rect 2186 3374 2198 3376
rect 2240 3414 2304 3806
rect 2506 3904 2518 3906
rect 2506 3896 2508 3904
rect 2516 3896 2518 3904
rect 2240 3406 2244 3414
rect 2252 3406 2256 3414
rect 2264 3406 2268 3414
rect 2276 3406 2280 3414
rect 2288 3406 2292 3414
rect 2300 3406 2304 3414
rect 2090 2996 2092 3004
rect 2100 2996 2102 3004
rect 2090 2994 2102 2996
rect 2240 3014 2304 3406
rect 2240 3006 2244 3014
rect 2252 3006 2256 3014
rect 2264 3006 2268 3014
rect 2276 3006 2280 3014
rect 2288 3006 2292 3014
rect 2300 3006 2304 3014
rect 2058 2636 2060 2644
rect 2068 2636 2070 2644
rect 2058 2634 2070 2636
rect 2240 2614 2304 3006
rect 2240 2606 2244 2614
rect 2252 2606 2256 2614
rect 2264 2606 2268 2614
rect 2276 2606 2280 2614
rect 2288 2606 2292 2614
rect 2300 2606 2304 2614
rect 2026 2376 2028 2384
rect 2036 2376 2038 2384
rect 2026 2374 2038 2376
rect 2122 2524 2134 2526
rect 2122 2516 2124 2524
rect 2132 2516 2134 2524
rect 1930 1996 1932 2004
rect 1940 1996 1942 2004
rect 1930 1994 1942 1996
rect 1994 2124 2006 2126
rect 1994 2116 1996 2124
rect 2004 2116 2006 2124
rect 1962 1964 1974 1966
rect 1962 1956 1964 1964
rect 1972 1956 1974 1964
rect 1834 1716 1836 1724
rect 1844 1716 1846 1724
rect 1674 1344 1686 1346
rect 1674 1336 1676 1344
rect 1684 1336 1686 1344
rect 1674 1304 1686 1336
rect 1834 1324 1846 1716
rect 1866 1884 1878 1886
rect 1866 1876 1868 1884
rect 1876 1876 1878 1884
rect 1866 1464 1878 1876
rect 1930 1864 1942 1866
rect 1930 1856 1932 1864
rect 1940 1856 1942 1864
rect 1930 1684 1942 1856
rect 1930 1676 1932 1684
rect 1940 1676 1942 1684
rect 1930 1674 1942 1676
rect 1866 1456 1868 1464
rect 1876 1456 1878 1464
rect 1866 1454 1878 1456
rect 1930 1464 1942 1466
rect 1930 1456 1932 1464
rect 1940 1456 1942 1464
rect 1834 1316 1836 1324
rect 1844 1316 1846 1324
rect 1834 1314 1846 1316
rect 1674 1296 1676 1304
rect 1684 1296 1686 1304
rect 1674 1294 1686 1296
rect 1898 1264 1910 1266
rect 1898 1256 1900 1264
rect 1908 1256 1910 1264
rect 1802 1124 1814 1126
rect 1802 1116 1804 1124
rect 1812 1116 1814 1124
rect 1642 916 1644 924
rect 1652 916 1654 924
rect 1642 914 1654 916
rect 1674 984 1686 986
rect 1674 976 1676 984
rect 1684 976 1686 984
rect 1546 716 1548 724
rect 1556 716 1558 724
rect 1546 714 1558 716
rect 1578 904 1590 906
rect 1578 896 1580 904
rect 1588 896 1590 904
rect 1578 724 1590 896
rect 1578 716 1580 724
rect 1588 716 1590 724
rect 1578 714 1590 716
rect 1642 744 1654 746
rect 1642 736 1644 744
rect 1652 736 1654 744
rect 1642 524 1654 736
rect 1674 604 1686 976
rect 1674 596 1676 604
rect 1684 596 1686 604
rect 1674 594 1686 596
rect 1642 516 1644 524
rect 1652 516 1654 524
rect 1642 514 1654 516
rect 1802 464 1814 1116
rect 1898 824 1910 1256
rect 1930 904 1942 1456
rect 1962 1344 1974 1956
rect 1994 1464 2006 2116
rect 2026 2004 2038 2006
rect 2026 1996 2028 2004
rect 2036 1996 2038 2004
rect 2026 1704 2038 1996
rect 2026 1696 2028 1704
rect 2036 1696 2038 1704
rect 2026 1694 2038 1696
rect 2090 1924 2102 1926
rect 2090 1916 2092 1924
rect 2100 1916 2102 1924
rect 2058 1684 2070 1686
rect 2058 1676 2060 1684
rect 2068 1676 2070 1684
rect 2058 1624 2070 1676
rect 2058 1616 2060 1624
rect 2068 1616 2070 1624
rect 2058 1614 2070 1616
rect 1994 1456 1996 1464
rect 2004 1456 2006 1464
rect 1994 1424 2006 1456
rect 1994 1416 1996 1424
rect 2004 1416 2006 1424
rect 1994 1414 2006 1416
rect 1962 1336 1964 1344
rect 1972 1336 1974 1344
rect 1962 1334 1974 1336
rect 2026 1384 2038 1386
rect 2026 1376 2028 1384
rect 2036 1376 2038 1384
rect 1994 1324 2006 1326
rect 1994 1316 1996 1324
rect 2004 1316 2006 1324
rect 1962 1244 1974 1246
rect 1962 1236 1964 1244
rect 1972 1236 1974 1244
rect 1962 1124 1974 1236
rect 1962 1116 1964 1124
rect 1972 1116 1974 1124
rect 1962 1114 1974 1116
rect 1930 896 1932 904
rect 1940 896 1942 904
rect 1930 894 1942 896
rect 1898 816 1900 824
rect 1908 816 1910 824
rect 1898 814 1910 816
rect 1930 824 1942 826
rect 1930 816 1932 824
rect 1940 816 1942 824
rect 1898 784 1910 786
rect 1898 776 1900 784
rect 1908 776 1910 784
rect 1834 724 1846 726
rect 1834 716 1836 724
rect 1844 716 1846 724
rect 1834 484 1846 716
rect 1898 624 1910 776
rect 1898 616 1900 624
rect 1908 616 1910 624
rect 1898 614 1910 616
rect 1930 564 1942 816
rect 1930 556 1932 564
rect 1940 556 1942 564
rect 1930 554 1942 556
rect 1994 544 2006 1316
rect 2026 1324 2038 1376
rect 2026 1316 2028 1324
rect 2036 1316 2038 1324
rect 2026 1314 2038 1316
rect 2090 1184 2102 1916
rect 2122 1724 2134 2516
rect 2122 1716 2124 1724
rect 2132 1716 2134 1724
rect 2122 1714 2134 1716
rect 2240 2214 2304 2606
rect 2240 2206 2244 2214
rect 2252 2206 2256 2214
rect 2264 2206 2268 2214
rect 2276 2206 2280 2214
rect 2288 2206 2292 2214
rect 2300 2206 2304 2214
rect 2240 1814 2304 2206
rect 2378 3664 2390 3666
rect 2378 3656 2380 3664
rect 2388 3656 2390 3664
rect 2378 2284 2390 3656
rect 2506 3384 2518 3896
rect 2538 3844 2550 4236
rect 2570 4044 2582 4576
rect 2570 4036 2572 4044
rect 2580 4036 2582 4044
rect 2570 4034 2582 4036
rect 2602 4424 2614 4426
rect 2602 4416 2604 4424
rect 2612 4416 2614 4424
rect 2538 3836 2540 3844
rect 2548 3836 2550 3844
rect 2538 3834 2550 3836
rect 2506 3376 2508 3384
rect 2516 3376 2518 3384
rect 2506 3374 2518 3376
rect 2602 3304 2614 4416
rect 2922 3884 2934 4976
rect 3744 4814 3808 5206
rect 4682 5144 4694 5146
rect 4682 5136 4684 5144
rect 4692 5136 4694 5144
rect 3978 5104 3990 5106
rect 3978 5096 3980 5104
rect 3988 5096 3990 5104
rect 3978 4884 3990 5096
rect 3978 4876 3980 4884
rect 3988 4876 3990 4884
rect 3978 4874 3990 4876
rect 3744 4806 3748 4814
rect 3756 4806 3760 4814
rect 3768 4806 3772 4814
rect 3780 4806 3784 4814
rect 3792 4806 3796 4814
rect 3804 4806 3808 4814
rect 3626 4804 3638 4806
rect 3626 4796 3628 4804
rect 3636 4796 3638 4804
rect 3402 4704 3414 4706
rect 3402 4696 3404 4704
rect 3412 4696 3414 4704
rect 3114 4684 3126 4686
rect 3114 4676 3116 4684
rect 3124 4676 3126 4684
rect 3082 4544 3094 4546
rect 3082 4536 3084 4544
rect 3092 4536 3094 4544
rect 2922 3876 2924 3884
rect 2932 3876 2934 3884
rect 2922 3874 2934 3876
rect 3018 4184 3030 4186
rect 3018 4176 3020 4184
rect 3028 4176 3030 4184
rect 2602 3296 2604 3304
rect 2612 3296 2614 3304
rect 2602 3294 2614 3296
rect 2762 3864 2774 3866
rect 2762 3856 2764 3864
rect 2772 3856 2774 3864
rect 2698 3264 2710 3266
rect 2698 3256 2700 3264
rect 2708 3256 2710 3264
rect 2634 3204 2646 3206
rect 2634 3196 2636 3204
rect 2644 3196 2646 3204
rect 2570 2784 2582 2786
rect 2570 2776 2572 2784
rect 2580 2776 2582 2784
rect 2378 2276 2380 2284
rect 2388 2276 2390 2284
rect 2378 2204 2390 2276
rect 2378 2196 2380 2204
rect 2388 2196 2390 2204
rect 2378 2194 2390 2196
rect 2506 2504 2518 2506
rect 2506 2496 2508 2504
rect 2516 2496 2518 2504
rect 2506 2264 2518 2496
rect 2506 2256 2508 2264
rect 2516 2256 2518 2264
rect 2378 2144 2390 2146
rect 2378 2136 2380 2144
rect 2388 2136 2390 2144
rect 2240 1806 2244 1814
rect 2252 1806 2256 1814
rect 2264 1806 2268 1814
rect 2276 1806 2280 1814
rect 2288 1806 2292 1814
rect 2300 1806 2304 1814
rect 2154 1464 2166 1466
rect 2154 1456 2156 1464
rect 2164 1456 2166 1464
rect 2090 1176 2092 1184
rect 2100 1176 2102 1184
rect 2090 1174 2102 1176
rect 2122 1184 2134 1186
rect 2122 1176 2124 1184
rect 2132 1176 2134 1184
rect 2122 1024 2134 1176
rect 2122 1016 2124 1024
rect 2132 1016 2134 1024
rect 2122 1014 2134 1016
rect 2154 1024 2166 1456
rect 2240 1414 2304 1806
rect 2346 1924 2358 1926
rect 2346 1916 2348 1924
rect 2356 1916 2358 1924
rect 2346 1704 2358 1916
rect 2346 1696 2348 1704
rect 2356 1696 2358 1704
rect 2346 1694 2358 1696
rect 2346 1644 2358 1646
rect 2346 1636 2348 1644
rect 2356 1636 2358 1644
rect 2346 1484 2358 1636
rect 2346 1476 2348 1484
rect 2356 1476 2358 1484
rect 2346 1474 2358 1476
rect 2240 1406 2244 1414
rect 2252 1406 2256 1414
rect 2264 1406 2268 1414
rect 2276 1406 2280 1414
rect 2288 1406 2292 1414
rect 2300 1406 2304 1414
rect 2186 1344 2198 1346
rect 2186 1336 2188 1344
rect 2196 1336 2198 1344
rect 2186 1164 2198 1336
rect 2186 1156 2188 1164
rect 2196 1156 2198 1164
rect 2186 1154 2198 1156
rect 2154 1016 2156 1024
rect 2164 1016 2166 1024
rect 2154 1014 2166 1016
rect 2240 1014 2304 1406
rect 2240 1006 2244 1014
rect 2252 1006 2256 1014
rect 2264 1006 2268 1014
rect 2276 1006 2280 1014
rect 2288 1006 2292 1014
rect 2300 1006 2304 1014
rect 2058 944 2070 946
rect 2058 936 2060 944
rect 2068 936 2070 944
rect 2058 904 2070 936
rect 2058 896 2060 904
rect 2068 896 2070 904
rect 2058 894 2070 896
rect 1994 536 1996 544
rect 2004 536 2006 544
rect 1994 534 2006 536
rect 2186 624 2198 626
rect 2186 616 2188 624
rect 2196 616 2198 624
rect 1834 476 1836 484
rect 1844 476 1846 484
rect 1834 474 1846 476
rect 1802 456 1804 464
rect 1812 456 1814 464
rect 1802 454 1814 456
rect 1962 444 1974 446
rect 1962 436 1964 444
rect 1972 436 1974 444
rect 1642 404 1654 406
rect 1642 396 1644 404
rect 1652 396 1654 404
rect 1226 244 1238 246
rect 1226 236 1228 244
rect 1236 236 1238 244
rect 1226 64 1238 236
rect 1226 56 1228 64
rect 1236 56 1238 64
rect 1226 54 1238 56
rect 1194 36 1196 44
rect 1204 36 1206 44
rect 1194 34 1206 36
rect 1642 44 1654 396
rect 1962 384 1974 436
rect 2186 444 2198 616
rect 2186 436 2188 444
rect 2196 436 2198 444
rect 2186 404 2198 436
rect 2186 396 2188 404
rect 2196 396 2198 404
rect 2186 394 2198 396
rect 2240 614 2304 1006
rect 2378 804 2390 2136
rect 2506 2064 2518 2256
rect 2570 2224 2582 2776
rect 2634 2784 2646 3196
rect 2634 2776 2636 2784
rect 2644 2776 2646 2784
rect 2634 2774 2646 2776
rect 2666 3204 2678 3206
rect 2666 3196 2668 3204
rect 2676 3196 2678 3204
rect 2666 2704 2678 3196
rect 2666 2696 2668 2704
rect 2676 2696 2678 2704
rect 2666 2694 2678 2696
rect 2666 2624 2678 2626
rect 2666 2616 2668 2624
rect 2676 2616 2678 2624
rect 2570 2216 2572 2224
rect 2580 2216 2582 2224
rect 2570 2214 2582 2216
rect 2634 2504 2646 2506
rect 2634 2496 2636 2504
rect 2644 2496 2646 2504
rect 2634 2144 2646 2496
rect 2634 2136 2636 2144
rect 2644 2136 2646 2144
rect 2634 2134 2646 2136
rect 2666 2104 2678 2616
rect 2698 2544 2710 3256
rect 2698 2536 2700 2544
rect 2708 2536 2710 2544
rect 2698 2534 2710 2536
rect 2666 2096 2668 2104
rect 2676 2096 2678 2104
rect 2666 2094 2678 2096
rect 2698 2504 2710 2506
rect 2698 2496 2700 2504
rect 2708 2496 2710 2504
rect 2698 2464 2710 2496
rect 2698 2456 2700 2464
rect 2708 2456 2710 2464
rect 2698 2104 2710 2456
rect 2698 2096 2700 2104
rect 2708 2096 2710 2104
rect 2698 2094 2710 2096
rect 2506 2056 2508 2064
rect 2516 2056 2518 2064
rect 2506 2054 2518 2056
rect 2762 2004 2774 3856
rect 2858 3444 2870 3446
rect 2858 3436 2860 3444
rect 2868 3436 2870 3444
rect 2858 3304 2870 3436
rect 2858 3296 2860 3304
rect 2868 3296 2870 3304
rect 2858 3294 2870 3296
rect 3018 3264 3030 4176
rect 3082 4164 3094 4536
rect 3114 4444 3126 4676
rect 3114 4436 3116 4444
rect 3124 4436 3126 4444
rect 3114 4434 3126 4436
rect 3082 4156 3084 4164
rect 3092 4156 3094 4164
rect 3082 4154 3094 4156
rect 3178 4324 3190 4326
rect 3178 4316 3180 4324
rect 3188 4316 3190 4324
rect 3146 4104 3158 4106
rect 3146 4096 3148 4104
rect 3156 4096 3158 4104
rect 3018 3256 3020 3264
rect 3028 3256 3030 3264
rect 3018 3254 3030 3256
rect 3082 3524 3094 3526
rect 3082 3516 3084 3524
rect 3092 3516 3094 3524
rect 2922 3184 2934 3186
rect 2922 3176 2924 3184
rect 2932 3176 2934 3184
rect 2890 3144 2902 3146
rect 2890 3136 2892 3144
rect 2900 3136 2902 3144
rect 2794 3084 2806 3086
rect 2794 3076 2796 3084
rect 2804 3076 2806 3084
rect 2794 2124 2806 3076
rect 2858 2964 2870 2966
rect 2858 2956 2860 2964
rect 2868 2956 2870 2964
rect 2858 2344 2870 2956
rect 2858 2336 2860 2344
rect 2868 2336 2870 2344
rect 2858 2334 2870 2336
rect 2890 2144 2902 3136
rect 2922 2804 2934 3176
rect 3082 2904 3094 3516
rect 3146 3084 3158 4096
rect 3178 3724 3190 4316
rect 3274 4184 3286 4186
rect 3274 4176 3276 4184
rect 3284 4176 3286 4184
rect 3274 3744 3286 4176
rect 3402 4044 3414 4696
rect 3402 4036 3404 4044
rect 3412 4036 3414 4044
rect 3274 3736 3276 3744
rect 3284 3736 3286 3744
rect 3274 3734 3286 3736
rect 3306 3824 3318 3826
rect 3306 3816 3308 3824
rect 3316 3816 3318 3824
rect 3178 3716 3180 3724
rect 3188 3716 3190 3724
rect 3178 3714 3190 3716
rect 3146 3076 3148 3084
rect 3156 3076 3158 3084
rect 3146 3074 3158 3076
rect 3178 3484 3190 3486
rect 3178 3476 3180 3484
rect 3188 3476 3190 3484
rect 3082 2896 3084 2904
rect 3092 2896 3094 2904
rect 3082 2894 3094 2896
rect 2922 2796 2924 2804
rect 2932 2796 2934 2804
rect 2922 2794 2934 2796
rect 3114 2584 3126 2586
rect 3114 2576 3116 2584
rect 3124 2576 3126 2584
rect 2890 2136 2892 2144
rect 2900 2136 2902 2144
rect 2890 2134 2902 2136
rect 3050 2544 3062 2546
rect 3050 2536 3052 2544
rect 3060 2536 3062 2544
rect 2794 2116 2796 2124
rect 2804 2116 2806 2124
rect 2794 2114 2806 2116
rect 3050 2124 3062 2536
rect 3050 2116 3052 2124
rect 3060 2116 3062 2124
rect 3050 2114 3062 2116
rect 2762 1996 2764 2004
rect 2772 1996 2774 2004
rect 2762 1994 2774 1996
rect 2858 1944 2870 1946
rect 2858 1936 2860 1944
rect 2868 1936 2870 1944
rect 2602 1864 2614 1866
rect 2602 1856 2604 1864
rect 2612 1856 2614 1864
rect 2442 1744 2454 1746
rect 2442 1736 2444 1744
rect 2452 1736 2454 1744
rect 2410 1344 2422 1346
rect 2410 1336 2412 1344
rect 2420 1336 2422 1344
rect 2410 1024 2422 1336
rect 2410 1016 2412 1024
rect 2420 1016 2422 1024
rect 2410 1014 2422 1016
rect 2442 1024 2454 1736
rect 2570 1744 2582 1746
rect 2570 1736 2572 1744
rect 2580 1736 2582 1744
rect 2506 1244 2518 1246
rect 2506 1236 2508 1244
rect 2516 1236 2518 1244
rect 2506 1184 2518 1236
rect 2506 1176 2508 1184
rect 2516 1176 2518 1184
rect 2506 1174 2518 1176
rect 2442 1016 2444 1024
rect 2452 1016 2454 1024
rect 2442 1014 2454 1016
rect 2474 1104 2486 1106
rect 2474 1096 2476 1104
rect 2484 1096 2486 1104
rect 2474 984 2486 1096
rect 2474 976 2476 984
rect 2484 976 2486 984
rect 2474 974 2486 976
rect 2378 796 2380 804
rect 2388 796 2390 804
rect 2378 794 2390 796
rect 2240 606 2244 614
rect 2252 606 2256 614
rect 2264 606 2268 614
rect 2276 606 2280 614
rect 2288 606 2292 614
rect 2300 606 2304 614
rect 1962 376 1964 384
rect 1972 376 1974 384
rect 1962 374 1974 376
rect 1738 364 1750 366
rect 1738 356 1740 364
rect 1748 356 1750 364
rect 1738 324 1750 356
rect 1738 316 1740 324
rect 1748 316 1750 324
rect 1738 314 1750 316
rect 1642 36 1644 44
rect 1652 36 1654 44
rect 1642 34 1654 36
rect 2240 214 2304 606
rect 2570 684 2582 1736
rect 2602 1224 2614 1856
rect 2762 1784 2774 1786
rect 2762 1776 2764 1784
rect 2772 1776 2774 1784
rect 2762 1766 2774 1776
rect 2762 1764 2790 1766
rect 2762 1756 2780 1764
rect 2788 1756 2790 1764
rect 2762 1754 2790 1756
rect 2762 1724 2774 1726
rect 2762 1716 2764 1724
rect 2772 1716 2774 1724
rect 2602 1216 2604 1224
rect 2612 1216 2614 1224
rect 2602 1214 2614 1216
rect 2730 1564 2742 1566
rect 2730 1556 2732 1564
rect 2740 1556 2742 1564
rect 2730 1184 2742 1556
rect 2762 1424 2774 1716
rect 2858 1724 2870 1936
rect 2858 1716 2860 1724
rect 2868 1716 2870 1724
rect 2858 1714 2870 1716
rect 3050 1884 3062 1886
rect 3050 1876 3052 1884
rect 3060 1876 3062 1884
rect 2762 1416 2764 1424
rect 2772 1416 2774 1424
rect 2762 1414 2774 1416
rect 3018 1424 3030 1426
rect 3018 1416 3020 1424
rect 3028 1416 3030 1424
rect 2730 1176 2732 1184
rect 2740 1176 2742 1184
rect 2730 1174 2742 1176
rect 2890 1104 2902 1106
rect 2890 1096 2892 1104
rect 2900 1096 2902 1104
rect 2858 1024 2870 1026
rect 2858 1016 2860 1024
rect 2868 1016 2870 1024
rect 2570 676 2572 684
rect 2580 676 2582 684
rect 2570 564 2582 676
rect 2570 556 2572 564
rect 2580 556 2582 564
rect 2570 554 2582 556
rect 2826 824 2838 826
rect 2826 816 2828 824
rect 2836 816 2838 824
rect 2240 206 2244 214
rect 2252 206 2256 214
rect 2264 206 2268 214
rect 2276 206 2280 214
rect 2288 206 2292 214
rect 2300 206 2304 214
rect 736 6 740 14
rect 748 6 752 14
rect 760 6 764 14
rect 772 6 776 14
rect 784 6 788 14
rect 796 6 800 14
rect 736 -10 800 6
rect 2240 -10 2304 206
rect 2730 344 2742 346
rect 2730 336 2732 344
rect 2740 336 2742 344
rect 2730 184 2742 336
rect 2826 324 2838 816
rect 2826 316 2828 324
rect 2836 316 2838 324
rect 2826 314 2838 316
rect 2858 284 2870 1016
rect 2890 804 2902 1096
rect 3018 1024 3030 1416
rect 3050 1384 3062 1876
rect 3050 1376 3052 1384
rect 3060 1376 3062 1384
rect 3050 1374 3062 1376
rect 3018 1016 3020 1024
rect 3028 1016 3030 1024
rect 3018 1014 3030 1016
rect 3082 1084 3094 1086
rect 3082 1076 3084 1084
rect 3092 1076 3094 1084
rect 3050 984 3062 986
rect 3050 976 3052 984
rect 3060 976 3062 984
rect 3050 944 3062 976
rect 3050 936 3052 944
rect 3060 936 3062 944
rect 3050 934 3062 936
rect 2890 796 2892 804
rect 2900 796 2902 804
rect 2890 794 2902 796
rect 3050 904 3062 906
rect 3050 896 3052 904
rect 3060 896 3062 904
rect 3050 344 3062 896
rect 3082 884 3094 1076
rect 3082 876 3084 884
rect 3092 876 3094 884
rect 3082 874 3094 876
rect 3114 884 3126 2576
rect 3146 2544 3158 2546
rect 3146 2536 3148 2544
rect 3156 2536 3158 2544
rect 3146 2144 3158 2536
rect 3146 2136 3148 2144
rect 3156 2136 3158 2144
rect 3146 2134 3158 2136
rect 3178 1864 3190 3476
rect 3210 3404 3222 3406
rect 3210 3396 3212 3404
rect 3220 3396 3222 3404
rect 3210 2604 3222 3396
rect 3306 3364 3318 3816
rect 3306 3356 3308 3364
rect 3316 3356 3318 3364
rect 3306 3354 3318 3356
rect 3402 3324 3414 4036
rect 3562 4104 3574 4106
rect 3562 4096 3564 4104
rect 3572 4096 3574 4104
rect 3562 3804 3574 4096
rect 3562 3796 3564 3804
rect 3572 3796 3574 3804
rect 3562 3794 3574 3796
rect 3626 3764 3638 4796
rect 3744 4414 3808 4806
rect 4362 4784 4374 4786
rect 4362 4776 4364 4784
rect 4372 4776 4374 4784
rect 3744 4406 3748 4414
rect 3756 4406 3760 4414
rect 3768 4406 3772 4414
rect 3780 4406 3784 4414
rect 3792 4406 3796 4414
rect 3804 4406 3808 4414
rect 3690 4124 3702 4126
rect 3690 4116 3692 4124
rect 3700 4116 3702 4124
rect 3626 3756 3628 3764
rect 3636 3756 3638 3764
rect 3626 3754 3638 3756
rect 3658 3764 3670 3766
rect 3658 3756 3660 3764
rect 3668 3756 3670 3764
rect 3402 3316 3404 3324
rect 3412 3316 3414 3324
rect 3402 3314 3414 3316
rect 3434 3604 3446 3606
rect 3434 3596 3436 3604
rect 3444 3596 3446 3604
rect 3338 3204 3350 3206
rect 3338 3196 3340 3204
rect 3348 3196 3350 3204
rect 3338 2984 3350 3196
rect 3338 2976 3340 2984
rect 3348 2976 3350 2984
rect 3338 2974 3350 2976
rect 3370 3084 3382 3086
rect 3370 3076 3372 3084
rect 3380 3076 3382 3084
rect 3370 2624 3382 3076
rect 3434 2724 3446 3596
rect 3498 3124 3510 3126
rect 3498 3116 3500 3124
rect 3508 3116 3510 3124
rect 3466 2964 3478 2966
rect 3466 2956 3468 2964
rect 3476 2956 3478 2964
rect 3466 2844 3478 2956
rect 3466 2836 3468 2844
rect 3476 2836 3478 2844
rect 3466 2834 3478 2836
rect 3498 2844 3510 3116
rect 3626 3044 3638 3046
rect 3626 3036 3628 3044
rect 3636 3036 3638 3044
rect 3626 2984 3638 3036
rect 3626 2976 3628 2984
rect 3636 2976 3638 2984
rect 3626 2974 3638 2976
rect 3658 2944 3670 3756
rect 3658 2936 3660 2944
rect 3668 2936 3670 2944
rect 3658 2934 3670 2936
rect 3498 2836 3500 2844
rect 3508 2836 3510 2844
rect 3498 2834 3510 2836
rect 3434 2716 3436 2724
rect 3444 2716 3446 2724
rect 3434 2714 3446 2716
rect 3690 2704 3702 4116
rect 3690 2696 3692 2704
rect 3700 2696 3702 2704
rect 3370 2616 3372 2624
rect 3380 2616 3382 2624
rect 3370 2614 3382 2616
rect 3466 2644 3478 2646
rect 3466 2636 3468 2644
rect 3476 2636 3478 2644
rect 3210 2596 3212 2604
rect 3220 2596 3222 2604
rect 3210 2594 3222 2596
rect 3274 2384 3286 2386
rect 3274 2376 3276 2384
rect 3284 2376 3286 2384
rect 3178 1856 3180 1864
rect 3188 1856 3190 1864
rect 3178 1854 3190 1856
rect 3210 2204 3222 2206
rect 3210 2196 3212 2204
rect 3220 2196 3222 2204
rect 3210 1604 3222 2196
rect 3242 1904 3254 1906
rect 3242 1896 3244 1904
rect 3252 1896 3254 1904
rect 3242 1764 3254 1896
rect 3242 1756 3244 1764
rect 3252 1756 3254 1764
rect 3242 1754 3254 1756
rect 3274 1704 3286 2376
rect 3466 2384 3478 2636
rect 3466 2376 3468 2384
rect 3476 2376 3478 2384
rect 3466 2374 3478 2376
rect 3594 2504 3606 2506
rect 3594 2496 3596 2504
rect 3604 2496 3606 2504
rect 3466 2344 3478 2346
rect 3466 2336 3468 2344
rect 3476 2336 3478 2344
rect 3434 2324 3446 2326
rect 3434 2316 3436 2324
rect 3444 2316 3446 2324
rect 3306 2284 3318 2286
rect 3306 2276 3308 2284
rect 3316 2276 3318 2284
rect 3306 2064 3318 2276
rect 3306 2056 3308 2064
rect 3316 2056 3318 2064
rect 3306 2054 3318 2056
rect 3402 2024 3414 2026
rect 3402 2016 3404 2024
rect 3412 2016 3414 2024
rect 3274 1696 3276 1704
rect 3284 1696 3286 1704
rect 3274 1694 3286 1696
rect 3306 1884 3318 1886
rect 3306 1876 3308 1884
rect 3316 1876 3318 1884
rect 3306 1644 3318 1876
rect 3402 1724 3414 2016
rect 3434 1984 3446 2316
rect 3434 1976 3436 1984
rect 3444 1976 3446 1984
rect 3434 1974 3446 1976
rect 3466 1944 3478 2336
rect 3530 2184 3542 2186
rect 3530 2176 3532 2184
rect 3540 2176 3542 2184
rect 3530 2144 3542 2176
rect 3530 2136 3532 2144
rect 3540 2136 3542 2144
rect 3530 2134 3542 2136
rect 3594 2104 3606 2496
rect 3690 2444 3702 2696
rect 3690 2436 3692 2444
rect 3700 2436 3702 2444
rect 3690 2434 3702 2436
rect 3744 4014 3808 4406
rect 3744 4006 3748 4014
rect 3756 4006 3760 4014
rect 3768 4006 3772 4014
rect 3780 4006 3784 4014
rect 3792 4006 3796 4014
rect 3804 4006 3808 4014
rect 3744 3614 3808 4006
rect 3946 4764 3958 4766
rect 3946 4756 3948 4764
rect 3956 4756 3958 4764
rect 3744 3606 3748 3614
rect 3756 3606 3760 3614
rect 3768 3606 3772 3614
rect 3780 3606 3784 3614
rect 3792 3606 3796 3614
rect 3804 3606 3808 3614
rect 3744 3214 3808 3606
rect 3744 3206 3748 3214
rect 3756 3206 3760 3214
rect 3768 3206 3772 3214
rect 3780 3206 3784 3214
rect 3792 3206 3796 3214
rect 3804 3206 3808 3214
rect 3744 2814 3808 3206
rect 3744 2806 3748 2814
rect 3756 2806 3760 2814
rect 3768 2806 3772 2814
rect 3780 2806 3784 2814
rect 3792 2806 3796 2814
rect 3804 2806 3808 2814
rect 3744 2414 3808 2806
rect 3744 2406 3748 2414
rect 3756 2406 3760 2414
rect 3768 2406 3772 2414
rect 3780 2406 3784 2414
rect 3792 2406 3796 2414
rect 3804 2406 3808 2414
rect 3626 2404 3638 2406
rect 3626 2396 3628 2404
rect 3636 2396 3638 2404
rect 3626 2124 3638 2396
rect 3626 2116 3628 2124
rect 3636 2116 3638 2124
rect 3626 2114 3638 2116
rect 3658 2224 3670 2226
rect 3658 2216 3660 2224
rect 3668 2216 3670 2224
rect 3594 2096 3596 2104
rect 3604 2096 3606 2104
rect 3594 2094 3606 2096
rect 3466 1936 3468 1944
rect 3476 1936 3478 1944
rect 3466 1934 3478 1936
rect 3562 2084 3574 2086
rect 3562 2076 3564 2084
rect 3572 2076 3574 2084
rect 3402 1716 3404 1724
rect 3412 1716 3414 1724
rect 3402 1714 3414 1716
rect 3306 1636 3308 1644
rect 3316 1636 3318 1644
rect 3306 1634 3318 1636
rect 3210 1596 3212 1604
rect 3220 1596 3222 1604
rect 3210 1594 3222 1596
rect 3530 1584 3542 1586
rect 3530 1576 3532 1584
rect 3540 1576 3542 1584
rect 3242 1504 3254 1506
rect 3242 1496 3244 1504
rect 3252 1496 3254 1504
rect 3210 1324 3222 1326
rect 3210 1316 3212 1324
rect 3220 1316 3222 1324
rect 3210 1284 3222 1316
rect 3210 1276 3212 1284
rect 3220 1276 3222 1284
rect 3210 1274 3222 1276
rect 3242 904 3254 1496
rect 3338 1484 3350 1486
rect 3338 1476 3340 1484
rect 3348 1476 3350 1484
rect 3274 1404 3286 1406
rect 3274 1396 3276 1404
rect 3284 1396 3286 1404
rect 3274 1264 3286 1396
rect 3274 1256 3276 1264
rect 3284 1256 3286 1264
rect 3274 1254 3286 1256
rect 3306 1144 3318 1146
rect 3306 1136 3308 1144
rect 3316 1136 3318 1144
rect 3306 984 3318 1136
rect 3306 976 3308 984
rect 3316 976 3318 984
rect 3306 974 3318 976
rect 3242 896 3244 904
rect 3252 896 3254 904
rect 3242 894 3254 896
rect 3114 876 3116 884
rect 3124 876 3126 884
rect 3082 724 3094 726
rect 3082 716 3084 724
rect 3092 716 3094 724
rect 3082 624 3094 716
rect 3082 616 3084 624
rect 3092 616 3094 624
rect 3082 614 3094 616
rect 3114 364 3126 876
rect 3306 844 3318 846
rect 3306 836 3308 844
rect 3316 836 3318 844
rect 3242 784 3254 786
rect 3242 776 3244 784
rect 3252 776 3254 784
rect 3242 584 3254 776
rect 3306 624 3318 836
rect 3338 824 3350 1476
rect 3402 1364 3414 1366
rect 3402 1356 3404 1364
rect 3412 1356 3414 1364
rect 3370 1224 3382 1226
rect 3370 1216 3372 1224
rect 3380 1216 3382 1224
rect 3370 1044 3382 1216
rect 3370 1036 3372 1044
rect 3380 1036 3382 1044
rect 3370 1034 3382 1036
rect 3338 816 3340 824
rect 3348 816 3350 824
rect 3338 814 3350 816
rect 3402 744 3414 1356
rect 3530 1044 3542 1576
rect 3562 1084 3574 2076
rect 3594 1984 3606 1986
rect 3594 1976 3596 1984
rect 3604 1976 3606 1984
rect 3594 1684 3606 1976
rect 3594 1676 3596 1684
rect 3604 1676 3606 1684
rect 3594 1674 3606 1676
rect 3658 1864 3670 2216
rect 3658 1856 3660 1864
rect 3668 1856 3670 1864
rect 3626 1584 3638 1586
rect 3626 1576 3628 1584
rect 3636 1576 3638 1584
rect 3626 1364 3638 1576
rect 3658 1464 3670 1856
rect 3658 1456 3660 1464
rect 3668 1456 3670 1464
rect 3658 1454 3670 1456
rect 3744 2014 3808 2406
rect 3744 2006 3748 2014
rect 3756 2006 3760 2014
rect 3768 2006 3772 2014
rect 3780 2006 3784 2014
rect 3792 2006 3796 2014
rect 3804 2006 3808 2014
rect 3744 1614 3808 2006
rect 3744 1606 3748 1614
rect 3756 1606 3760 1614
rect 3768 1606 3772 1614
rect 3780 1606 3784 1614
rect 3792 1606 3796 1614
rect 3804 1606 3808 1614
rect 3626 1356 3628 1364
rect 3636 1356 3638 1364
rect 3626 1354 3638 1356
rect 3690 1244 3702 1246
rect 3690 1236 3692 1244
rect 3700 1236 3702 1244
rect 3562 1076 3564 1084
rect 3572 1076 3574 1084
rect 3562 1074 3574 1076
rect 3626 1124 3638 1126
rect 3626 1116 3628 1124
rect 3636 1116 3638 1124
rect 3530 1036 3532 1044
rect 3540 1036 3542 1044
rect 3530 1034 3542 1036
rect 3498 984 3510 986
rect 3498 976 3500 984
rect 3508 976 3510 984
rect 3498 904 3510 976
rect 3498 896 3500 904
rect 3508 896 3510 904
rect 3498 894 3510 896
rect 3562 964 3574 966
rect 3562 956 3564 964
rect 3572 956 3574 964
rect 3402 736 3404 744
rect 3412 736 3414 744
rect 3402 734 3414 736
rect 3562 704 3574 956
rect 3626 724 3638 1116
rect 3690 904 3702 1236
rect 3690 896 3692 904
rect 3700 896 3702 904
rect 3690 894 3702 896
rect 3744 1214 3808 1606
rect 3744 1206 3748 1214
rect 3756 1206 3760 1214
rect 3768 1206 3772 1214
rect 3780 1206 3784 1214
rect 3792 1206 3796 1214
rect 3804 1206 3808 1214
rect 3626 716 3628 724
rect 3636 716 3638 724
rect 3626 714 3638 716
rect 3744 814 3808 1206
rect 3850 3964 3862 3966
rect 3850 3956 3852 3964
rect 3860 3956 3862 3964
rect 3850 1204 3862 3956
rect 3914 3864 3926 3866
rect 3914 3856 3916 3864
rect 3924 3856 3926 3864
rect 3882 3344 3894 3346
rect 3882 3336 3884 3344
rect 3892 3336 3894 3344
rect 3882 3244 3894 3336
rect 3882 3236 3884 3244
rect 3892 3236 3894 3244
rect 3882 3234 3894 3236
rect 3882 2804 3894 2806
rect 3882 2796 3884 2804
rect 3892 2796 3894 2804
rect 3882 2584 3894 2796
rect 3882 2576 3884 2584
rect 3892 2576 3894 2584
rect 3882 2574 3894 2576
rect 3882 2244 3894 2246
rect 3882 2236 3884 2244
rect 3892 2236 3894 2244
rect 3882 1564 3894 2236
rect 3882 1556 3884 1564
rect 3892 1556 3894 1564
rect 3882 1554 3894 1556
rect 3850 1196 3852 1204
rect 3860 1196 3862 1204
rect 3850 1194 3862 1196
rect 3914 1184 3926 3856
rect 3946 3524 3958 4756
rect 4106 4724 4118 4726
rect 4106 4716 4108 4724
rect 4116 4716 4118 4724
rect 4106 4686 4118 4716
rect 4170 4714 4214 4726
rect 4170 4686 4182 4714
rect 4202 4704 4214 4714
rect 4202 4696 4204 4704
rect 4212 4696 4214 4704
rect 4202 4694 4214 4696
rect 4106 4674 4182 4686
rect 4362 4284 4374 4776
rect 4586 4744 4598 4746
rect 4586 4736 4588 4744
rect 4596 4736 4598 4744
rect 4586 4524 4598 4736
rect 4586 4516 4588 4524
rect 4596 4516 4598 4524
rect 4586 4514 4598 4516
rect 4362 4276 4364 4284
rect 4372 4276 4374 4284
rect 4362 4274 4374 4276
rect 4426 4424 4438 4426
rect 4426 4416 4428 4424
rect 4436 4416 4438 4424
rect 4010 4164 4022 4166
rect 4010 4156 4012 4164
rect 4020 4156 4022 4164
rect 4010 3624 4022 4156
rect 4426 3924 4438 4416
rect 4682 4324 4694 5136
rect 4714 5064 4726 5066
rect 4714 5056 4716 5064
rect 4724 5056 4726 5064
rect 4714 4624 4726 5056
rect 4746 4764 4758 5216
rect 5002 5084 5014 5086
rect 5002 5076 5004 5084
rect 5012 5076 5014 5084
rect 4746 4756 4748 4764
rect 4756 4756 4758 4764
rect 4746 4754 4758 4756
rect 4906 4864 4918 4866
rect 4906 4856 4908 4864
rect 4916 4856 4918 4864
rect 4714 4616 4716 4624
rect 4724 4616 4726 4624
rect 4714 4614 4726 4616
rect 4746 4724 4758 4726
rect 4746 4716 4748 4724
rect 4756 4716 4758 4724
rect 4746 4364 4758 4716
rect 4778 4704 4790 4706
rect 4778 4696 4780 4704
rect 4788 4696 4790 4704
rect 4778 4504 4790 4696
rect 4778 4496 4780 4504
rect 4788 4496 4790 4504
rect 4778 4494 4790 4496
rect 4746 4356 4748 4364
rect 4756 4356 4758 4364
rect 4746 4354 4758 4356
rect 4874 4384 4886 4386
rect 4874 4376 4876 4384
rect 4884 4376 4886 4384
rect 4682 4316 4684 4324
rect 4692 4316 4694 4324
rect 4682 4314 4694 4316
rect 4426 3916 4428 3924
rect 4436 3916 4438 3924
rect 4426 3914 4438 3916
rect 4458 4284 4470 4286
rect 4458 4276 4460 4284
rect 4468 4276 4470 4284
rect 4458 3904 4470 4276
rect 4458 3896 4460 3904
rect 4468 3896 4470 3904
rect 4362 3784 4374 3786
rect 4362 3776 4364 3784
rect 4372 3776 4374 3784
rect 4010 3616 4012 3624
rect 4020 3616 4022 3624
rect 4010 3614 4022 3616
rect 4138 3664 4150 3666
rect 4138 3656 4140 3664
rect 4148 3656 4150 3664
rect 3946 3516 3948 3524
rect 3956 3516 3958 3524
rect 3946 3514 3958 3516
rect 4074 3204 4086 3206
rect 4074 3196 4076 3204
rect 4084 3196 4086 3204
rect 4010 3084 4022 3086
rect 4010 3076 4012 3084
rect 4020 3076 4022 3084
rect 4010 2724 4022 3076
rect 4010 2716 4012 2724
rect 4020 2716 4022 2724
rect 4010 2714 4022 2716
rect 4010 2544 4022 2546
rect 4010 2536 4012 2544
rect 4020 2536 4022 2544
rect 3946 2524 3958 2526
rect 3946 2516 3948 2524
rect 3956 2516 3958 2524
rect 3946 1944 3958 2516
rect 3946 1936 3948 1944
rect 3956 1936 3958 1944
rect 3946 1934 3958 1936
rect 4010 1704 4022 2536
rect 4074 2164 4086 3196
rect 4106 2964 4118 2966
rect 4106 2956 4108 2964
rect 4116 2956 4118 2964
rect 4106 2524 4118 2956
rect 4106 2516 4108 2524
rect 4116 2516 4118 2524
rect 4106 2514 4118 2516
rect 4074 2156 4076 2164
rect 4084 2156 4086 2164
rect 4074 2154 4086 2156
rect 4074 1964 4086 1966
rect 4074 1956 4076 1964
rect 4084 1956 4086 1964
rect 4074 1804 4086 1956
rect 4074 1796 4076 1804
rect 4084 1796 4086 1804
rect 4074 1794 4086 1796
rect 4138 1784 4150 3656
rect 4362 3524 4374 3776
rect 4458 3784 4470 3896
rect 4458 3776 4460 3784
rect 4468 3776 4470 3784
rect 4458 3774 4470 3776
rect 4490 3964 4502 3966
rect 4490 3956 4492 3964
rect 4500 3956 4502 3964
rect 4490 3764 4502 3956
rect 4874 3884 4886 4376
rect 4874 3876 4876 3884
rect 4884 3876 4886 3884
rect 4874 3874 4886 3876
rect 4906 3884 4918 4856
rect 5002 4684 5014 5076
rect 5194 5064 5206 5066
rect 5194 5056 5196 5064
rect 5204 5056 5206 5064
rect 5002 4676 5004 4684
rect 5012 4676 5014 4684
rect 5002 4674 5014 4676
rect 5162 4704 5174 4706
rect 5162 4696 5164 4704
rect 5172 4696 5174 4704
rect 5002 4564 5014 4566
rect 5002 4556 5004 4564
rect 5012 4556 5014 4564
rect 4970 4344 4982 4346
rect 4970 4336 4972 4344
rect 4980 4336 4982 4344
rect 4970 3984 4982 4336
rect 4970 3976 4972 3984
rect 4980 3976 4982 3984
rect 4970 3974 4982 3976
rect 5002 3904 5014 4556
rect 5130 4424 5142 4426
rect 5130 4416 5132 4424
rect 5140 4416 5142 4424
rect 5098 4304 5110 4306
rect 5098 4296 5100 4304
rect 5108 4296 5110 4304
rect 5002 3896 5004 3904
rect 5012 3896 5014 3904
rect 5002 3894 5014 3896
rect 5034 4184 5046 4186
rect 5034 4176 5036 4184
rect 5044 4176 5046 4184
rect 4906 3876 4908 3884
rect 4916 3876 4918 3884
rect 4906 3874 4918 3876
rect 4490 3756 4492 3764
rect 4500 3756 4502 3764
rect 4490 3754 4502 3756
rect 4586 3584 4598 3586
rect 4586 3576 4588 3584
rect 4596 3576 4598 3584
rect 4362 3516 4364 3524
rect 4372 3516 4374 3524
rect 4362 3514 4374 3516
rect 4426 3524 4438 3526
rect 4426 3516 4428 3524
rect 4436 3516 4438 3524
rect 4426 3324 4438 3516
rect 4522 3384 4534 3386
rect 4522 3376 4524 3384
rect 4532 3376 4534 3384
rect 4426 3316 4428 3324
rect 4436 3316 4438 3324
rect 4426 3314 4438 3316
rect 4490 3364 4502 3366
rect 4490 3356 4492 3364
rect 4500 3356 4502 3364
rect 4490 3284 4502 3356
rect 4490 3276 4492 3284
rect 4500 3276 4502 3284
rect 4490 3274 4502 3276
rect 4522 3124 4534 3376
rect 4522 3116 4524 3124
rect 4532 3116 4534 3124
rect 4522 3114 4534 3116
rect 4458 3064 4470 3066
rect 4458 3056 4460 3064
rect 4468 3056 4470 3064
rect 4426 2944 4438 2946
rect 4426 2936 4428 2944
rect 4436 2936 4438 2944
rect 4394 2704 4406 2706
rect 4394 2696 4396 2704
rect 4404 2696 4406 2704
rect 4362 2564 4374 2566
rect 4362 2556 4364 2564
rect 4372 2556 4374 2564
rect 4138 1776 4140 1784
rect 4148 1776 4150 1784
rect 4138 1774 4150 1776
rect 4202 2444 4214 2446
rect 4202 2436 4204 2444
rect 4212 2436 4214 2444
rect 4010 1696 4012 1704
rect 4020 1696 4022 1704
rect 4010 1694 4022 1696
rect 4170 1504 4182 1506
rect 4170 1496 4172 1504
rect 4180 1496 4182 1504
rect 3946 1324 3958 1326
rect 3946 1316 3948 1324
rect 3956 1316 3958 1324
rect 3946 1264 3958 1316
rect 4170 1304 4182 1496
rect 4202 1484 4214 2436
rect 4266 2324 4278 2326
rect 4266 2316 4268 2324
rect 4276 2316 4278 2324
rect 4266 1724 4278 2316
rect 4298 2064 4310 2066
rect 4298 2056 4300 2064
rect 4308 2056 4310 2064
rect 4298 1844 4310 2056
rect 4298 1836 4300 1844
rect 4308 1836 4310 1844
rect 4298 1834 4310 1836
rect 4330 1884 4342 1886
rect 4330 1876 4332 1884
rect 4340 1876 4342 1884
rect 4266 1716 4268 1724
rect 4276 1716 4278 1724
rect 4266 1714 4278 1716
rect 4202 1476 4204 1484
rect 4212 1476 4214 1484
rect 4202 1474 4214 1476
rect 4266 1684 4278 1686
rect 4266 1676 4268 1684
rect 4276 1676 4278 1684
rect 4234 1464 4246 1466
rect 4234 1456 4236 1464
rect 4244 1456 4246 1464
rect 4234 1324 4246 1456
rect 4234 1316 4236 1324
rect 4244 1316 4246 1324
rect 4234 1314 4246 1316
rect 4170 1296 4172 1304
rect 4180 1296 4182 1304
rect 4170 1294 4182 1296
rect 3946 1256 3948 1264
rect 3956 1256 3958 1264
rect 3946 1254 3958 1256
rect 3914 1176 3916 1184
rect 3924 1176 3926 1184
rect 3744 806 3748 814
rect 3756 806 3760 814
rect 3768 806 3772 814
rect 3780 806 3784 814
rect 3792 806 3796 814
rect 3804 806 3808 814
rect 3562 696 3564 704
rect 3572 696 3574 704
rect 3562 694 3574 696
rect 3306 616 3308 624
rect 3316 616 3318 624
rect 3306 614 3318 616
rect 3242 576 3244 584
rect 3252 576 3254 584
rect 3242 574 3254 576
rect 3402 604 3414 606
rect 3402 596 3404 604
rect 3412 596 3414 604
rect 3402 444 3414 596
rect 3402 436 3404 444
rect 3412 436 3414 444
rect 3402 434 3414 436
rect 3114 356 3116 364
rect 3124 356 3126 364
rect 3114 354 3126 356
rect 3744 414 3808 806
rect 3744 406 3748 414
rect 3756 406 3760 414
rect 3768 406 3772 414
rect 3780 406 3784 414
rect 3792 406 3796 414
rect 3804 406 3808 414
rect 3050 336 3052 344
rect 3060 336 3062 344
rect 3050 334 3062 336
rect 2858 276 2860 284
rect 2868 276 2870 284
rect 2858 274 2870 276
rect 2730 176 2732 184
rect 2740 176 2742 184
rect 2730 174 2742 176
rect 3744 14 3808 406
rect 3850 1084 3862 1086
rect 3850 1076 3852 1084
rect 3860 1076 3862 1084
rect 3850 344 3862 1076
rect 3850 336 3852 344
rect 3860 336 3862 344
rect 3850 334 3862 336
rect 3882 864 3894 866
rect 3882 856 3884 864
rect 3892 856 3894 864
rect 3882 344 3894 856
rect 3914 724 3926 1176
rect 3946 1164 3958 1166
rect 3946 1156 3948 1164
rect 3956 1156 3958 1164
rect 3946 904 3958 1156
rect 4266 1164 4278 1676
rect 4330 1624 4342 1876
rect 4330 1616 4332 1624
rect 4340 1616 4342 1624
rect 4330 1614 4342 1616
rect 4362 1504 4374 2556
rect 4394 1864 4406 2696
rect 4426 2524 4438 2936
rect 4458 2704 4470 3056
rect 4458 2696 4460 2704
rect 4468 2696 4470 2704
rect 4458 2694 4470 2696
rect 4522 3064 4534 3066
rect 4522 3056 4524 3064
rect 4532 3056 4534 3064
rect 4426 2516 4428 2524
rect 4436 2516 4438 2524
rect 4426 2514 4438 2516
rect 4426 2464 4438 2466
rect 4426 2456 4428 2464
rect 4436 2456 4438 2464
rect 4426 2064 4438 2456
rect 4522 2464 4534 3056
rect 4522 2456 4524 2464
rect 4532 2456 4534 2464
rect 4522 2454 4534 2456
rect 4522 2404 4534 2406
rect 4522 2396 4524 2404
rect 4532 2396 4534 2404
rect 4522 2144 4534 2396
rect 4586 2404 4598 3576
rect 4714 3564 4726 3566
rect 4714 3556 4716 3564
rect 4724 3556 4726 3564
rect 4586 2396 4588 2404
rect 4596 2396 4598 2404
rect 4586 2394 4598 2396
rect 4618 3504 4630 3506
rect 4618 3496 4620 3504
rect 4628 3496 4630 3504
rect 4618 3324 4630 3496
rect 4714 3344 4726 3556
rect 5034 3564 5046 4176
rect 5098 3884 5110 4296
rect 5130 3966 5142 4416
rect 5162 4304 5174 4696
rect 5194 4644 5206 5056
rect 5194 4636 5196 4644
rect 5204 4636 5206 4644
rect 5194 4634 5206 4636
rect 5248 5014 5312 5216
rect 6752 5214 6816 5216
rect 6752 5206 6756 5214
rect 6764 5206 6768 5214
rect 6776 5206 6780 5214
rect 6788 5206 6792 5214
rect 6800 5206 6804 5214
rect 6812 5206 6816 5214
rect 5248 5006 5252 5014
rect 5260 5006 5264 5014
rect 5272 5006 5276 5014
rect 5284 5006 5288 5014
rect 5296 5006 5300 5014
rect 5308 5006 5312 5014
rect 5162 4296 5164 4304
rect 5172 4296 5174 4304
rect 5162 4104 5174 4296
rect 5162 4096 5164 4104
rect 5172 4096 5174 4104
rect 5162 4094 5174 4096
rect 5248 4614 5312 5006
rect 6282 5024 6294 5026
rect 6282 5016 6284 5024
rect 6292 5016 6294 5024
rect 5738 4944 5750 4946
rect 5738 4936 5740 4944
rect 5748 4936 5750 4944
rect 5738 4926 5750 4936
rect 5610 4914 5750 4926
rect 5834 4944 5846 4946
rect 5834 4936 5836 4944
rect 5844 4936 5846 4944
rect 5610 4904 5622 4914
rect 5610 4896 5612 4904
rect 5620 4896 5622 4904
rect 5610 4894 5622 4896
rect 5248 4606 5252 4614
rect 5260 4606 5264 4614
rect 5272 4606 5276 4614
rect 5284 4606 5288 4614
rect 5296 4606 5300 4614
rect 5308 4606 5312 4614
rect 5248 4214 5312 4606
rect 5248 4206 5252 4214
rect 5260 4206 5264 4214
rect 5272 4206 5276 4214
rect 5284 4206 5288 4214
rect 5296 4206 5300 4214
rect 5308 4206 5312 4214
rect 5130 3954 5174 3966
rect 5098 3876 5100 3884
rect 5108 3876 5110 3884
rect 5098 3874 5110 3876
rect 5034 3556 5036 3564
rect 5044 3556 5046 3564
rect 4810 3504 4822 3506
rect 4810 3496 4812 3504
rect 4820 3496 4822 3504
rect 4714 3336 4716 3344
rect 4724 3336 4726 3344
rect 4714 3334 4726 3336
rect 4778 3384 4790 3386
rect 4778 3376 4780 3384
rect 4788 3376 4790 3384
rect 4618 3316 4620 3324
rect 4628 3316 4630 3324
rect 4618 2924 4630 3316
rect 4746 3324 4758 3326
rect 4746 3316 4748 3324
rect 4756 3316 4758 3324
rect 4618 2916 4620 2924
rect 4628 2916 4630 2924
rect 4522 2136 4524 2144
rect 4532 2136 4534 2144
rect 4522 2134 4534 2136
rect 4586 2364 4598 2366
rect 4586 2356 4588 2364
rect 4596 2356 4598 2364
rect 4554 2104 4566 2106
rect 4554 2096 4556 2104
rect 4564 2096 4566 2104
rect 4426 2056 4428 2064
rect 4436 2056 4438 2064
rect 4426 2054 4438 2056
rect 4490 2084 4502 2086
rect 4490 2076 4492 2084
rect 4500 2076 4502 2084
rect 4394 1856 4396 1864
rect 4404 1856 4406 1864
rect 4394 1854 4406 1856
rect 4458 1644 4470 1646
rect 4458 1636 4460 1644
rect 4468 1636 4470 1644
rect 4458 1544 4470 1636
rect 4458 1536 4460 1544
rect 4468 1536 4470 1544
rect 4458 1534 4470 1536
rect 4362 1496 4364 1504
rect 4372 1496 4374 1504
rect 4362 1494 4374 1496
rect 4394 1524 4406 1526
rect 4394 1516 4396 1524
rect 4404 1516 4406 1524
rect 4394 1484 4406 1516
rect 4394 1476 4396 1484
rect 4404 1476 4406 1484
rect 4394 1474 4406 1476
rect 4490 1364 4502 2076
rect 4522 1844 4534 1846
rect 4522 1836 4524 1844
rect 4532 1836 4534 1844
rect 4522 1504 4534 1836
rect 4554 1824 4566 2096
rect 4586 1904 4598 2356
rect 4618 2144 4630 2916
rect 4650 3224 4662 3226
rect 4650 3216 4652 3224
rect 4660 3216 4662 3224
rect 4650 2364 4662 3216
rect 4746 3204 4758 3316
rect 4746 3196 4748 3204
rect 4756 3196 4758 3204
rect 4746 3194 4758 3196
rect 4746 3044 4758 3046
rect 4746 3036 4748 3044
rect 4756 3036 4758 3044
rect 4746 2924 4758 3036
rect 4746 2916 4748 2924
rect 4756 2916 4758 2924
rect 4746 2704 4758 2916
rect 4778 2784 4790 3376
rect 4810 3364 4822 3496
rect 4810 3356 4812 3364
rect 4820 3356 4822 3364
rect 4810 3354 4822 3356
rect 4938 3504 4950 3506
rect 4938 3496 4940 3504
rect 4948 3496 4950 3504
rect 4938 3304 4950 3496
rect 4938 3296 4940 3304
rect 4948 3296 4950 3304
rect 4938 2904 4950 3296
rect 5034 3164 5046 3556
rect 5034 3156 5036 3164
rect 5044 3156 5046 3164
rect 5034 3154 5046 3156
rect 5098 3544 5110 3546
rect 5098 3536 5100 3544
rect 5108 3536 5110 3544
rect 5098 3144 5110 3536
rect 5130 3524 5142 3526
rect 5130 3516 5132 3524
rect 5140 3516 5142 3524
rect 5130 3404 5142 3516
rect 5162 3464 5174 3954
rect 5162 3456 5164 3464
rect 5172 3456 5174 3464
rect 5162 3454 5174 3456
rect 5248 3814 5312 4206
rect 5514 4824 5526 4826
rect 5514 4816 5516 4824
rect 5524 4816 5526 4824
rect 5248 3806 5252 3814
rect 5260 3806 5264 3814
rect 5272 3806 5276 3814
rect 5284 3806 5288 3814
rect 5296 3806 5300 3814
rect 5308 3806 5312 3814
rect 5248 3414 5312 3806
rect 5482 3924 5494 3926
rect 5482 3916 5484 3924
rect 5492 3916 5494 3924
rect 5418 3704 5430 3706
rect 5418 3696 5420 3704
rect 5428 3696 5430 3704
rect 5248 3406 5252 3414
rect 5260 3406 5264 3414
rect 5272 3406 5276 3414
rect 5284 3406 5288 3414
rect 5296 3406 5300 3414
rect 5308 3406 5312 3414
rect 5130 3396 5132 3404
rect 5140 3396 5142 3404
rect 5130 3394 5142 3396
rect 5162 3404 5174 3406
rect 5162 3396 5164 3404
rect 5172 3396 5174 3404
rect 5098 3136 5100 3144
rect 5108 3136 5110 3144
rect 5098 3134 5110 3136
rect 5130 3344 5142 3346
rect 5130 3336 5132 3344
rect 5140 3336 5142 3344
rect 5066 3084 5078 3086
rect 5066 3076 5068 3084
rect 5076 3076 5078 3084
rect 4938 2896 4940 2904
rect 4948 2896 4950 2904
rect 4938 2894 4950 2896
rect 4970 3064 4982 3066
rect 4970 3056 4972 3064
rect 4980 3056 4982 3064
rect 4778 2776 4780 2784
rect 4788 2776 4790 2784
rect 4778 2774 4790 2776
rect 4970 2784 4982 3056
rect 5034 2864 5046 2866
rect 5034 2856 5036 2864
rect 5044 2856 5046 2864
rect 5034 2824 5046 2856
rect 5034 2816 5036 2824
rect 5044 2816 5046 2824
rect 5034 2814 5046 2816
rect 5066 2844 5078 3076
rect 5066 2836 5068 2844
rect 5076 2836 5078 2844
rect 4970 2776 4972 2784
rect 4980 2776 4982 2784
rect 4970 2774 4982 2776
rect 4746 2696 4748 2704
rect 4756 2696 4758 2704
rect 4746 2694 4758 2696
rect 4714 2634 4758 2646
rect 4714 2624 4726 2634
rect 4714 2616 4716 2624
rect 4724 2616 4726 2624
rect 4714 2614 4726 2616
rect 4746 2604 4758 2634
rect 4746 2596 4748 2604
rect 4756 2596 4758 2604
rect 4746 2594 4758 2596
rect 5066 2564 5078 2836
rect 5130 3084 5142 3336
rect 5130 3076 5132 3084
rect 5140 3076 5142 3084
rect 5066 2556 5068 2564
rect 5076 2556 5078 2564
rect 5066 2554 5078 2556
rect 5098 2704 5110 2706
rect 5098 2696 5100 2704
rect 5108 2696 5110 2704
rect 4650 2356 4652 2364
rect 4660 2356 4662 2364
rect 4650 2354 4662 2356
rect 4682 2464 4694 2466
rect 4682 2456 4684 2464
rect 4692 2456 4694 2464
rect 4618 2136 4620 2144
rect 4628 2136 4630 2144
rect 4618 2134 4630 2136
rect 4586 1896 4588 1904
rect 4596 1896 4598 1904
rect 4586 1894 4598 1896
rect 4554 1816 4556 1824
rect 4564 1816 4566 1824
rect 4554 1814 4566 1816
rect 4618 1824 4630 1826
rect 4618 1816 4620 1824
rect 4628 1816 4630 1824
rect 4522 1496 4524 1504
rect 4532 1496 4534 1504
rect 4522 1494 4534 1496
rect 4554 1784 4566 1786
rect 4554 1776 4556 1784
rect 4564 1776 4566 1784
rect 4490 1356 4492 1364
rect 4500 1356 4502 1364
rect 4490 1354 4502 1356
rect 4554 1344 4566 1776
rect 4554 1336 4556 1344
rect 4564 1336 4566 1344
rect 4554 1334 4566 1336
rect 4266 1156 4268 1164
rect 4276 1156 4278 1164
rect 4266 1154 4278 1156
rect 4426 964 4438 966
rect 4426 956 4428 964
rect 4436 956 4438 964
rect 4298 944 4310 946
rect 4298 936 4300 944
rect 4308 936 4310 944
rect 4298 926 4310 936
rect 3946 896 3948 904
rect 3956 896 3958 904
rect 3946 894 3958 896
rect 4074 924 4086 926
rect 4074 916 4076 924
rect 4084 916 4086 924
rect 3914 716 3916 724
rect 3924 716 3926 724
rect 3914 714 3926 716
rect 3882 336 3884 344
rect 3892 336 3894 344
rect 3882 334 3894 336
rect 3914 444 3926 446
rect 3914 436 3916 444
rect 3924 436 3926 444
rect 3914 304 3926 436
rect 4074 424 4086 916
rect 4106 914 4310 926
rect 4426 926 4438 956
rect 4458 944 4470 946
rect 4458 936 4460 944
rect 4468 936 4470 944
rect 4458 926 4470 936
rect 4426 914 4470 926
rect 4106 904 4118 914
rect 4106 896 4108 904
rect 4116 896 4118 904
rect 4106 894 4118 896
rect 4618 904 4630 1816
rect 4682 1704 4694 2456
rect 5002 2364 5014 2366
rect 5002 2356 5004 2364
rect 5012 2356 5014 2364
rect 4874 2324 4886 2326
rect 4874 2316 4876 2324
rect 4884 2316 4886 2324
rect 4842 1904 4854 1906
rect 4842 1896 4844 1904
rect 4852 1896 4854 1904
rect 4842 1844 4854 1896
rect 4842 1836 4844 1844
rect 4852 1836 4854 1844
rect 4842 1834 4854 1836
rect 4682 1696 4684 1704
rect 4692 1696 4694 1704
rect 4682 1694 4694 1696
rect 4842 1644 4854 1646
rect 4842 1636 4844 1644
rect 4852 1636 4854 1644
rect 4778 1404 4790 1406
rect 4778 1396 4780 1404
rect 4788 1396 4790 1404
rect 4778 1224 4790 1396
rect 4778 1216 4780 1224
rect 4788 1216 4790 1224
rect 4778 1214 4790 1216
rect 4842 1104 4854 1636
rect 4874 1404 4886 2316
rect 4970 2244 4982 2246
rect 4970 2236 4972 2244
rect 4980 2236 4982 2244
rect 4970 2204 4982 2236
rect 4970 2196 4972 2204
rect 4980 2196 4982 2204
rect 4970 2194 4982 2196
rect 5002 2024 5014 2356
rect 5002 2016 5004 2024
rect 5012 2016 5014 2024
rect 5002 2014 5014 2016
rect 5066 2224 5078 2226
rect 5066 2216 5068 2224
rect 5076 2216 5078 2224
rect 5002 1884 5014 1886
rect 5002 1876 5004 1884
rect 5012 1876 5014 1884
rect 5002 1524 5014 1876
rect 5002 1516 5004 1524
rect 5012 1516 5014 1524
rect 5002 1514 5014 1516
rect 5034 1844 5046 1846
rect 5034 1836 5036 1844
rect 5044 1836 5046 1844
rect 4874 1396 4876 1404
rect 4884 1396 4886 1404
rect 4874 1394 4886 1396
rect 5034 1324 5046 1836
rect 5034 1316 5036 1324
rect 5044 1316 5046 1324
rect 5034 1314 5046 1316
rect 5066 1224 5078 2216
rect 5098 2024 5110 2696
rect 5130 2544 5142 3076
rect 5162 2824 5174 3396
rect 5248 3014 5312 3406
rect 5354 3464 5366 3466
rect 5354 3456 5356 3464
rect 5364 3456 5366 3464
rect 5354 3364 5366 3456
rect 5354 3356 5356 3364
rect 5364 3356 5366 3364
rect 5354 3354 5366 3356
rect 5418 3144 5430 3696
rect 5482 3524 5494 3916
rect 5482 3516 5484 3524
rect 5492 3516 5494 3524
rect 5482 3514 5494 3516
rect 5418 3136 5420 3144
rect 5428 3136 5430 3144
rect 5418 3134 5430 3136
rect 5450 3504 5462 3506
rect 5450 3496 5452 3504
rect 5460 3496 5462 3504
rect 5248 3006 5252 3014
rect 5260 3006 5264 3014
rect 5272 3006 5276 3014
rect 5284 3006 5288 3014
rect 5296 3006 5300 3014
rect 5308 3006 5312 3014
rect 5162 2816 5164 2824
rect 5172 2816 5174 2824
rect 5162 2814 5174 2816
rect 5194 2964 5206 2966
rect 5194 2956 5196 2964
rect 5204 2956 5206 2964
rect 5194 2824 5206 2956
rect 5194 2816 5196 2824
rect 5204 2816 5206 2824
rect 5194 2814 5206 2816
rect 5130 2536 5132 2544
rect 5140 2536 5142 2544
rect 5130 2534 5142 2536
rect 5194 2704 5206 2706
rect 5194 2696 5196 2704
rect 5204 2696 5206 2704
rect 5130 2324 5142 2326
rect 5130 2316 5132 2324
rect 5140 2316 5142 2324
rect 5130 2104 5142 2316
rect 5194 2324 5206 2696
rect 5194 2316 5196 2324
rect 5204 2316 5206 2324
rect 5194 2314 5206 2316
rect 5248 2614 5312 3006
rect 5450 2784 5462 3496
rect 5514 3504 5526 4816
rect 5802 4824 5814 4826
rect 5802 4816 5804 4824
rect 5812 4816 5814 4824
rect 5674 4804 5686 4806
rect 5674 4796 5676 4804
rect 5684 4796 5686 4804
rect 5610 4384 5622 4386
rect 5610 4376 5612 4384
rect 5620 4376 5622 4384
rect 5610 3844 5622 4376
rect 5610 3836 5612 3844
rect 5620 3836 5622 3844
rect 5610 3834 5622 3836
rect 5674 3544 5686 4796
rect 5802 4064 5814 4816
rect 5802 4056 5804 4064
rect 5812 4056 5814 4064
rect 5802 4054 5814 4056
rect 5674 3536 5676 3544
rect 5684 3536 5686 3544
rect 5674 3534 5686 3536
rect 5738 3544 5750 3546
rect 5738 3536 5740 3544
rect 5748 3536 5750 3544
rect 5514 3496 5516 3504
rect 5524 3496 5526 3504
rect 5514 3494 5526 3496
rect 5546 3484 5558 3486
rect 5546 3476 5548 3484
rect 5556 3476 5558 3484
rect 5514 3404 5526 3406
rect 5514 3396 5516 3404
rect 5524 3396 5526 3404
rect 5514 3204 5526 3396
rect 5514 3196 5516 3204
rect 5524 3196 5526 3204
rect 5450 2776 5452 2784
rect 5460 2776 5462 2784
rect 5450 2774 5462 2776
rect 5482 3124 5494 3126
rect 5482 3116 5484 3124
rect 5492 3116 5494 3124
rect 5482 2904 5494 3116
rect 5514 2924 5526 3196
rect 5546 2964 5558 3476
rect 5546 2956 5548 2964
rect 5556 2956 5558 2964
rect 5546 2954 5558 2956
rect 5610 3344 5622 3346
rect 5610 3336 5612 3344
rect 5620 3336 5622 3344
rect 5610 3064 5622 3336
rect 5706 3184 5718 3186
rect 5706 3176 5708 3184
rect 5716 3176 5718 3184
rect 5706 3126 5718 3176
rect 5738 3184 5750 3536
rect 5738 3176 5740 3184
rect 5748 3176 5750 3184
rect 5738 3174 5750 3176
rect 5770 3184 5782 3186
rect 5770 3176 5772 3184
rect 5780 3176 5782 3184
rect 5770 3126 5782 3176
rect 5610 3056 5612 3064
rect 5620 3056 5622 3064
rect 5514 2916 5516 2924
rect 5524 2916 5526 2924
rect 5514 2914 5526 2916
rect 5546 2924 5558 2926
rect 5546 2916 5548 2924
rect 5556 2916 5558 2924
rect 5482 2896 5484 2904
rect 5492 2896 5494 2904
rect 5354 2764 5366 2766
rect 5354 2756 5356 2764
rect 5364 2756 5366 2764
rect 5354 2624 5366 2756
rect 5354 2616 5356 2624
rect 5364 2616 5366 2624
rect 5354 2614 5366 2616
rect 5418 2724 5430 2726
rect 5418 2716 5420 2724
rect 5428 2716 5430 2724
rect 5248 2606 5252 2614
rect 5260 2606 5264 2614
rect 5272 2606 5276 2614
rect 5284 2606 5288 2614
rect 5296 2606 5300 2614
rect 5308 2606 5312 2614
rect 5248 2214 5312 2606
rect 5386 2604 5398 2606
rect 5386 2596 5388 2604
rect 5396 2596 5398 2604
rect 5386 2524 5398 2596
rect 5386 2516 5388 2524
rect 5396 2516 5398 2524
rect 5386 2514 5398 2516
rect 5354 2464 5366 2466
rect 5354 2456 5356 2464
rect 5364 2456 5366 2464
rect 5354 2344 5366 2456
rect 5418 2384 5430 2716
rect 5482 2504 5494 2896
rect 5546 2524 5558 2916
rect 5578 2924 5590 2926
rect 5578 2916 5580 2924
rect 5588 2916 5590 2924
rect 5578 2784 5590 2916
rect 5578 2776 5580 2784
rect 5588 2776 5590 2784
rect 5578 2644 5590 2776
rect 5578 2636 5580 2644
rect 5588 2636 5590 2644
rect 5578 2634 5590 2636
rect 5546 2516 5548 2524
rect 5556 2516 5558 2524
rect 5482 2496 5484 2504
rect 5492 2496 5494 2504
rect 5482 2494 5494 2496
rect 5514 2504 5526 2506
rect 5514 2496 5516 2504
rect 5524 2496 5526 2504
rect 5418 2376 5420 2384
rect 5428 2376 5430 2384
rect 5418 2374 5430 2376
rect 5354 2336 5356 2344
rect 5364 2336 5366 2344
rect 5354 2334 5366 2336
rect 5248 2206 5252 2214
rect 5260 2206 5264 2214
rect 5272 2206 5276 2214
rect 5284 2206 5288 2214
rect 5296 2206 5300 2214
rect 5308 2206 5312 2214
rect 5130 2096 5132 2104
rect 5140 2096 5142 2104
rect 5130 2094 5142 2096
rect 5194 2104 5206 2106
rect 5194 2096 5196 2104
rect 5204 2096 5206 2104
rect 5098 2016 5100 2024
rect 5108 2016 5110 2024
rect 5098 2014 5110 2016
rect 5098 1584 5110 1586
rect 5098 1576 5100 1584
rect 5108 1576 5110 1584
rect 5098 1524 5110 1576
rect 5098 1516 5100 1524
rect 5108 1516 5110 1524
rect 5098 1514 5110 1516
rect 5066 1216 5068 1224
rect 5076 1216 5078 1224
rect 5066 1214 5078 1216
rect 5162 1404 5174 1406
rect 5162 1396 5164 1404
rect 5172 1396 5174 1404
rect 4842 1096 4844 1104
rect 4852 1096 4854 1104
rect 4842 1094 4854 1096
rect 5002 1144 5014 1146
rect 5002 1136 5004 1144
rect 5012 1136 5014 1144
rect 4842 964 4854 966
rect 4842 956 4844 964
rect 4852 956 4854 964
rect 4618 896 4620 904
rect 4628 896 4630 904
rect 4330 864 4342 866
rect 4330 856 4332 864
rect 4340 856 4342 864
rect 4330 444 4342 856
rect 4330 436 4332 444
rect 4340 436 4342 444
rect 4330 434 4342 436
rect 4362 724 4374 726
rect 4362 716 4364 724
rect 4372 716 4374 724
rect 4362 544 4374 716
rect 4618 724 4630 896
rect 4618 716 4620 724
rect 4628 716 4630 724
rect 4618 714 4630 716
rect 4682 904 4694 906
rect 4682 896 4684 904
rect 4692 896 4694 904
rect 4362 536 4364 544
rect 4372 536 4374 544
rect 4074 416 4076 424
rect 4084 416 4086 424
rect 4074 414 4086 416
rect 3914 296 3916 304
rect 3924 296 3926 304
rect 3914 294 3926 296
rect 4362 144 4374 536
rect 4394 664 4406 666
rect 4394 656 4396 664
rect 4404 656 4406 664
rect 4394 164 4406 656
rect 4490 624 4502 626
rect 4490 616 4492 624
rect 4500 616 4502 624
rect 4490 224 4502 616
rect 4682 544 4694 896
rect 4842 664 4854 956
rect 5002 784 5014 1136
rect 5002 776 5004 784
rect 5012 776 5014 784
rect 5002 774 5014 776
rect 5162 724 5174 1396
rect 5194 1124 5206 2096
rect 5194 1116 5196 1124
rect 5204 1116 5206 1124
rect 5194 1114 5206 1116
rect 5248 1814 5312 2206
rect 5386 2284 5398 2286
rect 5386 2276 5388 2284
rect 5396 2276 5398 2284
rect 5354 2184 5366 2186
rect 5354 2176 5356 2184
rect 5364 2176 5366 2184
rect 5354 2044 5366 2176
rect 5354 2036 5356 2044
rect 5364 2036 5366 2044
rect 5354 2034 5366 2036
rect 5386 1964 5398 2276
rect 5386 1956 5388 1964
rect 5396 1956 5398 1964
rect 5386 1954 5398 1956
rect 5450 2224 5462 2226
rect 5450 2216 5452 2224
rect 5460 2216 5462 2224
rect 5248 1806 5252 1814
rect 5260 1806 5264 1814
rect 5272 1806 5276 1814
rect 5284 1806 5288 1814
rect 5296 1806 5300 1814
rect 5308 1806 5312 1814
rect 5248 1414 5312 1806
rect 5386 1824 5398 1826
rect 5386 1816 5388 1824
rect 5396 1816 5398 1824
rect 5386 1584 5398 1816
rect 5450 1764 5462 2216
rect 5450 1756 5452 1764
rect 5460 1756 5462 1764
rect 5450 1754 5462 1756
rect 5482 1924 5494 1926
rect 5482 1916 5484 1924
rect 5492 1916 5494 1924
rect 5482 1604 5494 1916
rect 5514 1924 5526 2496
rect 5514 1916 5516 1924
rect 5524 1916 5526 1924
rect 5514 1914 5526 1916
rect 5482 1596 5484 1604
rect 5492 1596 5494 1604
rect 5482 1594 5494 1596
rect 5386 1576 5388 1584
rect 5396 1576 5398 1584
rect 5386 1574 5398 1576
rect 5546 1504 5558 2516
rect 5610 2484 5622 3056
rect 5642 3124 5654 3126
rect 5642 3116 5644 3124
rect 5652 3116 5654 3124
rect 5642 2724 5654 3116
rect 5706 3114 5782 3126
rect 5642 2716 5644 2724
rect 5652 2716 5654 2724
rect 5642 2714 5654 2716
rect 5674 3104 5686 3106
rect 5674 3096 5676 3104
rect 5684 3096 5686 3104
rect 5674 2544 5686 3096
rect 5674 2536 5676 2544
rect 5684 2536 5686 2544
rect 5674 2534 5686 2536
rect 5610 2476 5612 2484
rect 5620 2476 5622 2484
rect 5610 2474 5622 2476
rect 5610 2384 5622 2386
rect 5610 2376 5612 2384
rect 5620 2376 5622 2384
rect 5610 2124 5622 2376
rect 5610 2116 5612 2124
rect 5620 2116 5622 2124
rect 5610 2114 5622 2116
rect 5834 2124 5846 4936
rect 6282 4684 6294 5016
rect 6666 4844 6678 4846
rect 6666 4836 6668 4844
rect 6676 4836 6678 4844
rect 6282 4676 6284 4684
rect 6292 4676 6294 4684
rect 6282 4674 6294 4676
rect 6314 4824 6326 4826
rect 6314 4816 6316 4824
rect 6324 4816 6326 4824
rect 6058 4584 6070 4586
rect 6058 4576 6060 4584
rect 6068 4576 6070 4584
rect 6058 4524 6070 4576
rect 6154 4544 6166 4546
rect 6154 4536 6156 4544
rect 6164 4536 6166 4544
rect 6058 4516 6060 4524
rect 6068 4516 6070 4524
rect 6058 4514 6070 4516
rect 6090 4524 6102 4526
rect 6090 4516 6092 4524
rect 6100 4516 6102 4524
rect 6090 4484 6102 4516
rect 6090 4476 6092 4484
rect 6100 4476 6102 4484
rect 6090 4474 6102 4476
rect 5866 4344 5878 4346
rect 5866 4336 5868 4344
rect 5876 4336 5878 4344
rect 5866 4124 5878 4336
rect 6026 4284 6038 4286
rect 6026 4276 6028 4284
rect 6036 4276 6038 4284
rect 5866 4116 5868 4124
rect 5876 4116 5878 4124
rect 5866 4114 5878 4116
rect 5930 4264 5942 4266
rect 5930 4256 5932 4264
rect 5940 4256 5942 4264
rect 5930 3884 5942 4256
rect 6026 4024 6038 4276
rect 6154 4224 6166 4536
rect 6314 4324 6326 4816
rect 6314 4316 6316 4324
rect 6324 4316 6326 4324
rect 6314 4314 6326 4316
rect 6346 4344 6358 4346
rect 6346 4336 6348 4344
rect 6356 4336 6358 4344
rect 6154 4216 6156 4224
rect 6164 4216 6166 4224
rect 6122 4184 6134 4186
rect 6122 4176 6124 4184
rect 6132 4176 6134 4184
rect 6122 4124 6134 4176
rect 6122 4116 6124 4124
rect 6132 4116 6134 4124
rect 6122 4114 6134 4116
rect 6026 4016 6028 4024
rect 6036 4016 6038 4024
rect 6026 4014 6038 4016
rect 6154 3944 6166 4216
rect 6154 3936 6156 3944
rect 6164 3936 6166 3944
rect 6154 3934 6166 3936
rect 6186 4264 6198 4266
rect 6186 4256 6188 4264
rect 6196 4256 6198 4264
rect 5930 3876 5932 3884
rect 5940 3876 5942 3884
rect 5930 3874 5942 3876
rect 5994 3784 6006 3786
rect 5994 3776 5996 3784
rect 6004 3776 6006 3784
rect 5930 3244 5942 3246
rect 5930 3236 5932 3244
rect 5940 3236 5942 3244
rect 5898 2984 5910 2986
rect 5898 2976 5900 2984
rect 5908 2976 5910 2984
rect 5898 2924 5910 2976
rect 5898 2916 5900 2924
rect 5908 2916 5910 2924
rect 5898 2914 5910 2916
rect 5930 2824 5942 3236
rect 5994 3084 6006 3776
rect 5994 3076 5996 3084
rect 6004 3076 6006 3084
rect 5994 3074 6006 3076
rect 6058 3284 6070 3286
rect 6058 3276 6060 3284
rect 6068 3276 6070 3284
rect 5930 2816 5932 2824
rect 5940 2816 5942 2824
rect 5930 2814 5942 2816
rect 6058 2464 6070 3276
rect 6186 2944 6198 4256
rect 6250 4204 6262 4206
rect 6250 4196 6252 4204
rect 6260 4196 6262 4204
rect 6218 4184 6230 4186
rect 6218 4176 6220 4184
rect 6228 4176 6230 4184
rect 6218 3124 6230 4176
rect 6250 3344 6262 4196
rect 6250 3336 6252 3344
rect 6260 3336 6262 3344
rect 6250 3334 6262 3336
rect 6314 3404 6326 3406
rect 6314 3396 6316 3404
rect 6324 3396 6326 3404
rect 6314 3144 6326 3396
rect 6346 3304 6358 4336
rect 6378 3844 6390 3846
rect 6378 3836 6380 3844
rect 6388 3836 6390 3844
rect 6378 3344 6390 3836
rect 6378 3336 6380 3344
rect 6388 3336 6390 3344
rect 6378 3334 6390 3336
rect 6410 3804 6422 3806
rect 6410 3796 6412 3804
rect 6420 3796 6422 3804
rect 6346 3296 6348 3304
rect 6356 3296 6358 3304
rect 6346 3294 6358 3296
rect 6314 3136 6316 3144
rect 6324 3136 6326 3144
rect 6314 3134 6326 3136
rect 6410 3204 6422 3796
rect 6666 3724 6678 4836
rect 6752 4814 6816 5206
rect 7338 5064 7350 5066
rect 7338 5056 7340 5064
rect 7348 5056 7350 5064
rect 6752 4806 6756 4814
rect 6764 4806 6768 4814
rect 6776 4806 6780 4814
rect 6788 4806 6792 4814
rect 6800 4806 6804 4814
rect 6812 4806 6816 4814
rect 6698 4544 6710 4546
rect 6698 4536 6700 4544
rect 6708 4536 6710 4544
rect 6698 4184 6710 4536
rect 6698 4176 6700 4184
rect 6708 4176 6710 4184
rect 6698 4174 6710 4176
rect 6752 4414 6816 4806
rect 6752 4406 6756 4414
rect 6764 4406 6768 4414
rect 6776 4406 6780 4414
rect 6788 4406 6792 4414
rect 6800 4406 6804 4414
rect 6812 4406 6816 4414
rect 6666 3716 6668 3724
rect 6676 3716 6678 3724
rect 6666 3714 6678 3716
rect 6752 4014 6816 4406
rect 6858 5044 6870 5046
rect 6858 5036 6860 5044
rect 6868 5036 6870 5044
rect 6858 4304 6870 5036
rect 7306 5004 7318 5006
rect 7306 4996 7308 5004
rect 7316 4996 7318 5004
rect 6858 4296 6860 4304
rect 6868 4296 6870 4304
rect 6858 4294 6870 4296
rect 6954 4804 6966 4806
rect 6954 4796 6956 4804
rect 6964 4796 6966 4804
rect 6752 4006 6756 4014
rect 6764 4006 6768 4014
rect 6776 4006 6780 4014
rect 6788 4006 6792 4014
rect 6800 4006 6804 4014
rect 6812 4006 6816 4014
rect 6570 3644 6582 3646
rect 6570 3636 6572 3644
rect 6580 3636 6582 3644
rect 6538 3544 6550 3546
rect 6538 3536 6540 3544
rect 6548 3536 6550 3544
rect 6442 3504 6454 3506
rect 6442 3496 6444 3504
rect 6452 3496 6454 3504
rect 6442 3444 6454 3496
rect 6442 3436 6444 3444
rect 6452 3436 6454 3444
rect 6442 3434 6454 3436
rect 6538 3344 6550 3536
rect 6538 3336 6540 3344
rect 6548 3336 6550 3344
rect 6538 3334 6550 3336
rect 6410 3196 6412 3204
rect 6420 3196 6422 3204
rect 6218 3116 6220 3124
rect 6228 3116 6230 3124
rect 6218 3114 6230 3116
rect 6186 2936 6188 2944
rect 6196 2936 6198 2944
rect 6186 2934 6198 2936
rect 6218 3084 6230 3086
rect 6218 3076 6220 3084
rect 6228 3076 6230 3084
rect 6058 2456 6060 2464
rect 6068 2456 6070 2464
rect 6058 2454 6070 2456
rect 6154 2684 6166 2686
rect 6154 2676 6156 2684
rect 6164 2676 6166 2684
rect 5834 2116 5836 2124
rect 5844 2116 5846 2124
rect 5834 2114 5846 2116
rect 5962 2204 5974 2206
rect 5962 2196 5964 2204
rect 5972 2196 5974 2204
rect 5962 2064 5974 2196
rect 5962 2056 5964 2064
rect 5972 2056 5974 2064
rect 5962 2054 5974 2056
rect 6154 1884 6166 2676
rect 6186 2224 6198 2226
rect 6186 2216 6188 2224
rect 6196 2216 6198 2224
rect 6186 2084 6198 2216
rect 6218 2224 6230 3076
rect 6314 3084 6326 3086
rect 6314 3076 6316 3084
rect 6324 3076 6326 3084
rect 6250 2564 6262 2566
rect 6250 2556 6252 2564
rect 6260 2556 6262 2564
rect 6250 2524 6262 2556
rect 6250 2516 6252 2524
rect 6260 2516 6262 2524
rect 6250 2514 6262 2516
rect 6218 2216 6220 2224
rect 6228 2216 6230 2224
rect 6218 2214 6230 2216
rect 6186 2076 6188 2084
rect 6196 2076 6198 2084
rect 6186 2074 6198 2076
rect 6282 2124 6294 2126
rect 6282 2116 6284 2124
rect 6292 2116 6294 2124
rect 6154 1876 6156 1884
rect 6164 1876 6166 1884
rect 6154 1874 6166 1876
rect 5834 1824 5846 1826
rect 5834 1816 5836 1824
rect 5844 1816 5846 1824
rect 5546 1496 5548 1504
rect 5556 1496 5558 1504
rect 5546 1494 5558 1496
rect 5674 1764 5686 1766
rect 5674 1756 5676 1764
rect 5684 1756 5686 1764
rect 5248 1406 5252 1414
rect 5260 1406 5264 1414
rect 5272 1406 5276 1414
rect 5284 1406 5288 1414
rect 5296 1406 5300 1414
rect 5308 1406 5312 1414
rect 5162 716 5164 724
rect 5172 716 5174 724
rect 5162 714 5174 716
rect 5248 1014 5312 1406
rect 5578 1284 5590 1286
rect 5578 1276 5580 1284
rect 5588 1276 5590 1284
rect 5248 1006 5252 1014
rect 5260 1006 5264 1014
rect 5272 1006 5276 1014
rect 5284 1006 5288 1014
rect 5296 1006 5300 1014
rect 5308 1006 5312 1014
rect 4842 656 4844 664
rect 4852 656 4854 664
rect 4842 654 4854 656
rect 4682 536 4684 544
rect 4692 536 4694 544
rect 4682 534 4694 536
rect 5248 614 5312 1006
rect 5248 606 5252 614
rect 5260 606 5264 614
rect 5272 606 5276 614
rect 5284 606 5288 614
rect 5296 606 5300 614
rect 5308 606 5312 614
rect 4938 524 4950 526
rect 4938 516 4940 524
rect 4948 516 4950 524
rect 4490 216 4492 224
rect 4500 216 4502 224
rect 4490 214 4502 216
rect 4810 364 4822 366
rect 4810 356 4812 364
rect 4820 356 4822 364
rect 4394 156 4396 164
rect 4404 156 4406 164
rect 4394 154 4406 156
rect 4362 136 4364 144
rect 4372 136 4374 144
rect 4362 134 4374 136
rect 4810 124 4822 356
rect 4810 116 4812 124
rect 4820 116 4822 124
rect 4810 114 4822 116
rect 4938 124 4950 516
rect 4938 116 4940 124
rect 4948 116 4950 124
rect 4938 114 4950 116
rect 5248 214 5312 606
rect 5418 1224 5430 1226
rect 5418 1216 5420 1224
rect 5428 1216 5430 1224
rect 5248 206 5252 214
rect 5260 206 5264 214
rect 5272 206 5276 214
rect 5284 206 5288 214
rect 5296 206 5300 214
rect 5308 206 5312 214
rect 3744 6 3748 14
rect 3756 6 3760 14
rect 3768 6 3772 14
rect 3780 6 3784 14
rect 3792 6 3796 14
rect 3804 6 3808 14
rect 3744 -10 3808 6
rect 5248 -10 5312 206
rect 5354 544 5366 546
rect 5354 536 5356 544
rect 5364 536 5366 544
rect 5354 184 5366 536
rect 5354 176 5356 184
rect 5364 176 5366 184
rect 5354 174 5366 176
rect 5386 524 5398 526
rect 5386 516 5388 524
rect 5396 516 5398 524
rect 5386 144 5398 516
rect 5418 464 5430 1216
rect 5578 1024 5590 1276
rect 5578 1016 5580 1024
rect 5588 1016 5590 1024
rect 5578 1014 5590 1016
rect 5610 1124 5622 1126
rect 5610 1116 5612 1124
rect 5620 1116 5622 1124
rect 5610 904 5622 1116
rect 5610 896 5612 904
rect 5620 896 5622 904
rect 5610 894 5622 896
rect 5674 844 5686 1756
rect 5738 1264 5750 1266
rect 5738 1256 5740 1264
rect 5748 1256 5750 1264
rect 5738 1024 5750 1256
rect 5834 1124 5846 1816
rect 6282 1584 6294 2116
rect 6314 2124 6326 3076
rect 6410 2964 6422 3196
rect 6538 3284 6550 3286
rect 6538 3276 6540 3284
rect 6548 3276 6550 3284
rect 6474 3144 6486 3146
rect 6474 3136 6476 3144
rect 6484 3136 6486 3144
rect 6474 3024 6486 3136
rect 6474 3016 6476 3024
rect 6484 3016 6486 3024
rect 6474 3014 6486 3016
rect 6410 2956 6412 2964
rect 6420 2956 6422 2964
rect 6410 2954 6422 2956
rect 6410 2924 6422 2926
rect 6410 2916 6412 2924
rect 6420 2916 6422 2924
rect 6410 2704 6422 2916
rect 6410 2696 6412 2704
rect 6420 2696 6422 2704
rect 6410 2694 6422 2696
rect 6474 2584 6486 2586
rect 6474 2576 6476 2584
rect 6484 2576 6486 2584
rect 6314 2116 6316 2124
rect 6324 2116 6326 2124
rect 6314 2114 6326 2116
rect 6410 2544 6422 2546
rect 6410 2536 6412 2544
rect 6420 2536 6422 2544
rect 6410 1804 6422 2536
rect 6474 2544 6486 2576
rect 6474 2536 6476 2544
rect 6484 2536 6486 2544
rect 6474 2534 6486 2536
rect 6538 2484 6550 3276
rect 6570 2944 6582 3636
rect 6752 3614 6816 4006
rect 6954 3624 6966 4796
rect 7178 4764 7190 4766
rect 7178 4756 7180 4764
rect 7188 4756 7190 4764
rect 7178 4584 7190 4756
rect 7274 4764 7286 4766
rect 7274 4756 7276 4764
rect 7284 4756 7286 4764
rect 7178 4576 7180 4584
rect 7188 4576 7190 4584
rect 7178 4574 7190 4576
rect 7210 4604 7222 4606
rect 7210 4596 7212 4604
rect 7220 4596 7222 4604
rect 7210 3664 7222 4596
rect 7210 3656 7212 3664
rect 7220 3656 7222 3664
rect 7210 3654 7222 3656
rect 6954 3616 6956 3624
rect 6964 3616 6966 3624
rect 6954 3614 6966 3616
rect 6752 3606 6756 3614
rect 6764 3606 6768 3614
rect 6776 3606 6780 3614
rect 6788 3606 6792 3614
rect 6800 3606 6804 3614
rect 6812 3606 6816 3614
rect 6698 3304 6710 3306
rect 6698 3296 6700 3304
rect 6708 3296 6710 3304
rect 6570 2936 6572 2944
rect 6580 2936 6582 2944
rect 6570 2934 6582 2936
rect 6602 3084 6614 3086
rect 6602 3076 6604 3084
rect 6612 3076 6614 3084
rect 6602 2944 6614 3076
rect 6698 3044 6710 3296
rect 6698 3036 6700 3044
rect 6708 3036 6710 3044
rect 6698 3034 6710 3036
rect 6752 3214 6816 3606
rect 7274 3584 7286 4756
rect 7306 4604 7318 4996
rect 7306 4596 7308 4604
rect 7316 4596 7318 4604
rect 7306 4594 7318 4596
rect 7274 3576 7276 3584
rect 7284 3576 7286 3584
rect 7274 3574 7286 3576
rect 7306 3884 7318 3886
rect 7306 3876 7308 3884
rect 7316 3876 7318 3884
rect 7082 3564 7094 3566
rect 7082 3556 7084 3564
rect 7092 3556 7094 3564
rect 6752 3206 6756 3214
rect 6764 3206 6768 3214
rect 6776 3206 6780 3214
rect 6788 3206 6792 3214
rect 6800 3206 6804 3214
rect 6812 3206 6816 3214
rect 6602 2936 6604 2944
rect 6612 2936 6614 2944
rect 6602 2934 6614 2936
rect 6634 3024 6646 3026
rect 6634 3016 6636 3024
rect 6644 3016 6646 3024
rect 6570 2904 6582 2906
rect 6570 2896 6572 2904
rect 6580 2896 6582 2904
rect 6570 2724 6582 2896
rect 6634 2904 6646 3016
rect 6634 2896 6636 2904
rect 6644 2896 6646 2904
rect 6634 2894 6646 2896
rect 6570 2716 6572 2724
rect 6580 2716 6582 2724
rect 6570 2714 6582 2716
rect 6602 2844 6614 2846
rect 6602 2836 6604 2844
rect 6612 2836 6614 2844
rect 6538 2476 6540 2484
rect 6548 2476 6550 2484
rect 6538 2474 6550 2476
rect 6570 2144 6582 2146
rect 6570 2136 6572 2144
rect 6580 2136 6582 2144
rect 6410 1796 6412 1804
rect 6420 1796 6422 1804
rect 6410 1794 6422 1796
rect 6474 2104 6486 2106
rect 6474 2096 6476 2104
rect 6484 2096 6486 2104
rect 6474 1726 6486 2096
rect 6474 1714 6518 1726
rect 6282 1576 6284 1584
rect 6292 1576 6294 1584
rect 6282 1574 6294 1576
rect 5834 1116 5836 1124
rect 5844 1116 5846 1124
rect 5834 1114 5846 1116
rect 5962 1324 5974 1326
rect 5962 1316 5964 1324
rect 5972 1316 5974 1324
rect 5738 1016 5740 1024
rect 5748 1016 5750 1024
rect 5738 1014 5750 1016
rect 5962 1044 5974 1316
rect 6250 1324 6262 1326
rect 6250 1316 6252 1324
rect 6260 1316 6262 1324
rect 5962 1036 5964 1044
rect 5972 1036 5974 1044
rect 5674 836 5676 844
rect 5684 836 5686 844
rect 5674 834 5686 836
rect 5770 864 5782 866
rect 5770 856 5772 864
rect 5780 856 5782 864
rect 5770 664 5782 856
rect 5770 656 5772 664
rect 5780 656 5782 664
rect 5770 654 5782 656
rect 5962 624 5974 1036
rect 6218 1104 6230 1106
rect 6218 1096 6220 1104
rect 6228 1096 6230 1104
rect 6090 964 6102 966
rect 6090 956 6092 964
rect 6100 956 6102 964
rect 6090 884 6102 956
rect 6090 876 6092 884
rect 6100 876 6102 884
rect 6090 874 6102 876
rect 6154 964 6166 966
rect 6154 956 6156 964
rect 6164 956 6166 964
rect 6154 704 6166 956
rect 6154 696 6156 704
rect 6164 696 6166 704
rect 6154 694 6166 696
rect 6218 744 6230 1096
rect 6250 1084 6262 1316
rect 6250 1076 6252 1084
rect 6260 1076 6262 1084
rect 6250 1074 6262 1076
rect 6506 764 6518 1714
rect 6570 1284 6582 2136
rect 6602 1784 6614 2836
rect 6666 2824 6678 2826
rect 6666 2816 6668 2824
rect 6676 2816 6678 2824
rect 6634 2644 6646 2646
rect 6634 2636 6636 2644
rect 6644 2636 6646 2644
rect 6634 2144 6646 2636
rect 6666 2444 6678 2816
rect 6666 2436 6668 2444
rect 6676 2436 6678 2444
rect 6666 2434 6678 2436
rect 6752 2814 6816 3206
rect 6858 3524 6870 3526
rect 6858 3516 6860 3524
rect 6868 3516 6870 3524
rect 6858 2944 6870 3516
rect 6986 3364 6998 3366
rect 6986 3356 6988 3364
rect 6996 3356 6998 3364
rect 6922 3224 6934 3226
rect 6922 3216 6924 3224
rect 6932 3216 6934 3224
rect 6922 3084 6934 3216
rect 6986 3204 6998 3356
rect 6986 3196 6988 3204
rect 6996 3196 6998 3204
rect 6986 3194 6998 3196
rect 6922 3076 6924 3084
rect 6932 3076 6934 3084
rect 6922 3074 6934 3076
rect 6954 3184 6966 3186
rect 6954 3176 6956 3184
rect 6964 3176 6966 3184
rect 6858 2936 6860 2944
rect 6868 2936 6870 2944
rect 6858 2934 6870 2936
rect 6890 3064 6902 3066
rect 6890 3056 6892 3064
rect 6900 3056 6902 3064
rect 6752 2806 6756 2814
rect 6764 2806 6768 2814
rect 6776 2806 6780 2814
rect 6788 2806 6792 2814
rect 6800 2806 6804 2814
rect 6812 2806 6816 2814
rect 6634 2136 6636 2144
rect 6644 2136 6646 2144
rect 6634 2134 6646 2136
rect 6752 2414 6816 2806
rect 6890 2704 6902 3056
rect 6954 2964 6966 3176
rect 6954 2956 6956 2964
rect 6964 2956 6966 2964
rect 6954 2954 6966 2956
rect 7018 3184 7030 3186
rect 7018 3176 7020 3184
rect 7028 3176 7030 3184
rect 6890 2696 6892 2704
rect 6900 2696 6902 2704
rect 6890 2694 6902 2696
rect 6752 2406 6756 2414
rect 6764 2406 6768 2414
rect 6776 2406 6780 2414
rect 6788 2406 6792 2414
rect 6800 2406 6804 2414
rect 6812 2406 6816 2414
rect 6602 1776 6604 1784
rect 6612 1776 6614 1784
rect 6602 1774 6614 1776
rect 6752 2014 6816 2406
rect 6890 2664 6902 2666
rect 6890 2656 6892 2664
rect 6900 2656 6902 2664
rect 6890 2044 6902 2656
rect 6986 2544 6998 2546
rect 6986 2536 6988 2544
rect 6996 2536 6998 2544
rect 6954 2524 6966 2526
rect 6954 2516 6956 2524
rect 6964 2516 6966 2524
rect 6890 2036 6892 2044
rect 6900 2036 6902 2044
rect 6890 2034 6902 2036
rect 6922 2264 6934 2266
rect 6922 2256 6924 2264
rect 6932 2256 6934 2264
rect 6752 2006 6756 2014
rect 6764 2006 6768 2014
rect 6776 2006 6780 2014
rect 6788 2006 6792 2014
rect 6800 2006 6804 2014
rect 6812 2006 6816 2014
rect 6752 1614 6816 2006
rect 6922 1964 6934 2256
rect 6922 1956 6924 1964
rect 6932 1956 6934 1964
rect 6922 1954 6934 1956
rect 6954 1864 6966 2516
rect 6986 1884 6998 2536
rect 7018 1964 7030 3176
rect 7082 3144 7094 3556
rect 7210 3444 7222 3446
rect 7210 3436 7212 3444
rect 7220 3436 7222 3444
rect 7082 3136 7084 3144
rect 7092 3136 7094 3144
rect 7082 3134 7094 3136
rect 7178 3344 7190 3346
rect 7178 3336 7180 3344
rect 7188 3336 7190 3344
rect 7178 3064 7190 3336
rect 7178 3056 7180 3064
rect 7188 3056 7190 3064
rect 7178 3054 7190 3056
rect 7114 3024 7126 3026
rect 7114 3016 7116 3024
rect 7124 3016 7126 3024
rect 7114 2964 7126 3016
rect 7114 2956 7116 2964
rect 7124 2956 7126 2964
rect 7114 2954 7126 2956
rect 7082 2844 7094 2846
rect 7082 2836 7084 2844
rect 7092 2836 7094 2844
rect 7050 2504 7062 2506
rect 7050 2496 7052 2504
rect 7060 2496 7062 2504
rect 7050 2104 7062 2496
rect 7082 2304 7094 2836
rect 7146 2804 7158 2806
rect 7146 2796 7148 2804
rect 7156 2796 7158 2804
rect 7146 2464 7158 2796
rect 7178 2744 7190 2746
rect 7178 2736 7180 2744
rect 7188 2736 7190 2744
rect 7178 2564 7190 2736
rect 7178 2556 7180 2564
rect 7188 2556 7190 2564
rect 7178 2554 7190 2556
rect 7146 2456 7148 2464
rect 7156 2456 7158 2464
rect 7146 2454 7158 2456
rect 7178 2464 7190 2466
rect 7178 2456 7180 2464
rect 7188 2456 7190 2464
rect 7082 2296 7084 2304
rect 7092 2296 7094 2304
rect 7082 2294 7094 2296
rect 7114 2324 7126 2326
rect 7114 2316 7116 2324
rect 7124 2316 7126 2324
rect 7050 2096 7052 2104
rect 7060 2096 7062 2104
rect 7050 2094 7062 2096
rect 7082 2264 7094 2266
rect 7082 2256 7084 2264
rect 7092 2256 7094 2264
rect 7018 1956 7020 1964
rect 7028 1956 7030 1964
rect 7018 1954 7030 1956
rect 6986 1876 6988 1884
rect 6996 1876 6998 1884
rect 6986 1874 6998 1876
rect 6954 1856 6956 1864
rect 6964 1856 6966 1864
rect 6752 1606 6756 1614
rect 6764 1606 6768 1614
rect 6776 1606 6780 1614
rect 6788 1606 6792 1614
rect 6800 1606 6804 1614
rect 6812 1606 6816 1614
rect 6570 1276 6572 1284
rect 6580 1276 6582 1284
rect 6570 1274 6582 1276
rect 6634 1284 6646 1286
rect 6634 1276 6636 1284
rect 6644 1276 6646 1284
rect 6506 756 6508 764
rect 6516 756 6518 764
rect 6506 754 6518 756
rect 6538 1204 6550 1206
rect 6538 1196 6540 1204
rect 6548 1196 6550 1204
rect 6218 736 6220 744
rect 6228 736 6230 744
rect 6218 704 6230 736
rect 6218 696 6220 704
rect 6228 696 6230 704
rect 6218 694 6230 696
rect 5962 616 5964 624
rect 5972 616 5974 624
rect 5962 614 5974 616
rect 5418 456 5420 464
rect 5428 456 5430 464
rect 5418 454 5430 456
rect 5610 544 5622 546
rect 5610 536 5612 544
rect 5620 536 5622 544
rect 5610 324 5622 536
rect 5610 316 5612 324
rect 5620 316 5622 324
rect 5610 314 5622 316
rect 5674 364 5686 366
rect 5674 356 5676 364
rect 5684 356 5686 364
rect 5386 136 5388 144
rect 5396 136 5398 144
rect 5386 134 5398 136
rect 5674 24 5686 356
rect 6538 304 6550 1196
rect 6634 564 6646 1276
rect 6752 1214 6816 1606
rect 6922 1704 6934 1706
rect 6922 1696 6924 1704
rect 6932 1696 6934 1704
rect 6922 1404 6934 1696
rect 6954 1444 6966 1856
rect 7050 1704 7062 1706
rect 7050 1696 7052 1704
rect 7060 1696 7062 1704
rect 6954 1436 6956 1444
rect 6964 1436 6966 1444
rect 6954 1434 6966 1436
rect 6986 1444 6998 1446
rect 6986 1436 6988 1444
rect 6996 1436 6998 1444
rect 6922 1396 6924 1404
rect 6932 1396 6934 1404
rect 6922 1394 6934 1396
rect 6954 1404 6966 1406
rect 6954 1396 6956 1404
rect 6964 1396 6966 1404
rect 6752 1206 6756 1214
rect 6764 1206 6768 1214
rect 6776 1206 6780 1214
rect 6788 1206 6792 1214
rect 6800 1206 6804 1214
rect 6812 1206 6816 1214
rect 6698 1084 6710 1086
rect 6698 1076 6700 1084
rect 6708 1076 6710 1084
rect 6698 1044 6710 1076
rect 6698 1036 6700 1044
rect 6708 1036 6710 1044
rect 6698 1034 6710 1036
rect 6698 984 6710 986
rect 6698 976 6700 984
rect 6708 976 6710 984
rect 6698 804 6710 976
rect 6698 796 6700 804
rect 6708 796 6710 804
rect 6698 794 6710 796
rect 6752 814 6816 1206
rect 6954 844 6966 1396
rect 6954 836 6956 844
rect 6964 836 6966 844
rect 6954 834 6966 836
rect 6752 806 6756 814
rect 6764 806 6768 814
rect 6776 806 6780 814
rect 6788 806 6792 814
rect 6800 806 6804 814
rect 6812 806 6816 814
rect 6634 556 6636 564
rect 6644 556 6646 564
rect 6634 554 6646 556
rect 6538 296 6540 304
rect 6548 296 6550 304
rect 6538 294 6550 296
rect 6752 414 6816 806
rect 6986 724 6998 1436
rect 7050 1444 7062 1696
rect 7050 1436 7052 1444
rect 7060 1436 7062 1444
rect 7050 1434 7062 1436
rect 7082 1284 7094 2256
rect 7114 2124 7126 2316
rect 7114 2116 7116 2124
rect 7124 2116 7126 2124
rect 7114 2114 7126 2116
rect 7146 2124 7158 2126
rect 7146 2116 7148 2124
rect 7156 2116 7158 2124
rect 7114 2084 7126 2086
rect 7114 2076 7116 2084
rect 7124 2076 7126 2084
rect 7114 1824 7126 2076
rect 7114 1816 7116 1824
rect 7124 1816 7126 1824
rect 7114 1814 7126 1816
rect 7114 1764 7126 1766
rect 7114 1756 7116 1764
rect 7124 1756 7126 1764
rect 7114 1464 7126 1756
rect 7114 1456 7116 1464
rect 7124 1456 7126 1464
rect 7114 1454 7126 1456
rect 7082 1276 7084 1284
rect 7092 1276 7094 1284
rect 7082 1274 7094 1276
rect 7082 1124 7094 1126
rect 7082 1116 7084 1124
rect 7092 1116 7094 1124
rect 7082 1024 7094 1116
rect 7082 1016 7084 1024
rect 7092 1016 7094 1024
rect 7082 1014 7094 1016
rect 6986 716 6988 724
rect 6996 716 6998 724
rect 6986 714 6998 716
rect 6752 406 6756 414
rect 6764 406 6768 414
rect 6776 406 6780 414
rect 6788 406 6792 414
rect 6800 406 6804 414
rect 6812 406 6816 414
rect 5674 16 5676 24
rect 5684 16 5686 24
rect 5674 14 5686 16
rect 6752 14 6816 406
rect 7146 284 7158 2116
rect 7178 1404 7190 2456
rect 7210 2224 7222 3436
rect 7274 3324 7286 3326
rect 7274 3316 7276 3324
rect 7284 3316 7286 3324
rect 7242 3304 7254 3306
rect 7242 3296 7244 3304
rect 7252 3296 7254 3304
rect 7242 2924 7254 3296
rect 7242 2916 7244 2924
rect 7252 2916 7254 2924
rect 7242 2914 7254 2916
rect 7274 2704 7286 3316
rect 7274 2696 7276 2704
rect 7284 2696 7286 2704
rect 7274 2694 7286 2696
rect 7210 2216 7212 2224
rect 7220 2216 7222 2224
rect 7210 2214 7222 2216
rect 7242 2684 7254 2686
rect 7242 2676 7244 2684
rect 7252 2676 7254 2684
rect 7242 2544 7254 2676
rect 7242 2536 7244 2544
rect 7252 2536 7254 2544
rect 7210 1884 7222 1886
rect 7210 1876 7212 1884
rect 7220 1876 7222 1884
rect 7210 1704 7222 1876
rect 7242 1764 7254 2536
rect 7274 2344 7286 2346
rect 7274 2336 7276 2344
rect 7284 2336 7286 2344
rect 7274 1904 7286 2336
rect 7274 1896 7276 1904
rect 7284 1896 7286 1904
rect 7274 1894 7286 1896
rect 7242 1756 7244 1764
rect 7252 1756 7254 1764
rect 7242 1754 7254 1756
rect 7210 1696 7212 1704
rect 7220 1696 7222 1704
rect 7210 1694 7222 1696
rect 7178 1396 7180 1404
rect 7188 1396 7190 1404
rect 7178 1394 7190 1396
rect 7274 1644 7286 1646
rect 7274 1636 7276 1644
rect 7284 1636 7286 1644
rect 7178 1364 7190 1366
rect 7178 1356 7180 1364
rect 7188 1356 7190 1364
rect 7178 1304 7190 1356
rect 7178 1296 7180 1304
rect 7188 1296 7190 1304
rect 7178 1294 7190 1296
rect 7242 944 7254 946
rect 7242 936 7244 944
rect 7252 936 7254 944
rect 7242 524 7254 936
rect 7274 884 7286 1636
rect 7306 1084 7318 3876
rect 7338 3624 7350 5056
rect 7530 5064 7542 5066
rect 7530 5056 7532 5064
rect 7540 5056 7542 5064
rect 7466 4924 7478 4926
rect 7466 4916 7468 4924
rect 7476 4916 7478 4924
rect 7402 4724 7414 4726
rect 7402 4716 7404 4724
rect 7412 4716 7414 4724
rect 7370 4324 7382 4326
rect 7370 4316 7372 4324
rect 7380 4316 7382 4324
rect 7370 3764 7382 4316
rect 7402 3944 7414 4716
rect 7434 4724 7446 4726
rect 7434 4716 7436 4724
rect 7444 4716 7446 4724
rect 7434 4164 7446 4716
rect 7434 4156 7436 4164
rect 7444 4156 7446 4164
rect 7434 4154 7446 4156
rect 7402 3936 7404 3944
rect 7412 3936 7414 3944
rect 7402 3934 7414 3936
rect 7434 3944 7446 3946
rect 7434 3936 7436 3944
rect 7444 3936 7446 3944
rect 7370 3756 7372 3764
rect 7380 3756 7382 3764
rect 7370 3754 7382 3756
rect 7402 3904 7414 3906
rect 7402 3896 7404 3904
rect 7412 3896 7414 3904
rect 7338 3616 7340 3624
rect 7348 3616 7350 3624
rect 7338 3614 7350 3616
rect 7370 3724 7382 3726
rect 7370 3716 7372 3724
rect 7380 3716 7382 3724
rect 7338 3364 7350 3366
rect 7338 3356 7340 3364
rect 7348 3356 7350 3364
rect 7338 2844 7350 3356
rect 7338 2836 7340 2844
rect 7348 2836 7350 2844
rect 7338 2834 7350 2836
rect 7370 2944 7382 3716
rect 7402 3704 7414 3896
rect 7402 3696 7404 3704
rect 7412 3696 7414 3704
rect 7402 3694 7414 3696
rect 7434 3684 7446 3936
rect 7434 3676 7436 3684
rect 7444 3676 7446 3684
rect 7434 3674 7446 3676
rect 7402 3664 7414 3666
rect 7402 3656 7404 3664
rect 7412 3656 7414 3664
rect 7402 3344 7414 3656
rect 7434 3644 7446 3646
rect 7434 3636 7436 3644
rect 7444 3636 7446 3644
rect 7434 3384 7446 3636
rect 7434 3376 7436 3384
rect 7444 3376 7446 3384
rect 7434 3374 7446 3376
rect 7402 3336 7404 3344
rect 7412 3336 7414 3344
rect 7402 3334 7414 3336
rect 7370 2936 7372 2944
rect 7380 2936 7382 2944
rect 7370 2584 7382 2936
rect 7402 3104 7414 3106
rect 7402 3096 7404 3104
rect 7412 3096 7414 3104
rect 7402 2604 7414 3096
rect 7402 2596 7404 2604
rect 7412 2596 7414 2604
rect 7402 2594 7414 2596
rect 7466 3084 7478 4916
rect 7498 4664 7510 4666
rect 7498 4656 7500 4664
rect 7508 4656 7510 4664
rect 7498 4184 7510 4656
rect 7498 4176 7500 4184
rect 7508 4176 7510 4184
rect 7498 4174 7510 4176
rect 7498 4044 7510 4046
rect 7498 4036 7500 4044
rect 7508 4036 7510 4044
rect 7498 3324 7510 4036
rect 7498 3316 7500 3324
rect 7508 3316 7510 3324
rect 7498 3314 7510 3316
rect 7466 3076 7468 3084
rect 7476 3076 7478 3084
rect 7466 2684 7478 3076
rect 7498 3184 7510 3186
rect 7498 3176 7500 3184
rect 7508 3176 7510 3184
rect 7498 2844 7510 3176
rect 7498 2836 7500 2844
rect 7508 2836 7510 2844
rect 7498 2834 7510 2836
rect 7466 2676 7468 2684
rect 7476 2676 7478 2684
rect 7370 2576 7372 2584
rect 7380 2576 7382 2584
rect 7306 1076 7308 1084
rect 7316 1076 7318 1084
rect 7306 1074 7318 1076
rect 7338 2564 7350 2566
rect 7338 2556 7340 2564
rect 7348 2556 7350 2564
rect 7338 1484 7350 2556
rect 7338 1476 7340 1484
rect 7348 1476 7350 1484
rect 7274 876 7276 884
rect 7284 876 7286 884
rect 7274 874 7286 876
rect 7242 516 7244 524
rect 7252 516 7254 524
rect 7242 514 7254 516
rect 7146 276 7148 284
rect 7156 276 7158 284
rect 7146 274 7158 276
rect 7338 124 7350 1476
rect 7370 1524 7382 2576
rect 7434 2544 7446 2546
rect 7434 2536 7436 2544
rect 7444 2536 7446 2544
rect 7434 1704 7446 2536
rect 7434 1696 7436 1704
rect 7444 1696 7446 1704
rect 7434 1694 7446 1696
rect 7466 2264 7478 2676
rect 7498 2764 7510 2766
rect 7498 2756 7500 2764
rect 7508 2756 7510 2764
rect 7498 2304 7510 2756
rect 7530 2684 7542 5056
rect 7530 2676 7532 2684
rect 7540 2676 7542 2684
rect 7530 2674 7542 2676
rect 7562 4964 7574 4966
rect 7562 4956 7564 4964
rect 7572 4956 7574 4964
rect 7530 2644 7542 2646
rect 7530 2636 7532 2644
rect 7540 2636 7542 2644
rect 7530 2524 7542 2636
rect 7562 2564 7574 4956
rect 7562 2556 7564 2564
rect 7572 2556 7574 2564
rect 7562 2554 7574 2556
rect 7530 2516 7532 2524
rect 7540 2516 7542 2524
rect 7530 2514 7542 2516
rect 7498 2296 7500 2304
rect 7508 2296 7510 2304
rect 7498 2294 7510 2296
rect 7530 2404 7542 2406
rect 7530 2396 7532 2404
rect 7540 2396 7542 2404
rect 7466 2256 7468 2264
rect 7476 2256 7478 2264
rect 7370 1516 7372 1524
rect 7380 1516 7382 1524
rect 7370 584 7382 1516
rect 7434 1104 7446 1106
rect 7434 1096 7436 1104
rect 7444 1096 7446 1104
rect 7434 744 7446 1096
rect 7434 736 7436 744
rect 7444 736 7446 744
rect 7434 734 7446 736
rect 7370 576 7372 584
rect 7380 576 7382 584
rect 7370 574 7382 576
rect 7466 144 7478 2256
rect 7498 2184 7510 2186
rect 7498 2176 7500 2184
rect 7508 2176 7510 2184
rect 7498 1724 7510 2176
rect 7530 1884 7542 2396
rect 7530 1876 7532 1884
rect 7540 1876 7542 1884
rect 7530 1874 7542 1876
rect 7562 1964 7574 1966
rect 7562 1956 7564 1964
rect 7572 1956 7574 1964
rect 7498 1716 7500 1724
rect 7508 1716 7510 1724
rect 7498 1714 7510 1716
rect 7530 1784 7542 1786
rect 7530 1776 7532 1784
rect 7540 1776 7542 1784
rect 7498 1684 7510 1686
rect 7498 1676 7500 1684
rect 7508 1676 7510 1684
rect 7498 544 7510 1676
rect 7530 1504 7542 1776
rect 7530 1496 7532 1504
rect 7540 1496 7542 1504
rect 7530 1494 7542 1496
rect 7562 1104 7574 1956
rect 7562 1096 7564 1104
rect 7572 1096 7574 1104
rect 7562 1094 7574 1096
rect 7498 536 7500 544
rect 7508 536 7510 544
rect 7498 534 7510 536
rect 7530 1004 7542 1006
rect 7530 996 7532 1004
rect 7540 996 7542 1004
rect 7466 136 7468 144
rect 7476 136 7478 144
rect 7466 134 7478 136
rect 7338 116 7340 124
rect 7348 116 7350 124
rect 7338 114 7350 116
rect 7530 124 7542 996
rect 7530 116 7532 124
rect 7540 116 7542 124
rect 7530 114 7542 116
rect 6752 6 6756 14
rect 6764 6 6768 14
rect 6776 6 6780 14
rect 6788 6 6792 14
rect 6800 6 6804 14
rect 6812 6 6816 14
rect 6752 -10 6816 6
use AOI21X1  _3496_
timestamp 1597059762
transform 1 0 8 0 -1 210
box -4 -6 68 206
use NAND2X1  _3495_
timestamp 1597059762
transform -1 0 120 0 -1 210
box -4 -6 52 206
use AOI21X1  _3457_
timestamp 1597059762
transform -1 0 184 0 -1 210
box -4 -6 68 206
use NAND2X1  _3455_
timestamp 1597059762
transform -1 0 232 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3508_
timestamp 1597059762
transform 1 0 8 0 1 210
box -4 -6 196 206
use DFFPOSX1  _3518_
timestamp 1597059762
transform 1 0 200 0 1 210
box -4 -6 196 206
use NAND2X1  _3456_
timestamp 1597059762
transform -1 0 280 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3512_
timestamp 1597059762
transform 1 0 280 0 -1 210
box -4 -6 196 206
use INVX8  _3960_
timestamp 1597059762
transform 1 0 392 0 1 210
box -4 -6 84 206
use DFFPOSX1  _3510_
timestamp 1597059762
transform 1 0 472 0 -1 210
box -4 -6 196 206
use INVX8  _3439_
timestamp 1597059762
transform -1 0 552 0 1 210
box -4 -6 84 206
use AOI21X1  _3472_
timestamp 1597059762
transform -1 0 616 0 1 210
box -4 -6 68 206
use NAND2X1  _3470_
timestamp 1597059762
transform -1 0 712 0 1 210
box -4 -6 52 206
use NAND2X1  _3471_
timestamp 1597059762
transform -1 0 664 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert132
timestamp 1597059762
transform -1 0 712 0 -1 210
box -4 -6 52 206
use FILL  SFILL8080x2100
timestamp 1597059762
transform 1 0 808 0 1 210
box -4 -6 20 206
use FILL  SFILL7920x2100
timestamp 1597059762
transform 1 0 792 0 1 210
box -4 -6 20 206
use FILL  SFILL7760x2100
timestamp 1597059762
transform 1 0 776 0 1 210
box -4 -6 20 206
use FILL  SFILL7600x2100
timestamp 1597059762
transform 1 0 760 0 1 210
box -4 -6 20 206
use FILL  SFILL7600x100
timestamp 1597059762
transform -1 0 776 0 -1 210
box -4 -6 20 206
use FILL  SFILL7440x100
timestamp 1597059762
transform -1 0 760 0 -1 210
box -4 -6 20 206
use FILL  SFILL7280x100
timestamp 1597059762
transform -1 0 744 0 -1 210
box -4 -6 20 206
use FILL  SFILL7120x100
timestamp 1597059762
transform -1 0 728 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_insert131
timestamp 1597059762
transform -1 0 760 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3509_
timestamp 1597059762
transform 1 0 776 0 -1 210
box -4 -6 196 206
use NAND2X1  _3476_
timestamp 1597059762
transform -1 0 1016 0 -1 210
box -4 -6 52 206
use AOI21X1  _3478_
timestamp 1597059762
transform -1 0 888 0 1 210
box -4 -6 68 206
use AOI21X1  _3469_
timestamp 1597059762
transform -1 0 952 0 1 210
box -4 -6 68 206
use NAND2X1  _3468_
timestamp 1597059762
transform 1 0 952 0 1 210
box -4 -6 52 206
use NAND2X1  _3477_
timestamp 1597059762
transform -1 0 1048 0 1 210
box -4 -6 52 206
use NAND2X1  _3467_
timestamp 1597059762
transform -1 0 1064 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert134
timestamp 1597059762
transform 1 0 1064 0 -1 210
box -4 -6 52 206
use AOI21X1  _3484_
timestamp 1597059762
transform 1 0 1112 0 -1 210
box -4 -6 68 206
use NAND2X1  _3482_
timestamp 1597059762
transform 1 0 1176 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert200
timestamp 1597059762
transform 1 0 1048 0 1 210
box -4 -6 52 206
use NAND2X1  _3483_
timestamp 1597059762
transform -1 0 1144 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3502_
timestamp 1597059762
transform 1 0 1144 0 1 210
box -4 -6 196 206
use NAND2X1  _3473_
timestamp 1597059762
transform 1 0 1224 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3294_
timestamp 1597059762
transform -1 0 1464 0 -1 210
box -4 -6 196 206
use INVX1  _3403_
timestamp 1597059762
transform 1 0 1336 0 1 210
box -4 -6 36 206
use INVX1  _3389_
timestamp 1597059762
transform 1 0 1368 0 1 210
box -4 -6 36 206
use INVX1  _3410_
timestamp 1597059762
transform 1 0 1400 0 1 210
box -4 -6 36 206
use NOR2X1  _3288_
timestamp 1597059762
transform -1 0 1512 0 -1 210
box -4 -6 52 206
use INVX1  _3255_
timestamp 1597059762
transform 1 0 1512 0 -1 210
box -4 -6 36 206
use BUFX2  _2048_
timestamp 1597059762
transform -1 0 1592 0 -1 210
box -4 -6 52 206
use OAI21X1  _3260_
timestamp 1597059762
transform -1 0 1656 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_insert133
timestamp 1597059762
transform 1 0 1432 0 1 210
box -4 -6 52 206
use INVX1  _3312_
timestamp 1597059762
transform 1 0 1480 0 1 210
box -4 -6 36 206
use INVX1  _3354_
timestamp 1597059762
transform 1 0 1512 0 1 210
box -4 -6 36 206
use AOI21X1  _3475_
timestamp 1597059762
transform -1 0 1608 0 1 210
box -4 -6 68 206
use NAND2X1  _3474_
timestamp 1597059762
transform -1 0 1656 0 1 210
box -4 -6 52 206
use NOR2X1  _3289_
timestamp 1597059762
transform 1 0 1656 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3291_
timestamp 1597059762
transform 1 0 1704 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _3511_
timestamp 1597059762
transform 1 0 1656 0 1 210
box -4 -6 196 206
use DFFPOSX1  _3293_
timestamp 1597059762
transform 1 0 1896 0 -1 210
box -4 -6 196 206
use INVX1  _3274_
timestamp 1597059762
transform -1 0 1880 0 1 210
box -4 -6 36 206
use DFFPOSX1  _3290_
timestamp 1597059762
transform 1 0 1880 0 1 210
box -4 -6 196 206
use INVX1  _3276_
timestamp 1597059762
transform -1 0 2120 0 -1 210
box -4 -6 36 206
use INVX1  _3270_
timestamp 1597059762
transform -1 0 2152 0 -1 210
box -4 -6 36 206
use OR2X2  _3271_
timestamp 1597059762
transform 1 0 2152 0 -1 210
box -4 -6 68 206
use OAI21X1  _3275_
timestamp 1597059762
transform -1 0 2136 0 1 210
box -4 -6 68 206
use OAI21X1  _3259_
timestamp 1597059762
transform 1 0 2136 0 1 210
box -4 -6 68 206
use NOR2X1  _3258_
timestamp 1597059762
transform 1 0 2200 0 1 210
box -4 -6 52 206
use FILL  SFILL22800x2100
timestamp 1597059762
transform 1 0 2280 0 1 210
box -4 -6 20 206
use FILL  SFILL22640x2100
timestamp 1597059762
transform 1 0 2264 0 1 210
box -4 -6 20 206
use FILL  SFILL22480x2100
timestamp 1597059762
transform 1 0 2248 0 1 210
box -4 -6 20 206
use FILL  SFILL22800x100
timestamp 1597059762
transform -1 0 2296 0 -1 210
box -4 -6 20 206
use NAND3X1  _3273_
timestamp 1597059762
transform 1 0 2216 0 -1 210
box -4 -6 68 206
use FILL  SFILL22960x2100
timestamp 1597059762
transform 1 0 2296 0 1 210
box -4 -6 20 206
use FILL  SFILL23280x100
timestamp 1597059762
transform -1 0 2344 0 -1 210
box -4 -6 20 206
use FILL  SFILL23120x100
timestamp 1597059762
transform -1 0 2328 0 -1 210
box -4 -6 20 206
use FILL  SFILL22960x100
timestamp 1597059762
transform -1 0 2312 0 -1 210
box -4 -6 20 206
use OAI21X1  _3272_
timestamp 1597059762
transform -1 0 2376 0 1 210
box -4 -6 68 206
use OAI21X1  _3269_
timestamp 1597059762
transform 1 0 2344 0 -1 210
box -4 -6 68 206
use NAND2X1  _3265_
timestamp 1597059762
transform -1 0 2456 0 1 210
box -4 -6 52 206
use INVX1  _3263_
timestamp 1597059762
transform -1 0 2408 0 1 210
box -4 -6 36 206
use INVX1  _3268_
timestamp 1597059762
transform -1 0 2440 0 -1 210
box -4 -6 36 206
use OR2X2  _3282_
timestamp 1597059762
transform 1 0 2440 0 -1 210
box -4 -6 68 206
use BUFX2  _2049_
timestamp 1597059762
transform -1 0 2552 0 -1 210
box -4 -6 52 206
use NAND2X1  _3257_
timestamp 1597059762
transform 1 0 2552 0 -1 210
box -4 -6 52 206
use INVX1  _3256_
timestamp 1597059762
transform -1 0 2632 0 -1 210
box -4 -6 36 206
use OAI21X1  _3266_
timestamp 1597059762
transform 1 0 2456 0 1 210
box -4 -6 68 206
use NOR2X1  _3287_
timestamp 1597059762
transform 1 0 2520 0 1 210
box -4 -6 52 206
use AND2X2  _3281_
timestamp 1597059762
transform -1 0 2632 0 1 210
box -4 -6 68 206
use AND2X2  _3284_
timestamp 1597059762
transform 1 0 2632 0 -1 210
box -4 -6 68 206
use INVX1  _4332_
timestamp 1597059762
transform 1 0 2696 0 -1 210
box -4 -6 36 206
use NOR2X1  _4338_
timestamp 1597059762
transform 1 0 2728 0 -1 210
box -4 -6 52 206
use INVX1  _4333_
timestamp 1597059762
transform -1 0 2808 0 -1 210
box -4 -6 36 206
use NOR2X1  _4334_
timestamp 1597059762
transform -1 0 2856 0 -1 210
box -4 -6 52 206
use AOI21X1  _3283_
timestamp 1597059762
transform 1 0 2632 0 1 210
box -4 -6 68 206
use NOR2X1  _3280_
timestamp 1597059762
transform -1 0 2744 0 1 210
box -4 -6 52 206
use INVX1  _3278_
timestamp 1597059762
transform -1 0 2776 0 1 210
box -4 -6 36 206
use NAND2X1  _3279_
timestamp 1597059762
transform -1 0 2824 0 1 210
box -4 -6 52 206
use NOR2X1  _4337_
timestamp 1597059762
transform 1 0 2856 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _4452_
timestamp 1597059762
transform 1 0 2904 0 -1 210
box -4 -6 196 206
use OR2X2  _3277_
timestamp 1597059762
transform -1 0 2888 0 1 210
box -4 -6 68 206
use AOI22X1  _4435_
timestamp 1597059762
transform 1 0 2888 0 1 210
box -4 -6 84 206
use AOI21X1  _4436_
timestamp 1597059762
transform 1 0 2968 0 1 210
box -4 -6 68 206
use INVX1  _4432_
timestamp 1597059762
transform 1 0 3096 0 -1 210
box -4 -6 36 206
use INVX1  _2095_
timestamp 1597059762
transform 1 0 3128 0 -1 210
box -4 -6 36 206
use OAI21X1  _2097_
timestamp 1597059762
transform 1 0 3160 0 -1 210
box -4 -6 68 206
use NAND3X1  _4434_
timestamp 1597059762
transform 1 0 3032 0 1 210
box -4 -6 68 206
use NAND3X1  _4431_
timestamp 1597059762
transform 1 0 3096 0 1 210
box -4 -6 68 206
use NAND2X1  _4433_
timestamp 1597059762
transform 1 0 3160 0 1 210
box -4 -6 52 206
use NAND2X1  _2096_
timestamp 1597059762
transform -1 0 3256 0 1 210
box -4 -6 52 206
use BUFX2  _2031_
timestamp 1597059762
transform 1 0 3224 0 -1 210
box -4 -6 52 206
use BUFX2  _2029_
timestamp 1597059762
transform 1 0 3272 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert186
timestamp 1597059762
transform 1 0 3320 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _4448_
timestamp 1597059762
transform 1 0 3368 0 -1 210
box -4 -6 196 206
use OAI21X1  _2091_
timestamp 1597059762
transform 1 0 3256 0 1 210
box -4 -6 68 206
use NAND2X1  _2090_
timestamp 1597059762
transform -1 0 3368 0 1 210
box -4 -6 52 206
use AOI21X1  _4410_
timestamp 1597059762
transform 1 0 3368 0 1 210
box -4 -6 68 206
use BUFX2  _2027_
timestamp 1597059762
transform -1 0 3608 0 -1 210
box -4 -6 52 206
use BUFX2  _2030_
timestamp 1597059762
transform 1 0 3608 0 -1 210
box -4 -6 52 206
use AOI22X1  _4409_
timestamp 1597059762
transform 1 0 3432 0 1 210
box -4 -6 84 206
use INVX1  _2092_
timestamp 1597059762
transform -1 0 3544 0 1 210
box -4 -6 36 206
use INVX1  _2083_
timestamp 1597059762
transform 1 0 3544 0 1 210
box -4 -6 36 206
use OAI21X1  _2085_
timestamp 1597059762
transform 1 0 3576 0 1 210
box -4 -6 68 206
use DFFPOSX1  _4446_
timestamp 1597059762
transform 1 0 3656 0 -1 210
box -4 -6 196 206
use OAI21X1  _2094_
timestamp 1597059762
transform 1 0 3640 0 1 210
box -4 -6 68 206
use INVX1  _4406_
timestamp 1597059762
transform -1 0 3736 0 1 210
box -4 -6 36 206
use AND2X2  _4398_
timestamp 1597059762
transform -1 0 3864 0 1 210
box -4 -6 68 206
use FILL  SFILL37360x2100
timestamp 1597059762
transform 1 0 3736 0 1 210
box -4 -6 20 206
use FILL  SFILL37520x2100
timestamp 1597059762
transform 1 0 3752 0 1 210
box -4 -6 20 206
use FILL  SFILL37680x2100
timestamp 1597059762
transform 1 0 3768 0 1 210
box -4 -6 20 206
use FILL  SFILL37840x2100
timestamp 1597059762
transform 1 0 3784 0 1 210
box -4 -6 20 206
use FILL  SFILL38800x100
timestamp 1597059762
transform -1 0 3896 0 -1 210
box -4 -6 20 206
use FILL  SFILL38640x100
timestamp 1597059762
transform -1 0 3880 0 -1 210
box -4 -6 20 206
use FILL  SFILL38480x100
timestamp 1597059762
transform -1 0 3864 0 -1 210
box -4 -6 20 206
use NAND3X1  _4405_
timestamp 1597059762
transform 1 0 3864 0 1 210
box -4 -6 68 206
use FILL  SFILL38960x100
timestamp 1597059762
transform -1 0 3912 0 -1 210
box -4 -6 20 206
use OAI21X1  _4397_
timestamp 1597059762
transform -1 0 3992 0 1 210
box -4 -6 68 206
use OAI21X1  _2079_
timestamp 1597059762
transform 1 0 3944 0 -1 210
box -4 -6 68 206
use INVX1  _2077_
timestamp 1597059762
transform 1 0 3912 0 -1 210
box -4 -6 36 206
use NAND2X1  _2078_
timestamp 1597059762
transform -1 0 4040 0 1 210
box -4 -6 52 206
use BUFX2  _2026_
timestamp 1597059762
transform 1 0 4008 0 -1 210
box -4 -6 52 206
use BUFX2  _2025_
timestamp 1597059762
transform 1 0 4056 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _4445_
timestamp 1597059762
transform 1 0 4104 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert187
timestamp 1597059762
transform -1 0 4088 0 1 210
box -4 -6 52 206
use OAI21X1  _4395_
timestamp 1597059762
transform -1 0 4152 0 1 210
box -4 -6 68 206
use NAND3X1  _4399_
timestamp 1597059762
transform 1 0 4152 0 1 210
box -4 -6 68 206
use INVX1  _4393_
timestamp 1597059762
transform 1 0 4216 0 1 210
box -4 -6 36 206
use AOI22X1  _4391_
timestamp 1597059762
transform 1 0 4296 0 -1 210
box -4 -6 84 206
use AOI21X1  _4392_
timestamp 1597059762
transform -1 0 4440 0 -1 210
box -4 -6 68 206
use OAI21X1  _4401_
timestamp 1597059762
transform 1 0 4248 0 1 210
box -4 -6 68 206
use INVX1  _4400_
timestamp 1597059762
transform -1 0 4344 0 1 210
box -4 -6 36 206
use NOR3X1  _4394_
timestamp 1597059762
transform 1 0 4344 0 1 210
box -4 -6 132 206
use INVX1  _4389_
timestamp 1597059762
transform 1 0 4440 0 -1 210
box -4 -6 36 206
use NAND3X1  _4390_
timestamp 1597059762
transform -1 0 4536 0 -1 210
box -4 -6 68 206
use OAI21X1  _4387_
timestamp 1597059762
transform -1 0 4600 0 -1 210
box -4 -6 68 206
use INVX1  _4380_
timestamp 1597059762
transform -1 0 4632 0 -1 210
box -4 -6 36 206
use NAND3X1  _4383_
timestamp 1597059762
transform 1 0 4472 0 1 210
box -4 -6 68 206
use NAND3X1  _4382_
timestamp 1597059762
transform -1 0 4600 0 1 210
box -4 -6 68 206
use OAI21X1  _4381_
timestamp 1597059762
transform -1 0 4664 0 1 210
box -4 -6 68 206
use NOR3X1  _4388_
timestamp 1597059762
transform 1 0 4632 0 -1 210
box -4 -6 132 206
use INVX1  _4386_
timestamp 1597059762
transform -1 0 4792 0 -1 210
box -4 -6 36 206
use INVX1  _2074_
timestamp 1597059762
transform 1 0 4792 0 -1 210
box -4 -6 36 206
use INVX1  _4374_
timestamp 1597059762
transform 1 0 4664 0 1 210
box -4 -6 36 206
use INVX1  _4370_
timestamp 1597059762
transform 1 0 4696 0 1 210
box -4 -6 36 206
use NAND3X1  _4371_
timestamp 1597059762
transform 1 0 4728 0 1 210
box -4 -6 68 206
use INVX1  _4367_
timestamp 1597059762
transform 1 0 4792 0 1 210
box -4 -6 36 206
use OAI21X1  _2076_
timestamp 1597059762
transform -1 0 4888 0 -1 210
box -4 -6 68 206
use BUFX2  _2024_
timestamp 1597059762
transform 1 0 4888 0 -1 210
box -4 -6 52 206
use AOI22X1  _4378_
timestamp 1597059762
transform 1 0 4936 0 -1 210
box -4 -6 84 206
use NAND3X1  _4377_
timestamp 1597059762
transform -1 0 5080 0 -1 210
box -4 -6 68 206
use OAI21X1  _4368_
timestamp 1597059762
transform -1 0 4888 0 1 210
box -4 -6 68 206
use NOR3X1  _4369_
timestamp 1597059762
transform 1 0 4888 0 1 210
box -4 -6 132 206
use OAI21X1  _4375_
timestamp 1597059762
transform -1 0 5080 0 1 210
box -4 -6 68 206
use AOI21X1  _4379_
timestamp 1597059762
transform 1 0 5080 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _4443_
timestamp 1597059762
transform 1 0 5144 0 -1 210
box -4 -6 196 206
use AOI22X1  _4365_
timestamp 1597059762
transform 1 0 5080 0 1 210
box -4 -6 84 206
use AOI21X1  _4366_
timestamp 1597059762
transform -1 0 5224 0 1 210
box -4 -6 68 206
use FILL  SFILL52880x2100
timestamp 1597059762
transform 1 0 5288 0 1 210
box -4 -6 20 206
use NAND3X1  _4364_
timestamp 1597059762
transform 1 0 5224 0 1 210
box -4 -6 68 206
use FILL  SFILL53360x2100
timestamp 1597059762
transform 1 0 5336 0 1 210
box -4 -6 20 206
use FILL  SFILL53200x2100
timestamp 1597059762
transform 1 0 5320 0 1 210
box -4 -6 20 206
use FILL  SFILL53040x2100
timestamp 1597059762
transform 1 0 5304 0 1 210
box -4 -6 20 206
use FILL  SFILL53520x100
timestamp 1597059762
transform -1 0 5368 0 -1 210
box -4 -6 20 206
use FILL  SFILL53360x100
timestamp 1597059762
transform -1 0 5352 0 -1 210
box -4 -6 20 206
use OAI21X1  _4361_
timestamp 1597059762
transform -1 0 5416 0 1 210
box -4 -6 68 206
use FILL  SFILL53840x100
timestamp 1597059762
transform -1 0 5400 0 -1 210
box -4 -6 20 206
use FILL  SFILL53680x100
timestamp 1597059762
transform -1 0 5384 0 -1 210
box -4 -6 20 206
use INVX1  _4363_
timestamp 1597059762
transform -1 0 5448 0 1 210
box -4 -6 36 206
use NAND3X1  _4376_
timestamp 1597059762
transform 1 0 5400 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _4441_
timestamp 1597059762
transform 1 0 5464 0 -1 210
box -4 -6 196 206
use NOR3X1  _4362_
timestamp 1597059762
transform 1 0 5448 0 1 210
box -4 -6 132 206
use INVX2  _4360_
timestamp 1597059762
transform -1 0 5608 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_insert185
timestamp 1597059762
transform -1 0 5656 0 1 210
box -4 -6 52 206
use BUFX2  _2028_
timestamp 1597059762
transform 1 0 5656 0 -1 210
box -4 -6 52 206
use BUFX2  _2019_
timestamp 1597059762
transform 1 0 5704 0 -1 210
box -4 -6 52 206
use BUFX2  _2017_
timestamp 1597059762
transform 1 0 5752 0 -1 210
box -4 -6 52 206
use BUFX2  _2016_
timestamp 1597059762
transform 1 0 5800 0 -1 210
box -4 -6 52 206
use INVX1  _2053_
timestamp 1597059762
transform 1 0 5656 0 1 210
box -4 -6 36 206
use OAI21X1  _2055_
timestamp 1597059762
transform -1 0 5752 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_insert183
timestamp 1597059762
transform 1 0 5752 0 1 210
box -4 -6 52 206
use INVX1  _3035_
timestamp 1597059762
transform -1 0 5832 0 1 210
box -4 -6 36 206
use INVX1  _2068_
timestamp 1597059762
transform 1 0 5848 0 -1 210
box -4 -6 36 206
use OAI21X1  _2070_
timestamp 1597059762
transform 1 0 5880 0 -1 210
box -4 -6 68 206
use INVX1  _2071_
timestamp 1597059762
transform 1 0 5944 0 -1 210
box -4 -6 36 206
use BUFX2  _2022_
timestamp 1597059762
transform 1 0 5976 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert184
timestamp 1597059762
transform 1 0 5832 0 1 210
box -4 -6 52 206
use NAND2X1  _2069_
timestamp 1597059762
transform 1 0 5880 0 1 210
box -4 -6 52 206
use NOR2X1  _2246_
timestamp 1597059762
transform 1 0 5928 0 1 210
box -4 -6 52 206
use NOR2X1  _2244_
timestamp 1597059762
transform -1 0 6024 0 1 210
box -4 -6 52 206
use INVX1  _2062_
timestamp 1597059762
transform 1 0 6024 0 -1 210
box -4 -6 36 206
use BUFX2  _2020_
timestamp 1597059762
transform -1 0 6104 0 -1 210
box -4 -6 52 206
use OAI21X1  _2064_
timestamp 1597059762
transform -1 0 6168 0 -1 210
box -4 -6 68 206
use OAI21X1  _2073_
timestamp 1597059762
transform -1 0 6232 0 -1 210
box -4 -6 68 206
use AND2X2  _2245_
timestamp 1597059762
transform -1 0 6088 0 1 210
box -4 -6 68 206
use NAND2X1  _2063_
timestamp 1597059762
transform -1 0 6136 0 1 210
box -4 -6 52 206
use INVX1  _2442_
timestamp 1597059762
transform -1 0 6168 0 1 210
box -4 -6 36 206
use NAND2X1  _2072_
timestamp 1597059762
transform -1 0 6216 0 1 210
box -4 -6 52 206
use INVX1  _2630_
timestamp 1597059762
transform 1 0 6216 0 1 210
box -4 -6 36 206
use INVX1  _2065_
timestamp 1597059762
transform 1 0 6232 0 -1 210
box -4 -6 36 206
use OAI21X1  _2067_
timestamp 1597059762
transform 1 0 6264 0 -1 210
box -4 -6 68 206
use BUFX2  _2023_
timestamp 1597059762
transform 1 0 6328 0 -1 210
box -4 -6 52 206
use BUFX2  _2021_
timestamp 1597059762
transform 1 0 6376 0 -1 210
box -4 -6 52 206
use NAND2X1  _2066_
timestamp 1597059762
transform 1 0 6248 0 1 210
box -4 -6 52 206
use XNOR2X1  _2435_
timestamp 1597059762
transform 1 0 6296 0 1 210
box -4 -6 116 206
use XNOR2X1  _2634_
timestamp 1597059762
transform 1 0 6408 0 1 210
box -4 -6 116 206
use BUFX2  _2037_
timestamp 1597059762
transform 1 0 6424 0 -1 210
box -4 -6 52 206
use XNOR2X1  _2635_
timestamp 1597059762
transform 1 0 6472 0 -1 210
box -4 -6 116 206
use BUFX2  _2036_
timestamp 1597059762
transform 1 0 6584 0 -1 210
box -4 -6 52 206
use NAND3X1  _2636_
timestamp 1597059762
transform 1 0 6520 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_insert147
timestamp 1597059762
transform 1 0 6584 0 1 210
box -4 -6 52 206
use INVX1  _2721_
timestamp 1597059762
transform 1 0 6712 0 1 210
box -4 -6 36 206
use INVX1  _2720_
timestamp 1597059762
transform 1 0 6680 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_insert137
timestamp 1597059762
transform 1 0 6632 0 1 210
box -4 -6 52 206
use AOI21X1  _2725_
timestamp 1597059762
transform 1 0 6712 0 -1 210
box -4 -6 68 206
use NAND2X1  _2746_
timestamp 1597059762
transform 1 0 6664 0 -1 210
box -4 -6 52 206
use INVX1  _2723_
timestamp 1597059762
transform 1 0 6632 0 -1 210
box -4 -6 36 206
use FILL  SFILL67920x2100
timestamp 1597059762
transform 1 0 6792 0 1 210
box -4 -6 20 206
use FILL  SFILL67760x2100
timestamp 1597059762
transform 1 0 6776 0 1 210
box -4 -6 20 206
use FILL  SFILL67600x2100
timestamp 1597059762
transform 1 0 6760 0 1 210
box -4 -6 20 206
use FILL  SFILL67440x2100
timestamp 1597059762
transform 1 0 6744 0 1 210
box -4 -6 20 206
use FILL  SFILL67920x100
timestamp 1597059762
transform -1 0 6808 0 -1 210
box -4 -6 20 206
use FILL  SFILL67760x100
timestamp 1597059762
transform -1 0 6792 0 -1 210
box -4 -6 20 206
use FILL  SFILL68240x100
timestamp 1597059762
transform -1 0 6840 0 -1 210
box -4 -6 20 206
use FILL  SFILL68080x100
timestamp 1597059762
transform -1 0 6824 0 -1 210
box -4 -6 20 206
use AOI22X1  _2722_
timestamp 1597059762
transform -1 0 6888 0 1 210
box -4 -6 84 206
use OAI21X1  _2747_
timestamp 1597059762
transform 1 0 6840 0 -1 210
box -4 -6 68 206
use AOI21X1  _2754_
timestamp 1597059762
transform 1 0 6904 0 -1 210
box -4 -6 68 206
use INVX1  _2748_
timestamp 1597059762
transform 1 0 6968 0 -1 210
box -4 -6 36 206
use NAND2X1  _2749_
timestamp 1597059762
transform -1 0 7048 0 -1 210
box -4 -6 52 206
use NOR2X1  _2724_
timestamp 1597059762
transform -1 0 6936 0 1 210
box -4 -6 52 206
use NAND2X1  _2745_
timestamp 1597059762
transform -1 0 6984 0 1 210
box -4 -6 52 206
use NAND3X1  _2726_
timestamp 1597059762
transform 1 0 6984 0 1 210
box -4 -6 68 206
use OAI21X1  _2753_
timestamp 1597059762
transform -1 0 7112 0 -1 210
box -4 -6 68 206
use NOR2X1  _2750_
timestamp 1597059762
transform -1 0 7160 0 -1 210
box -4 -6 52 206
use BUFX2  _2039_
timestamp 1597059762
transform -1 0 7208 0 -1 210
box -4 -6 52 206
use OR2X2  _2715_
timestamp 1597059762
transform 1 0 7208 0 -1 210
box -4 -6 68 206
use XNOR2X1  _2557_
timestamp 1597059762
transform 1 0 7048 0 1 210
box -4 -6 116 206
use NAND2X1  _2559_
timestamp 1597059762
transform 1 0 7160 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert135
timestamp 1597059762
transform 1 0 7208 0 1 210
box -4 -6 52 206
use NAND2X1  _2752_
timestamp 1597059762
transform -1 0 7320 0 -1 210
box -4 -6 52 206
use INVX1  _2751_
timestamp 1597059762
transform -1 0 7352 0 -1 210
box -4 -6 36 206
use XNOR2X1  _2558_
timestamp 1597059762
transform -1 0 7464 0 -1 210
box -4 -6 116 206
use NAND2X1  _2716_
timestamp 1597059762
transform 1 0 7256 0 1 210
box -4 -6 52 206
use AOI22X1  _2719_
timestamp 1597059762
transform 1 0 7304 0 1 210
box -4 -6 84 206
use NAND2X1  _2718_
timestamp 1597059762
transform -1 0 7432 0 1 210
box -4 -6 52 206
use AOI22X1  _2826_
timestamp 1597059762
transform -1 0 7544 0 -1 210
box -4 -6 84 206
use NOR2X1  _2829_
timestamp 1597059762
transform 1 0 7432 0 1 210
box -4 -6 52 206
use OR2X2  _2717_
timestamp 1597059762
transform -1 0 7544 0 1 210
box -4 -6 68 206
use FILL  FILL72240x100
timestamp 1597059762
transform -1 0 7560 0 -1 210
box -4 -6 20 206
use FILL  FILL72240x2100
timestamp 1597059762
transform 1 0 7544 0 1 210
box -4 -6 20 206
use DFFPOSX1  _3521_
timestamp 1597059762
transform 1 0 8 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _3505_
timestamp 1597059762
transform 1 0 200 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _3513_
timestamp 1597059762
transform -1 0 584 0 -1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert201
timestamp 1597059762
transform -1 0 632 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert20
timestamp 1597059762
transform -1 0 680 0 -1 610
box -4 -6 52 206
use NAND2X1  _3458_
timestamp 1597059762
transform 1 0 680 0 -1 610
box -4 -6 52 206
use NAND2X1  _3441_
timestamp 1597059762
transform -1 0 840 0 -1 610
box -4 -6 52 206
use FILL  SFILL7280x4100
timestamp 1597059762
transform -1 0 744 0 -1 610
box -4 -6 20 206
use FILL  SFILL7440x4100
timestamp 1597059762
transform -1 0 760 0 -1 610
box -4 -6 20 206
use FILL  SFILL7600x4100
timestamp 1597059762
transform -1 0 776 0 -1 610
box -4 -6 20 206
use FILL  SFILL7760x4100
timestamp 1597059762
transform -1 0 792 0 -1 610
box -4 -6 20 206
use AOI21X1  _3442_
timestamp 1597059762
transform 1 0 840 0 -1 610
box -4 -6 68 206
use AOI21X1  _3486_
timestamp 1597059762
transform 1 0 904 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _3503_
timestamp 1597059762
transform 1 0 968 0 -1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert18
timestamp 1597059762
transform 1 0 1160 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _3501_
timestamp 1597059762
transform 1 0 1208 0 -1 610
box -4 -6 196 206
use AOI21X1  _3481_
timestamp 1597059762
transform -1 0 1464 0 -1 610
box -4 -6 68 206
use NAND2X1  _3480_
timestamp 1597059762
transform -1 0 1512 0 -1 610
box -4 -6 52 206
use NAND2X1  _3479_
timestamp 1597059762
transform 1 0 1512 0 -1 610
box -4 -6 52 206
use NAND2X1  _3444_
timestamp 1597059762
transform 1 0 1560 0 -1 610
box -4 -6 52 206
use NAND2X1  _3497_
timestamp 1597059762
transform 1 0 1608 0 -1 610
box -4 -6 52 206
use AOI21X1  _3499_
timestamp 1597059762
transform -1 0 1720 0 -1 610
box -4 -6 68 206
use NAND2X1  _3498_
timestamp 1597059762
transform -1 0 1768 0 -1 610
box -4 -6 52 206
use AND2X2  _3437_
timestamp 1597059762
transform 1 0 1768 0 -1 610
box -4 -6 68 206
use INVX1  _3428_
timestamp 1597059762
transform 1 0 1832 0 -1 610
box -4 -6 36 206
use AND2X2  _3431_
timestamp 1597059762
transform 1 0 1864 0 -1 610
box -4 -6 68 206
use NAND2X1  _3261_
timestamp 1597059762
transform 1 0 1928 0 -1 610
box -4 -6 52 206
use OAI21X1  _3262_
timestamp 1597059762
transform 1 0 1976 0 -1 610
box -4 -6 68 206
use NOR2X1  _3285_
timestamp 1597059762
transform -1 0 2088 0 -1 610
box -4 -6 52 206
use NOR3X1  _3264_
timestamp 1597059762
transform -1 0 2216 0 -1 610
box -4 -6 132 206
use INVX1  _4498_
timestamp 1597059762
transform 1 0 2216 0 -1 610
box -4 -6 36 206
use OAI21X1  _3267_
timestamp 1597059762
transform -1 0 2376 0 -1 610
box -4 -6 68 206
use NOR3X1  _3286_
timestamp 1597059762
transform -1 0 2504 0 -1 610
box -4 -6 132 206
use FILL  SFILL22480x4100
timestamp 1597059762
transform -1 0 2264 0 -1 610
box -4 -6 20 206
use FILL  SFILL22640x4100
timestamp 1597059762
transform -1 0 2280 0 -1 610
box -4 -6 20 206
use FILL  SFILL22800x4100
timestamp 1597059762
transform -1 0 2296 0 -1 610
box -4 -6 20 206
use FILL  SFILL22960x4100
timestamp 1597059762
transform -1 0 2312 0 -1 610
box -4 -6 20 206
use DFFPOSX1  _3292_
timestamp 1597059762
transform 1 0 2504 0 -1 610
box -4 -6 196 206
use OAI21X1  _4500_
timestamp 1597059762
transform 1 0 2696 0 -1 610
box -4 -6 68 206
use NAND2X1  _4499_
timestamp 1597059762
transform 1 0 2760 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _4451_
timestamp 1597059762
transform 1 0 2808 0 -1 610
box -4 -6 196 206
use INVX1  _4425_
timestamp 1597059762
transform 1 0 3000 0 -1 610
box -4 -6 36 206
use INVX1  _4418_
timestamp 1597059762
transform 1 0 3032 0 -1 610
box -4 -6 36 206
use OAI21X1  _4427_
timestamp 1597059762
transform -1 0 3128 0 -1 610
box -4 -6 68 206
use NOR3X1  _4419_
timestamp 1597059762
transform 1 0 3128 0 -1 610
box -4 -6 132 206
use INVX1  _2089_
timestamp 1597059762
transform 1 0 3256 0 -1 610
box -4 -6 36 206
use INVX1  _4426_
timestamp 1597059762
transform -1 0 3320 0 -1 610
box -4 -6 36 206
use NAND3X1  _4408_
timestamp 1597059762
transform -1 0 3384 0 -1 610
box -4 -6 68 206
use NAND2X1  _4414_
timestamp 1597059762
transform 1 0 3384 0 -1 610
box -4 -6 52 206
use OAI21X1  _4413_
timestamp 1597059762
transform -1 0 3496 0 -1 610
box -4 -6 68 206
use NAND2X1  _4407_
timestamp 1597059762
transform 1 0 3496 0 -1 610
box -4 -6 52 206
use INVX1  _4411_
timestamp 1597059762
transform 1 0 3544 0 -1 610
box -4 -6 36 206
use NOR3X1  _4412_
timestamp 1597059762
transform 1 0 3576 0 -1 610
box -4 -6 132 206
use AOI22X1  _4396_
timestamp 1597059762
transform 1 0 3704 0 -1 610
box -4 -6 84 206
use FILL  SFILL37840x4100
timestamp 1597059762
transform -1 0 3800 0 -1 610
box -4 -6 20 206
use FILL  SFILL38000x4100
timestamp 1597059762
transform -1 0 3816 0 -1 610
box -4 -6 20 206
use FILL  SFILL38160x4100
timestamp 1597059762
transform -1 0 3832 0 -1 610
box -4 -6 20 206
use AOI22X1  _4403_
timestamp 1597059762
transform 1 0 3848 0 -1 610
box -4 -6 84 206
use INVX1  _2080_
timestamp 1597059762
transform 1 0 3928 0 -1 610
box -4 -6 36 206
use OAI21X1  _2082_
timestamp 1597059762
transform 1 0 3960 0 -1 610
box -4 -6 68 206
use FILL  SFILL38320x4100
timestamp 1597059762
transform -1 0 3848 0 -1 610
box -4 -6 20 206
use AOI21X1  _4404_
timestamp 1597059762
transform 1 0 4024 0 -1 610
box -4 -6 68 206
use NAND3X1  _4402_
timestamp 1597059762
transform 1 0 4088 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4447_
timestamp 1597059762
transform 1 0 4152 0 -1 610
box -4 -6 196 206
use AOI22X1  _4384_
timestamp 1597059762
transform 1 0 4344 0 -1 610
box -4 -6 84 206
use AOI21X1  _4385_
timestamp 1597059762
transform 1 0 4424 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4444_
timestamp 1597059762
transform 1 0 4488 0 -1 610
box -4 -6 196 206
use AOI22X1  _4372_
timestamp 1597059762
transform 1 0 4680 0 -1 610
box -4 -6 84 206
use AOI21X1  _4373_
timestamp 1597059762
transform 1 0 4760 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4442_
timestamp 1597059762
transform 1 0 4824 0 -1 610
box -4 -6 196 206
use INVX1  _4348_
timestamp 1597059762
transform 1 0 5016 0 -1 610
box -4 -6 36 206
use OAI21X1  _4355_
timestamp 1597059762
transform 1 0 5048 0 -1 610
box -4 -6 68 206
use INVX1  _4344_
timestamp 1597059762
transform -1 0 5144 0 -1 610
box -4 -6 36 206
use NAND3X1  _4356_
timestamp 1597059762
transform 1 0 5144 0 -1 610
box -4 -6 68 206
use INVX1  _2086_
timestamp 1597059762
transform 1 0 5208 0 -1 610
box -4 -6 36 206
use OAI21X1  _2088_
timestamp 1597059762
transform 1 0 5304 0 -1 610
box -4 -6 68 206
use OAI21X1  _2052_
timestamp 1597059762
transform -1 0 5432 0 -1 610
box -4 -6 68 206
use FILL  SFILL52400x4100
timestamp 1597059762
transform -1 0 5256 0 -1 610
box -4 -6 20 206
use FILL  SFILL52560x4100
timestamp 1597059762
transform -1 0 5272 0 -1 610
box -4 -6 20 206
use FILL  SFILL52720x4100
timestamp 1597059762
transform -1 0 5288 0 -1 610
box -4 -6 20 206
use FILL  SFILL52880x4100
timestamp 1597059762
transform -1 0 5304 0 -1 610
box -4 -6 20 206
use INVX1  _4354_
timestamp 1597059762
transform -1 0 5464 0 -1 610
box -4 -6 36 206
use INVX1  _2059_
timestamp 1597059762
transform 1 0 5464 0 -1 610
box -4 -6 36 206
use OAI21X1  _2061_
timestamp 1597059762
transform -1 0 5560 0 -1 610
box -4 -6 68 206
use INVX1  _2056_
timestamp 1597059762
transform 1 0 5560 0 -1 610
box -4 -6 36 206
use OAI21X1  _2058_
timestamp 1597059762
transform -1 0 5656 0 -1 610
box -4 -6 68 206
use BUFX2  _2018_
timestamp 1597059762
transform 1 0 5656 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert81
timestamp 1597059762
transform 1 0 5704 0 -1 610
box -4 -6 52 206
use XNOR2X1  _2436_
timestamp 1597059762
transform 1 0 5752 0 -1 610
box -4 -6 116 206
use XNOR2X1  _2428_
timestamp 1597059762
transform 1 0 5864 0 -1 610
box -4 -6 116 206
use NOR2X1  _2431_
timestamp 1597059762
transform 1 0 5976 0 -1 610
box -4 -6 52 206
use INVX1  _2430_
timestamp 1597059762
transform -1 0 6056 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert221
timestamp 1597059762
transform 1 0 6056 0 -1 610
box -4 -6 52 206
use NOR2X1  _2443_
timestamp 1597059762
transform -1 0 6152 0 -1 610
box -4 -6 52 206
use INVX1  _2631_
timestamp 1597059762
transform 1 0 6152 0 -1 610
box -4 -6 36 206
use OAI22X1  _2632_
timestamp 1597059762
transform -1 0 6264 0 -1 610
box -4 -6 84 206
use BUFX2  BUFX2_insert253
timestamp 1597059762
transform -1 0 6312 0 -1 610
box -4 -6 52 206
use INVX1  _2628_
timestamp 1597059762
transform 1 0 6312 0 -1 610
box -4 -6 36 206
use OAI22X1  _2629_
timestamp 1597059762
transform -1 0 6424 0 -1 610
box -4 -6 84 206
use NOR2X1  _2633_
timestamp 1597059762
transform -1 0 6472 0 -1 610
box -4 -6 52 206
use AOI22X1  _2664_
timestamp 1597059762
transform -1 0 6552 0 -1 610
box -4 -6 84 206
use NAND2X1  _2662_
timestamp 1597059762
transform 1 0 6552 0 -1 610
box -4 -6 52 206
use INVX1  _2661_
timestamp 1597059762
transform -1 0 6632 0 -1 610
box -4 -6 36 206
use INVX1  _2627_
timestamp 1597059762
transform -1 0 6664 0 -1 610
box -4 -6 36 206
use NAND2X1  _2657_
timestamp 1597059762
transform -1 0 6712 0 -1 610
box -4 -6 52 206
use XNOR2X1  _2211_
timestamp 1597059762
transform -1 0 6888 0 -1 610
box -4 -6 116 206
use FILL  SFILL67120x4100
timestamp 1597059762
transform -1 0 6728 0 -1 610
box -4 -6 20 206
use FILL  SFILL67280x4100
timestamp 1597059762
transform -1 0 6744 0 -1 610
box -4 -6 20 206
use FILL  SFILL67440x4100
timestamp 1597059762
transform -1 0 6760 0 -1 610
box -4 -6 20 206
use FILL  SFILL67600x4100
timestamp 1597059762
transform -1 0 6776 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert79
timestamp 1597059762
transform -1 0 6936 0 -1 610
box -4 -6 52 206
use NAND2X1  _2563_
timestamp 1597059762
transform 1 0 6936 0 -1 610
box -4 -6 52 206
use INVX1  _2562_
timestamp 1597059762
transform 1 0 6984 0 -1 610
box -4 -6 36 206
use NOR2X1  _2580_
timestamp 1597059762
transform -1 0 7064 0 -1 610
box -4 -6 52 206
use AOI21X1  _2212_
timestamp 1597059762
transform -1 0 7128 0 -1 610
box -4 -6 68 206
use OR2X2  _2209_
timestamp 1597059762
transform -1 0 7192 0 -1 610
box -4 -6 68 206
use NAND2X1  _2210_
timestamp 1597059762
transform 1 0 7192 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert251
timestamp 1597059762
transform 1 0 7240 0 -1 610
box -4 -6 52 206
use INVX1  _2208_
timestamp 1597059762
transform 1 0 7288 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert218
timestamp 1597059762
transform 1 0 7320 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert80
timestamp 1597059762
transform 1 0 7368 0 -1 610
box -4 -6 52 206
use NOR2X1  _2586_
timestamp 1597059762
transform 1 0 7416 0 -1 610
box -4 -6 52 206
use INVX1  _2585_
timestamp 1597059762
transform -1 0 7496 0 -1 610
box -4 -6 36 206
use INVX1  _2825_
timestamp 1597059762
transform 1 0 7496 0 -1 610
box -4 -6 36 206
use FILL  FILL72080x4100
timestamp 1597059762
transform -1 0 7544 0 -1 610
box -4 -6 20 206
use FILL  FILL72240x4100
timestamp 1597059762
transform -1 0 7560 0 -1 610
box -4 -6 20 206
use DFFPOSX1  _3514_
timestamp 1597059762
transform -1 0 200 0 1 610
box -4 -6 196 206
use AOI21X1  _3448_
timestamp 1597059762
transform 1 0 200 0 1 610
box -4 -6 68 206
use NAND2X1  _3446_
timestamp 1597059762
transform -1 0 312 0 1 610
box -4 -6 52 206
use AOI21X1  _3490_
timestamp 1597059762
transform -1 0 376 0 1 610
box -4 -6 68 206
use NAND2X1  _3447_
timestamp 1597059762
transform 1 0 376 0 1 610
box -4 -6 52 206
use NAND2X1  _3489_
timestamp 1597059762
transform -1 0 472 0 1 610
box -4 -6 52 206
use INVX8  _3746_
timestamp 1597059762
transform 1 0 472 0 1 610
box -4 -6 84 206
use BUFX2  BUFX2_insert203
timestamp 1597059762
transform -1 0 600 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert21
timestamp 1597059762
transform -1 0 648 0 1 610
box -4 -6 52 206
use NAND2X1  _3459_
timestamp 1597059762
transform 1 0 648 0 1 610
box -4 -6 52 206
use AOI21X1  _3460_
timestamp 1597059762
transform 1 0 696 0 1 610
box -4 -6 68 206
use FILL  SFILL7600x6100
timestamp 1597059762
transform 1 0 760 0 1 610
box -4 -6 20 206
use FILL  SFILL7760x6100
timestamp 1597059762
transform 1 0 776 0 1 610
box -4 -6 20 206
use FILL  SFILL7920x6100
timestamp 1597059762
transform 1 0 792 0 1 610
box -4 -6 20 206
use FILL  SFILL8080x6100
timestamp 1597059762
transform 1 0 808 0 1 610
box -4 -6 20 206
use NAND2X1  _3440_
timestamp 1597059762
transform -1 0 872 0 1 610
box -4 -6 52 206
use DFFPOSX1  _3519_
timestamp 1597059762
transform 1 0 872 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert202
timestamp 1597059762
transform 1 0 1064 0 1 610
box -4 -6 52 206
use NAND2X1  _3485_
timestamp 1597059762
transform -1 0 1160 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert19
timestamp 1597059762
transform 1 0 1160 0 1 610
box -4 -6 52 206
use INVX1  _3396_
timestamp 1597059762
transform 1 0 1208 0 1 610
box -4 -6 36 206
use INVX1  _3368_
timestamp 1597059762
transform 1 0 1240 0 1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert87
timestamp 1597059762
transform 1 0 1272 0 1 610
box -4 -6 52 206
use DFFPOSX1  _3504_
timestamp 1597059762
transform 1 0 1320 0 1 610
box -4 -6 196 206
use AOI21X1  _3488_
timestamp 1597059762
transform -1 0 1576 0 1 610
box -4 -6 68 206
use NAND2X1  _3487_
timestamp 1597059762
transform -1 0 1624 0 1 610
box -4 -6 52 206
use INVX1  _3319_
timestamp 1597059762
transform 1 0 1624 0 1 610
box -4 -6 36 206
use AOI21X1  _3445_
timestamp 1597059762
transform -1 0 1720 0 1 610
box -4 -6 68 206
use INVX8  _3438_
timestamp 1597059762
transform -1 0 1800 0 1 610
box -4 -6 84 206
use DFFPOSX1  _3500_
timestamp 1597059762
transform 1 0 1800 0 1 610
box -4 -6 196 206
use INVX1  _3361_
timestamp 1597059762
transform 1 0 1992 0 1 610
box -4 -6 36 206
use NAND3X1  _3411_
timestamp 1597059762
transform 1 0 2024 0 1 610
box -4 -6 68 206
use NAND3X1  _3355_
timestamp 1597059762
transform 1 0 2088 0 1 610
box -4 -6 68 206
use INVX1  _3326_
timestamp 1597059762
transform 1 0 2152 0 1 610
box -4 -6 36 206
use NAND3X1  _3327_
timestamp 1597059762
transform 1 0 2184 0 1 610
box -4 -6 68 206
use NAND3X1  _3362_
timestamp 1597059762
transform 1 0 2312 0 1 610
box -4 -6 68 206
use AND2X2  _3432_
timestamp 1597059762
transform 1 0 2376 0 1 610
box -4 -6 68 206
use FILL  SFILL22480x6100
timestamp 1597059762
transform 1 0 2248 0 1 610
box -4 -6 20 206
use FILL  SFILL22640x6100
timestamp 1597059762
transform 1 0 2264 0 1 610
box -4 -6 20 206
use FILL  SFILL22800x6100
timestamp 1597059762
transform 1 0 2280 0 1 610
box -4 -6 20 206
use FILL  SFILL22960x6100
timestamp 1597059762
transform 1 0 2296 0 1 610
box -4 -6 20 206
use INVX1  _3418_
timestamp 1597059762
transform 1 0 2440 0 1 610
box -4 -6 36 206
use NAND3X1  _3527_
timestamp 1597059762
transform -1 0 2536 0 1 610
box -4 -6 68 206
use INVX1  _3757_
timestamp 1597059762
transform -1 0 2568 0 1 610
box -4 -6 36 206
use NOR2X1  _3758_
timestamp 1597059762
transform 1 0 2568 0 1 610
box -4 -6 52 206
use INVX1  _4480_
timestamp 1597059762
transform 1 0 2616 0 1 610
box -4 -6 36 206
use INVX1  _3416_
timestamp 1597059762
transform 1 0 2648 0 1 610
box -4 -6 36 206
use DFFPOSX1  _4450_
timestamp 1597059762
transform 1 0 2680 0 1 610
box -4 -6 196 206
use AND2X2  _4423_
timestamp 1597059762
transform -1 0 2936 0 1 610
box -4 -6 68 206
use AOI22X1  _4421_
timestamp 1597059762
transform 1 0 2936 0 1 610
box -4 -6 84 206
use OAI21X1  _4422_
timestamp 1597059762
transform -1 0 3080 0 1 610
box -4 -6 68 206
use AOI21X1  _4430_
timestamp 1597059762
transform -1 0 3144 0 1 610
box -4 -6 68 206
use NAND3X1  _4428_
timestamp 1597059762
transform -1 0 3208 0 1 610
box -4 -6 68 206
use AOI22X1  _4429_
timestamp 1597059762
transform -1 0 3288 0 1 610
box -4 -6 84 206
use OAI21X1  _4420_
timestamp 1597059762
transform -1 0 3352 0 1 610
box -4 -6 68 206
use NAND3X1  _4424_
timestamp 1597059762
transform 1 0 3352 0 1 610
box -4 -6 68 206
use OAI21X1  _4416_
timestamp 1597059762
transform 1 0 3416 0 1 610
box -4 -6 68 206
use AOI22X1  _4415_
timestamp 1597059762
transform 1 0 3480 0 1 610
box -4 -6 84 206
use AND2X2  _4417_
timestamp 1597059762
transform 1 0 3560 0 1 610
box -4 -6 68 206
use NAND2X1  _2084_
timestamp 1597059762
transform -1 0 3672 0 1 610
box -4 -6 52 206
use NAND2X1  _2093_
timestamp 1597059762
transform -1 0 3720 0 1 610
box -4 -6 52 206
use INVX1  _4483_
timestamp 1597059762
transform 1 0 3720 0 1 610
box -4 -6 36 206
use OAI21X1  _4482_
timestamp 1597059762
transform -1 0 3880 0 1 610
box -4 -6 68 206
use FILL  SFILL37520x6100
timestamp 1597059762
transform 1 0 3752 0 1 610
box -4 -6 20 206
use FILL  SFILL37680x6100
timestamp 1597059762
transform 1 0 3768 0 1 610
box -4 -6 20 206
use FILL  SFILL37840x6100
timestamp 1597059762
transform 1 0 3784 0 1 610
box -4 -6 20 206
use FILL  SFILL38000x6100
timestamp 1597059762
transform 1 0 3800 0 1 610
box -4 -6 20 206
use OAI21X1  _4485_
timestamp 1597059762
transform -1 0 3944 0 1 610
box -4 -6 68 206
use NAND2X1  _4484_
timestamp 1597059762
transform 1 0 3944 0 1 610
box -4 -6 52 206
use NAND2X1  _2081_
timestamp 1597059762
transform -1 0 4040 0 1 610
box -4 -6 52 206
use DFFPOSX1  _4449_
timestamp 1597059762
transform 1 0 4040 0 1 610
box -4 -6 196 206
use AOI22X1  _4339_
timestamp 1597059762
transform -1 0 4312 0 1 610
box -4 -6 84 206
use AOI21X1  _4340_
timestamp 1597059762
transform 1 0 4312 0 1 610
box -4 -6 68 206
use NAND2X1  _4335_
timestamp 1597059762
transform -1 0 4424 0 1 610
box -4 -6 52 206
use DFFPOSX1  _4437_
timestamp 1597059762
transform 1 0 4424 0 1 610
box -4 -6 196 206
use INVX1  _4336_
timestamp 1597059762
transform 1 0 4616 0 1 610
box -4 -6 36 206
use NAND3X1  _4345_
timestamp 1597059762
transform 1 0 4648 0 1 610
box -4 -6 68 206
use NAND2X1  _4342_
timestamp 1597059762
transform 1 0 4712 0 1 610
box -4 -6 52 206
use INVX1  _4341_
timestamp 1597059762
transform 1 0 4760 0 1 610
box -4 -6 36 206
use NAND2X1  _2075_
timestamp 1597059762
transform -1 0 4840 0 1 610
box -4 -6 52 206
use OAI21X1  _4349_
timestamp 1597059762
transform 1 0 4840 0 1 610
box -4 -6 68 206
use NAND3X1  _4351_
timestamp 1597059762
transform -1 0 4968 0 1 610
box -4 -6 68 206
use NAND3X1  _4350_
timestamp 1597059762
transform -1 0 5032 0 1 610
box -4 -6 68 206
use NAND3X1  _4357_
timestamp 1597059762
transform 1 0 5032 0 1 610
box -4 -6 68 206
use AND2X2  _4343_
timestamp 1597059762
transform 1 0 5096 0 1 610
box -4 -6 68 206
use INVX1  _2050_
timestamp 1597059762
transform 1 0 5160 0 1 610
box -4 -6 36 206
use NAND2X1  _2087_
timestamp 1597059762
transform -1 0 5240 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert219
timestamp 1597059762
transform -1 0 5352 0 1 610
box -4 -6 52 206
use NAND2X1  _2051_
timestamp 1597059762
transform 1 0 5352 0 1 610
box -4 -6 52 206
use NAND2X1  _2057_
timestamp 1597059762
transform -1 0 5448 0 1 610
box -4 -6 52 206
use FILL  SFILL52400x6100
timestamp 1597059762
transform 1 0 5240 0 1 610
box -4 -6 20 206
use FILL  SFILL52560x6100
timestamp 1597059762
transform 1 0 5256 0 1 610
box -4 -6 20 206
use FILL  SFILL52720x6100
timestamp 1597059762
transform 1 0 5272 0 1 610
box -4 -6 20 206
use FILL  SFILL52880x6100
timestamp 1597059762
transform 1 0 5288 0 1 610
box -4 -6 20 206
use NAND2X1  _2060_
timestamp 1597059762
transform -1 0 5496 0 1 610
box -4 -6 52 206
use NAND2X1  _2054_
timestamp 1597059762
transform -1 0 5544 0 1 610
box -4 -6 52 206
use XNOR2X1  _2429_
timestamp 1597059762
transform 1 0 5544 0 1 610
box -4 -6 116 206
use XOR2X1  _2432_
timestamp 1597059762
transform -1 0 5768 0 1 610
box -4 -6 116 206
use NOR2X1  _2433_
timestamp 1597059762
transform 1 0 5768 0 1 610
box -4 -6 52 206
use NOR2X1  _2434_
timestamp 1597059762
transform -1 0 5864 0 1 610
box -4 -6 52 206
use NAND2X1  _2439_
timestamp 1597059762
transform 1 0 5864 0 1 610
box -4 -6 52 206
use OAI21X1  _2445_
timestamp 1597059762
transform 1 0 5912 0 1 610
box -4 -6 68 206
use AOI21X1  _2444_
timestamp 1597059762
transform 1 0 5976 0 1 610
box -4 -6 68 206
use OAI21X1  _2441_
timestamp 1597059762
transform -1 0 6104 0 1 610
box -4 -6 68 206
use INVX1  _2421_
timestamp 1597059762
transform -1 0 6136 0 1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert171
timestamp 1597059762
transform 1 0 6136 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert51
timestamp 1597059762
transform 1 0 6184 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert263
timestamp 1597059762
transform 1 0 6232 0 1 610
box -4 -6 52 206
use INVX1  _2658_
timestamp 1597059762
transform 1 0 6280 0 1 610
box -4 -6 36 206
use NAND2X1  _2659_
timestamp 1597059762
transform -1 0 6360 0 1 610
box -4 -6 52 206
use NOR2X1  _2660_
timestamp 1597059762
transform -1 0 6408 0 1 610
box -4 -6 52 206
use OAI21X1  _2663_
timestamp 1597059762
transform -1 0 6472 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert265
timestamp 1597059762
transform 1 0 6472 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert145
timestamp 1597059762
transform -1 0 6568 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert52
timestamp 1597059762
transform 1 0 6568 0 1 610
box -4 -6 52 206
use INVX1  _2560_
timestamp 1597059762
transform 1 0 6616 0 1 610
box -4 -6 36 206
use INVX1  _2564_
timestamp 1597059762
transform 1 0 6648 0 1 610
box -4 -6 36 206
use AOI22X1  _2565_
timestamp 1597059762
transform 1 0 6680 0 1 610
box -4 -6 84 206
use OR2X2  _2561_
timestamp 1597059762
transform 1 0 6824 0 1 610
box -4 -6 68 206
use FILL  SFILL67600x6100
timestamp 1597059762
transform 1 0 6760 0 1 610
box -4 -6 20 206
use FILL  SFILL67760x6100
timestamp 1597059762
transform 1 0 6776 0 1 610
box -4 -6 20 206
use FILL  SFILL67920x6100
timestamp 1597059762
transform 1 0 6792 0 1 610
box -4 -6 20 206
use FILL  SFILL68080x6100
timestamp 1597059762
transform 1 0 6808 0 1 610
box -4 -6 20 206
use NAND3X1  _2566_
timestamp 1597059762
transform -1 0 6952 0 1 610
box -4 -6 68 206
use NOR2X1  _2579_
timestamp 1597059762
transform -1 0 7000 0 1 610
box -4 -6 52 206
use AOI21X1  _2581_
timestamp 1597059762
transform 1 0 7000 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert173
timestamp 1597059762
transform -1 0 7112 0 1 610
box -4 -6 52 206
use NOR2X1  _2567_
timestamp 1597059762
transform 1 0 7112 0 1 610
box -4 -6 52 206
use OAI21X1  _2588_
timestamp 1597059762
transform 1 0 7160 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert249
timestamp 1597059762
transform 1 0 7224 0 1 610
box -4 -6 52 206
use NOR2X1  _2584_
timestamp 1597059762
transform 1 0 7272 0 1 610
box -4 -6 52 206
use AOI21X1  _2587_
timestamp 1597059762
transform -1 0 7384 0 1 610
box -4 -6 68 206
use NAND2X1  _2583_
timestamp 1597059762
transform -1 0 7432 0 1 610
box -4 -6 52 206
use XNOR2X1  _2811_
timestamp 1597059762
transform -1 0 7544 0 1 610
box -4 -6 116 206
use FILL  FILL72240x6100
timestamp 1597059762
transform 1 0 7544 0 1 610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert33
timestamp 1597059762
transform 1 0 8 0 -1 1010
box -4 -6 148 206
use NAND2X1  _3462_
timestamp 1597059762
transform 1 0 152 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3463_
timestamp 1597059762
transform 1 0 200 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3461_
timestamp 1597059762
transform -1 0 312 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3465_
timestamp 1597059762
transform 1 0 312 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3466_
timestamp 1597059762
transform 1 0 360 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3464_
timestamp 1597059762
transform 1 0 424 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3492_
timestamp 1597059762
transform -1 0 536 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3491_
timestamp 1597059762
transform -1 0 584 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3449_
timestamp 1597059762
transform -1 0 632 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3451_
timestamp 1597059762
transform 1 0 632 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _3516_
timestamp 1597059762
transform 1 0 760 0 -1 1010
box -4 -6 196 206
use FILL  SFILL6960x8100
timestamp 1597059762
transform -1 0 712 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7120x8100
timestamp 1597059762
transform -1 0 728 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7280x8100
timestamp 1597059762
transform -1 0 744 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7440x8100
timestamp 1597059762
transform -1 0 760 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  _3517_
timestamp 1597059762
transform -1 0 1144 0 -1 1010
box -4 -6 196 206
use NAND2X1  _3453_
timestamp 1597059762
transform 1 0 1144 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3454_
timestamp 1597059762
transform -1 0 1256 0 -1 1010
box -4 -6 68 206
use AOI21X1  _3494_
timestamp 1597059762
transform -1 0 1320 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3452_
timestamp 1597059762
transform -1 0 1368 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3493_
timestamp 1597059762
transform -1 0 1416 0 -1 1010
box -4 -6 52 206
use OAI21X1  _3623_
timestamp 1597059762
transform 1 0 1416 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3622_
timestamp 1597059762
transform -1 0 1528 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _4239_
timestamp 1597059762
transform 1 0 1528 0 -1 1010
box -4 -6 196 206
use NAND2X1  _3443_
timestamp 1597059762
transform -1 0 1768 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _3520_
timestamp 1597059762
transform 1 0 1768 0 -1 1010
box -4 -6 196 206
use BUFX2  BUFX2_insert166
timestamp 1597059762
transform -1 0 2008 0 -1 1010
box -4 -6 52 206
use NAND3X1  _3397_
timestamp 1597059762
transform 1 0 2008 0 -1 1010
box -4 -6 68 206
use NOR2X1  _3303_
timestamp 1597059762
transform 1 0 2072 0 -1 1010
box -4 -6 52 206
use INVX4  _3542_
timestamp 1597059762
transform -1 0 2168 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3407_
timestamp 1597059762
transform -1 0 2216 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3365_
timestamp 1597059762
transform -1 0 2264 0 -1 1010
box -4 -6 52 206
use NOR2X1  _3429_
timestamp 1597059762
transform -1 0 2376 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3351_
timestamp 1597059762
transform 1 0 2376 0 -1 1010
box -4 -6 52 206
use FILL  SFILL22640x8100
timestamp 1597059762
transform -1 0 2280 0 -1 1010
box -4 -6 20 206
use FILL  SFILL22800x8100
timestamp 1597059762
transform -1 0 2296 0 -1 1010
box -4 -6 20 206
use FILL  SFILL22960x8100
timestamp 1597059762
transform -1 0 2312 0 -1 1010
box -4 -6 20 206
use FILL  SFILL23120x8100
timestamp 1597059762
transform -1 0 2328 0 -1 1010
box -4 -6 20 206
use NAND2X1  _3372_
timestamp 1597059762
transform -1 0 2472 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert129
timestamp 1597059762
transform -1 0 2520 0 -1 1010
box -4 -6 52 206
use NOR2X1  _3419_
timestamp 1597059762
transform -1 0 2568 0 -1 1010
box -4 -6 52 206
use AND2X2  _3434_
timestamp 1597059762
transform 1 0 2568 0 -1 1010
box -4 -6 68 206
use INVX1  _3422_
timestamp 1597059762
transform 1 0 2632 0 -1 1010
box -4 -6 36 206
use NOR2X1  _3423_
timestamp 1597059762
transform -1 0 2712 0 -1 1010
box -4 -6 52 206
use NOR2X1  _3417_
timestamp 1597059762
transform -1 0 2760 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert164
timestamp 1597059762
transform 1 0 2760 0 -1 1010
box -4 -6 52 206
use INVX1  _4459_
timestamp 1597059762
transform 1 0 2808 0 -1 1010
box -4 -6 36 206
use AND2X2  _3433_
timestamp 1597059762
transform 1 0 2840 0 -1 1010
box -4 -6 68 206
use INVX1  _3420_
timestamp 1597059762
transform 1 0 2904 0 -1 1010
box -4 -6 36 206
use INVX1  _4492_
timestamp 1597059762
transform 1 0 2936 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4494_
timestamp 1597059762
transform 1 0 2968 0 -1 1010
box -4 -6 68 206
use NOR2X1  _3421_
timestamp 1597059762
transform -1 0 3080 0 -1 1010
box -4 -6 52 206
use INVX1  _4474_
timestamp 1597059762
transform 1 0 3080 0 -1 1010
box -4 -6 36 206
use INVX1  _4495_
timestamp 1597059762
transform 1 0 3112 0 -1 1010
box -4 -6 36 206
use NAND2X1  _4493_
timestamp 1597059762
transform 1 0 3144 0 -1 1010
box -4 -6 52 206
use INVX1  _4477_
timestamp 1597059762
transform 1 0 3192 0 -1 1010
box -4 -6 36 206
use INVX1  _4462_
timestamp 1597059762
transform 1 0 3224 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4497_
timestamp 1597059762
transform 1 0 3256 0 -1 1010
box -4 -6 68 206
use INVX1  _4453_
timestamp 1597059762
transform 1 0 3320 0 -1 1010
box -4 -6 36 206
use INVX1  _4465_
timestamp 1597059762
transform 1 0 3352 0 -1 1010
box -4 -6 36 206
use INVX1  _4489_
timestamp 1597059762
transform 1 0 3384 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4491_
timestamp 1597059762
transform 1 0 3416 0 -1 1010
box -4 -6 68 206
use NAND2X1  _4490_
timestamp 1597059762
transform 1 0 3480 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4455_
timestamp 1597059762
transform -1 0 3592 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert167
timestamp 1597059762
transform -1 0 3640 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4461_
timestamp 1597059762
transform 1 0 3640 0 -1 1010
box -4 -6 68 206
use NAND2X1  _4481_
timestamp 1597059762
transform 1 0 3704 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4464_
timestamp 1597059762
transform 1 0 3816 0 -1 1010
box -4 -6 68 206
use FILL  SFILL37520x8100
timestamp 1597059762
transform -1 0 3768 0 -1 1010
box -4 -6 20 206
use FILL  SFILL37680x8100
timestamp 1597059762
transform -1 0 3784 0 -1 1010
box -4 -6 20 206
use FILL  SFILL37840x8100
timestamp 1597059762
transform -1 0 3800 0 -1 1010
box -4 -6 20 206
use FILL  SFILL38000x8100
timestamp 1597059762
transform -1 0 3816 0 -1 1010
box -4 -6 20 206
use NAND2X1  _4463_
timestamp 1597059762
transform -1 0 3928 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4476_
timestamp 1597059762
transform 1 0 3928 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert162
timestamp 1597059762
transform 1 0 3992 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4479_
timestamp 1597059762
transform 1 0 4040 0 -1 1010
box -4 -6 68 206
use NAND2X1  _4478_
timestamp 1597059762
transform 1 0 4104 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4467_
timestamp 1597059762
transform 1 0 4152 0 -1 1010
box -4 -6 68 206
use INVX1  _4471_
timestamp 1597059762
transform 1 0 4216 0 -1 1010
box -4 -6 36 206
use OAI21X1  _4473_
timestamp 1597059762
transform 1 0 4248 0 -1 1010
box -4 -6 68 206
use AOI22X1  _4346_
timestamp 1597059762
transform 1 0 4312 0 -1 1010
box -4 -6 84 206
use AOI21X1  _4347_
timestamp 1597059762
transform -1 0 4456 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _4438_
timestamp 1597059762
transform 1 0 4456 0 -1 1010
box -4 -6 196 206
use AOI22X1  _4352_
timestamp 1597059762
transform 1 0 4648 0 -1 1010
box -4 -6 84 206
use AOI22X1  _4358_
timestamp 1597059762
transform 1 0 4728 0 -1 1010
box -4 -6 84 206
use AOI21X1  _4353_
timestamp 1597059762
transform 1 0 4808 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _4439_
timestamp 1597059762
transform 1 0 4872 0 -1 1010
box -4 -6 196 206
use AOI21X1  _4359_
timestamp 1597059762
transform 1 0 5064 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _4440_
timestamp 1597059762
transform 1 0 5128 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  _4303_
timestamp 1597059762
transform 1 0 5384 0 -1 1010
box -4 -6 196 206
use FILL  SFILL53200x8100
timestamp 1597059762
transform -1 0 5336 0 -1 1010
box -4 -6 20 206
use FILL  SFILL53360x8100
timestamp 1597059762
transform -1 0 5352 0 -1 1010
box -4 -6 20 206
use FILL  SFILL53520x8100
timestamp 1597059762
transform -1 0 5368 0 -1 1010
box -4 -6 20 206
use FILL  SFILL53680x8100
timestamp 1597059762
transform -1 0 5384 0 -1 1010
box -4 -6 20 206
use NAND2X1  _3043_
timestamp 1597059762
transform 1 0 5576 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2491_
timestamp 1597059762
transform -1 0 5672 0 -1 1010
box -4 -6 52 206
use NOR2X1  _2490_
timestamp 1597059762
transform 1 0 5672 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3065_
timestamp 1597059762
transform -1 0 5768 0 -1 1010
box -4 -6 52 206
use AOI22X1  _2427_
timestamp 1597059762
transform -1 0 5848 0 -1 1010
box -4 -6 84 206
use NOR2X1  _2440_
timestamp 1597059762
transform 1 0 5848 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2423_
timestamp 1597059762
transform 1 0 5896 0 -1 1010
box -4 -6 52 206
use OAI21X1  _2418_
timestamp 1597059762
transform -1 0 6008 0 -1 1010
box -4 -6 68 206
use OAI21X1  _2425_
timestamp 1597059762
transform 1 0 6008 0 -1 1010
box -4 -6 68 206
use NAND2X1  _2422_
timestamp 1597059762
transform -1 0 6120 0 -1 1010
box -4 -6 52 206
use INVX1  _2415_
timestamp 1597059762
transform -1 0 6152 0 -1 1010
box -4 -6 36 206
use XNOR2X1  _2416_
timestamp 1597059762
transform -1 0 6264 0 -1 1010
box -4 -6 116 206
use AND2X2  _2307_
timestamp 1597059762
transform -1 0 6328 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert148
timestamp 1597059762
transform 1 0 6328 0 -1 1010
box -4 -6 52 206
use AND2X2  _2130_
timestamp 1597059762
transform 1 0 6376 0 -1 1010
box -4 -6 68 206
use XNOR2X1  _2817_
timestamp 1597059762
transform -1 0 6552 0 -1 1010
box -4 -6 116 206
use NOR2X1  _2124_
timestamp 1597059762
transform 1 0 6552 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert49
timestamp 1597059762
transform 1 0 6600 0 -1 1010
box -4 -6 52 206
use OR2X2  _2126_
timestamp 1597059762
transform 1 0 6648 0 -1 1010
box -4 -6 68 206
use NAND2X1  _2128_
timestamp 1597059762
transform -1 0 6760 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2127_
timestamp 1597059762
transform 1 0 6824 0 -1 1010
box -4 -6 52 206
use FILL  SFILL67600x8100
timestamp 1597059762
transform -1 0 6776 0 -1 1010
box -4 -6 20 206
use FILL  SFILL67760x8100
timestamp 1597059762
transform -1 0 6792 0 -1 1010
box -4 -6 20 206
use FILL  SFILL67920x8100
timestamp 1597059762
transform -1 0 6808 0 -1 1010
box -4 -6 20 206
use FILL  SFILL68080x8100
timestamp 1597059762
transform -1 0 6824 0 -1 1010
box -4 -6 20 206
use AND2X2  _2131_
timestamp 1597059762
transform -1 0 6936 0 -1 1010
box -4 -6 68 206
use INVX1  _2814_
timestamp 1597059762
transform 1 0 6936 0 -1 1010
box -4 -6 36 206
use INVX1  _2836_
timestamp 1597059762
transform 1 0 6968 0 -1 1010
box -4 -6 36 206
use NOR2X1  _2837_
timestamp 1597059762
transform 1 0 7000 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2816_
timestamp 1597059762
transform -1 0 7096 0 -1 1010
box -4 -6 52 206
use NOR2X1  _2835_
timestamp 1597059762
transform 1 0 7096 0 -1 1010
box -4 -6 52 206
use AOI21X1  _2838_
timestamp 1597059762
transform -1 0 7208 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert139
timestamp 1597059762
transform 1 0 7208 0 -1 1010
box -4 -6 52 206
use NOR2X1  _2143_
timestamp 1597059762
transform -1 0 7304 0 -1 1010
box -4 -6 52 206
use AND2X2  _2144_
timestamp 1597059762
transform -1 0 7368 0 -1 1010
box -4 -6 68 206
use NAND2X1  _2813_
timestamp 1597059762
transform -1 0 7416 0 -1 1010
box -4 -6 52 206
use INVX1  _2839_
timestamp 1597059762
transform 1 0 7416 0 -1 1010
box -4 -6 36 206
use NOR2X1  _2840_
timestamp 1597059762
transform -1 0 7496 0 -1 1010
box -4 -6 52 206
use AOI21X1  _2843_
timestamp 1597059762
transform -1 0 7560 0 -1 1010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert29
timestamp 1597059762
transform 1 0 8 0 1 1010
box -4 -6 148 206
use DFFPOSX1  _3515_
timestamp 1597059762
transform -1 0 344 0 1 1010
box -4 -6 196 206
use INVX1  _3375_
timestamp 1597059762
transform 1 0 344 0 1 1010
box -4 -6 36 206
use INVX1  _3333_
timestamp 1597059762
transform -1 0 408 0 1 1010
box -4 -6 36 206
use DFFPOSX1  _3506_
timestamp 1597059762
transform 1 0 408 0 1 1010
box -4 -6 196 206
use NAND2X1  _3450_
timestamp 1597059762
transform 1 0 600 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert193
timestamp 1597059762
transform -1 0 696 0 1 1010
box -4 -6 52 206
use INVX1  _3340_
timestamp 1597059762
transform 1 0 696 0 1 1010
box -4 -6 36 206
use DFFPOSX1  _4223_
timestamp 1597059762
transform 1 0 792 0 1 1010
box -4 -6 196 206
use FILL  SFILL7280x10100
timestamp 1597059762
transform 1 0 728 0 1 1010
box -4 -6 20 206
use FILL  SFILL7440x10100
timestamp 1597059762
transform 1 0 744 0 1 1010
box -4 -6 20 206
use FILL  SFILL7600x10100
timestamp 1597059762
transform 1 0 760 0 1 1010
box -4 -6 20 206
use FILL  SFILL7760x10100
timestamp 1597059762
transform 1 0 776 0 1 1010
box -4 -6 20 206
use AOI21X1  _3723_
timestamp 1597059762
transform 1 0 984 0 1 1010
box -4 -6 68 206
use NOR2X1  _3722_
timestamp 1597059762
transform -1 0 1096 0 1 1010
box -4 -6 52 206
use OAI21X1  _4012_
timestamp 1597059762
transform 1 0 1096 0 1 1010
box -4 -6 68 206
use OAI21X1  _3800_
timestamp 1597059762
transform 1 0 1160 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _3507_
timestamp 1597059762
transform 1 0 1224 0 1 1010
box -4 -6 196 206
use MUX2X1  _4006_
timestamp 1597059762
transform 1 0 1416 0 1 1010
box -4 -6 100 206
use NOR2X1  _3655_
timestamp 1597059762
transform 1 0 1512 0 1 1010
box -4 -6 52 206
use AOI21X1  _3656_
timestamp 1597059762
transform -1 0 1624 0 1 1010
box -4 -6 68 206
use MUX2X1  _3794_
timestamp 1597059762
transform 1 0 1624 0 1 1010
box -4 -6 100 206
use DFFPOSX1  _4255_
timestamp 1597059762
transform -1 0 1912 0 1 1010
box -4 -6 196 206
use INVX1  _3302_
timestamp 1597059762
transform -1 0 1944 0 1 1010
box -4 -6 36 206
use INVX1  _3347_
timestamp 1597059762
transform -1 0 1976 0 1 1010
box -4 -6 36 206
use NAND3X1  _3320_
timestamp 1597059762
transform 1 0 1976 0 1 1010
box -4 -6 68 206
use NAND3X1  _3369_
timestamp 1597059762
transform 1 0 2040 0 1 1010
box -4 -6 68 206
use NAND3X1  _3334_
timestamp 1597059762
transform 1 0 2104 0 1 1010
box -4 -6 68 206
use NAND3X1  _3348_
timestamp 1597059762
transform 1 0 2168 0 1 1010
box -4 -6 68 206
use NAND2X1  _3336_
timestamp 1597059762
transform 1 0 2296 0 1 1010
box -4 -6 52 206
use NAND3X1  _3390_
timestamp 1597059762
transform 1 0 2344 0 1 1010
box -4 -6 68 206
use NAND3X1  _3404_
timestamp 1597059762
transform 1 0 2408 0 1 1010
box -4 -6 68 206
use FILL  SFILL22320x10100
timestamp 1597059762
transform 1 0 2232 0 1 1010
box -4 -6 20 206
use FILL  SFILL22480x10100
timestamp 1597059762
transform 1 0 2248 0 1 1010
box -4 -6 20 206
use FILL  SFILL22640x10100
timestamp 1597059762
transform 1 0 2264 0 1 1010
box -4 -6 20 206
use FILL  SFILL22800x10100
timestamp 1597059762
transform 1 0 2280 0 1 1010
box -4 -6 20 206
use NAND3X1  _3341_
timestamp 1597059762
transform 1 0 2472 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert130
timestamp 1597059762
transform 1 0 2536 0 1 1010
box -4 -6 52 206
use NAND2X1  _3330_
timestamp 1597059762
transform 1 0 2584 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert127
timestamp 1597059762
transform 1 0 2632 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert128
timestamp 1597059762
transform 1 0 2680 0 1 1010
box -4 -6 52 206
use AND2X2  _3435_
timestamp 1597059762
transform -1 0 2792 0 1 1010
box -4 -6 68 206
use INVX1  _3424_
timestamp 1597059762
transform 1 0 2792 0 1 1010
box -4 -6 36 206
use AND2X2  _3436_
timestamp 1597059762
transform 1 0 2824 0 1 1010
box -4 -6 68 206
use INVX1  _3426_
timestamp 1597059762
transform 1 0 2888 0 1 1010
box -4 -6 36 206
use NOR2X1  _3427_
timestamp 1597059762
transform -1 0 2968 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert168
timestamp 1597059762
transform -1 0 3016 0 1 1010
box -4 -6 52 206
use NOR2X1  _3425_
timestamp 1597059762
transform -1 0 3064 0 1 1010
box -4 -6 52 206
use AND2X2  _3430_
timestamp 1597059762
transform 1 0 3064 0 1 1010
box -4 -6 68 206
use INVX1  _3414_
timestamp 1597059762
transform 1 0 3128 0 1 1010
box -4 -6 36 206
use NOR2X1  _3415_
timestamp 1597059762
transform 1 0 3160 0 1 1010
box -4 -6 52 206
use INVX1  _4468_
timestamp 1597059762
transform 1 0 3208 0 1 1010
box -4 -6 36 206
use INVX1  _4486_
timestamp 1597059762
transform 1 0 3240 0 1 1010
box -4 -6 36 206
use NAND2X1  _4496_
timestamp 1597059762
transform 1 0 3272 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert165
timestamp 1597059762
transform -1 0 3368 0 1 1010
box -4 -6 52 206
use INVX1  _4456_
timestamp 1597059762
transform 1 0 3368 0 1 1010
box -4 -6 36 206
use OAI21X1  _4488_
timestamp 1597059762
transform 1 0 3400 0 1 1010
box -4 -6 68 206
use NAND2X1  _4487_
timestamp 1597059762
transform 1 0 3464 0 1 1010
box -4 -6 52 206
use NAND2X1  _4454_
timestamp 1597059762
transform -1 0 3560 0 1 1010
box -4 -6 52 206
use INVX4  _4331_
timestamp 1597059762
transform -1 0 3608 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert163
timestamp 1597059762
transform 1 0 3608 0 1 1010
box -4 -6 52 206
use NAND2X1  _4460_
timestamp 1597059762
transform 1 0 3656 0 1 1010
box -4 -6 52 206
use OAI21X1  _4458_
timestamp 1597059762
transform 1 0 3704 0 1 1010
box -4 -6 68 206
use FILL  SFILL37680x10100
timestamp 1597059762
transform 1 0 3768 0 1 1010
box -4 -6 20 206
use FILL  SFILL37840x10100
timestamp 1597059762
transform 1 0 3784 0 1 1010
box -4 -6 20 206
use FILL  SFILL38000x10100
timestamp 1597059762
transform 1 0 3800 0 1 1010
box -4 -6 20 206
use FILL  SFILL38160x10100
timestamp 1597059762
transform 1 0 3816 0 1 1010
box -4 -6 20 206
use NAND2X1  _4457_
timestamp 1597059762
transform 1 0 3832 0 1 1010
box -4 -6 52 206
use OAI21X1  _4470_
timestamp 1597059762
transform 1 0 3880 0 1 1010
box -4 -6 68 206
use NAND2X1  _4475_
timestamp 1597059762
transform 1 0 3944 0 1 1010
box -4 -6 52 206
use NAND2X1  _4469_
timestamp 1597059762
transform -1 0 4040 0 1 1010
box -4 -6 52 206
use AOI21X1  _4016_
timestamp 1597059762
transform 1 0 4040 0 1 1010
box -4 -6 68 206
use OAI21X1  _4015_
timestamp 1597059762
transform -1 0 4168 0 1 1010
box -4 -6 68 206
use NAND2X1  _4466_
timestamp 1597059762
transform 1 0 4168 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert169
timestamp 1597059762
transform 1 0 4216 0 1 1010
box -4 -6 52 206
use NAND2X1  _4472_
timestamp 1597059762
transform 1 0 4264 0 1 1010
box -4 -6 52 206
use AOI21X1  _3804_
timestamp 1597059762
transform 1 0 4312 0 1 1010
box -4 -6 68 206
use OAI21X1  _3803_
timestamp 1597059762
transform -1 0 4440 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _4305_
timestamp 1597059762
transform 1 0 4440 0 1 1010
box -4 -6 196 206
use DFFPOSX1  _4319_
timestamp 1597059762
transform 1 0 4632 0 1 1010
box -4 -6 196 206
use BUFX2  BUFX2_insert77
timestamp 1597059762
transform -1 0 4872 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert144
timestamp 1597059762
transform 1 0 4872 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2360_
timestamp 1597059762
transform 1 0 4920 0 1 1010
box -4 -6 116 206
use NAND2X1  _2999_
timestamp 1597059762
transform -1 0 5080 0 1 1010
box -4 -6 52 206
use XOR2X1  _2413_
timestamp 1597059762
transform -1 0 5192 0 1 1010
box -4 -6 116 206
use BUFX2  BUFX2_insert262
timestamp 1597059762
transform -1 0 5240 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2414_
timestamp 1597059762
transform -1 0 5416 0 1 1010
box -4 -6 116 206
use NOR2X1  _2426_
timestamp 1597059762
transform 1 0 5416 0 1 1010
box -4 -6 52 206
use FILL  SFILL52400x10100
timestamp 1597059762
transform 1 0 5240 0 1 1010
box -4 -6 20 206
use FILL  SFILL52560x10100
timestamp 1597059762
transform 1 0 5256 0 1 1010
box -4 -6 20 206
use FILL  SFILL52720x10100
timestamp 1597059762
transform 1 0 5272 0 1 1010
box -4 -6 20 206
use FILL  SFILL52880x10100
timestamp 1597059762
transform 1 0 5288 0 1 1010
box -4 -6 20 206
use NAND2X1  _3021_
timestamp 1597059762
transform -1 0 5512 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2424_
timestamp 1597059762
transform -1 0 5624 0 1 1010
box -4 -6 116 206
use BUFX2  BUFX2_insert138
timestamp 1597059762
transform 1 0 5624 0 1 1010
box -4 -6 52 206
use XOR2X1  _2489_
timestamp 1597059762
transform -1 0 5784 0 1 1010
box -4 -6 116 206
use NAND2X1  _2417_
timestamp 1597059762
transform -1 0 5832 0 1 1010
box -4 -6 52 206
use NAND2X1  _2438_
timestamp 1597059762
transform 1 0 5832 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert170
timestamp 1597059762
transform 1 0 5880 0 1 1010
box -4 -6 52 206
use INVX1  _2419_
timestamp 1597059762
transform 1 0 5928 0 1 1010
box -4 -6 36 206
use NAND2X1  _2420_
timestamp 1597059762
transform -1 0 6008 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2437_
timestamp 1597059762
transform -1 0 6120 0 1 1010
box -4 -6 116 206
use BUFX2  BUFX2_insert53
timestamp 1597059762
transform -1 0 6168 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert264
timestamp 1597059762
transform -1 0 6216 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert146
timestamp 1597059762
transform 1 0 6216 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert266
timestamp 1597059762
transform 1 0 6264 0 1 1010
box -4 -6 52 206
use NAND2X1  _2120_
timestamp 1597059762
transform 1 0 6312 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2129_
timestamp 1597059762
transform 1 0 6360 0 1 1010
box -4 -6 116 206
use OAI21X1  _2125_
timestamp 1597059762
transform -1 0 6536 0 1 1010
box -4 -6 68 206
use NOR2X1  _2133_
timestamp 1597059762
transform 1 0 6536 0 1 1010
box -4 -6 52 206
use NAND2X1  _2136_
timestamp 1597059762
transform 1 0 6584 0 1 1010
box -4 -6 52 206
use NOR2X1  _2135_
timestamp 1597059762
transform -1 0 6680 0 1 1010
box -4 -6 52 206
use AOI21X1  _2132_
timestamp 1597059762
transform 1 0 6680 0 1 1010
box -4 -6 68 206
use NOR2X1  _2134_
timestamp 1597059762
transform 1 0 6808 0 1 1010
box -4 -6 52 206
use FILL  SFILL67440x10100
timestamp 1597059762
transform 1 0 6744 0 1 1010
box -4 -6 20 206
use FILL  SFILL67600x10100
timestamp 1597059762
transform 1 0 6760 0 1 1010
box -4 -6 20 206
use FILL  SFILL67760x10100
timestamp 1597059762
transform 1 0 6776 0 1 1010
box -4 -6 20 206
use FILL  SFILL67920x10100
timestamp 1597059762
transform 1 0 6792 0 1 1010
box -4 -6 20 206
use BUFX2  BUFX2_insert172
timestamp 1597059762
transform -1 0 6904 0 1 1010
box -4 -6 52 206
use OR2X2  _2815_
timestamp 1597059762
transform -1 0 6968 0 1 1010
box -4 -6 68 206
use NAND3X1  _2818_
timestamp 1597059762
transform 1 0 6968 0 1 1010
box -4 -6 68 206
use NOR2X1  _2819_
timestamp 1597059762
transform -1 0 7080 0 1 1010
box -4 -6 52 206
use OAI21X1  _2844_
timestamp 1597059762
transform -1 0 7144 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert78
timestamp 1597059762
transform 1 0 7144 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert220
timestamp 1597059762
transform 1 0 7192 0 1 1010
box -4 -6 52 206
use NOR2X1  _2145_
timestamp 1597059762
transform -1 0 7288 0 1 1010
box -4 -6 52 206
use INVX1  _2841_
timestamp 1597059762
transform 1 0 7288 0 1 1010
box -4 -6 36 206
use NOR2X1  _2842_
timestamp 1597059762
transform -1 0 7368 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2812_
timestamp 1597059762
transform -1 0 7480 0 1 1010
box -4 -6 116 206
use NOR2X1  _2576_
timestamp 1597059762
transform -1 0 7528 0 1 1010
box -4 -6 52 206
use FILL  FILL72080x10100
timestamp 1597059762
transform 1 0 7528 0 1 1010
box -4 -6 20 206
use FILL  FILL72240x10100
timestamp 1597059762
transform 1 0 7544 0 1 1010
box -4 -6 20 206
use DFFPOSX1  _4271_
timestamp 1597059762
transform -1 0 200 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _4191_
timestamp 1597059762
transform 1 0 200 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _4287_
timestamp 1597059762
transform 1 0 392 0 -1 1410
box -4 -6 196 206
use MUX2X1  _4010_
timestamp 1597059762
transform -1 0 680 0 -1 1410
box -4 -6 100 206
use MUX2X1  _3798_
timestamp 1597059762
transform -1 0 776 0 -1 1410
box -4 -6 100 206
use FILL  SFILL7760x12100
timestamp 1597059762
transform -1 0 792 0 -1 1410
box -4 -6 20 206
use FILL  SFILL7920x12100
timestamp 1597059762
transform -1 0 808 0 -1 1410
box -4 -6 20 206
use FILL  SFILL8080x12100
timestamp 1597059762
transform -1 0 824 0 -1 1410
box -4 -6 20 206
use DFFPOSX1  _4273_
timestamp 1597059762
transform 1 0 840 0 -1 1410
box -4 -6 196 206
use FILL  SFILL8240x12100
timestamp 1597059762
transform -1 0 840 0 -1 1410
box -4 -6 20 206
use AOI21X1  _3652_
timestamp 1597059762
transform 1 0 1032 0 -1 1410
box -4 -6 68 206
use NOR2X1  _3651_
timestamp 1597059762
transform -1 0 1144 0 -1 1410
box -4 -6 52 206
use OAI22X1  _4013_
timestamp 1597059762
transform -1 0 1224 0 -1 1410
box -4 -6 84 206
use NOR2X1  _4011_
timestamp 1597059762
transform 1 0 1224 0 -1 1410
box -4 -6 52 206
use OAI22X1  _3801_
timestamp 1597059762
transform 1 0 1272 0 -1 1410
box -4 -6 84 206
use BUFX2  BUFX2_insert121
timestamp 1597059762
transform -1 0 1400 0 -1 1410
box -4 -6 52 206
use OAI21X1  _4008_
timestamp 1597059762
transform 1 0 1400 0 -1 1410
box -4 -6 68 206
use OAI22X1  _4009_
timestamp 1597059762
transform -1 0 1544 0 -1 1410
box -4 -6 84 206
use MUX2X1  _4014_
timestamp 1597059762
transform 1 0 1544 0 -1 1410
box -4 -6 100 206
use OAI21X1  _3796_
timestamp 1597059762
transform 1 0 1640 0 -1 1410
box -4 -6 68 206
use NOR2X1  _4007_
timestamp 1597059762
transform -1 0 1752 0 -1 1410
box -4 -6 52 206
use OAI22X1  _3797_
timestamp 1597059762
transform 1 0 1752 0 -1 1410
box -4 -6 84 206
use MUX2X1  _3802_
timestamp 1597059762
transform 1 0 1832 0 -1 1410
box -4 -6 100 206
use INVX4  _3536_
timestamp 1597059762
transform -1 0 1976 0 -1 1410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert28
timestamp 1597059762
transform 1 0 1976 0 -1 1410
box -4 -6 148 206
use NAND3X1  _3370_
timestamp 1597059762
transform -1 0 2184 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3371_
timestamp 1597059762
transform -1 0 2232 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3335_
timestamp 1597059762
transform -1 0 2360 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3357_
timestamp 1597059762
transform 1 0 2360 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3356_
timestamp 1597059762
transform -1 0 2472 0 -1 1410
box -4 -6 68 206
use FILL  SFILL22320x12100
timestamp 1597059762
transform -1 0 2248 0 -1 1410
box -4 -6 20 206
use FILL  SFILL22480x12100
timestamp 1597059762
transform -1 0 2264 0 -1 1410
box -4 -6 20 206
use FILL  SFILL22640x12100
timestamp 1597059762
transform -1 0 2280 0 -1 1410
box -4 -6 20 206
use FILL  SFILL22800x12100
timestamp 1597059762
transform -1 0 2296 0 -1 1410
box -4 -6 20 206
use NAND3X1  _3321_
timestamp 1597059762
transform -1 0 2536 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3322_
timestamp 1597059762
transform -1 0 2584 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3316_
timestamp 1597059762
transform -1 0 2632 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3386_
timestamp 1597059762
transform 1 0 2632 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3393_
timestamp 1597059762
transform 1 0 2680 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3309_
timestamp 1597059762
transform 1 0 2728 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3349_
timestamp 1597059762
transform -1 0 2840 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3350_
timestamp 1597059762
transform -1 0 2888 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3400_
timestamp 1597059762
transform -1 0 2936 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3344_
timestamp 1597059762
transform 1 0 2936 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3328_
timestamp 1597059762
transform -1 0 3048 0 -1 1410
box -4 -6 68 206
use NAND2X1  _3329_
timestamp 1597059762
transform -1 0 3096 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3323_
timestamp 1597059762
transform -1 0 3144 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3337_
timestamp 1597059762
transform 1 0 3144 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3358_
timestamp 1597059762
transform -1 0 3240 0 -1 1410
box -4 -6 52 206
use NAND2X1  _3295_
timestamp 1597059762
transform -1 0 3288 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3353_
timestamp 1597059762
transform 1 0 3288 0 -1 1410
box -4 -6 68 206
use OAI21X1  _3346_
timestamp 1597059762
transform 1 0 3352 0 -1 1410
box -4 -6 68 206
use OAI21X1  _3332_
timestamp 1597059762
transform 1 0 3416 0 -1 1410
box -4 -6 68 206
use OAI21X1  _3325_
timestamp 1597059762
transform 1 0 3480 0 -1 1410
box -4 -6 68 206
use INVX1  _3331_
timestamp 1597059762
transform -1 0 3576 0 -1 1410
box -4 -6 36 206
use INVX1  _3352_
timestamp 1597059762
transform -1 0 3608 0 -1 1410
box -4 -6 36 206
use INVX1  _3324_
timestamp 1597059762
transform -1 0 3640 0 -1 1410
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert23
timestamp 1597059762
transform 1 0 3640 0 -1 1410
box -4 -6 148 206
use FILL  SFILL37840x12100
timestamp 1597059762
transform -1 0 3800 0 -1 1410
box -4 -6 20 206
use FILL  SFILL38000x12100
timestamp 1597059762
transform -1 0 3816 0 -1 1410
box -4 -6 20 206
use FILL  SFILL38160x12100
timestamp 1597059762
transform -1 0 3832 0 -1 1410
box -4 -6 20 206
use BUFX2  BUFX2_insert102
timestamp 1597059762
transform 1 0 3848 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _4320_
timestamp 1597059762
transform 1 0 3896 0 -1 1410
box -4 -6 196 206
use FILL  SFILL38320x12100
timestamp 1597059762
transform -1 0 3848 0 -1 1410
box -4 -6 20 206
use INVX1  _2895_
timestamp 1597059762
transform 1 0 4088 0 -1 1410
box -4 -6 36 206
use NAND2X1  _2896_
timestamp 1597059762
transform 1 0 4120 0 -1 1410
box -4 -6 52 206
use NOR3X1  _2915_
timestamp 1597059762
transform 1 0 4168 0 -1 1410
box -4 -6 132 206
use INVX1  _3345_
timestamp 1597059762
transform -1 0 4328 0 -1 1410
box -4 -6 36 206
use NAND2X1  _2902_
timestamp 1597059762
transform -1 0 4376 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3814_
timestamp 1597059762
transform -1 0 4440 0 -1 1410
box -4 -6 68 206
use OR2X2  _2276_
timestamp 1597059762
transform 1 0 4440 0 -1 1410
box -4 -6 68 206
use AOI22X1  _2962_
timestamp 1597059762
transform -1 0 4584 0 -1 1410
box -4 -6 84 206
use AND2X2  _2292_
timestamp 1597059762
transform 1 0 4584 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert50
timestamp 1597059762
transform 1 0 4648 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2238_
timestamp 1597059762
transform 1 0 4696 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2240_
timestamp 1597059762
transform 1 0 4744 0 -1 1410
box -4 -6 52 206
use AND2X2  _2239_
timestamp 1597059762
transform -1 0 4856 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2243_
timestamp 1597059762
transform -1 0 4904 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2241_
timestamp 1597059762
transform 1 0 4904 0 -1 1410
box -4 -6 52 206
use NOR2X1  _3004_
timestamp 1597059762
transform 1 0 4952 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3000_
timestamp 1597059762
transform -1 0 5064 0 -1 1410
box -4 -6 68 206
use INVX1  _2998_
timestamp 1597059762
transform -1 0 5096 0 -1 1410
box -4 -6 36 206
use AND2X2  _2295_
timestamp 1597059762
transform 1 0 5096 0 -1 1410
box -4 -6 68 206
use NOR2X1  _3041_
timestamp 1597059762
transform -1 0 5208 0 -1 1410
box -4 -6 52 206
use INVX1  _3036_
timestamp 1597059762
transform 1 0 5208 0 -1 1410
box -4 -6 36 206
use OAI22X1  _3037_
timestamp 1597059762
transform -1 0 5384 0 -1 1410
box -4 -6 84 206
use NAND3X1  _3056_
timestamp 1597059762
transform 1 0 5384 0 -1 1410
box -4 -6 68 206
use FILL  SFILL52400x12100
timestamp 1597059762
transform -1 0 5256 0 -1 1410
box -4 -6 20 206
use FILL  SFILL52560x12100
timestamp 1597059762
transform -1 0 5272 0 -1 1410
box -4 -6 20 206
use FILL  SFILL52720x12100
timestamp 1597059762
transform -1 0 5288 0 -1 1410
box -4 -6 20 206
use FILL  SFILL52880x12100
timestamp 1597059762
transform -1 0 5304 0 -1 1410
box -4 -6 20 206
use NOR2X1  _3048_
timestamp 1597059762
transform -1 0 5496 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3022_
timestamp 1597059762
transform -1 0 5560 0 -1 1410
box -4 -6 68 206
use INVX1  _3020_
timestamp 1597059762
transform -1 0 5592 0 -1 1410
box -4 -6 36 206
use OAI21X1  _3044_
timestamp 1597059762
transform -1 0 5656 0 -1 1410
box -4 -6 68 206
use INVX1  _3042_
timestamp 1597059762
transform -1 0 5688 0 -1 1410
box -4 -6 36 206
use NOR2X1  _3070_
timestamp 1597059762
transform 1 0 5688 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3066_
timestamp 1597059762
transform -1 0 5800 0 -1 1410
box -4 -6 68 206
use INVX1  _3064_
timestamp 1597059762
transform 1 0 5800 0 -1 1410
box -4 -6 36 206
use BUFX2  BUFX2_insert252
timestamp 1597059762
transform -1 0 5880 0 -1 1410
box -4 -6 52 206
use AOI22X1  _3028_
timestamp 1597059762
transform 1 0 5880 0 -1 1410
box -4 -6 84 206
use OR2X2  _2279_
timestamp 1597059762
transform -1 0 6024 0 -1 1410
box -4 -6 68 206
use AND2X2  _2297_
timestamp 1597059762
transform 1 0 6024 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2308_
timestamp 1597059762
transform -1 0 6136 0 -1 1410
box -4 -6 52 206
use AND2X2  _2309_
timestamp 1597059762
transform 1 0 6136 0 -1 1410
box -4 -6 68 206
use OAI22X1  _2310_
timestamp 1597059762
transform -1 0 6280 0 -1 1410
box -4 -6 84 206
use NOR2X1  _2306_
timestamp 1597059762
transform 1 0 6280 0 -1 1410
box -4 -6 52 206
use AND2X2  _2294_
timestamp 1597059762
transform 1 0 6328 0 -1 1410
box -4 -6 68 206
use AOI22X1  _3006_
timestamp 1597059762
transform 1 0 6392 0 -1 1410
box -4 -6 84 206
use OR2X2  _2278_
timestamp 1597059762
transform -1 0 6536 0 -1 1410
box -4 -6 68 206
use OR2X2  _2119_
timestamp 1597059762
transform 1 0 6536 0 -1 1410
box -4 -6 68 206
use NAND2X1  _2121_
timestamp 1597059762
transform 1 0 6600 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2207_
timestamp 1597059762
transform -1 0 6696 0 -1 1410
box -4 -6 52 206
use XNOR2X1  _2122_
timestamp 1597059762
transform -1 0 6808 0 -1 1410
box -4 -6 116 206
use FILL  SFILL68080x12100
timestamp 1597059762
transform -1 0 6824 0 -1 1410
box -4 -6 20 206
use FILL  SFILL68240x12100
timestamp 1597059762
transform -1 0 6840 0 -1 1410
box -4 -6 20 206
use INVX1  _2123_
timestamp 1597059762
transform 1 0 6872 0 -1 1410
box -4 -6 36 206
use OAI21X1  _2137_
timestamp 1597059762
transform 1 0 6904 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2148_
timestamp 1597059762
transform 1 0 6968 0 -1 1410
box -4 -6 52 206
use AOI21X1  _2151_
timestamp 1597059762
transform 1 0 7016 0 -1 1410
box -4 -6 68 206
use FILL  SFILL68400x12100
timestamp 1597059762
transform -1 0 6856 0 -1 1410
box -4 -6 20 206
use FILL  SFILL68560x12100
timestamp 1597059762
transform -1 0 6872 0 -1 1410
box -4 -6 20 206
use NAND2X1  _2213_
timestamp 1597059762
transform 1 0 7080 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2150_
timestamp 1597059762
transform 1 0 7128 0 -1 1410
box -4 -6 68 206
use NAND2X1  _2147_
timestamp 1597059762
transform -1 0 7240 0 -1 1410
box -4 -6 52 206
use AOI21X1  _2149_
timestamp 1597059762
transform -1 0 7304 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2140_
timestamp 1597059762
transform -1 0 7352 0 -1 1410
box -4 -6 52 206
use AND2X2  _2138_
timestamp 1597059762
transform -1 0 7416 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2139_
timestamp 1597059762
transform 1 0 7416 0 -1 1410
box -4 -6 52 206
use INVX1  _2582_
timestamp 1597059762
transform -1 0 7496 0 -1 1410
box -4 -6 36 206
use BUFX2  _2038_
timestamp 1597059762
transform 1 0 7496 0 -1 1410
box -4 -6 52 206
use FILL  FILL72240x12100
timestamp 1597059762
transform -1 0 7560 0 -1 1410
box -4 -6 20 206
use NOR2X1  _3936_
timestamp 1597059762
transform 1 0 8 0 1 1410
box -4 -6 52 206
use AOI21X1  _3937_
timestamp 1597059762
transform -1 0 120 0 1 1410
box -4 -6 68 206
use OAI21X1  _3690_
timestamp 1597059762
transform 1 0 120 0 1 1410
box -4 -6 68 206
use NAND2X1  _3689_
timestamp 1597059762
transform 1 0 184 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _4289_
timestamp 1597059762
transform 1 0 232 0 1 1410
box -4 -6 196 206
use AOI21X1  _4148_
timestamp 1597059762
transform 1 0 424 0 1 1410
box -4 -6 68 206
use NOR2X1  _4147_
timestamp 1597059762
transform -1 0 536 0 1 1410
box -4 -6 52 206
use AOI21X1  _4152_
timestamp 1597059762
transform 1 0 536 0 1 1410
box -4 -6 68 206
use NOR2X1  _4151_
timestamp 1597059762
transform -1 0 648 0 1 1410
box -4 -6 52 206
use AOI21X1  _3941_
timestamp 1597059762
transform 1 0 648 0 1 1410
box -4 -6 68 206
use NOR2X1  _3940_
timestamp 1597059762
transform -1 0 760 0 1 1410
box -4 -6 52 206
use FILL  SFILL7600x14100
timestamp 1597059762
transform 1 0 760 0 1 1410
box -4 -6 20 206
use FILL  SFILL7760x14100
timestamp 1597059762
transform 1 0 776 0 1 1410
box -4 -6 20 206
use FILL  SFILL7920x14100
timestamp 1597059762
transform 1 0 792 0 1 1410
box -4 -6 20 206
use FILL  SFILL8080x14100
timestamp 1597059762
transform 1 0 808 0 1 1410
box -4 -6 20 206
use DFFPOSX1  _4253_
timestamp 1597059762
transform 1 0 824 0 1 1410
box -4 -6 196 206
use MUX2X1  _3772_
timestamp 1597059762
transform 1 0 1016 0 1 1410
box -4 -6 100 206
use MUX2X1  _3984_
timestamp 1597059762
transform 1 0 1112 0 1 1410
box -4 -6 100 206
use NOR2X1  _3799_
timestamp 1597059762
transform 1 0 1208 0 1 1410
box -4 -6 52 206
use MUX2X1  _4032_
timestamp 1597059762
transform 1 0 1256 0 1 1410
box -4 -6 100 206
use MUX2X1  _3820_
timestamp 1597059762
transform 1 0 1352 0 1 1410
box -4 -6 100 206
use NAND2X1  _3618_
timestamp 1597059762
transform 1 0 1448 0 1 1410
box -4 -6 52 206
use OAI21X1  _3619_
timestamp 1597059762
transform 1 0 1496 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _4237_
timestamp 1597059762
transform -1 0 1752 0 1 1410
box -4 -6 196 206
use NOR2X1  _3795_
timestamp 1597059762
transform -1 0 1800 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert255
timestamp 1597059762
transform 1 0 1800 0 1 1410
box -4 -6 52 206
use INVX4  _3551_
timestamp 1597059762
transform -1 0 1896 0 1 1410
box -4 -6 52 206
use INVX4  _3557_
timestamp 1597059762
transform -1 0 1944 0 1 1410
box -4 -6 52 206
use INVX1  _3304_
timestamp 1597059762
transform 1 0 1944 0 1 1410
box -4 -6 36 206
use NOR2X1  _3305_
timestamp 1597059762
transform -1 0 2024 0 1 1410
box -4 -6 52 206
use NAND3X1  _3376_
timestamp 1597059762
transform 1 0 2024 0 1 1410
box -4 -6 68 206
use NAND2X1  _3413_
timestamp 1597059762
transform -1 0 2136 0 1 1410
box -4 -6 52 206
use NAND3X1  _3412_
timestamp 1597059762
transform -1 0 2200 0 1 1410
box -4 -6 68 206
use NAND3X1  _3313_
timestamp 1597059762
transform 1 0 2200 0 1 1410
box -4 -6 68 206
use INVX1  _3382_
timestamp 1597059762
transform 1 0 2328 0 1 1410
box -4 -6 36 206
use NAND3X1  _3383_
timestamp 1597059762
transform 1 0 2360 0 1 1410
box -4 -6 68 206
use FILL  SFILL22640x14100
timestamp 1597059762
transform 1 0 2264 0 1 1410
box -4 -6 20 206
use FILL  SFILL22800x14100
timestamp 1597059762
transform 1 0 2280 0 1 1410
box -4 -6 20 206
use FILL  SFILL22960x14100
timestamp 1597059762
transform 1 0 2296 0 1 1410
box -4 -6 20 206
use FILL  SFILL23120x14100
timestamp 1597059762
transform 1 0 2312 0 1 1410
box -4 -6 20 206
use NAND3X1  _3306_
timestamp 1597059762
transform 1 0 2424 0 1 1410
box -4 -6 68 206
use NAND3X1  _3398_
timestamp 1597059762
transform -1 0 2552 0 1 1410
box -4 -6 68 206
use NAND2X1  _3399_
timestamp 1597059762
transform -1 0 2600 0 1 1410
box -4 -6 52 206
use INVX4  _3296_
timestamp 1597059762
transform -1 0 2648 0 1 1410
box -4 -6 52 206
use NAND3X1  _3405_
timestamp 1597059762
transform -1 0 2712 0 1 1410
box -4 -6 68 206
use INVX4  _3548_
timestamp 1597059762
transform -1 0 2760 0 1 1410
box -4 -6 52 206
use OAI21X1  _3318_
timestamp 1597059762
transform -1 0 2824 0 1 1410
box -4 -6 68 206
use OAI21X1  _3395_
timestamp 1597059762
transform 1 0 2824 0 1 1410
box -4 -6 68 206
use NAND2X1  _3379_
timestamp 1597059762
transform 1 0 2888 0 1 1410
box -4 -6 52 206
use OAI21X1  _3402_
timestamp 1597059762
transform 1 0 2936 0 1 1410
box -4 -6 68 206
use NAND3X1  _3342_
timestamp 1597059762
transform -1 0 3064 0 1 1410
box -4 -6 68 206
use OAI21X1  _3339_
timestamp 1597059762
transform 1 0 3064 0 1 1410
box -4 -6 68 206
use NAND2X1  _3343_
timestamp 1597059762
transform -1 0 3176 0 1 1410
box -4 -6 52 206
use INVX1  _3299_
timestamp 1597059762
transform 1 0 3176 0 1 1410
box -4 -6 36 206
use NAND2X1  _3300_
timestamp 1597059762
transform -1 0 3256 0 1 1410
box -4 -6 52 206
use INVX1  _3338_
timestamp 1597059762
transform -1 0 3288 0 1 1410
box -4 -6 36 206
use OR2X2  _3298_
timestamp 1597059762
transform -1 0 3352 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert270
timestamp 1597059762
transform 1 0 3352 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _4321_
timestamp 1597059762
transform 1 0 3400 0 1 1410
box -4 -6 196 206
use BUFX2  BUFX2_insert268
timestamp 1597059762
transform 1 0 3592 0 1 1410
box -4 -6 52 206
use NAND2X1  _2901_
timestamp 1597059762
transform 1 0 3640 0 1 1410
box -4 -6 52 206
use NOR2X1  _2876_
timestamp 1597059762
transform 1 0 3688 0 1 1410
box -4 -6 52 206
use INVX1  _2878_
timestamp 1597059762
transform 1 0 3736 0 1 1410
box -4 -6 36 206
use FILL  SFILL37680x14100
timestamp 1597059762
transform 1 0 3768 0 1 1410
box -4 -6 20 206
use FILL  SFILL37840x14100
timestamp 1597059762
transform 1 0 3784 0 1 1410
box -4 -6 20 206
use FILL  SFILL38000x14100
timestamp 1597059762
transform 1 0 3800 0 1 1410
box -4 -6 20 206
use FILL  SFILL38160x14100
timestamp 1597059762
transform 1 0 3816 0 1 1410
box -4 -6 20 206
use NAND2X1  _2879_
timestamp 1597059762
transform -1 0 3880 0 1 1410
box -4 -6 52 206
use AOI21X1  _3815_
timestamp 1597059762
transform 1 0 3880 0 1 1410
box -4 -6 68 206
use NOR3X1  _2916_
timestamp 1597059762
transform -1 0 4072 0 1 1410
box -4 -6 132 206
use NAND3X1  _2887_
timestamp 1597059762
transform -1 0 4136 0 1 1410
box -4 -6 68 206
use NOR2X1  _2903_
timestamp 1597059762
transform 1 0 4136 0 1 1410
box -4 -6 52 206
use NOR2X1  _2918_
timestamp 1597059762
transform -1 0 4232 0 1 1410
box -4 -6 52 206
use AND2X2  _2919_
timestamp 1597059762
transform 1 0 4232 0 1 1410
box -4 -6 68 206
use AOI21X1  _4038_
timestamp 1597059762
transform 1 0 4296 0 1 1410
box -4 -6 68 206
use OAI21X1  _4037_
timestamp 1597059762
transform -1 0 4424 0 1 1410
box -4 -6 68 206
use INVX1  _2992_
timestamp 1597059762
transform 1 0 4424 0 1 1410
box -4 -6 36 206
use OAI22X1  _2993_
timestamp 1597059762
transform -1 0 4536 0 1 1410
box -4 -6 84 206
use INVX1  _2991_
timestamp 1597059762
transform 1 0 4536 0 1 1410
box -4 -6 36 206
use NOR2X1  _2997_
timestamp 1597059762
transform -1 0 4616 0 1 1410
box -4 -6 52 206
use OAI21X1  _2996_
timestamp 1597059762
transform -1 0 4680 0 1 1410
box -4 -6 68 206
use INVX1  _2994_
timestamp 1597059762
transform -1 0 4712 0 1 1410
box -4 -6 36 206
use NAND3X1  _3012_
timestamp 1597059762
transform 1 0 4712 0 1 1410
box -4 -6 68 206
use AND2X2  _2242_
timestamp 1597059762
transform 1 0 4776 0 1 1410
box -4 -6 68 206
use INVX1  _3013_
timestamp 1597059762
transform 1 0 4840 0 1 1410
box -4 -6 36 206
use OAI22X1  _3015_
timestamp 1597059762
transform 1 0 4872 0 1 1410
box -4 -6 84 206
use INVX1  _3014_
timestamp 1597059762
transform -1 0 4984 0 1 1410
box -4 -6 36 206
use OAI21X1  _3003_
timestamp 1597059762
transform -1 0 5048 0 1 1410
box -4 -6 68 206
use INVX1  _3001_
timestamp 1597059762
transform -1 0 5080 0 1 1410
box -4 -6 36 206
use INVX1  _3038_
timestamp 1597059762
transform 1 0 5080 0 1 1410
box -4 -6 36 206
use OAI21X1  _3040_
timestamp 1597059762
transform -1 0 5176 0 1 1410
box -4 -6 68 206
use INVX1  _3060_
timestamp 1597059762
transform 1 0 5176 0 1 1410
box -4 -6 36 206
use OAI21X1  _3062_
timestamp 1597059762
transform 1 0 5208 0 1 1410
box -4 -6 68 206
use NOR2X1  _3063_
timestamp 1597059762
transform 1 0 5336 0 1 1410
box -4 -6 52 206
use NAND3X1  _3078_
timestamp 1597059762
transform -1 0 5448 0 1 1410
box -4 -6 68 206
use FILL  SFILL52720x14100
timestamp 1597059762
transform 1 0 5272 0 1 1410
box -4 -6 20 206
use FILL  SFILL52880x14100
timestamp 1597059762
transform 1 0 5288 0 1 1410
box -4 -6 20 206
use FILL  SFILL53040x14100
timestamp 1597059762
transform 1 0 5304 0 1 1410
box -4 -6 20 206
use FILL  SFILL53200x14100
timestamp 1597059762
transform 1 0 5320 0 1 1410
box -4 -6 20 206
use INVX1  _3058_
timestamp 1597059762
transform 1 0 5448 0 1 1410
box -4 -6 36 206
use OAI22X1  _3059_
timestamp 1597059762
transform -1 0 5560 0 1 1410
box -4 -6 84 206
use OAI21X1  _3047_
timestamp 1597059762
transform -1 0 5624 0 1 1410
box -4 -6 68 206
use INVX1  _3045_
timestamp 1597059762
transform 1 0 5624 0 1 1410
box -4 -6 36 206
use OAI21X1  _3069_
timestamp 1597059762
transform -1 0 5720 0 1 1410
box -4 -6 68 206
use INVX1  _3067_
timestamp 1597059762
transform -1 0 5752 0 1 1410
box -4 -6 36 206
use INVX1  _3057_
timestamp 1597059762
transform -1 0 5784 0 1 1410
box -4 -6 36 206
use NOR2X1  _2247_
timestamp 1597059762
transform 1 0 5784 0 1 1410
box -4 -6 52 206
use NOR2X1  _2249_
timestamp 1597059762
transform 1 0 5832 0 1 1410
box -4 -6 52 206
use AND2X2  _2248_
timestamp 1597059762
transform -1 0 5944 0 1 1410
box -4 -6 68 206
use NOR2X1  _3055_
timestamp 1597059762
transform -1 0 5992 0 1 1410
box -4 -6 52 206
use OR2X2  _2281_
timestamp 1597059762
transform 1 0 5992 0 1 1410
box -4 -6 68 206
use AOI22X1  _3072_
timestamp 1597059762
transform -1 0 6136 0 1 1410
box -4 -6 84 206
use NAND2X1  _3073_
timestamp 1597059762
transform -1 0 6184 0 1 1410
box -4 -6 52 206
use NOR2X1  _3077_
timestamp 1597059762
transform -1 0 6232 0 1 1410
box -4 -6 52 206
use NOR2X1  _3011_
timestamp 1597059762
transform -1 0 6280 0 1 1410
box -4 -6 52 206
use NAND2X1  _3007_
timestamp 1597059762
transform 1 0 6280 0 1 1410
box -4 -6 52 206
use NAND2X1  _3054_
timestamp 1597059762
transform -1 0 6376 0 1 1410
box -4 -6 52 206
use AOI22X1  _3052_
timestamp 1597059762
transform -1 0 6456 0 1 1410
box -4 -6 84 206
use NAND2X1  _3010_
timestamp 1597059762
transform -1 0 6504 0 1 1410
box -4 -6 52 206
use AOI22X1  _3008_
timestamp 1597059762
transform -1 0 6584 0 1 1410
box -4 -6 84 206
use AOI22X1  _3074_
timestamp 1597059762
transform 1 0 6584 0 1 1410
box -4 -6 84 206
use NAND2X1  _3076_
timestamp 1597059762
transform 1 0 6664 0 1 1410
box -4 -6 52 206
use AOI22X1  _3009_
timestamp 1597059762
transform -1 0 6792 0 1 1410
box -4 -6 84 206
use FILL  SFILL67920x14100
timestamp 1597059762
transform 1 0 6792 0 1 1410
box -4 -6 20 206
use FILL  SFILL68080x14100
timestamp 1597059762
transform 1 0 6808 0 1 1410
box -4 -6 20 206
use FILL  SFILL68240x14100
timestamp 1597059762
transform 1 0 6824 0 1 1410
box -4 -6 20 206
use AOI22X1  _3053_
timestamp 1597059762
transform 1 0 6856 0 1 1410
box -4 -6 84 206
use AOI22X1  _3075_
timestamp 1597059762
transform 1 0 6936 0 1 1410
box -4 -6 84 206
use XOR2X1  _2141_
timestamp 1597059762
transform 1 0 7016 0 1 1410
box -4 -6 116 206
use FILL  SFILL68400x14100
timestamp 1597059762
transform 1 0 6840 0 1 1410
box -4 -6 20 206
use NAND2X1  _2118_
timestamp 1597059762
transform -1 0 7176 0 1 1410
box -4 -6 52 206
use XNOR2X1  _2146_
timestamp 1597059762
transform -1 0 7288 0 1 1410
box -4 -6 116 206
use AOI21X1  _2142_
timestamp 1597059762
transform 1 0 7288 0 1 1410
box -4 -6 68 206
use XNOR2X1  _2371_
timestamp 1597059762
transform -1 0 7464 0 1 1410
box -4 -6 116 206
use NAND2X1  _2099_
timestamp 1597059762
transform -1 0 7512 0 1 1410
box -4 -6 52 206
use BUFX2  _2034_
timestamp 1597059762
transform 1 0 7512 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _4269_
timestamp 1597059762
transform -1 0 200 0 -1 1810
box -4 -6 196 206
use AOI21X1  _3933_
timestamp 1597059762
transform 1 0 200 0 -1 1810
box -4 -6 68 206
use NOR2X1  _3932_
timestamp 1597059762
transform -1 0 312 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert76
timestamp 1597059762
transform 1 0 312 0 -1 1810
box -4 -6 52 206
use AOI21X1  _4144_
timestamp 1597059762
transform 1 0 360 0 -1 1810
box -4 -6 68 206
use NOR2X1  _4143_
timestamp 1597059762
transform -1 0 472 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3693_
timestamp 1597059762
transform 1 0 472 0 -1 1810
box -4 -6 52 206
use OAI21X1  _3694_
timestamp 1597059762
transform -1 0 584 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  _4193_
timestamp 1597059762
transform -1 0 776 0 -1 1810
box -4 -6 196 206
use FILL  SFILL7760x16100
timestamp 1597059762
transform -1 0 792 0 -1 1810
box -4 -6 20 206
use FILL  SFILL7920x16100
timestamp 1597059762
transform -1 0 808 0 -1 1810
box -4 -6 20 206
use FILL  SFILL8080x16100
timestamp 1597059762
transform -1 0 824 0 -1 1810
box -4 -6 20 206
use OAI21X1  _3774_
timestamp 1597059762
transform 1 0 840 0 -1 1810
box -4 -6 68 206
use OAI22X1  _3775_
timestamp 1597059762
transform 1 0 904 0 -1 1810
box -4 -6 84 206
use OAI21X1  _3986_
timestamp 1597059762
transform 1 0 984 0 -1 1810
box -4 -6 68 206
use FILL  SFILL8240x16100
timestamp 1597059762
transform -1 0 840 0 -1 1810
box -4 -6 20 206
use OAI22X1  _3987_
timestamp 1597059762
transform 1 0 1048 0 -1 1810
box -4 -6 84 206
use MUX2X1  _3992_
timestamp 1597059762
transform 1 0 1128 0 -1 1810
box -4 -6 100 206
use NOR2X1  _3773_
timestamp 1597059762
transform -1 0 1272 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3985_
timestamp 1597059762
transform 1 0 1272 0 -1 1810
box -4 -6 52 206
use NOR2X1  _4033_
timestamp 1597059762
transform -1 0 1368 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3821_
timestamp 1597059762
transform 1 0 1368 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3823_
timestamp 1597059762
transform -1 0 1496 0 -1 1810
box -4 -6 84 206
use OAI22X1  _4035_
timestamp 1597059762
transform -1 0 1576 0 -1 1810
box -4 -6 84 206
use OAI21X1  _3822_
timestamp 1597059762
transform -1 0 1640 0 -1 1810
box -4 -6 68 206
use OAI21X1  _4034_
timestamp 1597059762
transform -1 0 1704 0 -1 1810
box -4 -6 68 206
use MUX2X1  _3824_
timestamp 1597059762
transform -1 0 1800 0 -1 1810
box -4 -6 100 206
use NOR2X1  _3817_
timestamp 1597059762
transform -1 0 1848 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3819_
timestamp 1597059762
transform 1 0 1848 0 -1 1810
box -4 -6 84 206
use OAI21X1  _3818_
timestamp 1597059762
transform -1 0 1992 0 -1 1810
box -4 -6 68 206
use NOR2X1  _4029_
timestamp 1597059762
transform -1 0 2040 0 -1 1810
box -4 -6 52 206
use OAI21X1  _4030_
timestamp 1597059762
transform 1 0 2040 0 -1 1810
box -4 -6 68 206
use OAI22X1  _4031_
timestamp 1597059762
transform 1 0 2104 0 -1 1810
box -4 -6 84 206
use MUX2X1  _4036_
timestamp 1597059762
transform 1 0 2184 0 -1 1810
box -4 -6 100 206
use NAND3X1  _3377_
timestamp 1597059762
transform -1 0 2408 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3378_
timestamp 1597059762
transform -1 0 2456 0 -1 1810
box -4 -6 52 206
use FILL  SFILL22800x16100
timestamp 1597059762
transform -1 0 2296 0 -1 1810
box -4 -6 20 206
use FILL  SFILL22960x16100
timestamp 1597059762
transform -1 0 2312 0 -1 1810
box -4 -6 20 206
use FILL  SFILL23120x16100
timestamp 1597059762
transform -1 0 2328 0 -1 1810
box -4 -6 20 206
use FILL  SFILL23280x16100
timestamp 1597059762
transform -1 0 2344 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  _4209_
timestamp 1597059762
transform -1 0 2648 0 -1 1810
box -4 -6 196 206
use NAND2X1  _3392_
timestamp 1597059762
transform 1 0 2648 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3391_
timestamp 1597059762
transform -1 0 2760 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3315_
timestamp 1597059762
transform 1 0 2760 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3314_
timestamp 1597059762
transform -1 0 2872 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3406_
timestamp 1597059762
transform -1 0 2920 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3385_
timestamp 1597059762
transform 1 0 2920 0 -1 1810
box -4 -6 52 206
use NAND3X1  _3384_
timestamp 1597059762
transform -1 0 3032 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3307_
timestamp 1597059762
transform -1 0 3096 0 -1 1810
box -4 -6 68 206
use NAND3X1  _3363_
timestamp 1597059762
transform 1 0 3096 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3364_
timestamp 1597059762
transform -1 0 3208 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3308_
timestamp 1597059762
transform -1 0 3256 0 -1 1810
box -4 -6 52 206
use OAI21X1  _3360_
timestamp 1597059762
transform 1 0 3256 0 -1 1810
box -4 -6 68 206
use INVX1  _3317_
timestamp 1597059762
transform -1 0 3352 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  _4306_
timestamp 1597059762
transform 1 0 3352 0 -1 1810
box -4 -6 196 206
use AOI21X1  _3826_
timestamp 1597059762
transform 1 0 3544 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert100
timestamp 1597059762
transform 1 0 3608 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert250
timestamp 1597059762
transform 1 0 3656 0 -1 1810
box -4 -6 52 206
use AOI21X1  _3994_
timestamp 1597059762
transform 1 0 3704 0 -1 1810
box -4 -6 68 206
use FILL  SFILL37680x16100
timestamp 1597059762
transform -1 0 3784 0 -1 1810
box -4 -6 20 206
use FILL  SFILL37840x16100
timestamp 1597059762
transform -1 0 3800 0 -1 1810
box -4 -6 20 206
use FILL  SFILL38000x16100
timestamp 1597059762
transform -1 0 3816 0 -1 1810
box -4 -6 20 206
use FILL  SFILL38160x16100
timestamp 1597059762
transform -1 0 3832 0 -1 1810
box -4 -6 20 206
use OAI21X1  _3993_
timestamp 1597059762
transform -1 0 3896 0 -1 1810
box -4 -6 68 206
use OAI21X1  _3825_
timestamp 1597059762
transform -1 0 3960 0 -1 1810
box -4 -6 68 206
use NOR3X1  _2912_
timestamp 1597059762
transform -1 0 4088 0 -1 1810
box -4 -6 132 206
use INVX1  _2891_
timestamp 1597059762
transform 1 0 4088 0 -1 1810
box -4 -6 36 206
use NAND2X1  _2892_
timestamp 1597059762
transform -1 0 4168 0 -1 1810
box -4 -6 52 206
use OR2X2  _2884_
timestamp 1597059762
transform 1 0 4168 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2885_
timestamp 1597059762
transform -1 0 4280 0 -1 1810
box -4 -6 52 206
use NOR2X1  _2909_
timestamp 1597059762
transform 1 0 4280 0 -1 1810
box -4 -6 52 206
use NOR3X1  _2908_
timestamp 1597059762
transform -1 0 4456 0 -1 1810
box -4 -6 132 206
use INVX1  _2873_
timestamp 1597059762
transform 1 0 4456 0 -1 1810
box -4 -6 36 206
use NAND2X1  _2874_
timestamp 1597059762
transform 1 0 4488 0 -1 1810
box -4 -6 52 206
use NOR3X1  _2920_
timestamp 1597059762
transform 1 0 4536 0 -1 1810
box -4 -6 132 206
use NAND2X1  _2995_
timestamp 1597059762
transform -1 0 4712 0 -1 1810
box -4 -6 52 206
use NAND2X1  _2963_
timestamp 1597059762
transform -1 0 4760 0 -1 1810
box -4 -6 52 206
use NAND2X1  _2958_
timestamp 1597059762
transform 1 0 4760 0 -1 1810
box -4 -6 52 206
use NAND2X1  _2973_
timestamp 1597059762
transform 1 0 4808 0 -1 1810
box -4 -6 52 206
use OAI21X1  _2974_
timestamp 1597059762
transform -1 0 4920 0 -1 1810
box -4 -6 68 206
use INVX1  _2972_
timestamp 1597059762
transform -1 0 4952 0 -1 1810
box -4 -6 36 206
use NOR2X1  _2975_
timestamp 1597059762
transform 1 0 4952 0 -1 1810
box -4 -6 52 206
use OAI22X1  _2971_
timestamp 1597059762
transform 1 0 5000 0 -1 1810
box -4 -6 84 206
use INVX1  _2970_
timestamp 1597059762
transform 1 0 5080 0 -1 1810
box -4 -6 36 206
use NAND2X1  _3002_
timestamp 1597059762
transform -1 0 5160 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3039_
timestamp 1597059762
transform -1 0 5208 0 -1 1810
box -4 -6 52 206
use NAND3X1  _2990_
timestamp 1597059762
transform 1 0 5208 0 -1 1810
box -4 -6 68 206
use INVX1  _3016_
timestamp 1597059762
transform 1 0 5336 0 -1 1810
box -4 -6 36 206
use NOR2X1  _3019_
timestamp 1597059762
transform -1 0 5416 0 -1 1810
box -4 -6 52 206
use OAI21X1  _3018_
timestamp 1597059762
transform 1 0 5416 0 -1 1810
box -4 -6 68 206
use FILL  SFILL52720x16100
timestamp 1597059762
transform -1 0 5288 0 -1 1810
box -4 -6 20 206
use FILL  SFILL52880x16100
timestamp 1597059762
transform -1 0 5304 0 -1 1810
box -4 -6 20 206
use FILL  SFILL53040x16100
timestamp 1597059762
transform -1 0 5320 0 -1 1810
box -4 -6 20 206
use FILL  SFILL53200x16100
timestamp 1597059762
transform -1 0 5336 0 -1 1810
box -4 -6 20 206
use NAND3X1  _3034_
timestamp 1597059762
transform 1 0 5480 0 -1 1810
box -4 -6 68 206
use NOR2X1  _3026_
timestamp 1597059762
transform -1 0 5592 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3046_
timestamp 1597059762
transform -1 0 5640 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3068_
timestamp 1597059762
transform 1 0 5640 0 -1 1810
box -4 -6 52 206
use OR2X2  _2280_
timestamp 1597059762
transform 1 0 5688 0 -1 1810
box -4 -6 68 206
use AOI22X1  _3050_
timestamp 1597059762
transform -1 0 5832 0 -1 1810
box -4 -6 84 206
use INVX1  _3023_
timestamp 1597059762
transform -1 0 5864 0 -1 1810
box -4 -6 36 206
use OAI21X1  _3025_
timestamp 1597059762
transform 1 0 5864 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3024_
timestamp 1597059762
transform -1 0 5976 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3051_
timestamp 1597059762
transform -1 0 6024 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3029_
timestamp 1597059762
transform -1 0 6072 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3033_
timestamp 1597059762
transform -1 0 6120 0 -1 1810
box -4 -6 52 206
use AOI22X1  _3027_
timestamp 1597059762
transform -1 0 6200 0 -1 1810
box -4 -6 84 206
use AOI22X1  _3071_
timestamp 1597059762
transform -1 0 6280 0 -1 1810
box -4 -6 84 206
use AOI22X1  _3005_
timestamp 1597059762
transform 1 0 6280 0 -1 1810
box -4 -6 84 206
use AOI22X1  _3030_
timestamp 1597059762
transform 1 0 6360 0 -1 1810
box -4 -6 84 206
use NAND2X1  _3032_
timestamp 1597059762
transform 1 0 6440 0 -1 1810
box -4 -6 52 206
use AOI22X1  _3031_
timestamp 1597059762
transform -1 0 6568 0 -1 1810
box -4 -6 84 206
use AOI22X1  _2984_
timestamp 1597059762
transform 1 0 6568 0 -1 1810
box -4 -6 84 206
use NAND2X1  _2985_
timestamp 1597059762
transform -1 0 6696 0 -1 1810
box -4 -6 52 206
use NOR2X1  _2989_
timestamp 1597059762
transform -1 0 6744 0 -1 1810
box -4 -6 52 206
use AOI22X1  _2983_
timestamp 1597059762
transform -1 0 6888 0 -1 1810
box -4 -6 84 206
use FILL  SFILL67440x16100
timestamp 1597059762
transform -1 0 6760 0 -1 1810
box -4 -6 20 206
use FILL  SFILL67600x16100
timestamp 1597059762
transform -1 0 6776 0 -1 1810
box -4 -6 20 206
use FILL  SFILL67760x16100
timestamp 1597059762
transform -1 0 6792 0 -1 1810
box -4 -6 20 206
use FILL  SFILL67920x16100
timestamp 1597059762
transform -1 0 6808 0 -1 1810
box -4 -6 20 206
use AOI22X1  _2986_
timestamp 1597059762
transform 1 0 6888 0 -1 1810
box -4 -6 84 206
use NAND2X1  _2988_
timestamp 1597059762
transform 1 0 6968 0 -1 1810
box -4 -6 52 206
use AOI22X1  _2987_
timestamp 1597059762
transform 1 0 7016 0 -1 1810
box -4 -6 84 206
use AOI21X1  _2214_
timestamp 1597059762
transform -1 0 7160 0 -1 1810
box -4 -6 68 206
use XNOR2X1  _2114_
timestamp 1597059762
transform 1 0 7160 0 -1 1810
box -4 -6 116 206
use NAND3X1  _2115_
timestamp 1597059762
transform 1 0 7272 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2113_
timestamp 1597059762
transform -1 0 7384 0 -1 1810
box -4 -6 52 206
use AOI21X1  _2117_
timestamp 1597059762
transform -1 0 7448 0 -1 1810
box -4 -6 68 206
use INVX1  _2116_
timestamp 1597059762
transform 1 0 7448 0 -1 1810
box -4 -6 36 206
use BUFX2  BUFX2_insert156
timestamp 1597059762
transform 1 0 7480 0 -1 1810
box -4 -6 52 206
use INVX1  _2824_
timestamp 1597059762
transform -1 0 7560 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  _4189_
timestamp 1597059762
transform -1 0 200 0 1 1810
box -4 -6 196 206
use OAI21X1  _3686_
timestamp 1597059762
transform 1 0 200 0 1 1810
box -4 -6 68 206
use NAND2X1  _3685_
timestamp 1597059762
transform -1 0 312 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _4285_
timestamp 1597059762
transform 1 0 312 0 1 1810
box -4 -6 196 206
use MUX2X1  _3776_
timestamp 1597059762
transform 1 0 504 0 1 1810
box -4 -6 100 206
use MUX2X1  _3988_
timestamp 1597059762
transform -1 0 696 0 1 1810
box -4 -6 100 206
use DFFPOSX1  _4205_
timestamp 1597059762
transform 1 0 760 0 1 1810
box -4 -6 196 206
use FILL  SFILL6960x18100
timestamp 1597059762
transform 1 0 696 0 1 1810
box -4 -6 20 206
use FILL  SFILL7120x18100
timestamp 1597059762
transform 1 0 712 0 1 1810
box -4 -6 20 206
use FILL  SFILL7280x18100
timestamp 1597059762
transform 1 0 728 0 1 1810
box -4 -6 20 206
use FILL  SFILL7440x18100
timestamp 1597059762
transform 1 0 744 0 1 1810
box -4 -6 20 206
use OAI21X1  _3585_
timestamp 1597059762
transform 1 0 952 0 1 1810
box -4 -6 68 206
use NAND2X1  _3584_
timestamp 1597059762
transform 1 0 1016 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _4207_
timestamp 1597059762
transform 1 0 1064 0 1 1810
box -4 -6 196 206
use OAI21X1  _3589_
timestamp 1597059762
transform -1 0 1320 0 1 1810
box -4 -6 68 206
use NAND2X1  _3588_
timestamp 1597059762
transform -1 0 1368 0 1 1810
box -4 -6 52 206
use OAI22X1  _3991_
timestamp 1597059762
transform -1 0 1448 0 1 1810
box -4 -6 84 206
use NOR2X1  _3989_
timestamp 1597059762
transform -1 0 1496 0 1 1810
box -4 -6 52 206
use NOR2X1  _3777_
timestamp 1597059762
transform 1 0 1496 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert259
timestamp 1597059762
transform -1 0 1592 0 1 1810
box -4 -6 52 206
use NOR2X1  _3726_
timestamp 1597059762
transform -1 0 1640 0 1 1810
box -4 -6 52 206
use AOI21X1  _3727_
timestamp 1597059762
transform -1 0 1704 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _4225_
timestamp 1597059762
transform -1 0 1896 0 1 1810
box -4 -6 196 206
use OAI21X1  _3627_
timestamp 1597059762
transform 1 0 1896 0 1 1810
box -4 -6 68 206
use NAND2X1  _3626_
timestamp 1597059762
transform -1 0 2008 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _4241_
timestamp 1597059762
transform 1 0 2008 0 1 1810
box -4 -6 196 206
use MUX2X1  _3816_
timestamp 1597059762
transform 1 0 2200 0 1 1810
box -4 -6 100 206
use MUX2X1  _4028_
timestamp 1597059762
transform -1 0 2456 0 1 1810
box -4 -6 100 206
use FILL  SFILL22960x18100
timestamp 1597059762
transform 1 0 2296 0 1 1810
box -4 -6 20 206
use FILL  SFILL23120x18100
timestamp 1597059762
transform 1 0 2312 0 1 1810
box -4 -6 20 206
use FILL  SFILL23280x18100
timestamp 1597059762
transform 1 0 2328 0 1 1810
box -4 -6 20 206
use FILL  SFILL23440x18100
timestamp 1597059762
transform 1 0 2344 0 1 1810
box -4 -6 20 206
use NOR2X1  _3659_
timestamp 1597059762
transform 1 0 2456 0 1 1810
box -4 -6 52 206
use AOI21X1  _3660_
timestamp 1597059762
transform -1 0 2568 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _4257_
timestamp 1597059762
transform 1 0 2568 0 1 1810
box -4 -6 196 206
use NAND2X1  _3592_
timestamp 1597059762
transform 1 0 2760 0 1 1810
box -4 -6 52 206
use OAI21X1  _3593_
timestamp 1597059762
transform -1 0 2872 0 1 1810
box -4 -6 68 206
use INVX4  _3533_
timestamp 1597059762
transform 1 0 2872 0 1 1810
box -4 -6 52 206
use INVX4  _3563_
timestamp 1597059762
transform -1 0 2968 0 1 1810
box -4 -6 52 206
use INVX4  _3572_
timestamp 1597059762
transform 1 0 2968 0 1 1810
box -4 -6 52 206
use INVX4  _3539_
timestamp 1597059762
transform -1 0 3064 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _4177_
timestamp 1597059762
transform -1 0 3256 0 1 1810
box -4 -6 196 206
use INVX4  _3522_
timestamp 1597059762
transform 1 0 3256 0 1 1810
box -4 -6 52 206
use OAI21X1  _3301_
timestamp 1597059762
transform 1 0 3304 0 1 1810
box -4 -6 68 206
use OAI21X1  _3367_
timestamp 1597059762
transform 1 0 3368 0 1 1810
box -4 -6 68 206
use OAI21X1  _3381_
timestamp 1597059762
transform 1 0 3432 0 1 1810
box -4 -6 68 206
use OAI21X1  _3374_
timestamp 1597059762
transform 1 0 3496 0 1 1810
box -4 -6 68 206
use OAI21X1  _3388_
timestamp 1597059762
transform 1 0 3560 0 1 1810
box -4 -6 68 206
use OAI21X1  _3311_
timestamp 1597059762
transform 1 0 3624 0 1 1810
box -4 -6 68 206
use OAI21X1  _3409_
timestamp 1597059762
transform 1 0 3688 0 1 1810
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert24
timestamp 1597059762
transform -1 0 3960 0 1 1810
box -4 -6 148 206
use FILL  SFILL37520x18100
timestamp 1597059762
transform 1 0 3752 0 1 1810
box -4 -6 20 206
use FILL  SFILL37680x18100
timestamp 1597059762
transform 1 0 3768 0 1 1810
box -4 -6 20 206
use FILL  SFILL37840x18100
timestamp 1597059762
transform 1 0 3784 0 1 1810
box -4 -6 20 206
use FILL  SFILL38000x18100
timestamp 1597059762
transform 1 0 3800 0 1 1810
box -4 -6 20 206
use DFFPOSX1  _4301_
timestamp 1597059762
transform 1 0 3960 0 1 1810
box -4 -6 196 206
use BUFX2  BUFX2_insert90
timestamp 1597059762
transform -1 0 4200 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert136
timestamp 1597059762
transform 1 0 4200 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert178
timestamp 1597059762
transform -1 0 4296 0 1 1810
box -4 -6 52 206
use INVX1  _2880_
timestamp 1597059762
transform 1 0 4296 0 1 1810
box -4 -6 36 206
use NOR2X1  _2897_
timestamp 1597059762
transform 1 0 4328 0 1 1810
box -4 -6 52 206
use INVX1  _2893_
timestamp 1597059762
transform 1 0 4376 0 1 1810
box -4 -6 36 206
use NAND2X1  _2905_
timestamp 1597059762
transform -1 0 4456 0 1 1810
box -4 -6 52 206
use NAND2X1  _2894_
timestamp 1597059762
transform -1 0 4504 0 1 1810
box -4 -6 52 206
use NOR2X1  _2911_
timestamp 1597059762
transform 1 0 4504 0 1 1810
box -4 -6 52 206
use NAND2X1  _2877_
timestamp 1597059762
transform 1 0 4552 0 1 1810
box -4 -6 52 206
use INVX1  _2875_
timestamp 1597059762
transform 1 0 4600 0 1 1810
box -4 -6 36 206
use NAND2X1  _2881_
timestamp 1597059762
transform 1 0 4632 0 1 1810
box -4 -6 52 206
use NAND3X1  _2968_
timestamp 1597059762
transform 1 0 4680 0 1 1810
box -4 -6 68 206
use NOR2X1  _2967_
timestamp 1597059762
transform -1 0 4792 0 1 1810
box -4 -6 52 206
use AOI22X1  _2961_
timestamp 1597059762
transform -1 0 4872 0 1 1810
box -4 -6 84 206
use OAI21X1  _2959_
timestamp 1597059762
transform -1 0 4936 0 1 1810
box -4 -6 68 206
use INVX1  _2957_
timestamp 1597059762
transform -1 0 4968 0 1 1810
box -4 -6 36 206
use NOR2X1  _2960_
timestamp 1597059762
transform 1 0 4968 0 1 1810
box -4 -6 52 206
use OAI21X1  _2956_
timestamp 1597059762
transform -1 0 5080 0 1 1810
box -4 -6 68 206
use INVX1  _2954_
timestamp 1597059762
transform 1 0 5080 0 1 1810
box -4 -6 36 206
use XNOR2X1  _2359_
timestamp 1597059762
transform -1 0 5224 0 1 1810
box -4 -6 116 206
use INVX1  _2979_
timestamp 1597059762
transform 1 0 5224 0 1 1810
box -4 -6 36 206
use OAI21X1  _2981_
timestamp 1597059762
transform 1 0 5320 0 1 1810
box -4 -6 68 206
use NOR2X1  _2982_
timestamp 1597059762
transform 1 0 5384 0 1 1810
box -4 -6 52 206
use FILL  SFILL52560x18100
timestamp 1597059762
transform 1 0 5256 0 1 1810
box -4 -6 20 206
use FILL  SFILL52720x18100
timestamp 1597059762
transform 1 0 5272 0 1 1810
box -4 -6 20 206
use FILL  SFILL52880x18100
timestamp 1597059762
transform 1 0 5288 0 1 1810
box -4 -6 20 206
use FILL  SFILL53040x18100
timestamp 1597059762
transform 1 0 5304 0 1 1810
box -4 -6 20 206
use OAI21X1  _2978_
timestamp 1597059762
transform -1 0 5496 0 1 1810
box -4 -6 68 206
use INVX1  _2976_
timestamp 1597059762
transform -1 0 5528 0 1 1810
box -4 -6 36 206
use NAND2X1  _2980_
timestamp 1597059762
transform -1 0 5576 0 1 1810
box -4 -6 52 206
use NAND2X1  _3061_
timestamp 1597059762
transform 1 0 5576 0 1 1810
box -4 -6 52 206
use NAND2X1  _3017_
timestamp 1597059762
transform -1 0 5672 0 1 1810
box -4 -6 52 206
use AND2X2  _2296_
timestamp 1597059762
transform 1 0 5672 0 1 1810
box -4 -6 68 206
use NOR2X1  _2329_
timestamp 1597059762
transform -1 0 5784 0 1 1810
box -4 -6 52 206
use AND2X2  _2330_
timestamp 1597059762
transform 1 0 5784 0 1 1810
box -4 -6 68 206
use AOI21X1  _2446_
timestamp 1597059762
transform 1 0 5848 0 1 1810
box -4 -6 68 206
use OAI22X1  _2333_
timestamp 1597059762
transform 1 0 5912 0 1 1810
box -4 -6 84 206
use NOR2X1  _2331_
timestamp 1597059762
transform -1 0 6040 0 1 1810
box -4 -6 52 206
use AND2X2  _2332_
timestamp 1597059762
transform 1 0 6040 0 1 1810
box -4 -6 68 206
use AOI22X1  _3049_
timestamp 1597059762
transform -1 0 6184 0 1 1810
box -4 -6 84 206
use NOR2X1  _2311_
timestamp 1597059762
transform 1 0 6184 0 1 1810
box -4 -6 52 206
use AND2X2  _2312_
timestamp 1597059762
transform 1 0 6232 0 1 1810
box -4 -6 68 206
use NOR2X1  _2316_
timestamp 1597059762
transform 1 0 6296 0 1 1810
box -4 -6 52 206
use OAI22X1  _2315_
timestamp 1597059762
transform 1 0 6344 0 1 1810
box -4 -6 84 206
use BUFX2  BUFX2_insert177
timestamp 1597059762
transform -1 0 6472 0 1 1810
box -4 -6 52 206
use NOR2X1  _2313_
timestamp 1597059762
transform 1 0 6472 0 1 1810
box -4 -6 52 206
use AND2X2  _2293_
timestamp 1597059762
transform 1 0 6520 0 1 1810
box -4 -6 68 206
use OR2X2  _2277_
timestamp 1597059762
transform 1 0 6584 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert91
timestamp 1597059762
transform 1 0 6648 0 1 1810
box -4 -6 52 206
use NAND2X1  _2966_
timestamp 1597059762
transform -1 0 6744 0 1 1810
box -4 -6 52 206
use AOI22X1  _2964_
timestamp 1597059762
transform -1 0 6888 0 1 1810
box -4 -6 84 206
use FILL  SFILL67440x18100
timestamp 1597059762
transform 1 0 6744 0 1 1810
box -4 -6 20 206
use FILL  SFILL67600x18100
timestamp 1597059762
transform 1 0 6760 0 1 1810
box -4 -6 20 206
use FILL  SFILL67760x18100
timestamp 1597059762
transform 1 0 6776 0 1 1810
box -4 -6 20 206
use FILL  SFILL67920x18100
timestamp 1597059762
transform 1 0 6792 0 1 1810
box -4 -6 20 206
use OAI21X1  _2755_
timestamp 1597059762
transform 1 0 6888 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert176
timestamp 1597059762
transform 1 0 6952 0 1 1810
box -4 -6 52 206
use AOI22X1  _2965_
timestamp 1597059762
transform 1 0 7000 0 1 1810
box -4 -6 84 206
use XOR2X1  _2109_
timestamp 1597059762
transform 1 0 7080 0 1 1810
box -4 -6 116 206
use AOI21X1  _2110_
timestamp 1597059762
transform 1 0 7192 0 1 1810
box -4 -6 68 206
use NOR2X1  _2108_
timestamp 1597059762
transform -1 0 7304 0 1 1810
box -4 -6 52 206
use NOR2X1  _2107_
timestamp 1597059762
transform -1 0 7352 0 1 1810
box -4 -6 52 206
use AND2X2  _2112_
timestamp 1597059762
transform -1 0 7416 0 1 1810
box -4 -6 68 206
use NOR2X1  _2111_
timestamp 1597059762
transform 1 0 7416 0 1 1810
box -4 -6 52 206
use INVX1  _2828_
timestamp 1597059762
transform -1 0 7496 0 1 1810
box -4 -6 36 206
use AND2X2  _2106_
timestamp 1597059762
transform 1 0 7496 0 1 1810
box -4 -6 68 206
use INVX1  _3524_
timestamp 1597059762
transform 1 0 8 0 -1 2210
box -4 -6 36 206
use NOR2X1  _3612_
timestamp 1597059762
transform 1 0 40 0 -1 2210
box -4 -6 52 206
use NOR2X1  _3525_
timestamp 1597059762
transform -1 0 136 0 -1 2210
box -4 -6 52 206
use INVX1  _3523_
timestamp 1597059762
transform -1 0 168 0 -1 2210
box -4 -6 36 206
use NOR2X1  _3679_
timestamp 1597059762
transform -1 0 216 0 -1 2210
box -4 -6 52 206
use AND2X2  _3713_
timestamp 1597059762
transform -1 0 280 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3680_
timestamp 1597059762
transform 1 0 280 0 -1 2210
box -4 -6 52 206
use AND2X2  _3646_
timestamp 1597059762
transform 1 0 328 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3613_
timestamp 1597059762
transform 1 0 392 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3529_
timestamp 1597059762
transform -1 0 488 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3579_
timestamp 1597059762
transform 1 0 488 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3530_
timestamp 1597059762
transform -1 0 584 0 -1 2210
box -4 -6 52 206
use OAI21X1  _3603_
timestamp 1597059762
transform 1 0 584 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3602_
timestamp 1597059762
transform -1 0 696 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert8
timestamp 1597059762
transform 1 0 696 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert13
timestamp 1597059762
transform 1 0 808 0 -1 2210
box -4 -6 52 206
use FILL  SFILL7440x20100
timestamp 1597059762
transform -1 0 760 0 -1 2210
box -4 -6 20 206
use FILL  SFILL7600x20100
timestamp 1597059762
transform -1 0 776 0 -1 2210
box -4 -6 20 206
use FILL  SFILL7760x20100
timestamp 1597059762
transform -1 0 792 0 -1 2210
box -4 -6 20 206
use FILL  SFILL7920x20100
timestamp 1597059762
transform -1 0 808 0 -1 2210
box -4 -6 20 206
use MUX2X1  _3780_
timestamp 1597059762
transform 1 0 856 0 -1 2210
box -4 -6 100 206
use OAI22X1  _3779_
timestamp 1597059762
transform -1 0 1032 0 -1 2210
box -4 -6 84 206
use OAI21X1  _3778_
timestamp 1597059762
transform -1 0 1096 0 -1 2210
box -4 -6 68 206
use NOR2X1  _3718_
timestamp 1597059762
transform 1 0 1096 0 -1 2210
box -4 -6 52 206
use AOI21X1  _3719_
timestamp 1597059762
transform -1 0 1208 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4221_
timestamp 1597059762
transform 1 0 1208 0 -1 2210
box -4 -6 196 206
use OAI21X1  _3990_
timestamp 1597059762
transform 1 0 1400 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4173_
timestamp 1597059762
transform -1 0 1656 0 -1 2210
box -4 -6 196 206
use OAI21X1  _3537_
timestamp 1597059762
transform -1 0 1720 0 -1 2210
box -4 -6 68 206
use OAI21X1  _3538_
timestamp 1597059762
transform -1 0 1784 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert207
timestamp 1597059762
transform -1 0 1832 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert228
timestamp 1597059762
transform 1 0 1832 0 -1 2210
box -4 -6 52 206
use OAI21X1  _3543_
timestamp 1597059762
transform 1 0 1880 0 -1 2210
box -4 -6 68 206
use OAI21X1  _3544_
timestamp 1597059762
transform -1 0 2008 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4175_
timestamp 1597059762
transform -1 0 2200 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_insert85
timestamp 1597059762
transform -1 0 2248 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4246_
timestamp 1597059762
transform 1 0 2312 0 -1 2210
box -4 -6 196 206
use FILL  SFILL22480x20100
timestamp 1597059762
transform -1 0 2264 0 -1 2210
box -4 -6 20 206
use FILL  SFILL22640x20100
timestamp 1597059762
transform -1 0 2280 0 -1 2210
box -4 -6 20 206
use FILL  SFILL22800x20100
timestamp 1597059762
transform -1 0 2296 0 -1 2210
box -4 -6 20 206
use FILL  SFILL22960x20100
timestamp 1597059762
transform -1 0 2312 0 -1 2210
box -4 -6 20 206
use NAND2X1  _3636_
timestamp 1597059762
transform 1 0 2504 0 -1 2210
box -4 -6 52 206
use OAI21X1  _3637_
timestamp 1597059762
transform -1 0 2616 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert124
timestamp 1597059762
transform -1 0 2664 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert109
timestamp 1597059762
transform 1 0 2664 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert226
timestamp 1597059762
transform 1 0 2712 0 -1 2210
box -4 -6 52 206
use OAI21X1  _3549_
timestamp 1597059762
transform 1 0 2760 0 -1 2210
box -4 -6 68 206
use OAI21X1  _3550_
timestamp 1597059762
transform -1 0 2888 0 -1 2210
box -4 -6 68 206
use NOR2X1  _3669_
timestamp 1597059762
transform 1 0 2888 0 -1 2210
box -4 -6 52 206
use AOI21X1  _3670_
timestamp 1597059762
transform 1 0 2936 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert15
timestamp 1597059762
transform -1 0 3048 0 -1 2210
box -4 -6 52 206
use AOI21X1  _3648_
timestamp 1597059762
transform 1 0 3048 0 -1 2210
box -4 -6 68 206
use NOR2X1  _3647_
timestamp 1597059762
transform -1 0 3160 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4251_
timestamp 1597059762
transform 1 0 3160 0 -1 2210
box -4 -6 196 206
use AOI21X1  _4049_
timestamp 1597059762
transform 1 0 3352 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4322_
timestamp 1597059762
transform 1 0 3416 0 -1 2210
box -4 -6 196 206
use OAI21X1  _4048_
timestamp 1597059762
transform -1 0 3672 0 -1 2210
box -4 -6 68 206
use AOI21X1  _3782_
timestamp 1597059762
transform 1 0 3672 0 -1 2210
box -4 -6 68 206
use OAI21X1  _3781_
timestamp 1597059762
transform -1 0 3864 0 -1 2210
box -4 -6 68 206
use FILL  SFILL37360x20100
timestamp 1597059762
transform -1 0 3752 0 -1 2210
box -4 -6 20 206
use FILL  SFILL37520x20100
timestamp 1597059762
transform -1 0 3768 0 -1 2210
box -4 -6 20 206
use FILL  SFILL37680x20100
timestamp 1597059762
transform -1 0 3784 0 -1 2210
box -4 -6 20 206
use FILL  SFILL37840x20100
timestamp 1597059762
transform -1 0 3800 0 -1 2210
box -4 -6 20 206
use DFFPOSX1  _4302_
timestamp 1597059762
transform 1 0 3864 0 -1 2210
box -4 -6 196 206
use INVX1  _3401_
timestamp 1597059762
transform -1 0 4088 0 -1 2210
box -4 -6 36 206
use DFFPOSX1  _4304_
timestamp 1597059762
transform 1 0 4088 0 -1 2210
box -4 -6 196 206
use DFFPOSX1  _4317_
timestamp 1597059762
transform 1 0 4280 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_insert61
timestamp 1597059762
transform -1 0 4520 0 -1 2210
box -4 -6 52 206
use NOR2X1  _2953_
timestamp 1597059762
transform 1 0 4520 0 -1 2210
box -4 -6 52 206
use INVX1  _2948_
timestamp 1597059762
transform 1 0 4568 0 -1 2210
box -4 -6 36 206
use OAI22X1  _2949_
timestamp 1597059762
transform -1 0 4680 0 -1 2210
box -4 -6 84 206
use INVX1  _2402_
timestamp 1597059762
transform -1 0 4712 0 -1 2210
box -4 -6 36 206
use INVX1  _2947_
timestamp 1597059762
transform -1 0 4744 0 -1 2210
box -4 -6 36 206
use NOR2X1  _2232_
timestamp 1597059762
transform 1 0 4744 0 -1 2210
box -4 -6 52 206
use NOR2X1  _2234_
timestamp 1597059762
transform 1 0 4792 0 -1 2210
box -4 -6 52 206
use AND2X2  _2233_
timestamp 1597059762
transform 1 0 4840 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert174
timestamp 1597059762
transform -1 0 4952 0 -1 2210
box -4 -6 52 206
use INVX1  _2969_
timestamp 1597059762
transform 1 0 4952 0 -1 2210
box -4 -6 36 206
use OR2X2  _2396_
timestamp 1597059762
transform 1 0 4984 0 -1 2210
box -4 -6 68 206
use NAND2X1  _2397_
timestamp 1597059762
transform -1 0 5096 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2395_
timestamp 1597059762
transform -1 0 5144 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2955_
timestamp 1597059762
transform -1 0 5192 0 -1 2210
box -4 -6 52 206
use INVX1  _3310_
timestamp 1597059762
transform -1 0 5224 0 -1 2210
box -4 -6 36 206
use XNOR2X1  _2398_
timestamp 1597059762
transform -1 0 5400 0 -1 2210
box -4 -6 116 206
use NAND2X1  _2407_
timestamp 1597059762
transform 1 0 5400 0 -1 2210
box -4 -6 52 206
use FILL  SFILL52240x20100
timestamp 1597059762
transform -1 0 5240 0 -1 2210
box -4 -6 20 206
use FILL  SFILL52400x20100
timestamp 1597059762
transform -1 0 5256 0 -1 2210
box -4 -6 20 206
use FILL  SFILL52560x20100
timestamp 1597059762
transform -1 0 5272 0 -1 2210
box -4 -6 20 206
use FILL  SFILL52720x20100
timestamp 1597059762
transform -1 0 5288 0 -1 2210
box -4 -6 20 206
use OAI21X1  _2412_
timestamp 1597059762
transform 1 0 5448 0 -1 2210
box -4 -6 68 206
use INVX1  _2928_
timestamp 1597059762
transform 1 0 5512 0 -1 2210
box -4 -6 36 206
use OAI21X1  _2930_
timestamp 1597059762
transform 1 0 5544 0 -1 2210
box -4 -6 68 206
use NAND2X1  _2929_
timestamp 1597059762
transform -1 0 5656 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3127_
timestamp 1597059762
transform -1 0 5704 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2936_
timestamp 1597059762
transform 1 0 5704 0 -1 2210
box -4 -6 52 206
use OAI21X1  _2937_
timestamp 1597059762
transform -1 0 5816 0 -1 2210
box -4 -6 68 206
use INVX1  _2935_
timestamp 1597059762
transform -1 0 5848 0 -1 2210
box -4 -6 36 206
use NAND2X1  _2374_
timestamp 1597059762
transform -1 0 5896 0 -1 2210
box -4 -6 52 206
use XNOR2X1  _2405_
timestamp 1597059762
transform -1 0 6008 0 -1 2210
box -4 -6 116 206
use AND2X2  _2314_
timestamp 1597059762
transform 1 0 6008 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert59
timestamp 1597059762
transform 1 0 6072 0 -1 2210
box -4 -6 52 206
use XNOR2X1  _2372_
timestamp 1597059762
transform 1 0 6120 0 -1 2210
box -4 -6 116 206
use NAND2X1  _2373_
timestamp 1597059762
transform -1 0 6280 0 -1 2210
box -4 -6 52 206
use INVX1  _2639_
timestamp 1597059762
transform 1 0 6280 0 -1 2210
box -4 -6 36 206
use OAI22X1  _2640_
timestamp 1597059762
transform -1 0 6392 0 -1 2210
box -4 -6 84 206
use INVX1  _2638_
timestamp 1597059762
transform -1 0 6424 0 -1 2210
box -4 -6 36 206
use NAND2X1  _2728_
timestamp 1597059762
transform -1 0 6472 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert60
timestamp 1597059762
transform 1 0 6472 0 -1 2210
box -4 -6 52 206
use OAI21X1  _2665_
timestamp 1597059762
transform -1 0 6584 0 -1 2210
box -4 -6 68 206
use INVX1  _2738_
timestamp 1597059762
transform 1 0 6584 0 -1 2210
box -4 -6 36 206
use NAND2X1  _2739_
timestamp 1597059762
transform -1 0 6664 0 -1 2210
box -4 -6 52 206
use NOR2X1  _2740_
timestamp 1597059762
transform -1 0 6712 0 -1 2210
box -4 -6 52 206
use OAI21X1  _2743_
timestamp 1597059762
transform -1 0 6776 0 -1 2210
box -4 -6 68 206
use FILL  SFILL67760x20100
timestamp 1597059762
transform -1 0 6792 0 -1 2210
box -4 -6 20 206
use FILL  SFILL67920x20100
timestamp 1597059762
transform -1 0 6808 0 -1 2210
box -4 -6 20 206
use FILL  SFILL68080x20100
timestamp 1597059762
transform -1 0 6824 0 -1 2210
box -4 -6 20 206
use FILL  SFILL68240x20100
timestamp 1597059762
transform -1 0 6840 0 -1 2210
box -4 -6 20 206
use NAND2X1  _2742_
timestamp 1597059762
transform 1 0 6840 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert175
timestamp 1597059762
transform -1 0 6936 0 -1 2210
box -4 -6 52 206
use INVX1  _2741_
timestamp 1597059762
transform -1 0 6968 0 -1 2210
box -4 -6 36 206
use NOR2X1  _2536_
timestamp 1597059762
transform 1 0 6968 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert58
timestamp 1597059762
transform 1 0 7016 0 -1 2210
box -4 -6 52 206
use INVX1  _2530_
timestamp 1597059762
transform 1 0 7064 0 -1 2210
box -4 -6 36 206
use INVX1  _2534_
timestamp 1597059762
transform 1 0 7096 0 -1 2210
box -4 -6 36 206
use AOI21X1  _2537_
timestamp 1597059762
transform 1 0 7128 0 -1 2210
box -4 -6 68 206
use NOR2X1  _2535_
timestamp 1597059762
transform 1 0 7192 0 -1 2210
box -4 -6 52 206
use INVX1  _2831_
timestamp 1597059762
transform 1 0 7240 0 -1 2210
box -4 -6 36 206
use NOR2X1  _2832_
timestamp 1597059762
transform -1 0 7320 0 -1 2210
box -4 -6 52 206
use AOI21X1  _2833_
timestamp 1597059762
transform 1 0 7320 0 -1 2210
box -4 -6 68 206
use NAND2X1  _2830_
timestamp 1597059762
transform -1 0 7432 0 -1 2210
box -4 -6 52 206
use XNOR2X1  _2821_
timestamp 1597059762
transform -1 0 7544 0 -1 2210
box -4 -6 116 206
use FILL  FILL72240x20100
timestamp 1597059762
transform -1 0 7560 0 -1 2210
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert27
timestamp 1597059762
transform 1 0 8 0 1 2210
box -4 -6 148 206
use NOR2X1  _3926_
timestamp 1597059762
transform -1 0 200 0 1 2210
box -4 -6 52 206
use AND2X2  _4138_
timestamp 1597059762
transform -1 0 264 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert232
timestamp 1597059762
transform -1 0 312 0 1 2210
box -4 -6 52 206
use AND2X2  _3927_
timestamp 1597059762
transform 1 0 312 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert36
timestamp 1597059762
transform 1 0 376 0 1 2210
box -4 -6 52 206
use INVX1  _3526_
timestamp 1597059762
transform 1 0 424 0 1 2210
box -4 -6 36 206
use NOR2X1  _3528_
timestamp 1597059762
transform 1 0 456 0 1 2210
box -4 -6 52 206
use NOR2X1  _3578_
timestamp 1597059762
transform -1 0 552 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _4214_
timestamp 1597059762
transform 1 0 552 0 1 2210
box -4 -6 196 206
use OAI21X1  _3704_
timestamp 1597059762
transform 1 0 808 0 1 2210
box -4 -6 68 206
use FILL  SFILL7440x22100
timestamp 1597059762
transform 1 0 744 0 1 2210
box -4 -6 20 206
use FILL  SFILL7600x22100
timestamp 1597059762
transform 1 0 760 0 1 2210
box -4 -6 20 206
use FILL  SFILL7760x22100
timestamp 1597059762
transform 1 0 776 0 1 2210
box -4 -6 20 206
use FILL  SFILL7920x22100
timestamp 1597059762
transform 1 0 792 0 1 2210
box -4 -6 20 206
use DFFPOSX1  _4198_
timestamp 1597059762
transform 1 0 872 0 1 2210
box -4 -6 196 206
use BUFX2  BUFX2_insert69
timestamp 1597059762
transform -1 0 1112 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _4182_
timestamp 1597059762
transform 1 0 1112 0 1 2210
box -4 -6 196 206
use OAI21X1  _3565_
timestamp 1597059762
transform 1 0 1304 0 1 2210
box -4 -6 68 206
use OAI21X1  _3564_
timestamp 1597059762
transform -1 0 1432 0 1 2210
box -4 -6 68 206
use INVX4  _3560_
timestamp 1597059762
transform -1 0 1480 0 1 2210
box -4 -6 52 206
use OAI21X1  _3873_
timestamp 1597059762
transform 1 0 1480 0 1 2210
box -4 -6 68 206
use OAI22X1  _3874_
timestamp 1597059762
transform -1 0 1624 0 1 2210
box -4 -6 84 206
use NOR2X1  _3872_
timestamp 1597059762
transform 1 0 1624 0 1 2210
box -4 -6 52 206
use NOR2X1  _4084_
timestamp 1597059762
transform 1 0 1672 0 1 2210
box -4 -6 52 206
use OAI21X1  _4085_
timestamp 1597059762
transform 1 0 1720 0 1 2210
box -4 -6 68 206
use OAI22X1  _4086_
timestamp 1597059762
transform 1 0 1784 0 1 2210
box -4 -6 84 206
use MUX2X1  _4091_
timestamp 1597059762
transform 1 0 1864 0 1 2210
box -4 -6 100 206
use BUFX2  BUFX2_insert199
timestamp 1597059762
transform -1 0 2008 0 1 2210
box -4 -6 52 206
use INVX8  _3748_
timestamp 1597059762
transform 1 0 2008 0 1 2210
box -4 -6 84 206
use MUX2X1  _3871_
timestamp 1597059762
transform -1 0 2184 0 1 2210
box -4 -6 100 206
use MUX2X1  _4083_
timestamp 1597059762
transform -1 0 2280 0 1 2210
box -4 -6 100 206
use INVX4  _3569_
timestamp 1597059762
transform -1 0 2392 0 1 2210
box -4 -6 52 206
use NAND2X1  _3586_
timestamp 1597059762
transform 1 0 2392 0 1 2210
box -4 -6 52 206
use FILL  SFILL22800x22100
timestamp 1597059762
transform 1 0 2280 0 1 2210
box -4 -6 20 206
use FILL  SFILL22960x22100
timestamp 1597059762
transform 1 0 2296 0 1 2210
box -4 -6 20 206
use FILL  SFILL23120x22100
timestamp 1597059762
transform 1 0 2312 0 1 2210
box -4 -6 20 206
use FILL  SFILL23280x22100
timestamp 1597059762
transform 1 0 2328 0 1 2210
box -4 -6 20 206
use OAI21X1  _3587_
timestamp 1597059762
transform -1 0 2504 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4206_
timestamp 1597059762
transform -1 0 2696 0 1 2210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert26
timestamp 1597059762
transform -1 0 2840 0 1 2210
box -4 -6 148 206
use DFFPOSX1  _4262_
timestamp 1597059762
transform -1 0 3032 0 1 2210
box -4 -6 196 206
use DFFPOSX1  _4240_
timestamp 1597059762
transform 1 0 3032 0 1 2210
box -4 -6 196 206
use AOI21X1  _3837_
timestamp 1597059762
transform 1 0 3224 0 1 2210
box -4 -6 68 206
use OAI21X1  _3836_
timestamp 1597059762
transform 1 0 3288 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert272
timestamp 1597059762
transform -1 0 3400 0 1 2210
box -4 -6 52 206
use AOI21X1  _3793_
timestamp 1597059762
transform 1 0 3400 0 1 2210
box -4 -6 68 206
use OAI21X1  _3792_
timestamp 1597059762
transform -1 0 3528 0 1 2210
box -4 -6 68 206
use AOI21X1  _4005_
timestamp 1597059762
transform 1 0 3528 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert101
timestamp 1597059762
transform 1 0 3592 0 1 2210
box -4 -6 52 206
use OAI21X1  _4004_
timestamp 1597059762
transform -1 0 3704 0 1 2210
box -4 -6 68 206
use AOI21X1  _4027_
timestamp 1597059762
transform 1 0 3704 0 1 2210
box -4 -6 68 206
use FILL  SFILL37680x22100
timestamp 1597059762
transform 1 0 3768 0 1 2210
box -4 -6 20 206
use FILL  SFILL37840x22100
timestamp 1597059762
transform 1 0 3784 0 1 2210
box -4 -6 20 206
use FILL  SFILL38000x22100
timestamp 1597059762
transform 1 0 3800 0 1 2210
box -4 -6 20 206
use FILL  SFILL38160x22100
timestamp 1597059762
transform 1 0 3816 0 1 2210
box -4 -6 20 206
use OAI21X1  _4026_
timestamp 1597059762
transform -1 0 3896 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4318_
timestamp 1597059762
transform 1 0 3896 0 1 2210
box -4 -6 196 206
use BUFX2  BUFX2_insert238
timestamp 1597059762
transform -1 0 4136 0 1 2210
box -4 -6 52 206
use NAND2X1  _3244_
timestamp 1597059762
transform 1 0 4136 0 1 2210
box -4 -6 52 206
use INVX1  _2950_
timestamp 1597059762
transform 1 0 4184 0 1 2210
box -4 -6 36 206
use OAI21X1  _2952_
timestamp 1597059762
transform 1 0 4216 0 1 2210
box -4 -6 68 206
use NAND2X1  _2951_
timestamp 1597059762
transform -1 0 4328 0 1 2210
box -4 -6 52 206
use AND2X2  _2236_
timestamp 1597059762
transform 1 0 4328 0 1 2210
box -4 -6 68 206
use NOR2X1  _2237_
timestamp 1597059762
transform -1 0 4440 0 1 2210
box -4 -6 52 206
use NOR2X1  _2235_
timestamp 1597059762
transform 1 0 4440 0 1 2210
box -4 -6 52 206
use NAND2X1  _2409_
timestamp 1597059762
transform 1 0 4488 0 1 2210
box -4 -6 52 206
use NOR2X1  _2410_
timestamp 1597059762
transform 1 0 4536 0 1 2210
box -4 -6 52 206
use INVX1  _2408_
timestamp 1597059762
transform -1 0 4616 0 1 2210
box -4 -6 36 206
use AOI21X1  _2411_
timestamp 1597059762
transform -1 0 4680 0 1 2210
box -4 -6 68 206
use NOR2X1  _2403_
timestamp 1597059762
transform -1 0 4728 0 1 2210
box -4 -6 52 206
use AOI21X1  _2404_
timestamp 1597059762
transform -1 0 4792 0 1 2210
box -4 -6 68 206
use XNOR2X1  _2406_
timestamp 1597059762
transform 1 0 4792 0 1 2210
box -4 -6 116 206
use NAND2X1  _2977_
timestamp 1597059762
transform 1 0 4904 0 1 2210
box -4 -6 52 206
use NAND3X1  _2488_
timestamp 1597059762
transform -1 0 5016 0 1 2210
box -4 -6 68 206
use AOI21X1  _2492_
timestamp 1597059762
transform 1 0 5016 0 1 2210
box -4 -6 68 206
use INVX1  _2932_
timestamp 1597059762
transform 1 0 5080 0 1 2210
box -4 -6 36 206
use OAI21X1  _2934_
timestamp 1597059762
transform 1 0 5112 0 1 2210
box -4 -6 68 206
use NOR2X1  _2938_
timestamp 1597059762
transform -1 0 5224 0 1 2210
box -4 -6 52 206
use OAI21X1  _2494_
timestamp 1597059762
transform 1 0 5224 0 1 2210
box -4 -6 68 206
use OR2X2  _2375_
timestamp 1597059762
transform 1 0 5352 0 1 2210
box -4 -6 68 206
use NAND3X1  _2946_
timestamp 1597059762
transform 1 0 5416 0 1 2210
box -4 -6 68 206
use FILL  SFILL52880x22100
timestamp 1597059762
transform 1 0 5288 0 1 2210
box -4 -6 20 206
use FILL  SFILL53040x22100
timestamp 1597059762
transform 1 0 5304 0 1 2210
box -4 -6 20 206
use FILL  SFILL53200x22100
timestamp 1597059762
transform 1 0 5320 0 1 2210
box -4 -6 20 206
use FILL  SFILL53360x22100
timestamp 1597059762
transform 1 0 5336 0 1 2210
box -4 -6 20 206
use NOR2X1  _2931_
timestamp 1597059762
transform 1 0 5480 0 1 2210
box -4 -6 52 206
use AOI22X1  _2378_
timestamp 1597059762
transform 1 0 5528 0 1 2210
box -4 -6 84 206
use OR2X2  _2377_
timestamp 1597059762
transform -1 0 5672 0 1 2210
box -4 -6 68 206
use NAND2X1  _2376_
timestamp 1597059762
transform -1 0 5720 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert93
timestamp 1597059762
transform -1 0 5768 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert240
timestamp 1597059762
transform -1 0 5816 0 1 2210
box -4 -6 52 206
use INVX1  _2641_
timestamp 1597059762
transform 1 0 5816 0 1 2210
box -4 -6 36 206
use OAI22X1  _2643_
timestamp 1597059762
transform 1 0 5848 0 1 2210
box -4 -6 84 206
use INVX1  _2642_
timestamp 1597059762
transform -1 0 5960 0 1 2210
box -4 -6 36 206
use NOR2X1  _2644_
timestamp 1597059762
transform -1 0 6008 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert92
timestamp 1597059762
transform 1 0 6008 0 1 2210
box -4 -6 52 206
use NAND2X1  _2654_
timestamp 1597059762
transform 1 0 6056 0 1 2210
box -4 -6 52 206
use AOI22X1  _2656_
timestamp 1597059762
transform 1 0 6104 0 1 2210
box -4 -6 84 206
use BUFX2  BUFX2_insert236
timestamp 1597059762
transform 1 0 6184 0 1 2210
box -4 -6 52 206
use OR2X2  _2727_
timestamp 1597059762
transform 1 0 6232 0 1 2210
box -4 -6 68 206
use AOI22X1  _2731_
timestamp 1597059762
transform 1 0 6296 0 1 2210
box -4 -6 84 206
use OR2X2  _2729_
timestamp 1597059762
transform -1 0 6440 0 1 2210
box -4 -6 68 206
use NAND2X1  _2730_
timestamp 1597059762
transform -1 0 6488 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert239
timestamp 1597059762
transform 1 0 6488 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert237
timestamp 1597059762
transform 1 0 6536 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert94
timestamp 1597059762
transform 1 0 6584 0 1 2210
box -4 -6 52 206
use NAND2X1  _2532_
timestamp 1597059762
transform 1 0 6632 0 1 2210
box -4 -6 52 206
use OR2X2  _2531_
timestamp 1597059762
transform 1 0 6680 0 1 2210
box -4 -6 68 206
use NAND3X1  _2533_
timestamp 1597059762
transform -1 0 6872 0 1 2210
box -4 -6 68 206
use FILL  SFILL67440x22100
timestamp 1597059762
transform 1 0 6744 0 1 2210
box -4 -6 20 206
use FILL  SFILL67600x22100
timestamp 1597059762
transform 1 0 6760 0 1 2210
box -4 -6 20 206
use FILL  SFILL67760x22100
timestamp 1597059762
transform 1 0 6776 0 1 2210
box -4 -6 20 206
use FILL  SFILL67920x22100
timestamp 1597059762
transform 1 0 6792 0 1 2210
box -4 -6 20 206
use AOI21X1  _2744_
timestamp 1597059762
transform -1 0 6936 0 1 2210
box -4 -6 68 206
use XNOR2X1  _2529_
timestamp 1597059762
transform -1 0 7048 0 1 2210
box -4 -6 116 206
use AOI21X1  _2845_
timestamp 1597059762
transform -1 0 7112 0 1 2210
box -4 -6 68 206
use NAND3X1  _2868_
timestamp 1597059762
transform -1 0 7176 0 1 2210
box -4 -6 68 206
use INVX1  _2864_
timestamp 1597059762
transform -1 0 7208 0 1 2210
box -4 -6 36 206
use OAI21X1  _2834_
timestamp 1597059762
transform -1 0 7272 0 1 2210
box -4 -6 68 206
use NAND2X1  _2822_
timestamp 1597059762
transform -1 0 7320 0 1 2210
box -4 -6 52 206
use XNOR2X1  _2820_
timestamp 1597059762
transform -1 0 7432 0 1 2210
box -4 -6 116 206
use BUFX2  _2035_
timestamp 1597059762
transform 1 0 7432 0 1 2210
box -4 -6 52 206
use NOR2X1  _2100_
timestamp 1597059762
transform 1 0 7480 0 1 2210
box -4 -6 52 206
use INVX1  _2823_
timestamp 1597059762
transform -1 0 7560 0 1 2210
box -4 -6 36 206
use DFFPOSX1  _4294_
timestamp 1597059762
transform -1 0 200 0 -1 2610
box -4 -6 196 206
use AOI21X1  _3951_
timestamp 1597059762
transform -1 0 264 0 -1 2610
box -4 -6 68 206
use AOI21X1  _4162_
timestamp 1597059762
transform 1 0 264 0 -1 2610
box -4 -6 68 206
use NOR2X1  _4161_
timestamp 1597059762
transform -1 0 376 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _4222_
timestamp 1597059762
transform 1 0 376 0 -1 2610
box -4 -6 196 206
use AOI21X1  _3737_
timestamp 1597059762
transform 1 0 568 0 -1 2610
box -4 -6 68 206
use NOR2X1  _3736_
timestamp 1597059762
transform -1 0 680 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _4226_
timestamp 1597059762
transform 1 0 744 0 -1 2610
box -4 -6 196 206
use FILL  SFILL6800x24100
timestamp 1597059762
transform -1 0 696 0 -1 2610
box -4 -6 20 206
use FILL  SFILL6960x24100
timestamp 1597059762
transform -1 0 712 0 -1 2610
box -4 -6 20 206
use FILL  SFILL7120x24100
timestamp 1597059762
transform -1 0 728 0 -1 2610
box -4 -6 20 206
use FILL  SFILL7280x24100
timestamp 1597059762
transform -1 0 744 0 -1 2610
box -4 -6 20 206
use NOR2X1  _3728_
timestamp 1597059762
transform 1 0 936 0 -1 2610
box -4 -6 52 206
use AOI21X1  _3729_
timestamp 1597059762
transform -1 0 1048 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3553_
timestamp 1597059762
transform 1 0 1048 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3552_
timestamp 1597059762
transform 1 0 1112 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4178_
timestamp 1597059762
transform 1 0 1176 0 -1 2610
box -4 -6 196 206
use OAI21X1  _3789_
timestamp 1597059762
transform 1 0 1368 0 -1 2610
box -4 -6 68 206
use OAI22X1  _3790_
timestamp 1597059762
transform 1 0 1432 0 -1 2610
box -4 -6 84 206
use NOR2X1  _3788_
timestamp 1597059762
transform -1 0 1560 0 -1 2610
box -4 -6 52 206
use MUX2X1  _4047_
timestamp 1597059762
transform 1 0 1560 0 -1 2610
box -4 -6 100 206
use DFFPOSX1  _4194_
timestamp 1597059762
transform -1 0 1848 0 -1 2610
box -4 -6 196 206
use OAI21X1  _3696_
timestamp 1597059762
transform 1 0 1848 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3695_
timestamp 1597059762
transform 1 0 1912 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert209
timestamp 1597059762
transform -1 0 2008 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert235
timestamp 1597059762
transform -1 0 2056 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3687_
timestamp 1597059762
transform 1 0 2056 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3688_
timestamp 1597059762
transform -1 0 2168 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3682_
timestamp 1597059762
transform 1 0 2168 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3681_
timestamp 1597059762
transform -1 0 2344 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert6
timestamp 1597059762
transform 1 0 2344 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert82
timestamp 1597059762
transform 1 0 2392 0 -1 2610
box -4 -6 52 206
use FILL  SFILL22320x24100
timestamp 1597059762
transform -1 0 2248 0 -1 2610
box -4 -6 20 206
use FILL  SFILL22480x24100
timestamp 1597059762
transform -1 0 2264 0 -1 2610
box -4 -6 20 206
use FILL  SFILL22640x24100
timestamp 1597059762
transform -1 0 2280 0 -1 2610
box -4 -6 20 206
use FILL  SFILL22800x24100
timestamp 1597059762
transform -1 0 2296 0 -1 2610
box -4 -6 20 206
use OAI21X1  _3997_
timestamp 1597059762
transform 1 0 2440 0 -1 2610
box -4 -6 68 206
use MUX2X1  _4003_
timestamp 1597059762
transform -1 0 2600 0 -1 2610
box -4 -6 100 206
use MUX2X1  _3791_
timestamp 1597059762
transform -1 0 2696 0 -1 2610
box -4 -6 100 206
use OAI21X1  _3621_
timestamp 1597059762
transform 1 0 2696 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3620_
timestamp 1597059762
transform -1 0 2808 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _4238_
timestamp 1597059762
transform 1 0 2808 0 -1 2610
box -4 -6 196 206
use OAI21X1  _3581_
timestamp 1597059762
transform 1 0 3000 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3580_
timestamp 1597059762
transform -1 0 3112 0 -1 2610
box -4 -6 52 206
use INVX4  _3545_
timestamp 1597059762
transform -1 0 3160 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3625_
timestamp 1597059762
transform 1 0 3160 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3624_
timestamp 1597059762
transform -1 0 3272 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert104
timestamp 1597059762
transform -1 0 3320 0 -1 2610
box -4 -6 52 206
use INVX1  _3394_
timestamp 1597059762
transform -1 0 3352 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3615_
timestamp 1597059762
transform 1 0 3352 0 -1 2610
box -4 -6 68 206
use INVX1  _3366_
timestamp 1597059762
transform -1 0 3448 0 -1 2610
box -4 -6 36 206
use INVX1  _3297_
timestamp 1597059762
transform 1 0 3448 0 -1 2610
box -4 -6 36 206
use AOI21X1  _4093_
timestamp 1597059762
transform 1 0 3480 0 -1 2610
box -4 -6 68 206
use OAI21X1  _4092_
timestamp 1597059762
transform -1 0 3608 0 -1 2610
box -4 -6 68 206
use INVX1  _3380_
timestamp 1597059762
transform -1 0 3640 0 -1 2610
box -4 -6 36 206
use INVX1  _3387_
timestamp 1597059762
transform -1 0 3672 0 -1 2610
box -4 -6 36 206
use INVX1  _3373_
timestamp 1597059762
transform 1 0 3672 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  _4299_
timestamp 1597059762
transform 1 0 3768 0 -1 2610
box -4 -6 196 206
use FILL  SFILL37040x24100
timestamp 1597059762
transform -1 0 3720 0 -1 2610
box -4 -6 20 206
use FILL  SFILL37200x24100
timestamp 1597059762
transform -1 0 3736 0 -1 2610
box -4 -6 20 206
use FILL  SFILL37360x24100
timestamp 1597059762
transform -1 0 3752 0 -1 2610
box -4 -6 20 206
use FILL  SFILL37520x24100
timestamp 1597059762
transform -1 0 3768 0 -1 2610
box -4 -6 20 206
use INVX1  _3408_
timestamp 1597059762
transform -1 0 3992 0 -1 2610
box -4 -6 36 206
use BUFX2  BUFX2_insert111
timestamp 1597059762
transform 1 0 3992 0 -1 2610
box -4 -6 52 206
use INVX1  _3359_
timestamp 1597059762
transform -1 0 4072 0 -1 2610
box -4 -6 36 206
use AOI21X1  _3760_
timestamp 1597059762
transform 1 0 4072 0 -1 2610
box -4 -6 68 206
use OAI21X1  _3759_
timestamp 1597059762
transform -1 0 4200 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4315_
timestamp 1597059762
transform 1 0 4200 0 -1 2610
box -4 -6 196 206
use OAI21X1  _3245_
timestamp 1597059762
transform -1 0 4456 0 -1 2610
box -4 -6 68 206
use INVX1  _3243_
timestamp 1597059762
transform -1 0 4488 0 -1 2610
box -4 -6 36 206
use INVX1  _3082_
timestamp 1597059762
transform 1 0 4488 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3084_
timestamp 1597059762
transform 1 0 4520 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3083_
timestamp 1597059762
transform -1 0 4632 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert246
timestamp 1597059762
transform 1 0 4632 0 -1 2610
box -4 -6 52 206
use NOR2X1  _2226_
timestamp 1597059762
transform 1 0 4680 0 -1 2610
box -4 -6 52 206
use NOR2X1  _2228_
timestamp 1597059762
transform 1 0 4728 0 -1 2610
box -4 -6 52 206
use AND2X2  _2227_
timestamp 1597059762
transform -1 0 4840 0 -1 2610
box -4 -6 68 206
use INVX1  _2385_
timestamp 1597059762
transform 1 0 4840 0 -1 2610
box -4 -6 36 206
use NAND2X1  _2386_
timestamp 1597059762
transform 1 0 4872 0 -1 2610
box -4 -6 52 206
use AND2X2  _2399_
timestamp 1597059762
transform 1 0 4920 0 -1 2610
box -4 -6 68 206
use OAI21X1  _2401_
timestamp 1597059762
transform 1 0 4984 0 -1 2610
box -4 -6 68 206
use INVX1  _2387_
timestamp 1597059762
transform 1 0 5048 0 -1 2610
box -4 -6 36 206
use NAND2X1  _2388_
timestamp 1597059762
transform -1 0 5128 0 -1 2610
box -4 -6 52 206
use NOR2X1  _2393_
timestamp 1597059762
transform -1 0 5176 0 -1 2610
box -4 -6 52 206
use AOI21X1  _2394_
timestamp 1597059762
transform -1 0 5240 0 -1 2610
box -4 -6 68 206
use NAND2X1  _2391_
timestamp 1597059762
transform 1 0 5304 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3134_
timestamp 1597059762
transform 1 0 5352 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3135_
timestamp 1597059762
transform -1 0 5464 0 -1 2610
box -4 -6 68 206
use FILL  SFILL52400x24100
timestamp 1597059762
transform -1 0 5256 0 -1 2610
box -4 -6 20 206
use FILL  SFILL52560x24100
timestamp 1597059762
transform -1 0 5272 0 -1 2610
box -4 -6 20 206
use FILL  SFILL52720x24100
timestamp 1597059762
transform -1 0 5288 0 -1 2610
box -4 -6 20 206
use FILL  SFILL52880x24100
timestamp 1597059762
transform -1 0 5304 0 -1 2610
box -4 -6 20 206
use INVX1  _3133_
timestamp 1597059762
transform -1 0 5496 0 -1 2610
box -4 -6 36 206
use INVX1  _3126_
timestamp 1597059762
transform 1 0 5496 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3128_
timestamp 1597059762
transform 1 0 5528 0 -1 2610
box -4 -6 68 206
use INVX1  _2926_
timestamp 1597059762
transform 1 0 5592 0 -1 2610
box -4 -6 36 206
use OAI22X1  _2927_
timestamp 1597059762
transform -1 0 5704 0 -1 2610
box -4 -6 84 206
use INVX1  _2925_
timestamp 1597059762
transform -1 0 5736 0 -1 2610
box -4 -6 36 206
use NOR2X1  _2231_
timestamp 1597059762
transform -1 0 5784 0 -1 2610
box -4 -6 52 206
use NOR2X1  _2229_
timestamp 1597059762
transform -1 0 5832 0 -1 2610
box -4 -6 52 206
use XOR2X1  _2384_
timestamp 1597059762
transform 1 0 5832 0 -1 2610
box -4 -6 116 206
use INVX1  _2646_
timestamp 1597059762
transform 1 0 5944 0 -1 2610
box -4 -6 36 206
use OAI22X1  _2647_
timestamp 1597059762
transform 1 0 5976 0 -1 2610
box -4 -6 84 206
use INVX1  _2645_
timestamp 1597059762
transform -1 0 6088 0 -1 2610
box -4 -6 36 206
use NAND2X1  _2649_
timestamp 1597059762
transform -1 0 6136 0 -1 2610
box -4 -6 52 206
use OAI21X1  _2650_
timestamp 1597059762
transform -1 0 6200 0 -1 2610
box -4 -6 68 206
use INVX1  _2648_
timestamp 1597059762
transform -1 0 6232 0 -1 2610
box -4 -6 36 206
use OAI21X1  _2655_
timestamp 1597059762
transform 1 0 6232 0 -1 2610
box -4 -6 68 206
use NOR2X1  _2651_
timestamp 1597059762
transform 1 0 6296 0 -1 2610
box -4 -6 52 206
use AND2X2  _2652_
timestamp 1597059762
transform 1 0 6344 0 -1 2610
box -4 -6 68 206
use AOI22X1  _2939_
timestamp 1597059762
transform 1 0 6408 0 -1 2610
box -4 -6 84 206
use NAND2X1  _2941_
timestamp 1597059762
transform 1 0 6488 0 -1 2610
box -4 -6 52 206
use NOR2X1  _2945_
timestamp 1597059762
transform -1 0 6584 0 -1 2610
box -4 -6 52 206
use AOI22X1  _2942_
timestamp 1597059762
transform 1 0 6584 0 -1 2610
box -4 -6 84 206
use NAND2X1  _2944_
timestamp 1597059762
transform 1 0 6664 0 -1 2610
box -4 -6 52 206
use AOI22X1  _2943_
timestamp 1597059762
transform 1 0 6712 0 -1 2610
box -4 -6 84 206
use FILL  SFILL67920x24100
timestamp 1597059762
transform -1 0 6808 0 -1 2610
box -4 -6 20 206
use FILL  SFILL68080x24100
timestamp 1597059762
transform -1 0 6824 0 -1 2610
box -4 -6 20 206
use FILL  SFILL68240x24100
timestamp 1597059762
transform -1 0 6840 0 -1 2610
box -4 -6 20 206
use NOR3X1  _2784_
timestamp 1597059762
transform -1 0 6984 0 -1 2610
box -4 -6 132 206
use OAI21X1  _2781_
timestamp 1597059762
transform -1 0 7048 0 -1 2610
box -4 -6 68 206
use FILL  SFILL68400x24100
timestamp 1597059762
transform -1 0 6856 0 -1 2610
box -4 -6 20 206
use NOR2X1  _2736_
timestamp 1597059762
transform 1 0 7048 0 -1 2610
box -4 -6 52 206
use OAI21X1  _2737_
timestamp 1597059762
transform 1 0 7096 0 -1 2610
box -4 -6 68 206
use NAND2X1  _2733_
timestamp 1597059762
transform -1 0 7208 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert247
timestamp 1597059762
transform 1 0 7208 0 -1 2610
box -4 -6 52 206
use INVX1  _2865_
timestamp 1597059762
transform 1 0 7256 0 -1 2610
box -4 -6 36 206
use AOI21X1  _2867_
timestamp 1597059762
transform 1 0 7288 0 -1 2610
box -4 -6 68 206
use XNOR2X1  _2104_
timestamp 1597059762
transform 1 0 7352 0 -1 2610
box -4 -6 116 206
use OAI21X1  _2105_
timestamp 1597059762
transform 1 0 7464 0 -1 2610
box -4 -6 68 206
use FILL  FILL72080x24100
timestamp 1597059762
transform -1 0 7544 0 -1 2610
box -4 -6 20 206
use FILL  FILL72240x24100
timestamp 1597059762
transform -1 0 7560 0 -1 2610
box -4 -6 20 206
use DFFPOSX1  _4278_
timestamp 1597059762
transform -1 0 200 0 1 2610
box -4 -6 196 206
use NOR2X1  _3950_
timestamp 1597059762
transform 1 0 200 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert70
timestamp 1597059762
transform 1 0 248 0 1 2610
box -4 -6 52 206
use AOI21X1  _3721_
timestamp 1597059762
transform 1 0 296 0 1 2610
box -4 -6 68 206
use NOR2X1  _3720_
timestamp 1597059762
transform -1 0 408 0 1 2610
box -4 -6 52 206
use MUX2X1  _3875_
timestamp 1597059762
transform -1 0 504 0 1 2610
box -4 -6 100 206
use MUX2X1  _4087_
timestamp 1597059762
transform -1 0 600 0 1 2610
box -4 -6 100 206
use DFFPOSX1  _4230_
timestamp 1597059762
transform 1 0 600 0 1 2610
box -4 -6 196 206
use FILL  SFILL7920x26100
timestamp 1597059762
transform 1 0 792 0 1 2610
box -4 -6 20 206
use FILL  SFILL8080x26100
timestamp 1597059762
transform 1 0 808 0 1 2610
box -4 -6 20 206
use NAND2X1  _3703_
timestamp 1597059762
transform -1 0 904 0 1 2610
box -4 -6 52 206
use NOR2X1  _3876_
timestamp 1597059762
transform -1 0 952 0 1 2610
box -4 -6 52 206
use OAI21X1  _4089_
timestamp 1597059762
transform 1 0 952 0 1 2610
box -4 -6 68 206
use FILL  SFILL8240x26100
timestamp 1597059762
transform 1 0 824 0 1 2610
box -4 -6 20 206
use FILL  SFILL8400x26100
timestamp 1597059762
transform 1 0 840 0 1 2610
box -4 -6 20 206
use NOR2X1  _4088_
timestamp 1597059762
transform 1 0 1016 0 1 2610
box -4 -6 52 206
use OAI22X1  _4090_
timestamp 1597059762
transform 1 0 1064 0 1 2610
box -4 -6 84 206
use BUFX2  BUFX2_insert125
timestamp 1597059762
transform 1 0 1144 0 1 2610
box -4 -6 52 206
use OAI21X1  _4041_
timestamp 1597059762
transform 1 0 1192 0 1 2610
box -4 -6 68 206
use NOR2X1  _4040_
timestamp 1597059762
transform 1 0 1256 0 1 2610
box -4 -6 52 206
use OAI22X1  _4042_
timestamp 1597059762
transform 1 0 1304 0 1 2610
box -4 -6 84 206
use OAI21X1  _4001_
timestamp 1597059762
transform 1 0 1384 0 1 2610
box -4 -6 68 206
use NOR2X1  _3828_
timestamp 1597059762
transform 1 0 1448 0 1 2610
box -4 -6 52 206
use OAI22X1  _3830_
timestamp 1597059762
transform 1 0 1496 0 1 2610
box -4 -6 84 206
use OAI22X1  _4002_
timestamp 1597059762
transform 1 0 1576 0 1 2610
box -4 -6 84 206
use NOR2X1  _4000_
timestamp 1597059762
transform 1 0 1656 0 1 2610
box -4 -6 52 206
use OAI22X1  _4046_
timestamp 1597059762
transform -1 0 1784 0 1 2610
box -4 -6 84 206
use OAI21X1  _4045_
timestamp 1597059762
transform -1 0 1848 0 1 2610
box -4 -6 68 206
use NOR2X1  _4044_
timestamp 1597059762
transform 1 0 1848 0 1 2610
box -4 -6 52 206
use NOR2X1  _3832_
timestamp 1597059762
transform -1 0 1944 0 1 2610
box -4 -6 52 206
use OAI22X1  _3834_
timestamp 1597059762
transform -1 0 2024 0 1 2610
box -4 -6 84 206
use OAI21X1  _3833_
timestamp 1597059762
transform 1 0 2024 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert107
timestamp 1597059762
transform 1 0 2088 0 1 2610
box -4 -6 52 206
use MUX2X1  _3835_
timestamp 1597059762
transform 1 0 2136 0 1 2610
box -4 -6 100 206
use DFFPOSX1  _4190_
timestamp 1597059762
transform -1 0 2488 0 1 2610
box -4 -6 196 206
use FILL  SFILL22320x26100
timestamp 1597059762
transform 1 0 2232 0 1 2610
box -4 -6 20 206
use FILL  SFILL22480x26100
timestamp 1597059762
transform 1 0 2248 0 1 2610
box -4 -6 20 206
use FILL  SFILL22640x26100
timestamp 1597059762
transform 1 0 2264 0 1 2610
box -4 -6 20 206
use FILL  SFILL22800x26100
timestamp 1597059762
transform 1 0 2280 0 1 2610
box -4 -6 20 206
use DFFPOSX1  _4187_
timestamp 1597059762
transform 1 0 2488 0 1 2610
box -4 -6 196 206
use BUFX2  BUFX2_insert256
timestamp 1597059762
transform 1 0 2680 0 1 2610
box -4 -6 52 206
use OAI21X1  _3785_
timestamp 1597059762
transform 1 0 2728 0 1 2610
box -4 -6 68 206
use OAI22X1  _3786_
timestamp 1597059762
transform -1 0 2872 0 1 2610
box -4 -6 84 206
use OAI22X1  _3998_
timestamp 1597059762
transform 1 0 2872 0 1 2610
box -4 -6 84 206
use MUX2X1  _3995_
timestamp 1597059762
transform -1 0 3048 0 1 2610
box -4 -6 100 206
use MUX2X1  _3783_
timestamp 1597059762
transform -1 0 3144 0 1 2610
box -4 -6 100 206
use DFFPOSX1  _4254_
timestamp 1597059762
transform -1 0 3336 0 1 2610
box -4 -6 196 206
use NOR2X1  _3653_
timestamp 1597059762
transform 1 0 3336 0 1 2610
box -4 -6 52 206
use AOI21X1  _3654_
timestamp 1597059762
transform -1 0 3448 0 1 2610
box -4 -6 68 206
use NAND2X1  _3614_
timestamp 1597059762
transform -1 0 3496 0 1 2610
box -4 -6 52 206
use MUX2X1  _3747_
timestamp 1597059762
transform 1 0 3496 0 1 2610
box -4 -6 100 206
use MUX2X1  _3961_
timestamp 1597059762
transform 1 0 3592 0 1 2610
box -4 -6 100 206
use AOI21X1  _3972_
timestamp 1597059762
transform 1 0 3688 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4203_
timestamp 1597059762
transform 1 0 3816 0 1 2610
box -4 -6 196 206
use FILL  SFILL37520x26100
timestamp 1597059762
transform 1 0 3752 0 1 2610
box -4 -6 20 206
use FILL  SFILL37680x26100
timestamp 1597059762
transform 1 0 3768 0 1 2610
box -4 -6 20 206
use FILL  SFILL37840x26100
timestamp 1597059762
transform 1 0 3784 0 1 2610
box -4 -6 20 206
use FILL  SFILL38000x26100
timestamp 1597059762
transform 1 0 3800 0 1 2610
box -4 -6 20 206
use BUFX2  BUFX2_insert267
timestamp 1597059762
transform 1 0 4008 0 1 2610
box -4 -6 52 206
use OAI21X1  _3971_
timestamp 1597059762
transform -1 0 4120 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4235_
timestamp 1597059762
transform -1 0 4312 0 1 2610
box -4 -6 196 206
use OAI21X1  _3982_
timestamp 1597059762
transform -1 0 4376 0 1 2610
box -4 -6 68 206
use AOI21X1  _3983_
timestamp 1597059762
transform 1 0 4376 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4300_
timestamp 1597059762
transform 1 0 4440 0 1 2610
box -4 -6 196 206
use OAI21X1  _3216_
timestamp 1597059762
transform -1 0 4696 0 1 2610
box -4 -6 68 206
use INVX1  _3214_
timestamp 1597059762
transform -1 0 4728 0 1 2610
box -4 -6 36 206
use NOR2X1  _3246_
timestamp 1597059762
transform 1 0 4728 0 1 2610
box -4 -6 52 206
use NAND2X1  _3215_
timestamp 1597059762
transform -1 0 4824 0 1 2610
box -4 -6 52 206
use INVX1  _3240_
timestamp 1597059762
transform 1 0 4824 0 1 2610
box -4 -6 36 206
use OAI21X1  _3242_
timestamp 1597059762
transform -1 0 4920 0 1 2610
box -4 -6 68 206
use NOR2X1  _3085_
timestamp 1597059762
transform 1 0 4920 0 1 2610
box -4 -6 52 206
use NAND3X1  _3100_
timestamp 1597059762
transform 1 0 4968 0 1 2610
box -4 -6 68 206
use NOR2X1  _3092_
timestamp 1597059762
transform -1 0 5080 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert273
timestamp 1597059762
transform -1 0 5128 0 1 2610
box -4 -6 52 206
use NAND3X1  _2366_
timestamp 1597059762
transform 1 0 5128 0 1 2610
box -4 -6 68 206
use NAND2X1  _3090_
timestamp 1597059762
transform 1 0 5192 0 1 2610
box -4 -6 52 206
use OAI21X1  _3091_
timestamp 1597059762
transform -1 0 5368 0 1 2610
box -4 -6 68 206
use INVX1  _3089_
timestamp 1597059762
transform 1 0 5368 0 1 2610
box -4 -6 36 206
use NAND2X1  _3105_
timestamp 1597059762
transform 1 0 5400 0 1 2610
box -4 -6 52 206
use FILL  SFILL52400x26100
timestamp 1597059762
transform 1 0 5240 0 1 2610
box -4 -6 20 206
use FILL  SFILL52560x26100
timestamp 1597059762
transform 1 0 5256 0 1 2610
box -4 -6 20 206
use FILL  SFILL52720x26100
timestamp 1597059762
transform 1 0 5272 0 1 2610
box -4 -6 20 206
use FILL  SFILL52880x26100
timestamp 1597059762
transform 1 0 5288 0 1 2610
box -4 -6 20 206
use NAND2X1  _2390_
timestamp 1597059762
transform 1 0 5448 0 1 2610
box -4 -6 52 206
use NOR2X1  _2400_
timestamp 1597059762
transform 1 0 5496 0 1 2610
box -4 -6 52 206
use INVX1  _2871_
timestamp 1597059762
transform 1 0 5544 0 1 2610
box -4 -6 36 206
use INVX1  _2389_
timestamp 1597059762
transform -1 0 5608 0 1 2610
box -4 -6 36 206
use XNOR2X1  _2392_
timestamp 1597059762
transform -1 0 5720 0 1 2610
box -4 -6 116 206
use NAND2X1  _2933_
timestamp 1597059762
transform 1 0 5720 0 1 2610
box -4 -6 52 206
use NOR2X1  _3136_
timestamp 1597059762
transform 1 0 5768 0 1 2610
box -4 -6 52 206
use NAND3X1  _3144_
timestamp 1597059762
transform -1 0 5880 0 1 2610
box -4 -6 68 206
use NOR2X1  _3129_
timestamp 1597059762
transform 1 0 5880 0 1 2610
box -4 -6 52 206
use OAI22X1  _3125_
timestamp 1597059762
transform 1 0 5928 0 1 2610
box -4 -6 84 206
use NAND2X1  _2898_
timestamp 1597059762
transform 1 0 6008 0 1 2610
box -4 -6 52 206
use AND2X2  _2230_
timestamp 1597059762
transform 1 0 6056 0 1 2610
box -4 -6 68 206
use INVX1  _3124_
timestamp 1597059762
transform 1 0 6120 0 1 2610
box -4 -6 36 206
use BUFX2  BUFX2_insert114
timestamp 1597059762
transform -1 0 6200 0 1 2610
box -4 -6 52 206
use NOR2X1  _2339_
timestamp 1597059762
transform 1 0 6200 0 1 2610
box -4 -6 52 206
use NOR2X1  _2336_
timestamp 1597059762
transform -1 0 6296 0 1 2610
box -4 -6 52 206
use OAI22X1  _2338_
timestamp 1597059762
transform -1 0 6376 0 1 2610
box -4 -6 84 206
use NOR2X1  _2334_
timestamp 1597059762
transform 1 0 6376 0 1 2610
box -4 -6 52 206
use AND2X2  _2335_
timestamp 1597059762
transform -1 0 6488 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert245
timestamp 1597059762
transform -1 0 6536 0 1 2610
box -4 -6 52 206
use AND2X2  _2337_
timestamp 1597059762
transform -1 0 6600 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert274
timestamp 1597059762
transform -1 0 6648 0 1 2610
box -4 -6 52 206
use INVX1  _2637_
timestamp 1597059762
transform 1 0 6648 0 1 2610
box -4 -6 36 206
use NAND3X1  _2653_
timestamp 1597059762
transform 1 0 6680 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert154
timestamp 1597059762
transform -1 0 6856 0 1 2610
box -4 -6 52 206
use FILL  SFILL67440x26100
timestamp 1597059762
transform 1 0 6744 0 1 2610
box -4 -6 20 206
use FILL  SFILL67600x26100
timestamp 1597059762
transform 1 0 6760 0 1 2610
box -4 -6 20 206
use FILL  SFILL67760x26100
timestamp 1597059762
transform 1 0 6776 0 1 2610
box -4 -6 20 206
use FILL  SFILL67920x26100
timestamp 1597059762
transform 1 0 6792 0 1 2610
box -4 -6 20 206
use OR2X2  _2275_
timestamp 1597059762
transform 1 0 6856 0 1 2610
box -4 -6 68 206
use AOI22X1  _2940_
timestamp 1597059762
transform -1 0 7000 0 1 2610
box -4 -6 84 206
use AND2X2  _2291_
timestamp 1597059762
transform -1 0 7064 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert112
timestamp 1597059762
transform 1 0 7064 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert275
timestamp 1597059762
transform -1 0 7160 0 1 2610
box -4 -6 52 206
use OAI21X1  _2783_
timestamp 1597059762
transform -1 0 7224 0 1 2610
box -4 -6 68 206
use INVX1  _2782_
timestamp 1597059762
transform -1 0 7256 0 1 2610
box -4 -6 36 206
use BUFX2  BUFX2_insert248
timestamp 1597059762
transform 1 0 7256 0 1 2610
box -4 -6 52 206
use AOI21X1  _2780_
timestamp 1597059762
transform 1 0 7304 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert276
timestamp 1597059762
transform 1 0 7368 0 1 2610
box -4 -6 52 206
use INVX2  _2732_
timestamp 1597059762
transform -1 0 7448 0 1 2610
box -4 -6 36 206
use NOR2X1  _2735_
timestamp 1597059762
transform 1 0 7448 0 1 2610
box -4 -6 52 206
use INVX1  _2734_
timestamp 1597059762
transform -1 0 7528 0 1 2610
box -4 -6 36 206
use FILL  FILL72080x26100
timestamp 1597059762
transform 1 0 7528 0 1 2610
box -4 -6 20 206
use FILL  FILL72240x26100
timestamp 1597059762
transform 1 0 7544 0 1 2610
box -4 -6 20 206
use DFFPOSX1  _4286_
timestamp 1597059762
transform -1 0 200 0 -1 3010
box -4 -6 196 206
use AOI21X1  _3935_
timestamp 1597059762
transform 1 0 200 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3934_
timestamp 1597059762
transform -1 0 312 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert40
timestamp 1597059762
transform -1 0 360 0 -1 3010
box -4 -6 52 206
use MUX2X1  _3787_
timestamp 1597059762
transform -1 0 456 0 -1 3010
box -4 -6 100 206
use MUX2X1  _3999_
timestamp 1597059762
transform -1 0 552 0 -1 3010
box -4 -6 100 206
use DFFPOSX1  _4264_
timestamp 1597059762
transform 1 0 552 0 -1 3010
box -4 -6 196 206
use NOR2X1  _4106_
timestamp 1597059762
transform 1 0 808 0 -1 3010
box -4 -6 52 206
use FILL  SFILL7440x28100
timestamp 1597059762
transform -1 0 760 0 -1 3010
box -4 -6 20 206
use FILL  SFILL7600x28100
timestamp 1597059762
transform -1 0 776 0 -1 3010
box -4 -6 20 206
use FILL  SFILL7760x28100
timestamp 1597059762
transform -1 0 792 0 -1 3010
box -4 -6 20 206
use FILL  SFILL7920x28100
timestamp 1597059762
transform -1 0 808 0 -1 3010
box -4 -6 20 206
use OAI22X1  _3878_
timestamp 1597059762
transform -1 0 936 0 -1 3010
box -4 -6 84 206
use OAI21X1  _3877_
timestamp 1597059762
transform 1 0 936 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3894_
timestamp 1597059762
transform 1 0 1000 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4210_
timestamp 1597059762
transform 1 0 1048 0 -1 3010
box -4 -6 196 206
use MUX2X1  _3879_
timestamp 1597059762
transform -1 0 1336 0 -1 3010
box -4 -6 100 206
use OAI21X1  _3829_
timestamp 1597059762
transform 1 0 1336 0 -1 3010
box -4 -6 68 206
use AOI21X1  _3943_
timestamp 1597059762
transform 1 0 1400 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3942_
timestamp 1597059762
transform -1 0 1512 0 -1 3010
box -4 -6 52 206
use MUX2X1  _4043_
timestamp 1597059762
transform 1 0 1512 0 -1 3010
box -4 -6 100 206
use MUX2X1  _3831_
timestamp 1597059762
transform -1 0 1704 0 -1 3010
box -4 -6 100 206
use NOR2X1  _4153_
timestamp 1597059762
transform -1 0 1752 0 -1 3010
box -4 -6 52 206
use AOI21X1  _4154_
timestamp 1597059762
transform -1 0 1816 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert208
timestamp 1597059762
transform 1 0 1816 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4290_
timestamp 1597059762
transform -1 0 2056 0 -1 3010
box -4 -6 196 206
use AOI21X1  _3929_
timestamp 1597059762
transform 1 0 2056 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3928_
timestamp 1597059762
transform -1 0 2168 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert212
timestamp 1597059762
transform 1 0 2168 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4283_
timestamp 1597059762
transform 1 0 2280 0 -1 3010
box -4 -6 196 206
use FILL  SFILL22160x28100
timestamp 1597059762
transform -1 0 2232 0 -1 3010
box -4 -6 20 206
use FILL  SFILL22320x28100
timestamp 1597059762
transform -1 0 2248 0 -1 3010
box -4 -6 20 206
use FILL  SFILL22480x28100
timestamp 1597059762
transform -1 0 2264 0 -1 3010
box -4 -6 20 206
use FILL  SFILL22640x28100
timestamp 1597059762
transform -1 0 2280 0 -1 3010
box -4 -6 20 206
use MUX2X1  _3752_
timestamp 1597059762
transform 1 0 2472 0 -1 3010
box -4 -6 100 206
use NOR2X1  _3967_
timestamp 1597059762
transform -1 0 2616 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert194
timestamp 1597059762
transform 1 0 2616 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3753_
timestamp 1597059762
transform 1 0 2664 0 -1 3010
box -4 -6 52 206
use OAI22X1  _3755_
timestamp 1597059762
transform -1 0 2792 0 -1 3010
box -4 -6 84 206
use OAI21X1  _3754_
timestamp 1597059762
transform -1 0 2856 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3784_
timestamp 1597059762
transform -1 0 2904 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3541_
timestamp 1597059762
transform -1 0 2968 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _4174_
timestamp 1597059762
transform -1 0 3160 0 -1 3010
box -4 -6 196 206
use BUFX2  BUFX2_insert16
timestamp 1597059762
transform 1 0 3160 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3750_
timestamp 1597059762
transform -1 0 3272 0 -1 3010
box -4 -6 68 206
use OAI22X1  _3751_
timestamp 1597059762
transform 1 0 3272 0 -1 3010
box -4 -6 84 206
use MUX2X1  _3756_
timestamp 1597059762
transform 1 0 3352 0 -1 3010
box -4 -6 100 206
use MUX2X1  _3970_
timestamp 1597059762
transform -1 0 3544 0 -1 3010
box -4 -6 100 206
use OAI21X1  _3964_
timestamp 1597059762
transform 1 0 3544 0 -1 3010
box -4 -6 68 206
use OAI22X1  _3965_
timestamp 1597059762
transform 1 0 3608 0 -1 3010
box -4 -6 84 206
use AOI21X1  _3658_
timestamp 1597059762
transform 1 0 3688 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _4256_
timestamp 1597059762
transform -1 0 4008 0 -1 3010
box -4 -6 196 206
use FILL  SFILL37520x28100
timestamp 1597059762
transform -1 0 3768 0 -1 3010
box -4 -6 20 206
use FILL  SFILL37680x28100
timestamp 1597059762
transform -1 0 3784 0 -1 3010
box -4 -6 20 206
use FILL  SFILL37840x28100
timestamp 1597059762
transform -1 0 3800 0 -1 3010
box -4 -6 20 206
use FILL  SFILL38000x28100
timestamp 1597059762
transform -1 0 3816 0 -1 3010
box -4 -6 20 206
use DFFPOSX1  _4316_
timestamp 1597059762
transform 1 0 4008 0 -1 3010
box -4 -6 196 206
use OAI22X1  _3103_
timestamp 1597059762
transform 1 0 4200 0 -1 3010
box -4 -6 84 206
use BUFX2  BUFX2_insert157
timestamp 1597059762
transform 1 0 4280 0 -1 3010
box -4 -6 52 206
use INVX1  _3102_
timestamp 1597059762
transform 1 0 4328 0 -1 3010
box -4 -6 36 206
use INVX1  _3199_
timestamp 1597059762
transform 1 0 4360 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3201_
timestamp 1597059762
transform 1 0 4392 0 -1 3010
box -4 -6 68 206
use INVX1  _3192_
timestamp 1597059762
transform -1 0 4488 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3193_
timestamp 1597059762
transform -1 0 4536 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3200_
timestamp 1597059762
transform 1 0 4536 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3254_
timestamp 1597059762
transform -1 0 4648 0 -1 3010
box -4 -6 68 206
use INVX1  _3221_
timestamp 1597059762
transform -1 0 4680 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3223_
timestamp 1597059762
transform 1 0 4680 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3222_
timestamp 1597059762
transform 1 0 4744 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3237_
timestamp 1597059762
transform -1 0 4840 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3099_
timestamp 1597059762
transform -1 0 4888 0 -1 3010
box -4 -6 52 206
use INVX1  _3086_
timestamp 1597059762
transform 1 0 4888 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3088_
timestamp 1597059762
transform 1 0 4920 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3107_
timestamp 1597059762
transform -1 0 5032 0 -1 3010
box -4 -6 52 206
use INVX1  _3104_
timestamp 1597059762
transform 1 0 5032 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3106_
timestamp 1597059762
transform 1 0 5064 0 -1 3010
box -4 -6 68 206
use NAND3X1  _3122_
timestamp 1597059762
transform 1 0 5128 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3115_
timestamp 1597059762
transform 1 0 5192 0 -1 3010
box -4 -6 84 206
use NOR2X1  _3114_
timestamp 1597059762
transform -1 0 5384 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3113_
timestamp 1597059762
transform 1 0 5384 0 -1 3010
box -4 -6 68 206
use FILL  SFILL52720x28100
timestamp 1597059762
transform -1 0 5288 0 -1 3010
box -4 -6 20 206
use FILL  SFILL52880x28100
timestamp 1597059762
transform -1 0 5304 0 -1 3010
box -4 -6 20 206
use FILL  SFILL53040x28100
timestamp 1597059762
transform -1 0 5320 0 -1 3010
box -4 -6 20 206
use FILL  SFILL53200x28100
timestamp 1597059762
transform -1 0 5336 0 -1 3010
box -4 -6 20 206
use INVX1  _3111_
timestamp 1597059762
transform -1 0 5480 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3156_
timestamp 1597059762
transform 1 0 5480 0 -1 3010
box -4 -6 52 206
use OAI22X1  _2882_
timestamp 1597059762
transform 1 0 5528 0 -1 3010
box -4 -6 84 206
use INVX1  _2872_
timestamp 1597059762
transform 1 0 5608 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3098_
timestamp 1597059762
transform -1 0 5688 0 -1 3010
box -4 -6 52 206
use AOI22X1  _3096_
timestamp 1597059762
transform -1 0 5768 0 -1 3010
box -4 -6 84 206
use NOR2X1  _2889_
timestamp 1597059762
transform 1 0 5768 0 -1 3010
box -4 -6 52 206
use NAND3X1  _2924_
timestamp 1597059762
transform 1 0 5816 0 -1 3010
box -4 -6 68 206
use INVX1  _3123_
timestamp 1597059762
transform 1 0 5880 0 -1 3010
box -4 -6 36 206
use NOR2X1  _2907_
timestamp 1597059762
transform 1 0 5912 0 -1 3010
box -4 -6 52 206
use OAI21X1  _2906_
timestamp 1597059762
transform -1 0 6024 0 -1 3010
box -4 -6 68 206
use OAI21X1  _2899_
timestamp 1597059762
transform -1 0 6088 0 -1 3010
box -4 -6 68 206
use INVX1  _2890_
timestamp 1597059762
transform -1 0 6120 0 -1 3010
box -4 -6 36 206
use NAND2X1  _2383_
timestamp 1597059762
transform -1 0 6168 0 -1 3010
box -4 -6 52 206
use INVX1  _2900_
timestamp 1597059762
transform -1 0 6200 0 -1 3010
box -4 -6 36 206
use NOR2X1  _2352_
timestamp 1597059762
transform -1 0 6248 0 -1 3010
box -4 -6 52 206
use NOR3X1  _2367_
timestamp 1597059762
transform 1 0 6248 0 -1 3010
box -4 -6 132 206
use AND2X2  _2290_
timestamp 1597059762
transform 1 0 6376 0 -1 3010
box -4 -6 68 206
use AOI22X1  _2913_
timestamp 1597059762
transform 1 0 6440 0 -1 3010
box -4 -6 84 206
use NAND2X1  _2914_
timestamp 1597059762
transform 1 0 6520 0 -1 3010
box -4 -6 52 206
use NOR2X1  _2923_
timestamp 1597059762
transform -1 0 6616 0 -1 3010
box -4 -6 52 206
use NAND2X1  _2922_
timestamp 1597059762
transform 1 0 6616 0 -1 3010
box -4 -6 52 206
use AOI22X1  _2910_
timestamp 1597059762
transform -1 0 6744 0 -1 3010
box -4 -6 84 206
use OR2X2  _2274_
timestamp 1597059762
transform -1 0 6872 0 -1 3010
box -4 -6 68 206
use FILL  SFILL67440x28100
timestamp 1597059762
transform -1 0 6760 0 -1 3010
box -4 -6 20 206
use FILL  SFILL67600x28100
timestamp 1597059762
transform -1 0 6776 0 -1 3010
box -4 -6 20 206
use FILL  SFILL67760x28100
timestamp 1597059762
transform -1 0 6792 0 -1 3010
box -4 -6 20 206
use FILL  SFILL67920x28100
timestamp 1597059762
transform -1 0 6808 0 -1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert113
timestamp 1597059762
transform 1 0 6872 0 -1 3010
box -4 -6 52 206
use NOR3X1  _2597_
timestamp 1597059762
transform -1 0 7048 0 -1 3010
box -4 -6 132 206
use AOI21X1  _2594_
timestamp 1597059762
transform 1 0 7048 0 -1 3010
box -4 -6 68 206
use NAND2X1  _2595_
timestamp 1597059762
transform -1 0 7160 0 -1 3010
box -4 -6 52 206
use OAI21X1  _2544_
timestamp 1597059762
transform -1 0 7224 0 -1 3010
box -4 -6 68 206
use XNOR2X1  _2354_
timestamp 1597059762
transform 1 0 7224 0 -1 3010
box -4 -6 116 206
use NAND2X1  _2355_
timestamp 1597059762
transform -1 0 7384 0 -1 3010
box -4 -6 52 206
use XNOR2X1  _2353_
timestamp 1597059762
transform -1 0 7496 0 -1 3010
box -4 -6 116 206
use BUFX2  BUFX2_insert155
timestamp 1597059762
transform -1 0 7544 0 -1 3010
box -4 -6 52 206
use FILL  FILL72240x28100
timestamp 1597059762
transform -1 0 7560 0 -1 3010
box -4 -6 20 206
use NOR2X1  _4145_
timestamp 1597059762
transform 1 0 8 0 1 3010
box -4 -6 52 206
use AOI21X1  _4146_
timestamp 1597059762
transform -1 0 120 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert73
timestamp 1597059762
transform -1 0 168 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4270_
timestamp 1597059762
transform 1 0 168 0 1 3010
box -4 -6 196 206
use DFFPOSX1  _4184_
timestamp 1597059762
transform 1 0 360 0 1 3010
box -4 -6 196 206
use OAI21X1  _3571_
timestamp 1597059762
transform 1 0 552 0 1 3010
box -4 -6 68 206
use OAI21X1  _3570_
timestamp 1597059762
transform 1 0 616 0 1 3010
box -4 -6 68 206
use AOI21X1  _3674_
timestamp 1597059762
transform 1 0 680 0 1 3010
box -4 -6 68 206
use NOR2X1  _3673_
timestamp 1597059762
transform 1 0 808 0 1 3010
box -4 -6 52 206
use FILL  SFILL7440x30100
timestamp 1597059762
transform 1 0 744 0 1 3010
box -4 -6 20 206
use FILL  SFILL7600x30100
timestamp 1597059762
transform 1 0 760 0 1 3010
box -4 -6 20 206
use FILL  SFILL7760x30100
timestamp 1597059762
transform 1 0 776 0 1 3010
box -4 -6 20 206
use FILL  SFILL7920x30100
timestamp 1597059762
transform 1 0 792 0 1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert198
timestamp 1597059762
transform 1 0 856 0 1 3010
box -4 -6 52 206
use NOR2X1  _3661_
timestamp 1597059762
transform -1 0 952 0 1 3010
box -4 -6 52 206
use AOI21X1  _3662_
timestamp 1597059762
transform -1 0 1016 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4258_
timestamp 1597059762
transform 1 0 1016 0 1 3010
box -4 -6 196 206
use NAND2X1  _3594_
timestamp 1597059762
transform 1 0 1208 0 1 3010
box -4 -6 52 206
use OAI21X1  _3595_
timestamp 1597059762
transform -1 0 1320 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert254
timestamp 1597059762
transform 1 0 1320 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4274_
timestamp 1597059762
transform 1 0 1368 0 1 3010
box -4 -6 196 206
use BUFX2  BUFX2_insert7
timestamp 1597059762
transform 1 0 1560 0 1 3010
box -4 -6 52 206
use INVX4  _3575_
timestamp 1597059762
transform -1 0 1656 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert75
timestamp 1597059762
transform 1 0 1656 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4267_
timestamp 1597059762
transform 1 0 1704 0 1 3010
box -4 -6 196 206
use NOR2X1  _4139_
timestamp 1597059762
transform -1 0 1944 0 1 3010
box -4 -6 52 206
use AOI21X1  _4140_
timestamp 1597059762
transform -1 0 2008 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert108
timestamp 1597059762
transform -1 0 2056 0 1 3010
box -4 -6 52 206
use MUX2X1  _3966_
timestamp 1597059762
transform -1 0 2152 0 1 3010
box -4 -6 100 206
use NOR2X1  _3714_
timestamp 1597059762
transform -1 0 2200 0 1 3010
box -4 -6 52 206
use AOI21X1  _3715_
timestamp 1597059762
transform -1 0 2264 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4219_
timestamp 1597059762
transform 1 0 2328 0 1 3010
box -4 -6 196 206
use FILL  SFILL22640x30100
timestamp 1597059762
transform 1 0 2264 0 1 3010
box -4 -6 20 206
use FILL  SFILL22800x30100
timestamp 1597059762
transform 1 0 2280 0 1 3010
box -4 -6 20 206
use FILL  SFILL22960x30100
timestamp 1597059762
transform 1 0 2296 0 1 3010
box -4 -6 20 206
use FILL  SFILL23120x30100
timestamp 1597059762
transform 1 0 2312 0 1 3010
box -4 -6 20 206
use OAI21X1  _3968_
timestamp 1597059762
transform 1 0 2520 0 1 3010
box -4 -6 68 206
use OAI22X1  _3969_
timestamp 1597059762
transform 1 0 2584 0 1 3010
box -4 -6 84 206
use BUFX2  BUFX2_insert110
timestamp 1597059762
transform 1 0 2664 0 1 3010
box -4 -6 52 206
use OAI21X1  _3534_
timestamp 1597059762
transform 1 0 2712 0 1 3010
box -4 -6 68 206
use OAI21X1  _3540_
timestamp 1597059762
transform 1 0 2776 0 1 3010
box -4 -6 68 206
use NOR2X1  _3996_
timestamp 1597059762
transform 1 0 2840 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4176_
timestamp 1597059762
transform 1 0 2888 0 1 3010
box -4 -6 196 206
use OAI21X1  _3547_
timestamp 1597059762
transform 1 0 3080 0 1 3010
box -4 -6 68 206
use OAI21X1  _3546_
timestamp 1597059762
transform -1 0 3208 0 1 3010
box -4 -6 68 206
use OAI21X1  _3531_
timestamp 1597059762
transform 1 0 3208 0 1 3010
box -4 -6 68 206
use NOR2X1  _3749_
timestamp 1597059762
transform -1 0 3320 0 1 3010
box -4 -6 52 206
use OAI21X1  _3532_
timestamp 1597059762
transform -1 0 3384 0 1 3010
box -4 -6 68 206
use MUX2X1  _3805_
timestamp 1597059762
transform -1 0 3480 0 1 3010
box -4 -6 100 206
use MUX2X1  _4017_
timestamp 1597059762
transform -1 0 3576 0 1 3010
box -4 -6 100 206
use NOR2X1  _3963_
timestamp 1597059762
transform -1 0 3624 0 1 3010
box -4 -6 52 206
use NOR2X1  _3657_
timestamp 1597059762
transform 1 0 3624 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4171_
timestamp 1597059762
transform -1 0 3928 0 1 3010
box -4 -6 196 206
use FILL  SFILL36720x30100
timestamp 1597059762
transform 1 0 3672 0 1 3010
box -4 -6 20 206
use FILL  SFILL36880x30100
timestamp 1597059762
transform 1 0 3688 0 1 3010
box -4 -6 20 206
use FILL  SFILL37040x30100
timestamp 1597059762
transform 1 0 3704 0 1 3010
box -4 -6 20 206
use FILL  SFILL37200x30100
timestamp 1597059762
transform 1 0 3720 0 1 3010
box -4 -6 20 206
use AOI21X1  _3771_
timestamp 1597059762
transform 1 0 3928 0 1 3010
box -4 -6 68 206
use OAI21X1  _3770_
timestamp 1597059762
transform -1 0 4056 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert103
timestamp 1597059762
transform -1 0 4104 0 1 3010
box -4 -6 52 206
use INVX1  _3101_
timestamp 1597059762
transform 1 0 4104 0 1 3010
box -4 -6 36 206
use INVX1  _3190_
timestamp 1597059762
transform 1 0 4136 0 1 3010
box -4 -6 36 206
use OAI22X1  _3191_
timestamp 1597059762
transform -1 0 4248 0 1 3010
box -4 -6 84 206
use NOR2X1  _3195_
timestamp 1597059762
transform -1 0 4296 0 1 3010
box -4 -6 52 206
use NAND3X1  _3210_
timestamp 1597059762
transform 1 0 4296 0 1 3010
box -4 -6 68 206
use NOR2X1  _3202_
timestamp 1597059762
transform -1 0 4408 0 1 3010
box -4 -6 52 206
use OAI21X1  _3194_
timestamp 1597059762
transform -1 0 4472 0 1 3010
box -4 -6 68 206
use AOI22X1  _3093_
timestamp 1597059762
transform 1 0 4472 0 1 3010
box -4 -6 84 206
use NAND2X1  _3095_
timestamp 1597059762
transform 1 0 4552 0 1 3010
box -4 -6 52 206
use NOR2X1  _3253_
timestamp 1597059762
transform -1 0 4648 0 1 3010
box -4 -6 52 206
use NOR2X1  _3239_
timestamp 1597059762
transform -1 0 4696 0 1 3010
box -4 -6 52 206
use INVX1  _3236_
timestamp 1597059762
transform 1 0 4696 0 1 3010
box -4 -6 36 206
use OAI21X1  _3238_
timestamp 1597059762
transform 1 0 4728 0 1 3010
box -4 -6 68 206
use NAND2X1  _3171_
timestamp 1597059762
transform -1 0 4840 0 1 3010
box -4 -6 52 206
use OAI21X1  _3172_
timestamp 1597059762
transform -1 0 4904 0 1 3010
box -4 -6 68 206
use INVX1  _3170_
timestamp 1597059762
transform -1 0 4936 0 1 3010
box -4 -6 36 206
use INVX1  _3177_
timestamp 1597059762
transform 1 0 4936 0 1 3010
box -4 -6 36 206
use OAI21X1  _3179_
timestamp 1597059762
transform 1 0 4968 0 1 3010
box -4 -6 68 206
use NAND2X1  _3178_
timestamp 1597059762
transform -1 0 5080 0 1 3010
box -4 -6 52 206
use AOI22X1  _3250_
timestamp 1597059762
transform 1 0 5080 0 1 3010
box -4 -6 84 206
use NAND2X1  _3252_
timestamp 1597059762
transform 1 0 5160 0 1 3010
box -4 -6 52 206
use NAND2X1  _3117_
timestamp 1597059762
transform -1 0 5256 0 1 3010
box -4 -6 52 206
use NOR2X1  _3121_
timestamp 1597059762
transform -1 0 5368 0 1 3010
box -4 -6 52 206
use OAI21X1  _3110_
timestamp 1597059762
transform -1 0 5432 0 1 3010
box -4 -6 68 206
use FILL  SFILL52560x30100
timestamp 1597059762
transform 1 0 5256 0 1 3010
box -4 -6 20 206
use FILL  SFILL52720x30100
timestamp 1597059762
transform 1 0 5272 0 1 3010
box -4 -6 20 206
use FILL  SFILL52880x30100
timestamp 1597059762
transform 1 0 5288 0 1 3010
box -4 -6 20 206
use FILL  SFILL53040x30100
timestamp 1597059762
transform 1 0 5304 0 1 3010
box -4 -6 20 206
use INVX1  _3108_
timestamp 1597059762
transform -1 0 5464 0 1 3010
box -4 -6 36 206
use NAND2X1  _3112_
timestamp 1597059762
transform 1 0 5464 0 1 3010
box -4 -6 52 206
use OAI21X1  _3157_
timestamp 1597059762
transform -1 0 5576 0 1 3010
box -4 -6 68 206
use INVX1  _3155_
timestamp 1597059762
transform 1 0 5576 0 1 3010
box -4 -6 36 206
use NAND2X1  _3149_
timestamp 1597059762
transform 1 0 5608 0 1 3010
box -4 -6 52 206
use OAI21X1  _3150_
timestamp 1597059762
transform -1 0 5720 0 1 3010
box -4 -6 68 206
use INVX1  _3148_
timestamp 1597059762
transform -1 0 5752 0 1 3010
box -4 -6 36 206
use OAI21X1  _2888_
timestamp 1597059762
transform 1 0 5752 0 1 3010
box -4 -6 68 206
use NAND2X1  _2886_
timestamp 1597059762
transform -1 0 5864 0 1 3010
box -4 -6 52 206
use OAI21X1  _3132_
timestamp 1597059762
transform -1 0 5928 0 1 3010
box -4 -6 68 206
use INVX1  _3130_
timestamp 1597059762
transform -1 0 5960 0 1 3010
box -4 -6 36 206
use NAND2X1  _2904_
timestamp 1597059762
transform -1 0 6008 0 1 3010
box -4 -6 52 206
use AOI22X1  _3251_
timestamp 1597059762
transform 1 0 6008 0 1 3010
box -4 -6 84 206
use NOR3X1  _2382_
timestamp 1597059762
transform 1 0 6088 0 1 3010
box -4 -6 132 206
use NAND2X1  _2351_
timestamp 1597059762
transform -1 0 6264 0 1 3010
box -4 -6 52 206
use NAND2X1  _2328_
timestamp 1597059762
transform -1 0 6312 0 1 3010
box -4 -6 52 206
use AOI22X1  _3097_
timestamp 1597059762
transform 1 0 6312 0 1 3010
box -4 -6 84 206
use OAI21X1  _2863_
timestamp 1597059762
transform -1 0 6456 0 1 3010
box -4 -6 68 206
use NAND2X1  _2870_
timestamp 1597059762
transform -1 0 6504 0 1 3010
box -4 -6 52 206
use OR2X2  _2869_
timestamp 1597059762
transform -1 0 6568 0 1 3010
box -4 -6 68 206
use AOI22X1  _2917_
timestamp 1597059762
transform 1 0 6568 0 1 3010
box -4 -6 84 206
use AOI22X1  _2921_
timestamp 1597059762
transform 1 0 6648 0 1 3010
box -4 -6 84 206
use XOR2X1  _2098_
timestamp 1597059762
transform 1 0 6792 0 1 3010
box -4 -6 116 206
use FILL  SFILL67280x30100
timestamp 1597059762
transform 1 0 6728 0 1 3010
box -4 -6 20 206
use FILL  SFILL67440x30100
timestamp 1597059762
transform 1 0 6744 0 1 3010
box -4 -6 20 206
use FILL  SFILL67600x30100
timestamp 1597059762
transform 1 0 6760 0 1 3010
box -4 -6 20 206
use FILL  SFILL67760x30100
timestamp 1597059762
transform 1 0 6776 0 1 3010
box -4 -6 20 206
use NAND2X1  _3120_
timestamp 1597059762
transform -1 0 6952 0 1 3010
box -4 -6 52 206
use AOI22X1  _3118_
timestamp 1597059762
transform -1 0 7032 0 1 3010
box -4 -6 84 206
use OAI21X1  _2596_
timestamp 1597059762
transform 1 0 7032 0 1 3010
box -4 -6 68 206
use NAND2X1  _2542_
timestamp 1597059762
transform 1 0 7096 0 1 3010
box -4 -6 52 206
use INVX1  _2541_
timestamp 1597059762
transform -1 0 7176 0 1 3010
box -4 -6 36 206
use AOI21X1  _2543_
timestamp 1597059762
transform 1 0 7176 0 1 3010
box -4 -6 68 206
use XNOR2X1  _2157_
timestamp 1597059762
transform -1 0 7352 0 1 3010
box -4 -6 116 206
use NAND2X1  _2539_
timestamp 1597059762
transform 1 0 7352 0 1 3010
box -4 -6 52 206
use NOR2X1  _2540_
timestamp 1597059762
transform 1 0 7400 0 1 3010
box -4 -6 52 206
use INVX1  _2538_
timestamp 1597059762
transform -1 0 7480 0 1 3010
box -4 -6 36 206
use NAND2X1  _2101_
timestamp 1597059762
transform -1 0 7528 0 1 3010
box -4 -6 52 206
use FILL  FILL72080x30100
timestamp 1597059762
transform 1 0 7528 0 1 3010
box -4 -6 20 206
use FILL  FILL72240x30100
timestamp 1597059762
transform 1 0 7544 0 1 3010
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert34
timestamp 1597059762
transform 1 0 8 0 -1 3410
box -4 -6 148 206
use NOR2X1  _4165_
timestamp 1597059762
transform -1 0 200 0 -1 3410
box -4 -6 52 206
use AOI21X1  _4166_
timestamp 1597059762
transform -1 0 264 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4280_
timestamp 1597059762
transform 1 0 264 0 -1 3410
box -4 -6 196 206
use BUFX2  BUFX2_insert39
timestamp 1597059762
transform -1 0 504 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4248_
timestamp 1597059762
transform 1 0 504 0 -1 3410
box -4 -6 196 206
use MUX2X1  _4105_
timestamp 1597059762
transform 1 0 696 0 -1 3410
box -4 -6 100 206
use FILL  SFILL7920x32100
timestamp 1597059762
transform -1 0 808 0 -1 3410
box -4 -6 20 206
use FILL  SFILL8080x32100
timestamp 1597059762
transform -1 0 824 0 -1 3410
box -4 -6 20 206
use MUX2X1  _3893_
timestamp 1597059762
transform 1 0 856 0 -1 3410
box -4 -6 100 206
use OAI22X1  _3896_
timestamp 1597059762
transform -1 0 1032 0 -1 3410
box -4 -6 84 206
use FILL  SFILL8240x32100
timestamp 1597059762
transform -1 0 840 0 -1 3410
box -4 -6 20 206
use FILL  SFILL8400x32100
timestamp 1597059762
transform -1 0 856 0 -1 3410
box -4 -6 20 206
use NAND2X1  _3640_
timestamp 1597059762
transform 1 0 1032 0 -1 3410
box -4 -6 52 206
use OAI21X1  _3641_
timestamp 1597059762
transform -1 0 1144 0 -1 3410
box -4 -6 68 206
use OAI21X1  _3629_
timestamp 1597059762
transform 1 0 1144 0 -1 3410
box -4 -6 68 206
use NAND2X1  _3628_
timestamp 1597059762
transform -1 0 1256 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4242_
timestamp 1597059762
transform 1 0 1256 0 -1 3410
box -4 -6 196 206
use MUX2X1  _4039_
timestamp 1597059762
transform 1 0 1448 0 -1 3410
box -4 -6 100 206
use MUX2X1  _3827_
timestamp 1597059762
transform -1 0 1640 0 -1 3410
box -4 -6 100 206
use NOR2X1  _3930_
timestamp 1597059762
transform 1 0 1640 0 -1 3410
box -4 -6 52 206
use AOI21X1  _3931_
timestamp 1597059762
transform -1 0 1752 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4284_
timestamp 1597059762
transform -1 0 1944 0 -1 3410
box -4 -6 196 206
use NOR2X1  _4141_
timestamp 1597059762
transform 1 0 1944 0 -1 3410
box -4 -6 52 206
use AOI21X1  _4142_
timestamp 1597059762
transform -1 0 2056 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4220_
timestamp 1597059762
transform -1 0 2248 0 -1 3410
box -4 -6 196 206
use BUFX2  BUFX2_insert204
timestamp 1597059762
transform 1 0 2312 0 -1 3410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert31
timestamp 1597059762
transform 1 0 2360 0 -1 3410
box -4 -6 148 206
use FILL  SFILL22480x32100
timestamp 1597059762
transform -1 0 2264 0 -1 3410
box -4 -6 20 206
use FILL  SFILL22640x32100
timestamp 1597059762
transform -1 0 2280 0 -1 3410
box -4 -6 20 206
use FILL  SFILL22800x32100
timestamp 1597059762
transform -1 0 2296 0 -1 3410
box -4 -6 20 206
use FILL  SFILL22960x32100
timestamp 1597059762
transform -1 0 2312 0 -1 3410
box -4 -6 20 206
use BUFX2  BUFX2_insert119
timestamp 1597059762
transform 1 0 2504 0 -1 3410
box -4 -6 52 206
use MUX2X1  _3769_
timestamp 1597059762
transform -1 0 2648 0 -1 3410
box -4 -6 100 206
use BUFX2  BUFX2_insert257
timestamp 1597059762
transform 1 0 2648 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert89
timestamp 1597059762
transform 1 0 2696 0 -1 3410
box -4 -6 52 206
use OAI21X1  _3535_
timestamp 1597059762
transform 1 0 2744 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4172_
timestamp 1597059762
transform 1 0 2808 0 -1 3410
box -4 -6 196 206
use MUX2X1  _3981_
timestamp 1597059762
transform 1 0 3000 0 -1 3410
box -4 -6 100 206
use NOR2X1  _3806_
timestamp 1597059762
transform -1 0 3144 0 -1 3410
box -4 -6 52 206
use OAI22X1  _3808_
timestamp 1597059762
transform 1 0 3144 0 -1 3410
box -4 -6 84 206
use MUX2X1  _3813_
timestamp 1597059762
transform 1 0 3224 0 -1 3410
box -4 -6 100 206
use NOR2X1  _4018_
timestamp 1597059762
transform 1 0 3320 0 -1 3410
box -4 -6 52 206
use OAI21X1  _4019_
timestamp 1597059762
transform 1 0 3368 0 -1 3410
box -4 -6 68 206
use OAI22X1  _4020_
timestamp 1597059762
transform 1 0 3432 0 -1 3410
box -4 -6 84 206
use MUX2X1  _4025_
timestamp 1597059762
transform 1 0 3512 0 -1 3410
box -4 -6 100 206
use OAI21X1  _4114_
timestamp 1597059762
transform 1 0 3608 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4310_
timestamp 1597059762
transform 1 0 3736 0 -1 3410
box -4 -6 196 206
use FILL  SFILL36720x32100
timestamp 1597059762
transform -1 0 3688 0 -1 3410
box -4 -6 20 206
use FILL  SFILL36880x32100
timestamp 1597059762
transform -1 0 3704 0 -1 3410
box -4 -6 20 206
use FILL  SFILL37040x32100
timestamp 1597059762
transform -1 0 3720 0 -1 3410
box -4 -6 20 206
use FILL  SFILL37200x32100
timestamp 1597059762
transform -1 0 3736 0 -1 3410
box -4 -6 20 206
use AOI21X1  _3881_
timestamp 1597059762
transform 1 0 3928 0 -1 3410
box -4 -6 68 206
use OAI21X1  _3880_
timestamp 1597059762
transform -1 0 4056 0 -1 3410
box -4 -6 68 206
use OAI22X1  _3213_
timestamp 1597059762
transform 1 0 4056 0 -1 3410
box -4 -6 84 206
use INVX1  _3212_
timestamp 1597059762
transform 1 0 4136 0 -1 3410
box -4 -6 36 206
use INVX1  _3189_
timestamp 1597059762
transform 1 0 4168 0 -1 3410
box -4 -6 36 206
use NOR2X1  _3217_
timestamp 1597059762
transform -1 0 4248 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3232_
timestamp 1597059762
transform 1 0 4248 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3209_
timestamp 1597059762
transform -1 0 4360 0 -1 3410
box -4 -6 52 206
use INVX1  _3218_
timestamp 1597059762
transform 1 0 4360 0 -1 3410
box -4 -6 36 206
use OAI21X1  _3220_
timestamp 1597059762
transform 1 0 4392 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3224_
timestamp 1597059762
transform -1 0 4504 0 -1 3410
box -4 -6 52 206
use AOI22X1  _3225_
timestamp 1597059762
transform 1 0 4504 0 -1 3410
box -4 -6 84 206
use NOR2X1  _3231_
timestamp 1597059762
transform -1 0 4632 0 -1 3410
box -4 -6 52 206
use INVX1  _3080_
timestamp 1597059762
transform 1 0 4632 0 -1 3410
box -4 -6 36 206
use OAI22X1  _3081_
timestamp 1597059762
transform -1 0 4744 0 -1 3410
box -4 -6 84 206
use NOR2X1  _3173_
timestamp 1597059762
transform -1 0 4792 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3188_
timestamp 1597059762
transform 1 0 4792 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3187_
timestamp 1597059762
transform -1 0 4904 0 -1 3410
box -4 -6 52 206
use NOR2X1  _3180_
timestamp 1597059762
transform -1 0 4952 0 -1 3410
box -4 -6 52 206
use AOI22X1  _3206_
timestamp 1597059762
transform 1 0 4952 0 -1 3410
box -4 -6 84 206
use NAND2X1  _3208_
timestamp 1597059762
transform 1 0 5032 0 -1 3410
box -4 -6 52 206
use AOI22X1  _3228_
timestamp 1597059762
transform 1 0 5080 0 -1 3410
box -4 -6 84 206
use NAND2X1  _3230_
timestamp 1597059762
transform 1 0 5160 0 -1 3410
box -4 -6 52 206
use AND2X2  _2348_
timestamp 1597059762
transform -1 0 5272 0 -1 3410
box -4 -6 68 206
use NAND2X1  _3186_
timestamp 1597059762
transform -1 0 5384 0 -1 3410
box -4 -6 52 206
use AOI22X1  _3184_
timestamp 1597059762
transform -1 0 5464 0 -1 3410
box -4 -6 84 206
use FILL  SFILL52720x32100
timestamp 1597059762
transform -1 0 5288 0 -1 3410
box -4 -6 20 206
use FILL  SFILL52880x32100
timestamp 1597059762
transform -1 0 5304 0 -1 3410
box -4 -6 20 206
use FILL  SFILL53040x32100
timestamp 1597059762
transform -1 0 5320 0 -1 3410
box -4 -6 20 206
use FILL  SFILL53200x32100
timestamp 1597059762
transform -1 0 5336 0 -1 3410
box -4 -6 20 206
use NAND3X1  _3166_
timestamp 1597059762
transform 1 0 5464 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3151_
timestamp 1597059762
transform -1 0 5576 0 -1 3410
box -4 -6 52 206
use AOI22X1  _3185_
timestamp 1597059762
transform 1 0 5576 0 -1 3410
box -4 -6 84 206
use AOI22X1  _3229_
timestamp 1597059762
transform 1 0 5656 0 -1 3410
box -4 -6 84 206
use AOI22X1  _3207_
timestamp 1597059762
transform 1 0 5736 0 -1 3410
box -4 -6 84 206
use NOR2X1  _2256_
timestamp 1597059762
transform 1 0 5816 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2258_
timestamp 1597059762
transform 1 0 5864 0 -1 3410
box -4 -6 52 206
use AND2X2  _2257_
timestamp 1597059762
transform -1 0 5976 0 -1 3410
box -4 -6 68 206
use XNOR2X1  _2380_
timestamp 1597059762
transform 1 0 5976 0 -1 3410
box -4 -6 116 206
use NAND3X1  _2381_
timestamp 1597059762
transform -1 0 6152 0 -1 3410
box -4 -6 68 206
use XNOR2X1  _2379_
timestamp 1597059762
transform -1 0 6264 0 -1 3410
box -4 -6 116 206
use XNOR2X1  _2206_
timestamp 1597059762
transform 1 0 6264 0 -1 3410
box -4 -6 116 206
use AND2X2  _2205_
timestamp 1597059762
transform -1 0 6440 0 -1 3410
box -4 -6 68 206
use OR2X2  _2203_
timestamp 1597059762
transform -1 0 6504 0 -1 3410
box -4 -6 68 206
use INVX1  _2606_
timestamp 1597059762
transform 1 0 6504 0 -1 3410
box -4 -6 36 206
use NAND2X1  _2666_
timestamp 1597059762
transform -1 0 6584 0 -1 3410
box -4 -6 52 206
use NAND3X1  _2690_
timestamp 1597059762
transform 1 0 6584 0 -1 3410
box -4 -6 68 206
use INVX1  _2592_
timestamp 1597059762
transform 1 0 6648 0 -1 3410
box -4 -6 36 206
use AOI22X1  _2598_
timestamp 1597059762
transform 1 0 6680 0 -1 3410
box -4 -6 84 206
use NOR2X1  _3143_
timestamp 1597059762
transform -1 0 6872 0 -1 3410
box -4 -6 52 206
use FILL  SFILL67600x32100
timestamp 1597059762
transform -1 0 6776 0 -1 3410
box -4 -6 20 206
use FILL  SFILL67760x32100
timestamp 1597059762
transform -1 0 6792 0 -1 3410
box -4 -6 20 206
use FILL  SFILL67920x32100
timestamp 1597059762
transform -1 0 6808 0 -1 3410
box -4 -6 20 206
use FILL  SFILL68080x32100
timestamp 1597059762
transform -1 0 6824 0 -1 3410
box -4 -6 20 206
use NAND2X1  _3142_
timestamp 1597059762
transform -1 0 6920 0 -1 3410
box -4 -6 52 206
use AOI22X1  _3140_
timestamp 1597059762
transform -1 0 7000 0 -1 3410
box -4 -6 84 206
use AOI22X1  _3162_
timestamp 1597059762
transform 1 0 7000 0 -1 3410
box -4 -6 84 206
use NOR2X1  _3165_
timestamp 1597059762
transform -1 0 7128 0 -1 3410
box -4 -6 52 206
use NAND2X1  _3164_
timestamp 1597059762
transform 1 0 7128 0 -1 3410
box -4 -6 52 206
use INVX1  _2156_
timestamp 1597059762
transform 1 0 7176 0 -1 3410
box -4 -6 36 206
use AOI22X1  _3163_
timestamp 1597059762
transform 1 0 7208 0 -1 3410
box -4 -6 84 206
use AND2X2  _2593_
timestamp 1597059762
transform -1 0 7352 0 -1 3410
box -4 -6 68 206
use NAND3X1  _2568_
timestamp 1597059762
transform -1 0 7416 0 -1 3410
box -4 -6 68 206
use AOI21X1  _2589_
timestamp 1597059762
transform 1 0 7416 0 -1 3410
box -4 -6 68 206
use AOI21X1  _2827_
timestamp 1597059762
transform -1 0 7544 0 -1 3410
box -4 -6 68 206
use FILL  FILL72240x32100
timestamp 1597059762
transform -1 0 7560 0 -1 3410
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert25
timestamp 1597059762
transform 1 0 8 0 1 3410
box -4 -6 148 206
use DFFPOSX1  _4296_
timestamp 1597059762
transform 1 0 152 0 1 3410
box -4 -6 196 206
use DFFPOSX1  _4232_
timestamp 1597059762
transform 1 0 8 0 -1 3810
box -4 -6 196 206
use NOR2X1  _3740_
timestamp 1597059762
transform 1 0 200 0 -1 3810
box -4 -6 52 206
use AOI21X1  _3955_
timestamp 1597059762
transform 1 0 344 0 1 3410
box -4 -6 68 206
use NOR2X1  _3954_
timestamp 1597059762
transform -1 0 456 0 1 3410
box -4 -6 52 206
use AOI21X1  _3741_
timestamp 1597059762
transform -1 0 312 0 -1 3810
box -4 -6 68 206
use AOI21X1  _4170_
timestamp 1597059762
transform 1 0 312 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert231
timestamp 1597059762
transform 1 0 376 0 -1 3810
box -4 -6 52 206
use MUX2X1  _4109_
timestamp 1597059762
transform 1 0 456 0 1 3410
box -4 -6 100 206
use MUX2X1  _3897_
timestamp 1597059762
transform -1 0 648 0 1 3410
box -4 -6 100 206
use OAI21X1  _3708_
timestamp 1597059762
transform 1 0 424 0 -1 3810
box -4 -6 68 206
use NAND2X1  _3707_
timestamp 1597059762
transform -1 0 536 0 -1 3810
box -4 -6 52 206
use DFFPOSX1  _4200_
timestamp 1597059762
transform 1 0 536 0 -1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert5
timestamp 1597059762
transform 1 0 696 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert14
timestamp 1597059762
transform 1 0 648 0 1 3410
box -4 -6 52 206
use FILL  SFILL7760x36100
timestamp 1597059762
transform -1 0 792 0 -1 3810
box -4 -6 20 206
use FILL  SFILL7600x36100
timestamp 1597059762
transform -1 0 776 0 -1 3810
box -4 -6 20 206
use FILL  SFILL7440x36100
timestamp 1597059762
transform -1 0 760 0 -1 3810
box -4 -6 20 206
use FILL  SFILL7280x36100
timestamp 1597059762
transform -1 0 744 0 -1 3810
box -4 -6 20 206
use FILL  SFILL7760x34100
timestamp 1597059762
transform 1 0 776 0 1 3410
box -4 -6 20 206
use FILL  SFILL7600x34100
timestamp 1597059762
transform 1 0 760 0 1 3410
box -4 -6 20 206
use FILL  SFILL7440x34100
timestamp 1597059762
transform 1 0 744 0 1 3410
box -4 -6 20 206
use FILL  SFILL7920x34100
timestamp 1597059762
transform 1 0 792 0 1 3410
box -4 -6 20 206
use OAI21X1  _3899_
timestamp 1597059762
transform 1 0 792 0 -1 3810
box -4 -6 68 206
use OAI22X1  _4108_
timestamp 1597059762
transform 1 0 808 0 1 3410
box -4 -6 84 206
use MUX2X1  _4113_
timestamp 1597059762
transform 1 0 888 0 1 3410
box -4 -6 100 206
use OAI21X1  _4107_
timestamp 1597059762
transform -1 0 1048 0 1 3410
box -4 -6 68 206
use OAI22X1  _3900_
timestamp 1597059762
transform 1 0 856 0 -1 3810
box -4 -6 84 206
use OAI22X1  _4112_
timestamp 1597059762
transform -1 0 1016 0 -1 3810
box -4 -6 84 206
use OAI21X1  _3895_
timestamp 1597059762
transform -1 0 1112 0 1 3410
box -4 -6 68 206
use DFFPOSX1  _4216_
timestamp 1597059762
transform -1 0 1304 0 1 3410
box -4 -6 196 206
use OAI21X1  _4111_
timestamp 1597059762
transform 1 0 1016 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert229
timestamp 1597059762
transform 1 0 1080 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3633_
timestamp 1597059762
transform 1 0 1128 0 -1 3810
box -4 -6 68 206
use NAND2X1  _3632_
timestamp 1597059762
transform -1 0 1240 0 -1 3810
box -4 -6 52 206
use NAND2X1  _3606_
timestamp 1597059762
transform 1 0 1304 0 1 3410
box -4 -6 52 206
use OAI21X1  _3607_
timestamp 1597059762
transform -1 0 1416 0 1 3410
box -4 -6 68 206
use DFFPOSX1  _4244_
timestamp 1597059762
transform 1 0 1240 0 -1 3810
box -4 -6 196 206
use OAI21X1  _3576_
timestamp 1597059762
transform 1 0 1416 0 1 3410
box -4 -6 68 206
use DFFPOSX1  _4268_
timestamp 1597059762
transform 1 0 1480 0 1 3410
box -4 -6 196 206
use OAI21X1  _3577_
timestamp 1597059762
transform -1 0 1496 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4186_
timestamp 1597059762
transform -1 0 1688 0 -1 3810
box -4 -6 196 206
use MUX2X1  _3765_
timestamp 1597059762
transform 1 0 1672 0 1 3410
box -4 -6 100 206
use MUX2X1  _3977_
timestamp 1597059762
transform -1 0 1864 0 1 3410
box -4 -6 100 206
use BUFX2  BUFX2_insert234
timestamp 1597059762
transform -1 0 1736 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert123
timestamp 1597059762
transform 1 0 1736 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert197
timestamp 1597059762
transform 1 0 1784 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3767_
timestamp 1597059762
transform -1 0 1928 0 1 3410
box -4 -6 68 206
use OAI22X1  _3768_
timestamp 1597059762
transform -1 0 2008 0 1 3410
box -4 -6 84 206
use OAI22X1  _3980_
timestamp 1597059762
transform -1 0 2088 0 1 3410
box -4 -6 84 206
use NAND2X1  _3598_
timestamp 1597059762
transform 1 0 1832 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3599_
timestamp 1597059762
transform -1 0 1944 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert213
timestamp 1597059762
transform 1 0 1944 0 -1 3810
box -4 -6 52 206
use NOR2X1  _3766_
timestamp 1597059762
transform 1 0 1992 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3979_
timestamp 1597059762
transform -1 0 2152 0 1 3410
box -4 -6 68 206
use AOI21X1  _3717_
timestamp 1597059762
transform 1 0 2152 0 1 3410
box -4 -6 68 206
use NOR2X1  _3978_
timestamp 1597059762
transform -1 0 2088 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert233
timestamp 1597059762
transform 1 0 2088 0 -1 3810
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert30
timestamp 1597059762
transform 1 0 2136 0 -1 3810
box -4 -6 148 206
use FILL  SFILL22800x36100
timestamp 1597059762
transform -1 0 2296 0 -1 3810
box -4 -6 20 206
use FILL  SFILL22800x34100
timestamp 1597059762
transform 1 0 2280 0 1 3410
box -4 -6 20 206
use FILL  SFILL22640x34100
timestamp 1597059762
transform 1 0 2264 0 1 3410
box -4 -6 20 206
use NOR2X1  _3716_
timestamp 1597059762
transform -1 0 2264 0 1 3410
box -4 -6 52 206
use FILL  SFILL23280x36100
timestamp 1597059762
transform -1 0 2344 0 -1 3810
box -4 -6 20 206
use FILL  SFILL23120x36100
timestamp 1597059762
transform -1 0 2328 0 -1 3810
box -4 -6 20 206
use FILL  SFILL22960x36100
timestamp 1597059762
transform -1 0 2312 0 -1 3810
box -4 -6 20 206
use FILL  SFILL23120x34100
timestamp 1597059762
transform 1 0 2312 0 1 3410
box -4 -6 20 206
use FILL  SFILL22960x34100
timestamp 1597059762
transform 1 0 2296 0 1 3410
box -4 -6 20 206
use OAI21X1  _3617_
timestamp 1597059762
transform 1 0 2344 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert4
timestamp 1597059762
transform 1 0 2328 0 1 3410
box -4 -6 52 206
use NAND2X1  _3616_
timestamp 1597059762
transform -1 0 2456 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3583_
timestamp 1597059762
transform 1 0 2376 0 1 3410
box -4 -6 68 206
use NAND2X1  _3582_
timestamp 1597059762
transform -1 0 2488 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4204_
timestamp 1597059762
transform 1 0 2488 0 1 3410
box -4 -6 196 206
use DFFPOSX1  _4236_
timestamp 1597059762
transform 1 0 2456 0 -1 3810
box -4 -6 196 206
use INVX4  _3566_
timestamp 1597059762
transform 1 0 2680 0 1 3410
box -4 -6 52 206
use OAI22X1  _3764_
timestamp 1597059762
transform -1 0 2808 0 1 3410
box -4 -6 84 206
use NOR2X1  _3762_
timestamp 1597059762
transform 1 0 2808 0 1 3410
box -4 -6 52 206
use MUX2X1  _3761_
timestamp 1597059762
transform -1 0 2744 0 -1 3810
box -4 -6 100 206
use MUX2X1  _3973_
timestamp 1597059762
transform -1 0 2840 0 -1 3810
box -4 -6 100 206
use OAI21X1  _3763_
timestamp 1597059762
transform -1 0 2920 0 1 3410
box -4 -6 68 206
use NOR2X1  _3974_
timestamp 1597059762
transform 1 0 2920 0 1 3410
box -4 -6 52 206
use OAI22X1  _3976_
timestamp 1597059762
transform -1 0 3048 0 1 3410
box -4 -6 84 206
use NAND2X1  _3691_
timestamp 1597059762
transform -1 0 2888 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3692_
timestamp 1597059762
transform -1 0 2952 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4192_
timestamp 1597059762
transform 1 0 2952 0 -1 3810
box -4 -6 196 206
use OAI21X1  _3975_
timestamp 1597059762
transform 1 0 3048 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert17
timestamp 1597059762
transform 1 0 3112 0 1 3410
box -4 -6 52 206
use INVX4  _3554_
timestamp 1597059762
transform 1 0 3160 0 1 3410
box -4 -6 52 206
use OAI21X1  _3807_
timestamp 1597059762
transform -1 0 3272 0 1 3410
box -4 -6 68 206
use OAI21X1  _3811_
timestamp 1597059762
transform 1 0 3144 0 -1 3810
box -4 -6 68 206
use NOR2X1  _3810_
timestamp 1597059762
transform 1 0 3208 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3631_
timestamp 1597059762
transform 1 0 3272 0 1 3410
box -4 -6 68 206
use NAND2X1  _3630_
timestamp 1597059762
transform -1 0 3384 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4243_
timestamp 1597059762
transform 1 0 3384 0 1 3410
box -4 -6 196 206
use OAI22X1  _3812_
timestamp 1597059762
transform 1 0 3256 0 -1 3810
box -4 -6 84 206
use NOR2X1  _4022_
timestamp 1597059762
transform 1 0 3336 0 -1 3810
box -4 -6 52 206
use AOI21X1  _3650_
timestamp 1597059762
transform 1 0 3384 0 -1 3810
box -4 -6 68 206
use AOI21X1  _4115_
timestamp 1597059762
transform 1 0 3576 0 1 3410
box -4 -6 68 206
use NOR2X1  _3649_
timestamp 1597059762
transform 1 0 3448 0 -1 3810
box -4 -6 52 206
use NAND2X1  _3590_
timestamp 1597059762
transform 1 0 3496 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3591_
timestamp 1597059762
transform -1 0 3608 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4208_
timestamp 1597059762
transform -1 0 3800 0 -1 3810
box -4 -6 196 206
use DFFPOSX1  _4312_
timestamp 1597059762
transform 1 0 3640 0 1 3410
box -4 -6 196 206
use FILL  SFILL38000x36100
timestamp 1597059762
transform -1 0 3816 0 -1 3810
box -4 -6 20 206
use FILL  SFILL38160x36100
timestamp 1597059762
transform -1 0 3832 0 -1 3810
box -4 -6 20 206
use FILL  SFILL38480x36100
timestamp 1597059762
transform -1 0 3864 0 -1 3810
box -4 -6 20 206
use FILL  SFILL38320x36100
timestamp 1597059762
transform -1 0 3848 0 -1 3810
box -4 -6 20 206
use FILL  SFILL38800x34100
timestamp 1597059762
transform 1 0 3880 0 1 3410
box -4 -6 20 206
use FILL  SFILL38640x34100
timestamp 1597059762
transform 1 0 3864 0 1 3410
box -4 -6 20 206
use FILL  SFILL38480x34100
timestamp 1597059762
transform 1 0 3848 0 1 3410
box -4 -6 20 206
use FILL  SFILL38320x34100
timestamp 1597059762
transform 1 0 3832 0 1 3410
box -4 -6 20 206
use BUFX2  BUFX2_insert225
timestamp 1597059762
transform -1 0 3912 0 -1 3810
box -4 -6 52 206
use AND2X2  _2254_
timestamp 1597059762
transform -1 0 3960 0 1 3410
box -4 -6 68 206
use NOR2X1  _2253_
timestamp 1597059762
transform -1 0 4056 0 1 3410
box -4 -6 52 206
use NOR2X1  _2255_
timestamp 1597059762
transform -1 0 4008 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4326_
timestamp 1597059762
transform 1 0 3912 0 -1 3810
box -4 -6 196 206
use NOR2X1  _2265_
timestamp 1597059762
transform -1 0 4104 0 1 3410
box -4 -6 52 206
use NOR2X1  _2267_
timestamp 1597059762
transform 1 0 4104 0 1 3410
box -4 -6 52 206
use INVX1  _3196_
timestamp 1597059762
transform 1 0 4152 0 1 3410
box -4 -6 36 206
use OAI21X1  _3198_
timestamp 1597059762
transform 1 0 4184 0 1 3410
box -4 -6 68 206
use INVX1  _3211_
timestamp 1597059762
transform -1 0 4136 0 -1 3810
box -4 -6 36 206
use NOR2X1  _2268_
timestamp 1597059762
transform -1 0 4184 0 -1 3810
box -4 -6 52 206
use NOR2X1  _2270_
timestamp 1597059762
transform 1 0 4184 0 -1 3810
box -4 -6 52 206
use AOI22X1  _3203_
timestamp 1597059762
transform -1 0 4328 0 1 3410
box -4 -6 84 206
use NAND2X1  _3205_
timestamp 1597059762
transform -1 0 4376 0 1 3410
box -4 -6 52 206
use NAND2X1  _3249_
timestamp 1597059762
transform -1 0 4424 0 1 3410
box -4 -6 52 206
use AND2X2  _2269_
timestamp 1597059762
transform -1 0 4296 0 -1 3810
box -4 -6 68 206
use AND2X2  _2266_
timestamp 1597059762
transform -1 0 4360 0 -1 3810
box -4 -6 68 206
use OR2X2  _2287_
timestamp 1597059762
transform 1 0 4360 0 -1 3810
box -4 -6 68 206
use AOI22X1  _3247_
timestamp 1597059762
transform -1 0 4504 0 1 3410
box -4 -6 84 206
use INVX1  _3234_
timestamp 1597059762
transform 1 0 4504 0 1 3410
box -4 -6 36 206
use NAND2X1  _3227_
timestamp 1597059762
transform 1 0 4536 0 1 3410
box -4 -6 52 206
use OAI22X1  _3235_
timestamp 1597059762
transform -1 0 4664 0 1 3410
box -4 -6 84 206
use AOI22X1  _3204_
timestamp 1597059762
transform -1 0 4504 0 -1 3810
box -4 -6 84 206
use AOI22X1  _3094_
timestamp 1597059762
transform 1 0 4504 0 -1 3810
box -4 -6 84 206
use OR2X2  _2282_
timestamp 1597059762
transform -1 0 4648 0 -1 3810
box -4 -6 68 206
use OAI22X1  _3169_
timestamp 1597059762
transform 1 0 4664 0 1 3410
box -4 -6 84 206
use INVX1  _3168_
timestamp 1597059762
transform -1 0 4776 0 1 3410
box -4 -6 36 206
use AOI22X1  _3181_
timestamp 1597059762
transform 1 0 4776 0 1 3410
box -4 -6 84 206
use INVX1  _3167_
timestamp 1597059762
transform -1 0 4680 0 -1 3810
box -4 -6 36 206
use INVX1  _3079_
timestamp 1597059762
transform 1 0 4680 0 -1 3810
box -4 -6 36 206
use OR2X2  _2286_
timestamp 1597059762
transform 1 0 4712 0 -1 3810
box -4 -6 68 206
use AOI22X1  _3182_
timestamp 1597059762
transform -1 0 4856 0 -1 3810
box -4 -6 84 206
use NAND2X1  _3183_
timestamp 1597059762
transform -1 0 4904 0 1 3410
box -4 -6 52 206
use OAI21X1  _3176_
timestamp 1597059762
transform -1 0 4968 0 1 3410
box -4 -6 68 206
use INVX1  _3174_
timestamp 1597059762
transform -1 0 5000 0 1 3410
box -4 -6 36 206
use NOR2X1  _2345_
timestamp 1597059762
transform 1 0 5000 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert149
timestamp 1597059762
transform -1 0 4904 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert190
timestamp 1597059762
transform -1 0 4952 0 -1 3810
box -4 -6 52 206
use OR2X2  _2283_
timestamp 1597059762
transform 1 0 4952 0 -1 3810
box -4 -6 68 206
use AOI22X1  _3116_
timestamp 1597059762
transform -1 0 5096 0 -1 3810
box -4 -6 84 206
use AND2X2  _2346_
timestamp 1597059762
transform 1 0 5048 0 1 3410
box -4 -6 68 206
use OAI22X1  _2349_
timestamp 1597059762
transform 1 0 5112 0 1 3410
box -4 -6 84 206
use NOR2X1  _2350_
timestamp 1597059762
transform -1 0 5240 0 1 3410
box -4 -6 52 206
use NAND2X1  _2363_
timestamp 1597059762
transform 1 0 5096 0 -1 3810
box -4 -6 52 206
use OR2X2  _2364_
timestamp 1597059762
transform 1 0 5144 0 -1 3810
box -4 -6 68 206
use AOI22X1  _2365_
timestamp 1597059762
transform -1 0 5288 0 -1 3810
box -4 -6 84 206
use FILL  SFILL52880x36100
timestamp 1597059762
transform -1 0 5304 0 -1 3810
box -4 -6 20 206
use FILL  SFILL52880x34100
timestamp 1597059762
transform 1 0 5288 0 1 3410
box -4 -6 20 206
use FILL  SFILL52720x34100
timestamp 1597059762
transform 1 0 5272 0 1 3410
box -4 -6 20 206
use FILL  SFILL52560x34100
timestamp 1597059762
transform 1 0 5256 0 1 3410
box -4 -6 20 206
use FILL  SFILL52400x34100
timestamp 1597059762
transform 1 0 5240 0 1 3410
box -4 -6 20 206
use FILL  SFILL53360x36100
timestamp 1597059762
transform -1 0 5352 0 -1 3810
box -4 -6 20 206
use FILL  SFILL53200x36100
timestamp 1597059762
transform -1 0 5336 0 -1 3810
box -4 -6 20 206
use FILL  SFILL53040x36100
timestamp 1597059762
transform -1 0 5320 0 -1 3810
box -4 -6 20 206
use OR2X2  _2362_
timestamp 1597059762
transform -1 0 5416 0 -1 3810
box -4 -6 68 206
use INVX1  _3152_
timestamp 1597059762
transform 1 0 5352 0 1 3410
box -4 -6 36 206
use NOR2X1  _2347_
timestamp 1597059762
transform -1 0 5352 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert10
timestamp 1597059762
transform -1 0 5464 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3154_
timestamp 1597059762
transform 1 0 5384 0 1 3410
box -4 -6 68 206
use NOR2X1  _3158_
timestamp 1597059762
transform -1 0 5496 0 1 3410
box -4 -6 52 206
use OAI22X1  _3147_
timestamp 1597059762
transform 1 0 5496 0 1 3410
box -4 -6 84 206
use INVX1  _3146_
timestamp 1597059762
transform -1 0 5608 0 1 3410
box -4 -6 36 206
use XOR2X1  _2191_
timestamp 1597059762
transform -1 0 5720 0 1 3410
box -4 -6 116 206
use INVX1  _2187_
timestamp 1597059762
transform 1 0 5464 0 -1 3810
box -4 -6 36 206
use NOR2X1  _2189_
timestamp 1597059762
transform 1 0 5496 0 -1 3810
box -4 -6 52 206
use INVX1  _2188_
timestamp 1597059762
transform -1 0 5576 0 -1 3810
box -4 -6 36 206
use NOR2X1  _2190_
timestamp 1597059762
transform 1 0 5576 0 -1 3810
box -4 -6 52 206
use NAND2X1  _3131_
timestamp 1597059762
transform 1 0 5720 0 1 3410
box -4 -6 52 206
use AOI21X1  _2192_
timestamp 1597059762
transform 1 0 5768 0 1 3410
box -4 -6 68 206
use AOI22X1  _2603_
timestamp 1597059762
transform -1 0 5704 0 -1 3810
box -4 -6 84 206
use INVX1  _2520_
timestamp 1597059762
transform -1 0 5736 0 -1 3810
box -4 -6 36 206
use INVX1  _2883_
timestamp 1597059762
transform 1 0 5736 0 -1 3810
box -4 -6 36 206
use XNOR2X1  _2607_
timestamp 1597059762
transform -1 0 5880 0 -1 3810
box -4 -6 116 206
use XNOR2X1  _2197_
timestamp 1597059762
transform 1 0 5832 0 1 3410
box -4 -6 116 206
use NAND2X1  _2198_
timestamp 1597059762
transform -1 0 5992 0 1 3410
box -4 -6 52 206
use INVX1  _2200_
timestamp 1597059762
transform 1 0 5992 0 1 3410
box -4 -6 36 206
use XNOR2X1  _2219_
timestamp 1597059762
transform 1 0 5880 0 -1 3810
box -4 -6 116 206
use INVX1  _2522_
timestamp 1597059762
transform 1 0 5992 0 -1 3810
box -4 -6 36 206
use NAND2X1  _2194_
timestamp 1597059762
transform 1 0 6072 0 -1 3810
box -4 -6 52 206
use NOR2X1  _2193_
timestamp 1597059762
transform 1 0 6024 0 -1 3810
box -4 -6 52 206
use INVX1  _2195_
timestamp 1597059762
transform 1 0 6072 0 1 3410
box -4 -6 36 206
use NOR2X1  _2196_
timestamp 1597059762
transform 1 0 6024 0 1 3410
box -4 -6 52 206
use NAND2X1  _2525_
timestamp 1597059762
transform 1 0 6152 0 -1 3810
box -4 -6 52 206
use INVX1  _2521_
timestamp 1597059762
transform 1 0 6120 0 -1 3810
box -4 -6 36 206
use OAI21X1  _2201_
timestamp 1597059762
transform 1 0 6104 0 1 3410
box -4 -6 68 206
use OAI21X1  _2524_
timestamp 1597059762
transform 1 0 6200 0 -1 3810
box -4 -6 68 206
use NAND2X1  _2225_
timestamp 1597059762
transform -1 0 6264 0 1 3410
box -4 -6 52 206
use NAND2X1  _2224_
timestamp 1597059762
transform 1 0 6168 0 1 3410
box -4 -6 52 206
use INVX1  _2220_
timestamp 1597059762
transform 1 0 6264 0 1 3410
box -4 -6 36 206
use NAND3X1  _2221_
timestamp 1597059762
transform 1 0 6296 0 1 3410
box -4 -6 68 206
use OAI21X1  _2218_
timestamp 1597059762
transform -1 0 6424 0 1 3410
box -4 -6 68 206
use NAND2X1  _2523_
timestamp 1597059762
transform -1 0 6312 0 -1 3810
box -4 -6 52 206
use OAI21X1  _2526_
timestamp 1597059762
transform 1 0 6312 0 -1 3810
box -4 -6 68 206
use NOR2X1  _2527_
timestamp 1597059762
transform -1 0 6424 0 -1 3810
box -4 -6 52 206
use INVX1  _2222_
timestamp 1597059762
transform 1 0 6424 0 1 3410
box -4 -6 36 206
use OAI21X1  _2223_
timestamp 1597059762
transform 1 0 6456 0 1 3410
box -4 -6 68 206
use NAND2X1  _2204_
timestamp 1597059762
transform -1 0 6568 0 1 3410
box -4 -6 52 206
use AOI21X1  _2202_
timestamp 1597059762
transform -1 0 6632 0 1 3410
box -4 -6 68 206
use AND2X2  _2591_
timestamp 1597059762
transform 1 0 6424 0 -1 3810
box -4 -6 68 206
use NAND3X1  _2689_
timestamp 1597059762
transform 1 0 6488 0 -1 3810
box -4 -6 68 206
use OAI21X1  _2599_
timestamp 1597059762
transform 1 0 6552 0 -1 3810
box -4 -6 68 206
use AOI22X1  _3160_
timestamp 1597059762
transform 1 0 6616 0 -1 3810
box -4 -6 84 206
use AND2X2  _2301_
timestamp 1597059762
transform -1 0 6760 0 -1 3810
box -4 -6 68 206
use AOI22X1  _2785_
timestamp 1597059762
transform -1 0 6744 0 1 3410
box -4 -6 84 206
use INVX1  _2199_
timestamp 1597059762
transform -1 0 6664 0 1 3410
box -4 -6 36 206
use FILL  SFILL67920x36100
timestamp 1597059762
transform -1 0 6808 0 -1 3810
box -4 -6 20 206
use FILL  SFILL67760x36100
timestamp 1597059762
transform -1 0 6792 0 -1 3810
box -4 -6 20 206
use FILL  SFILL67600x36100
timestamp 1597059762
transform -1 0 6776 0 -1 3810
box -4 -6 20 206
use FILL  SFILL67920x34100
timestamp 1597059762
transform 1 0 6792 0 1 3410
box -4 -6 20 206
use FILL  SFILL67760x34100
timestamp 1597059762
transform 1 0 6776 0 1 3410
box -4 -6 20 206
use FILL  SFILL67600x34100
timestamp 1597059762
transform 1 0 6760 0 1 3410
box -4 -6 20 206
use FILL  SFILL67440x34100
timestamp 1597059762
transform 1 0 6744 0 1 3410
box -4 -6 20 206
use FILL  SFILL68080x36100
timestamp 1597059762
transform -1 0 6824 0 -1 3810
box -4 -6 20 206
use OR2X2  _2285_
timestamp 1597059762
transform -1 0 6888 0 -1 3810
box -4 -6 68 206
use NAND2X1  _2756_
timestamp 1597059762
transform 1 0 6808 0 1 3410
box -4 -6 52 206
use NAND2X1  _3139_
timestamp 1597059762
transform -1 0 6904 0 1 3410
box -4 -6 52 206
use INVX1  _3145_
timestamp 1597059762
transform -1 0 6936 0 1 3410
box -4 -6 36 206
use AOI22X1  _3137_
timestamp 1597059762
transform -1 0 7016 0 1 3410
box -4 -6 84 206
use AOI22X1  _3159_
timestamp 1597059762
transform 1 0 7016 0 1 3410
box -4 -6 84 206
use NOR2X1  _2259_
timestamp 1597059762
transform 1 0 6888 0 -1 3810
box -4 -6 52 206
use NOR2X1  _2261_
timestamp 1597059762
transform 1 0 6936 0 -1 3810
box -4 -6 52 206
use AND2X2  _2260_
timestamp 1597059762
transform 1 0 6984 0 -1 3810
box -4 -6 68 206
use NAND2X1  _3161_
timestamp 1597059762
transform -1 0 7144 0 1 3410
box -4 -6 52 206
use AOI22X1  _3141_
timestamp 1597059762
transform -1 0 7224 0 1 3410
box -4 -6 84 206
use AOI22X1  _3119_
timestamp 1597059762
transform -1 0 7304 0 1 3410
box -4 -6 84 206
use XNOR2X1  _2174_
timestamp 1597059762
transform 1 0 7048 0 -1 3810
box -4 -6 116 206
use NOR2X1  _2181_
timestamp 1597059762
transform -1 0 7208 0 -1 3810
box -4 -6 52 206
use AOI21X1  _2184_
timestamp 1597059762
transform 1 0 7208 0 -1 3810
box -4 -6 68 206
use OAI21X1  _2185_
timestamp 1597059762
transform -1 0 7368 0 1 3410
box -4 -6 68 206
use AOI21X1  _2217_
timestamp 1597059762
transform -1 0 7432 0 1 3410
box -4 -6 68 206
use XNOR2X1  _2180_
timestamp 1597059762
transform 1 0 7272 0 -1 3810
box -4 -6 116 206
use NAND2X1  _2182_
timestamp 1597059762
transform -1 0 7432 0 -1 3810
box -4 -6 52 206
use OAI21X1  _2216_
timestamp 1597059762
transform 1 0 7432 0 1 3410
box -4 -6 68 206
use INVX1  _2528_
timestamp 1597059762
transform 1 0 7496 0 1 3410
box -4 -6 36 206
use AND2X2  _2215_
timestamp 1597059762
transform 1 0 7432 0 -1 3810
box -4 -6 68 206
use BUFX2  _2032_
timestamp 1597059762
transform 1 0 7496 0 -1 3810
box -4 -6 52 206
use FILL  FILL72080x34100
timestamp 1597059762
transform 1 0 7528 0 1 3410
box -4 -6 20 206
use FILL  FILL72240x34100
timestamp 1597059762
transform 1 0 7544 0 1 3410
box -4 -6 20 206
use FILL  FILL72240x36100
timestamp 1597059762
transform -1 0 7560 0 -1 3810
box -4 -6 20 206
use DFFPOSX1  _4202_
timestamp 1597059762
transform 1 0 8 0 1 3810
box -4 -6 196 206
use NAND2X1  _3711_
timestamp 1597059762
transform 1 0 200 0 1 3810
box -4 -6 52 206
use OAI21X1  _3712_
timestamp 1597059762
transform -1 0 312 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4298_
timestamp 1597059762
transform 1 0 312 0 1 3810
box -4 -6 196 206
use OAI21X1  _3700_
timestamp 1597059762
transform 1 0 504 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4196_
timestamp 1597059762
transform 1 0 568 0 1 3810
box -4 -6 196 206
use FILL  SFILL7600x38100
timestamp 1597059762
transform 1 0 760 0 1 3810
box -4 -6 20 206
use FILL  SFILL7760x38100
timestamp 1597059762
transform 1 0 776 0 1 3810
box -4 -6 20 206
use FILL  SFILL7920x38100
timestamp 1597059762
transform 1 0 792 0 1 3810
box -4 -6 20 206
use FILL  SFILL8080x38100
timestamp 1597059762
transform 1 0 808 0 1 3810
box -4 -6 20 206
use NAND2X1  _3699_
timestamp 1597059762
transform 1 0 824 0 1 3810
box -4 -6 52 206
use NOR2X1  _3898_
timestamp 1597059762
transform 1 0 872 0 1 3810
box -4 -6 52 206
use NOR2X1  _4110_
timestamp 1597059762
transform 1 0 920 0 1 3810
box -4 -6 52 206
use MUX2X1  _3901_
timestamp 1597059762
transform 1 0 968 0 1 3810
box -4 -6 100 206
use BUFX2  BUFX2_insert230
timestamp 1597059762
transform -1 0 1112 0 1 3810
box -4 -6 52 206
use NOR2X1  _3744_
timestamp 1597059762
transform -1 0 1160 0 1 3810
box -4 -6 52 206
use DFFPOSX1  _4234_
timestamp 1597059762
transform -1 0 1352 0 1 3810
box -4 -6 196 206
use AOI21X1  _3745_
timestamp 1597059762
transform -1 0 1416 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert88
timestamp 1597059762
transform 1 0 1416 0 1 3810
box -4 -6 52 206
use OAI21X1  _3559_
timestamp 1597059762
transform 1 0 1464 0 1 3810
box -4 -6 68 206
use OAI21X1  _3558_
timestamp 1597059762
transform 1 0 1528 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4180_
timestamp 1597059762
transform 1 0 1592 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert205
timestamp 1597059762
transform -1 0 1832 0 1 3810
box -4 -6 52 206
use MUX2X1  _3849_
timestamp 1597059762
transform -1 0 1928 0 1 3810
box -4 -6 100 206
use MUX2X1  _4061_
timestamp 1597059762
transform -1 0 2024 0 1 3810
box -4 -6 100 206
use DFFPOSX1  _4212_
timestamp 1597059762
transform -1 0 2216 0 1 3810
box -4 -6 196 206
use NAND2X1  _3683_
timestamp 1597059762
transform 1 0 2216 0 1 3810
box -4 -6 52 206
use OAI21X1  _3684_
timestamp 1597059762
transform -1 0 2392 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4188_
timestamp 1597059762
transform -1 0 2584 0 1 3810
box -4 -6 196 206
use FILL  SFILL22640x38100
timestamp 1597059762
transform 1 0 2264 0 1 3810
box -4 -6 20 206
use FILL  SFILL22800x38100
timestamp 1597059762
transform 1 0 2280 0 1 3810
box -4 -6 20 206
use FILL  SFILL22960x38100
timestamp 1597059762
transform 1 0 2296 0 1 3810
box -4 -6 20 206
use FILL  SFILL23120x38100
timestamp 1597059762
transform 1 0 2312 0 1 3810
box -4 -6 20 206
use BUFX2  BUFX2_insert227
timestamp 1597059762
transform 1 0 2584 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert122
timestamp 1597059762
transform 1 0 2632 0 1 3810
box -4 -6 52 206
use NAND2X1  _3642_
timestamp 1597059762
transform 1 0 2680 0 1 3810
box -4 -6 52 206
use OAI21X1  _3643_
timestamp 1597059762
transform -1 0 2792 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4249_
timestamp 1597059762
transform 1 0 2792 0 1 3810
box -4 -6 196 206
use OAI21X1  _4023_
timestamp 1597059762
transform 1 0 2984 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4179_
timestamp 1597059762
transform -1 0 3240 0 1 3810
box -4 -6 196 206
use OAI22X1  _4024_
timestamp 1597059762
transform -1 0 3320 0 1 3810
box -4 -6 84 206
use DFFPOSX1  _4252_
timestamp 1597059762
transform -1 0 3512 0 1 3810
box -4 -6 196 206
use AOI21X1  _4126_
timestamp 1597059762
transform 1 0 3512 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4313_
timestamp 1597059762
transform 1 0 3576 0 1 3810
box -4 -6 196 206
use FILL  SFILL37680x38100
timestamp 1597059762
transform 1 0 3768 0 1 3810
box -4 -6 20 206
use FILL  SFILL37840x38100
timestamp 1597059762
transform 1 0 3784 0 1 3810
box -4 -6 20 206
use FILL  SFILL38000x38100
timestamp 1597059762
transform 1 0 3800 0 1 3810
box -4 -6 20 206
use FILL  SFILL38160x38100
timestamp 1597059762
transform 1 0 3816 0 1 3810
box -4 -6 20 206
use OAI21X1  _4125_
timestamp 1597059762
transform 1 0 3832 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4314_
timestamp 1597059762
transform 1 0 3896 0 1 3810
box -4 -6 196 206
use BUFX2  BUFX2_insert143
timestamp 1597059762
transform -1 0 4136 0 1 3810
box -4 -6 52 206
use OR2X2  _2288_
timestamp 1597059762
transform 1 0 4136 0 1 3810
box -4 -6 68 206
use AND2X2  _2305_
timestamp 1597059762
transform -1 0 4264 0 1 3810
box -4 -6 68 206
use OR2X2  _2289_
timestamp 1597059762
transform 1 0 4264 0 1 3810
box -4 -6 68 206
use AOI22X1  _3248_
timestamp 1597059762
transform -1 0 4408 0 1 3810
box -4 -6 84 206
use NAND2X1  _3219_
timestamp 1597059762
transform 1 0 4408 0 1 3810
box -4 -6 52 206
use AND2X2  _2298_
timestamp 1597059762
transform 1 0 4456 0 1 3810
box -4 -6 68 206
use AOI22X1  _3226_
timestamp 1597059762
transform -1 0 4600 0 1 3810
box -4 -6 84 206
use AND2X2  _2304_
timestamp 1597059762
transform -1 0 4664 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert140
timestamp 1597059762
transform 1 0 4664 0 1 3810
box -4 -6 52 206
use AND2X2  _2302_
timestamp 1597059762
transform 1 0 4712 0 1 3810
box -4 -6 68 206
use NAND2X1  _3241_
timestamp 1597059762
transform 1 0 4776 0 1 3810
box -4 -6 52 206
use NAND2X1  _3197_
timestamp 1597059762
transform -1 0 4872 0 1 3810
box -4 -6 52 206
use NAND2X1  _3175_
timestamp 1597059762
transform -1 0 4920 0 1 3810
box -4 -6 52 206
use NAND2X1  _3087_
timestamp 1597059762
transform -1 0 4968 0 1 3810
box -4 -6 52 206
use AND2X2  _2299_
timestamp 1597059762
transform 1 0 4968 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert47
timestamp 1597059762
transform 1 0 5032 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert48
timestamp 1597059762
transform 1 0 5080 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert151
timestamp 1597059762
transform 1 0 5128 0 1 3810
box -4 -6 52 206
use NAND2X1  _2361_
timestamp 1597059762
transform 1 0 5176 0 1 3810
box -4 -6 52 206
use XNOR2X1  _2608_
timestamp 1597059762
transform -1 0 5400 0 1 3810
box -4 -6 116 206
use NAND2X1  _3153_
timestamp 1597059762
transform 1 0 5400 0 1 3810
box -4 -6 52 206
use FILL  SFILL52240x38100
timestamp 1597059762
transform 1 0 5224 0 1 3810
box -4 -6 20 206
use FILL  SFILL52400x38100
timestamp 1597059762
transform 1 0 5240 0 1 3810
box -4 -6 20 206
use FILL  SFILL52560x38100
timestamp 1597059762
transform 1 0 5256 0 1 3810
box -4 -6 20 206
use FILL  SFILL52720x38100
timestamp 1597059762
transform 1 0 5272 0 1 3810
box -4 -6 20 206
use NAND2X1  _3109_
timestamp 1597059762
transform -1 0 5496 0 1 3810
box -4 -6 52 206
use NOR2X1  _2186_
timestamp 1597059762
transform 1 0 5496 0 1 3810
box -4 -6 52 206
use INVX1  _2600_
timestamp 1597059762
transform 1 0 5544 0 1 3810
box -4 -6 36 206
use AOI22X1  _2602_
timestamp 1597059762
transform 1 0 5576 0 1 3810
box -4 -6 84 206
use BUFX2  BUFX2_insert141
timestamp 1597059762
transform -1 0 5704 0 1 3810
box -4 -6 52 206
use INVX1  _2601_
timestamp 1597059762
transform -1 0 5736 0 1 3810
box -4 -6 36 206
use BUFX2  BUFX2_insert142
timestamp 1597059762
transform 1 0 5736 0 1 3810
box -4 -6 52 206
use NAND3X1  _2614_
timestamp 1597059762
transform -1 0 5848 0 1 3810
box -4 -6 68 206
use NAND2X1  _2668_
timestamp 1597059762
transform 1 0 5848 0 1 3810
box -4 -6 52 206
use OAI21X1  _2677_
timestamp 1597059762
transform 1 0 5896 0 1 3810
box -4 -6 68 206
use NAND2X1  _2370_
timestamp 1597059762
transform -1 0 6008 0 1 3810
box -4 -6 52 206
use XNOR2X1  _2368_
timestamp 1597059762
transform -1 0 6120 0 1 3810
box -4 -6 116 206
use INVX1  _2604_
timestamp 1597059762
transform 1 0 6120 0 1 3810
box -4 -6 36 206
use NOR2X1  _2605_
timestamp 1597059762
transform -1 0 6200 0 1 3810
box -4 -6 52 206
use AOI21X1  _2676_
timestamp 1597059762
transform -1 0 6264 0 1 3810
box -4 -6 68 206
use NOR2X1  _2675_
timestamp 1597059762
transform 1 0 6264 0 1 3810
box -4 -6 52 206
use INVX1  _2674_
timestamp 1597059762
transform 1 0 6312 0 1 3810
box -4 -6 36 206
use INVX1  _2667_
timestamp 1597059762
transform 1 0 6344 0 1 3810
box -4 -6 36 206
use AOI21X1  _2688_
timestamp 1597059762
transform -1 0 6440 0 1 3810
box -4 -6 68 206
use NOR2X1  _2626_
timestamp 1597059762
transform 1 0 6440 0 1 3810
box -4 -6 52 206
use OR2X2  _2284_
timestamp 1597059762
transform 1 0 6488 0 1 3810
box -4 -6 68 206
use AOI22X1  _3138_
timestamp 1597059762
transform -1 0 6632 0 1 3810
box -4 -6 84 206
use AND2X2  _2300_
timestamp 1597059762
transform -1 0 6696 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert11
timestamp 1597059762
transform -1 0 6744 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert191
timestamp 1597059762
transform 1 0 6808 0 1 3810
box -4 -6 52 206
use FILL  SFILL67440x38100
timestamp 1597059762
transform 1 0 6744 0 1 3810
box -4 -6 20 206
use FILL  SFILL67600x38100
timestamp 1597059762
transform 1 0 6760 0 1 3810
box -4 -6 20 206
use FILL  SFILL67760x38100
timestamp 1597059762
transform 1 0 6776 0 1 3810
box -4 -6 20 206
use FILL  SFILL67920x38100
timestamp 1597059762
transform 1 0 6792 0 1 3810
box -4 -6 20 206
use BUFX2  BUFX2_insert153
timestamp 1597059762
transform -1 0 6904 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert150
timestamp 1597059762
transform -1 0 6952 0 1 3810
box -4 -6 52 206
use NAND2X1  _2177_
timestamp 1597059762
transform 1 0 6952 0 1 3810
box -4 -6 52 206
use NOR2X1  _2166_
timestamp 1597059762
transform 1 0 7000 0 1 3810
box -4 -6 52 206
use INVX1  _2167_
timestamp 1597059762
transform 1 0 7048 0 1 3810
box -4 -6 36 206
use OAI21X1  _2168_
timestamp 1597059762
transform 1 0 7080 0 1 3810
box -4 -6 68 206
use INVX1  _2165_
timestamp 1597059762
transform -1 0 7176 0 1 3810
box -4 -6 36 206
use NAND2X1  _2173_
timestamp 1597059762
transform -1 0 7224 0 1 3810
box -4 -6 52 206
use NAND3X1  _2175_
timestamp 1597059762
transform -1 0 7288 0 1 3810
box -4 -6 68 206
use OAI21X1  _2183_
timestamp 1597059762
transform 1 0 7288 0 1 3810
box -4 -6 68 206
use NAND2X1  _2179_
timestamp 1597059762
transform 1 0 7352 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert152
timestamp 1597059762
transform 1 0 7400 0 1 3810
box -4 -6 52 206
use OR2X2  _2178_
timestamp 1597059762
transform -1 0 7512 0 1 3810
box -4 -6 68 206
use BUFX2  _2043_
timestamp 1597059762
transform 1 0 7512 0 1 3810
box -4 -6 52 206
use DFFPOSX1  _4276_
timestamp 1597059762
transform 1 0 8 0 -1 4210
box -4 -6 196 206
use AOI21X1  _3947_
timestamp 1597059762
transform 1 0 200 0 -1 4210
box -4 -6 68 206
use NOR2X1  _3946_
timestamp 1597059762
transform 1 0 264 0 -1 4210
box -4 -6 52 206
use NOR2X1  _4169_
timestamp 1597059762
transform -1 0 360 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4197_
timestamp 1597059762
transform -1 0 552 0 -1 4210
box -4 -6 196 206
use OAI21X1  _3702_
timestamp 1597059762
transform 1 0 552 0 -1 4210
box -4 -6 68 206
use NAND2X1  _3701_
timestamp 1597059762
transform -1 0 664 0 -1 4210
box -4 -6 52 206
use MUX2X1  _4131_
timestamp 1597059762
transform 1 0 664 0 -1 4210
box -4 -6 100 206
use FILL  SFILL7600x40100
timestamp 1597059762
transform -1 0 776 0 -1 4210
box -4 -6 20 206
use FILL  SFILL7760x40100
timestamp 1597059762
transform -1 0 792 0 -1 4210
box -4 -6 20 206
use FILL  SFILL7920x40100
timestamp 1597059762
transform -1 0 808 0 -1 4210
box -4 -6 20 206
use FILL  SFILL8080x40100
timestamp 1597059762
transform -1 0 824 0 -1 4210
box -4 -6 20 206
use NOR2X1  _4132_
timestamp 1597059762
transform 1 0 824 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4134_
timestamp 1597059762
transform -1 0 952 0 -1 4210
box -4 -6 84 206
use BUFX2  BUFX2_insert126
timestamp 1597059762
transform -1 0 1000 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4133_
timestamp 1597059762
transform -1 0 1064 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4181_
timestamp 1597059762
transform -1 0 1256 0 -1 4210
box -4 -6 196 206
use OAI21X1  _3562_
timestamp 1597059762
transform 1 0 1256 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3561_
timestamp 1597059762
transform -1 0 1384 0 -1 4210
box -4 -6 68 206
use MUX2X1  _4135_
timestamp 1597059762
transform 1 0 1384 0 -1 4210
box -4 -6 100 206
use BUFX2  BUFX2_insert258
timestamp 1597059762
transform -1 0 1528 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert210
timestamp 1597059762
transform -1 0 1576 0 -1 4210
box -4 -6 52 206
use NOR2X1  _4062_
timestamp 1597059762
transform -1 0 1624 0 -1 4210
box -4 -6 52 206
use NOR2X1  _3850_
timestamp 1597059762
transform -1 0 1672 0 -1 4210
box -4 -6 52 206
use OAI22X1  _3852_
timestamp 1597059762
transform 1 0 1672 0 -1 4210
box -4 -6 84 206
use OAI21X1  _3851_
timestamp 1597059762
transform -1 0 1816 0 -1 4210
box -4 -6 68 206
use OAI22X1  _4064_
timestamp 1597059762
transform 1 0 1816 0 -1 4210
box -4 -6 84 206
use OAI21X1  _4063_
timestamp 1597059762
transform -1 0 1960 0 -1 4210
box -4 -6 68 206
use INVX8  _3962_
timestamp 1597059762
transform -1 0 2040 0 -1 4210
box -4 -6 84 206
use OAI21X1  _3567_
timestamp 1597059762
transform 1 0 2040 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3568_
timestamp 1597059762
transform -1 0 2168 0 -1 4210
box -4 -6 68 206
use FILL  SFILL21680x40100
timestamp 1597059762
transform -1 0 2184 0 -1 4210
box -4 -6 20 206
use FILL  SFILL21840x40100
timestamp 1597059762
transform -1 0 2200 0 -1 4210
box -4 -6 20 206
use FILL  SFILL22000x40100
timestamp 1597059762
transform -1 0 2216 0 -1 4210
box -4 -6 20 206
use DFFPOSX1  _4183_
timestamp 1597059762
transform -1 0 2424 0 -1 4210
box -4 -6 196 206
use FILL  SFILL22160x40100
timestamp 1597059762
transform -1 0 2232 0 -1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert120
timestamp 1597059762
transform -1 0 2472 0 -1 4210
box -4 -6 52 206
use NAND2X1  _3608_
timestamp 1597059762
transform 1 0 2472 0 -1 4210
box -4 -6 52 206
use OAI21X1  _3609_
timestamp 1597059762
transform -1 0 2584 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4217_
timestamp 1597059762
transform -1 0 2776 0 -1 4210
box -4 -6 196 206
use BUFX2  BUFX2_insert83
timestamp 1597059762
transform 1 0 2776 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4185_
timestamp 1597059762
transform -1 0 3016 0 -1 4210
box -4 -6 196 206
use OAI21X1  _3574_
timestamp 1597059762
transform 1 0 3016 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3573_
timestamp 1597059762
transform -1 0 3144 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3555_
timestamp 1597059762
transform 1 0 3144 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3556_
timestamp 1597059762
transform -1 0 3272 0 -1 4210
box -4 -6 68 206
use AOI21X1  _3664_
timestamp 1597059762
transform 1 0 3272 0 -1 4210
box -4 -6 68 206
use NOR2X1  _3663_
timestamp 1597059762
transform -1 0 3384 0 -1 4210
box -4 -6 52 206
use MUX2X1  _4124_
timestamp 1597059762
transform 1 0 3384 0 -1 4210
box -4 -6 100 206
use OAI21X1  _3597_
timestamp 1597059762
transform 1 0 3480 0 -1 4210
box -4 -6 68 206
use NAND2X1  _3596_
timestamp 1597059762
transform -1 0 3592 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4211_
timestamp 1597059762
transform 1 0 3592 0 -1 4210
box -4 -6 196 206
use FILL  SFILL37840x40100
timestamp 1597059762
transform -1 0 3800 0 -1 4210
box -4 -6 20 206
use FILL  SFILL38000x40100
timestamp 1597059762
transform -1 0 3816 0 -1 4210
box -4 -6 20 206
use FILL  SFILL38160x40100
timestamp 1597059762
transform -1 0 3832 0 -1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert269
timestamp 1597059762
transform 1 0 3848 0 -1 4210
box -4 -6 52 206
use AOI21X1  _4137_
timestamp 1597059762
transform 1 0 3896 0 -1 4210
box -4 -6 68 206
use OAI21X1  _4136_
timestamp 1597059762
transform -1 0 4024 0 -1 4210
box -4 -6 68 206
use FILL  SFILL38320x40100
timestamp 1597059762
transform -1 0 3848 0 -1 4210
box -4 -6 20 206
use AOI21X1  _3903_
timestamp 1597059762
transform 1 0 4024 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert106
timestamp 1597059762
transform 1 0 4088 0 -1 4210
box -4 -6 52 206
use OAI21X1  _3902_
timestamp 1597059762
transform -1 0 4200 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert45
timestamp 1597059762
transform -1 0 4248 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert2
timestamp 1597059762
transform 1 0 4248 0 -1 4210
box -4 -6 52 206
use OAI21X1  _3913_
timestamp 1597059762
transform -1 0 4360 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2271_
timestamp 1597059762
transform -1 0 4408 0 -1 4210
box -4 -6 52 206
use AND2X2  _2303_
timestamp 1597059762
transform 1 0 4408 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert179
timestamp 1597059762
transform -1 0 4520 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2262_
timestamp 1597059762
transform 1 0 4520 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2264_
timestamp 1597059762
transform 1 0 4568 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2250_
timestamp 1597059762
transform 1 0 4616 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2252_
timestamp 1597059762
transform 1 0 4664 0 -1 4210
box -4 -6 52 206
use INVX1  _3233_
timestamp 1597059762
transform -1 0 4744 0 -1 4210
box -4 -6 36 206
use NOR2X1  _2273_
timestamp 1597059762
transform 1 0 4744 0 -1 4210
box -4 -6 52 206
use AND2X2  _2272_
timestamp 1597059762
transform -1 0 4856 0 -1 4210
box -4 -6 68 206
use XOR2X1  _2513_
timestamp 1597059762
transform -1 0 4968 0 -1 4210
box -4 -6 116 206
use BUFX2  BUFX2_insert46
timestamp 1597059762
transform -1 0 5016 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert55
timestamp 1597059762
transform -1 0 5064 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert96
timestamp 1597059762
transform -1 0 5112 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert54
timestamp 1597059762
transform 1 0 5112 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert180
timestamp 1597059762
transform 1 0 5160 0 -1 4210
box -4 -6 52 206
use AND2X2  _2320_
timestamp 1597059762
transform 1 0 5208 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert97
timestamp 1597059762
transform 1 0 5336 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert95
timestamp 1597059762
transform 1 0 5384 0 -1 4210
box -4 -6 52 206
use FILL  SFILL52720x40100
timestamp 1597059762
transform -1 0 5288 0 -1 4210
box -4 -6 20 206
use FILL  SFILL52880x40100
timestamp 1597059762
transform -1 0 5304 0 -1 4210
box -4 -6 20 206
use FILL  SFILL53040x40100
timestamp 1597059762
transform -1 0 5320 0 -1 4210
box -4 -6 20 206
use FILL  SFILL53200x40100
timestamp 1597059762
transform -1 0 5336 0 -1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert222
timestamp 1597059762
transform 1 0 5432 0 -1 4210
box -4 -6 52 206
use OR2X2  _2692_
timestamp 1597059762
transform 1 0 5480 0 -1 4210
box -4 -6 68 206
use NAND2X1  _2693_
timestamp 1597059762
transform 1 0 5544 0 -1 4210
box -4 -6 52 206
use AOI22X1  _2694_
timestamp 1597059762
transform -1 0 5672 0 -1 4210
box -4 -6 84 206
use INVX1  _2691_
timestamp 1597059762
transform -1 0 5704 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2695_
timestamp 1597059762
transform -1 0 5768 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert0
timestamp 1597059762
transform 1 0 5768 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2765_
timestamp 1597059762
transform -1 0 5864 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert181
timestamp 1597059762
transform 1 0 5864 0 -1 4210
box -4 -6 52 206
use XNOR2X1  _2369_
timestamp 1597059762
transform -1 0 6024 0 -1 4210
box -4 -6 116 206
use XNOR2X1  _2700_
timestamp 1597059762
transform -1 0 6136 0 -1 4210
box -4 -6 116 206
use OAI21X1  _2767_
timestamp 1597059762
transform -1 0 6200 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert188
timestamp 1597059762
transform -1 0 6248 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2757_
timestamp 1597059762
transform 1 0 6248 0 -1 4210
box -4 -6 52 206
use AOI21X1  _2779_
timestamp 1597059762
transform -1 0 6360 0 -1 4210
box -4 -6 68 206
use NOR3X1  _2714_
timestamp 1597059762
transform 1 0 6360 0 -1 4210
box -4 -6 132 206
use INVX1  _2709_
timestamp 1597059762
transform 1 0 6488 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2710_
timestamp 1597059762
transform -1 0 6568 0 -1 4210
box -4 -6 52 206
use XNOR2X1  _2712_
timestamp 1597059762
transform 1 0 6568 0 -1 4210
box -4 -6 116 206
use BUFX2  BUFX2_insert189
timestamp 1597059762
transform 1 0 6680 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert9
timestamp 1597059762
transform 1 0 6728 0 -1 4210
box -4 -6 52 206
use FILL  SFILL67760x40100
timestamp 1597059762
transform -1 0 6792 0 -1 4210
box -4 -6 20 206
use FILL  SFILL67920x40100
timestamp 1597059762
transform -1 0 6808 0 -1 4210
box -4 -6 20 206
use FILL  SFILL68080x40100
timestamp 1597059762
transform -1 0 6824 0 -1 4210
box -4 -6 20 206
use FILL  SFILL68240x40100
timestamp 1597059762
transform -1 0 6840 0 -1 4210
box -4 -6 20 206
use OAI21X1  _2687_
timestamp 1597059762
transform 1 0 6840 0 -1 4210
box -4 -6 68 206
use OR2X2  _2155_
timestamp 1597059762
transform -1 0 6968 0 -1 4210
box -4 -6 68 206
use INVX1  _2153_
timestamp 1597059762
transform -1 0 7000 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2158_
timestamp 1597059762
transform 1 0 7000 0 -1 4210
box -4 -6 68 206
use XNOR2X1  _2163_
timestamp 1597059762
transform 1 0 7064 0 -1 4210
box -4 -6 116 206
use INVX1  _2171_
timestamp 1597059762
transform 1 0 7176 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2172_
timestamp 1597059762
transform -1 0 7256 0 -1 4210
box -4 -6 52 206
use OAI21X1  _2176_
timestamp 1597059762
transform -1 0 7320 0 -1 4210
box -4 -6 68 206
use INVX1  _2170_
timestamp 1597059762
transform -1 0 7352 0 -1 4210
box -4 -6 36 206
use AND2X2  _2546_
timestamp 1597059762
transform 1 0 7352 0 -1 4210
box -4 -6 68 206
use INVX1  _2572_
timestamp 1597059762
transform 1 0 7416 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2574_
timestamp 1597059762
transform 1 0 7448 0 -1 4210
box -4 -6 52 206
use NOR2X1  _2573_
timestamp 1597059762
transform 1 0 7496 0 -1 4210
box -4 -6 52 206
use FILL  FILL72240x40100
timestamp 1597059762
transform -1 0 7560 0 -1 4210
box -4 -6 20 206
use DFFPOSX1  _4292_
timestamp 1597059762
transform 1 0 8 0 1 4210
box -4 -6 196 206
use AOI21X1  _4158_
timestamp 1597059762
transform 1 0 200 0 1 4210
box -4 -6 68 206
use NOR2X1  _4157_
timestamp 1597059762
transform 1 0 264 0 1 4210
box -4 -6 52 206
use MUX2X1  _3853_
timestamp 1597059762
transform -1 0 408 0 1 4210
box -4 -6 100 206
use MUX2X1  _4065_
timestamp 1597059762
transform 1 0 408 0 1 4210
box -4 -6 100 206
use OAI22X1  _3856_
timestamp 1597059762
transform -1 0 584 0 1 4210
box -4 -6 84 206
use NOR2X1  _3854_
timestamp 1597059762
transform -1 0 632 0 1 4210
box -4 -6 52 206
use MUX2X1  _3919_
timestamp 1597059762
transform 1 0 632 0 1 4210
box -4 -6 100 206
use OAI22X1  _4068_
timestamp 1597059762
transform -1 0 872 0 1 4210
box -4 -6 84 206
use FILL  SFILL7280x42100
timestamp 1597059762
transform 1 0 728 0 1 4210
box -4 -6 20 206
use FILL  SFILL7440x42100
timestamp 1597059762
transform 1 0 744 0 1 4210
box -4 -6 20 206
use FILL  SFILL7600x42100
timestamp 1597059762
transform 1 0 760 0 1 4210
box -4 -6 20 206
use FILL  SFILL7760x42100
timestamp 1597059762
transform 1 0 776 0 1 4210
box -4 -6 20 206
use NOR2X1  _4066_
timestamp 1597059762
transform 1 0 872 0 1 4210
box -4 -6 52 206
use NOR2X1  _3920_
timestamp 1597059762
transform 1 0 920 0 1 4210
box -4 -6 52 206
use OAI22X1  _3922_
timestamp 1597059762
transform 1 0 968 0 1 4210
box -4 -6 84 206
use OAI21X1  _3921_
timestamp 1597059762
transform -1 0 1112 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert84
timestamp 1597059762
transform -1 0 1160 0 1 4210
box -4 -6 52 206
use OAI21X1  _4129_
timestamp 1597059762
transform 1 0 1160 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert260
timestamp 1597059762
transform -1 0 1272 0 1 4210
box -4 -6 52 206
use OAI22X1  _4130_
timestamp 1597059762
transform -1 0 1352 0 1 4210
box -4 -6 84 206
use NOR2X1  _4128_
timestamp 1597059762
transform -1 0 1400 0 1 4210
box -4 -6 52 206
use OAI21X1  _3917_
timestamp 1597059762
transform 1 0 1400 0 1 4210
box -4 -6 68 206
use OAI22X1  _3918_
timestamp 1597059762
transform -1 0 1544 0 1 4210
box -4 -6 84 206
use NOR2X1  _3916_
timestamp 1597059762
transform 1 0 1544 0 1 4210
box -4 -6 52 206
use MUX2X1  _3923_
timestamp 1597059762
transform 1 0 1592 0 1 4210
box -4 -6 100 206
use MUX2X1  _3857_
timestamp 1597059762
transform 1 0 1688 0 1 4210
box -4 -6 100 206
use MUX2X1  _4069_
timestamp 1597059762
transform -1 0 1880 0 1 4210
box -4 -6 100 206
use DFFPOSX1  _4260_
timestamp 1597059762
transform -1 0 2072 0 1 4210
box -4 -6 196 206
use AOI21X1  _3666_
timestamp 1597059762
transform 1 0 2072 0 1 4210
box -4 -6 68 206
use NOR2X1  _3665_
timestamp 1597059762
transform 1 0 2136 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert211
timestamp 1597059762
transform 1 0 2184 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert206
timestamp 1597059762
transform 1 0 2296 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert86
timestamp 1597059762
transform -1 0 2392 0 1 4210
box -4 -6 52 206
use OAI21X1  _4118_
timestamp 1597059762
transform -1 0 2456 0 1 4210
box -4 -6 68 206
use FILL  SFILL22320x42100
timestamp 1597059762
transform 1 0 2232 0 1 4210
box -4 -6 20 206
use FILL  SFILL22480x42100
timestamp 1597059762
transform 1 0 2248 0 1 4210
box -4 -6 20 206
use FILL  SFILL22640x42100
timestamp 1597059762
transform 1 0 2264 0 1 4210
box -4 -6 20 206
use FILL  SFILL22800x42100
timestamp 1597059762
transform 1 0 2280 0 1 4210
box -4 -6 20 206
use OAI22X1  _4119_
timestamp 1597059762
transform -1 0 2536 0 1 4210
box -4 -6 84 206
use NOR2X1  _4117_
timestamp 1597059762
transform -1 0 2584 0 1 4210
box -4 -6 52 206
use MUX2X1  _4116_
timestamp 1597059762
transform -1 0 2680 0 1 4210
box -4 -6 100 206
use BUFX2  BUFX2_insert261
timestamp 1597059762
transform 1 0 2680 0 1 4210
box -4 -6 52 206
use OAI21X1  _3906_
timestamp 1597059762
transform 1 0 2728 0 1 4210
box -4 -6 68 206
use NOR2X1  _3905_
timestamp 1597059762
transform 1 0 2792 0 1 4210
box -4 -6 52 206
use OAI22X1  _3907_
timestamp 1597059762
transform 1 0 2840 0 1 4210
box -4 -6 84 206
use MUX2X1  _3904_
timestamp 1597059762
transform -1 0 3016 0 1 4210
box -4 -6 100 206
use MUX2X1  _3912_
timestamp 1597059762
transform 1 0 3016 0 1 4210
box -4 -6 100 206
use NOR2X1  _4051_
timestamp 1597059762
transform -1 0 3160 0 1 4210
box -4 -6 52 206
use NOR2X1  _3839_
timestamp 1597059762
transform 1 0 3160 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4259_
timestamp 1597059762
transform 1 0 3208 0 1 4210
box -4 -6 196 206
use MUX2X1  _4050_
timestamp 1597059762
transform 1 0 3400 0 1 4210
box -4 -6 100 206
use MUX2X1  _3838_
timestamp 1597059762
transform 1 0 3496 0 1 4210
box -4 -6 100 206
use OAI21X1  _3840_
timestamp 1597059762
transform 1 0 3592 0 1 4210
box -4 -6 68 206
use OAI22X1  _3841_
timestamp 1597059762
transform -1 0 3736 0 1 4210
box -4 -6 84 206
use MUX2X1  _3846_
timestamp 1597059762
transform 1 0 3800 0 1 4210
box -4 -6 100 206
use FILL  SFILL37360x42100
timestamp 1597059762
transform 1 0 3736 0 1 4210
box -4 -6 20 206
use FILL  SFILL37520x42100
timestamp 1597059762
transform 1 0 3752 0 1 4210
box -4 -6 20 206
use FILL  SFILL37680x42100
timestamp 1597059762
transform 1 0 3768 0 1 4210
box -4 -6 20 206
use FILL  SFILL37840x42100
timestamp 1597059762
transform 1 0 3784 0 1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert99
timestamp 1597059762
transform 1 0 3896 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert105
timestamp 1597059762
transform 1 0 3944 0 1 4210
box -4 -6 52 206
use OAI21X1  _3858_
timestamp 1597059762
transform -1 0 4056 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4328_
timestamp 1597059762
transform 1 0 4056 0 1 4210
box -4 -6 196 206
use OAI21X1  _3891_
timestamp 1597059762
transform -1 0 4312 0 1 4210
box -4 -6 68 206
use AOI21X1  _3914_
timestamp 1597059762
transform 1 0 4312 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4329_
timestamp 1597059762
transform 1 0 4376 0 1 4210
box -4 -6 196 206
use AND2X2  _2263_
timestamp 1597059762
transform 1 0 4568 0 1 4210
box -4 -6 68 206
use AND2X2  _2251_
timestamp 1597059762
transform 1 0 4632 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert118
timestamp 1597059762
transform -1 0 4744 0 1 4210
box -4 -6 52 206
use NAND2X1  _2519_
timestamp 1597059762
transform 1 0 4744 0 1 4210
box -4 -6 52 206
use NAND3X1  _2515_
timestamp 1597059762
transform -1 0 4856 0 1 4210
box -4 -6 68 206
use NAND2X1  _2518_
timestamp 1597059762
transform -1 0 4904 0 1 4210
box -4 -6 52 206
use INVX1  _2514_
timestamp 1597059762
transform 1 0 4904 0 1 4210
box -4 -6 36 206
use BUFX2  BUFX2_insert243
timestamp 1597059762
transform 1 0 4936 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert182
timestamp 1597059762
transform 1 0 4984 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert224
timestamp 1597059762
transform -1 0 5080 0 1 4210
box -4 -6 52 206
use AND2X2  _2318_
timestamp 1597059762
transform 1 0 5080 0 1 4210
box -4 -6 68 206
use NOR2X1  _2317_
timestamp 1597059762
transform -1 0 5192 0 1 4210
box -4 -6 52 206
use OAI22X1  _2321_
timestamp 1597059762
transform 1 0 5192 0 1 4210
box -4 -6 84 206
use NOR2X1  _2319_
timestamp 1597059762
transform -1 0 5384 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert115
timestamp 1597059762
transform 1 0 5384 0 1 4210
box -4 -6 52 206
use FILL  SFILL52720x42100
timestamp 1597059762
transform 1 0 5272 0 1 4210
box -4 -6 20 206
use FILL  SFILL52880x42100
timestamp 1597059762
transform 1 0 5288 0 1 4210
box -4 -6 20 206
use FILL  SFILL53040x42100
timestamp 1597059762
transform 1 0 5304 0 1 4210
box -4 -6 20 206
use FILL  SFILL53200x42100
timestamp 1597059762
transform 1 0 5320 0 1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert223
timestamp 1597059762
transform 1 0 5432 0 1 4210
box -4 -6 52 206
use XNOR2X1  _2786_
timestamp 1597059762
transform -1 0 5592 0 1 4210
box -4 -6 116 206
use NOR2X1  _2851_
timestamp 1597059762
transform 1 0 5592 0 1 4210
box -4 -6 52 206
use INVX1  _2850_
timestamp 1597059762
transform 1 0 5640 0 1 4210
box -4 -6 36 206
use AOI21X1  _2853_
timestamp 1597059762
transform -1 0 5736 0 1 4210
box -4 -6 68 206
use NOR2X1  _2852_
timestamp 1597059762
transform 1 0 5736 0 1 4210
box -4 -6 52 206
use INVX1  _2787_
timestamp 1597059762
transform 1 0 5784 0 1 4210
box -4 -6 36 206
use NAND2X1  _2789_
timestamp 1597059762
transform 1 0 5816 0 1 4210
box -4 -6 52 206
use OR2X2  _2788_
timestamp 1597059762
transform 1 0 5864 0 1 4210
box -4 -6 68 206
use NAND3X1  _2790_
timestamp 1597059762
transform 1 0 5928 0 1 4210
box -4 -6 68 206
use INVX1  _2762_
timestamp 1597059762
transform 1 0 5992 0 1 4210
box -4 -6 36 206
use NAND2X1  _2764_
timestamp 1597059762
transform 1 0 6024 0 1 4210
box -4 -6 52 206
use AOI21X1  _2766_
timestamp 1597059762
transform 1 0 6072 0 1 4210
box -4 -6 68 206
use NOR2X1  _2763_
timestamp 1597059762
transform -1 0 6184 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert241
timestamp 1597059762
transform -1 0 6232 0 1 4210
box -4 -6 52 206
use NOR2X1  _2327_
timestamp 1597059762
transform 1 0 6232 0 1 4210
box -4 -6 52 206
use INVX1  _2707_
timestamp 1597059762
transform 1 0 6280 0 1 4210
box -4 -6 36 206
use NAND2X1  _2708_
timestamp 1597059762
transform -1 0 6360 0 1 4210
box -4 -6 52 206
use INVX1  _2806_
timestamp 1597059762
transform 1 0 6360 0 1 4210
box -4 -6 36 206
use AOI22X1  _2807_
timestamp 1597059762
transform 1 0 6392 0 1 4210
box -4 -6 84 206
use INVX1  _2804_
timestamp 1597059762
transform 1 0 6472 0 1 4210
box -4 -6 36 206
use INVX1  _2775_
timestamp 1597059762
transform 1 0 6504 0 1 4210
box -4 -6 36 206
use NAND3X1  _2776_
timestamp 1597059762
transform 1 0 6536 0 1 4210
box -4 -6 68 206
use AND2X2  _2711_
timestamp 1597059762
transform 1 0 6600 0 1 4210
box -4 -6 68 206
use NOR2X1  _2623_
timestamp 1597059762
transform 1 0 6664 0 1 4210
box -4 -6 52 206
use INVX1  _2619_
timestamp 1597059762
transform 1 0 6712 0 1 4210
box -4 -6 36 206
use NAND2X1  _2685_
timestamp 1597059762
transform 1 0 6808 0 1 4210
box -4 -6 52 206
use FILL  SFILL67440x42100
timestamp 1597059762
transform 1 0 6744 0 1 4210
box -4 -6 20 206
use FILL  SFILL67600x42100
timestamp 1597059762
transform 1 0 6760 0 1 4210
box -4 -6 20 206
use FILL  SFILL67760x42100
timestamp 1597059762
transform 1 0 6776 0 1 4210
box -4 -6 20 206
use FILL  SFILL67920x42100
timestamp 1597059762
transform 1 0 6792 0 1 4210
box -4 -6 20 206
use AOI21X1  _2686_
timestamp 1597059762
transform -1 0 6920 0 1 4210
box -4 -6 68 206
use AOI22X1  _2621_
timestamp 1597059762
transform 1 0 6920 0 1 4210
box -4 -6 84 206
use NAND2X1  _2678_
timestamp 1597059762
transform 1 0 7000 0 1 4210
box -4 -6 52 206
use NOR2X1  _2624_
timestamp 1597059762
transform -1 0 7096 0 1 4210
box -4 -6 52 206
use INVX1  _2620_
timestamp 1597059762
transform -1 0 7128 0 1 4210
box -4 -6 36 206
use NOR2X1  _2622_
timestamp 1597059762
transform -1 0 7176 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert242
timestamp 1597059762
transform 1 0 7176 0 1 4210
box -4 -6 52 206
use NAND2X1  _2169_
timestamp 1597059762
transform -1 0 7272 0 1 4210
box -4 -6 52 206
use AND2X2  _2548_
timestamp 1597059762
transform 1 0 7272 0 1 4210
box -4 -6 68 206
use NOR2X1  _2547_
timestamp 1597059762
transform 1 0 7336 0 1 4210
box -4 -6 52 206
use OAI22X1  _2549_
timestamp 1597059762
transform -1 0 7464 0 1 4210
box -4 -6 84 206
use AOI21X1  _2577_
timestamp 1597059762
transform -1 0 7528 0 1 4210
box -4 -6 68 206
use FILL  FILL72080x42100
timestamp 1597059762
transform 1 0 7528 0 1 4210
box -4 -6 20 206
use FILL  FILL72240x42100
timestamp 1597059762
transform 1 0 7544 0 1 4210
box -4 -6 20 206
use NOR2X1  _3734_
timestamp 1597059762
transform 1 0 8 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3735_
timestamp 1597059762
transform -1 0 120 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert67
timestamp 1597059762
transform -1 0 168 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert74
timestamp 1597059762
transform 1 0 168 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3733_
timestamp 1597059762
transform 1 0 216 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3732_
timestamp 1597059762
transform -1 0 328 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3855_
timestamp 1597059762
transform 1 0 328 0 -1 4610
box -4 -6 68 206
use OAI21X1  _4067_
timestamp 1597059762
transform 1 0 392 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3865_
timestamp 1597059762
transform 1 0 456 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert196
timestamp 1597059762
transform -1 0 552 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert192
timestamp 1597059762
transform -1 0 600 0 -1 4610
box -4 -6 52 206
use NOR2X1  _4077_
timestamp 1597059762
transform 1 0 600 0 -1 4610
box -4 -6 52 206
use OAI21X1  _4074_
timestamp 1597059762
transform 1 0 648 0 -1 4610
box -4 -6 68 206
use OAI22X1  _4075_
timestamp 1597059762
transform 1 0 776 0 -1 4610
box -4 -6 84 206
use FILL  SFILL7120x44100
timestamp 1597059762
transform -1 0 728 0 -1 4610
box -4 -6 20 206
use FILL  SFILL7280x44100
timestamp 1597059762
transform -1 0 744 0 -1 4610
box -4 -6 20 206
use FILL  SFILL7440x44100
timestamp 1597059762
transform -1 0 760 0 -1 4610
box -4 -6 20 206
use FILL  SFILL7600x44100
timestamp 1597059762
transform -1 0 776 0 -1 4610
box -4 -6 20 206
use NOR2X1  _4073_
timestamp 1597059762
transform -1 0 904 0 -1 4610
box -4 -6 52 206
use NOR2X1  _3861_
timestamp 1597059762
transform 1 0 904 0 -1 4610
box -4 -6 52 206
use DFFPOSX1  _4218_
timestamp 1597059762
transform -1 0 1144 0 -1 4610
box -4 -6 196 206
use OAI21X1  _3611_
timestamp 1597059762
transform 1 0 1144 0 -1 4610
box -4 -6 68 206
use NAND2X1  _3610_
timestamp 1597059762
transform 1 0 1208 0 -1 4610
box -4 -6 52 206
use MUX2X1  _4127_
timestamp 1597059762
transform -1 0 1352 0 -1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert71
timestamp 1597059762
transform 1 0 1352 0 -1 4610
box -4 -6 52 206
use MUX2X1  _3915_
timestamp 1597059762
transform -1 0 1496 0 -1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert68
timestamp 1597059762
transform 1 0 1496 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3739_
timestamp 1597059762
transform 1 0 1544 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3738_
timestamp 1597059762
transform -1 0 1656 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3884_
timestamp 1597059762
transform 1 0 1656 0 -1 4610
box -4 -6 68 206
use OAI22X1  _3885_
timestamp 1597059762
transform -1 0 1800 0 -1 4610
box -4 -6 84 206
use MUX2X1  _3890_
timestamp 1597059762
transform 1 0 1800 0 -1 4610
box -4 -6 100 206
use OAI21X1  _3888_
timestamp 1597059762
transform -1 0 1960 0 -1 4610
box -4 -6 68 206
use OAI22X1  _3889_
timestamp 1597059762
transform -1 0 2040 0 -1 4610
box -4 -6 84 206
use NOR2X1  _3883_
timestamp 1597059762
transform 1 0 2040 0 -1 4610
box -4 -6 52 206
use NOR2X1  _3887_
timestamp 1597059762
transform -1 0 2136 0 -1 4610
box -4 -6 52 206
use NAND2X1  _3705_
timestamp 1597059762
transform 1 0 2136 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3706_
timestamp 1597059762
transform -1 0 2248 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4199_
timestamp 1597059762
transform -1 0 2504 0 -1 4610
box -4 -6 196 206
use FILL  SFILL22480x44100
timestamp 1597059762
transform -1 0 2264 0 -1 4610
box -4 -6 20 206
use FILL  SFILL22640x44100
timestamp 1597059762
transform -1 0 2280 0 -1 4610
box -4 -6 20 206
use FILL  SFILL22800x44100
timestamp 1597059762
transform -1 0 2296 0 -1 4610
box -4 -6 20 206
use FILL  SFILL22960x44100
timestamp 1597059762
transform -1 0 2312 0 -1 4610
box -4 -6 20 206
use OAI21X1  _3710_
timestamp 1597059762
transform 1 0 2504 0 -1 4610
box -4 -6 68 206
use NAND2X1  _3709_
timestamp 1597059762
transform -1 0 2616 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert195
timestamp 1597059762
transform 1 0 2616 0 -1 4610
box -4 -6 52 206
use NOR2X1  _3909_
timestamp 1597059762
transform 1 0 2664 0 -1 4610
box -4 -6 52 206
use OAI22X1  _3911_
timestamp 1597059762
transform -1 0 2792 0 -1 4610
box -4 -6 84 206
use OAI21X1  _3910_
timestamp 1597059762
transform -1 0 2856 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4233_
timestamp 1597059762
transform -1 0 3048 0 -1 4610
box -4 -6 196 206
use OAI21X1  _3698_
timestamp 1597059762
transform 1 0 3048 0 -1 4610
box -4 -6 68 206
use NAND2X1  _3697_
timestamp 1597059762
transform -1 0 3160 0 -1 4610
box -4 -6 52 206
use NOR2X1  _3843_
timestamp 1597059762
transform -1 0 3208 0 -1 4610
box -4 -6 52 206
use OAI21X1  _3844_
timestamp 1597059762
transform 1 0 3208 0 -1 4610
box -4 -6 68 206
use OAI22X1  _3845_
timestamp 1597059762
transform 1 0 3272 0 -1 4610
box -4 -6 84 206
use OAI22X1  _4053_
timestamp 1597059762
transform 1 0 3352 0 -1 4610
box -4 -6 84 206
use OAI21X1  _4052_
timestamp 1597059762
transform -1 0 3496 0 -1 4610
box -4 -6 68 206
use NOR2X1  _3730_
timestamp 1597059762
transform -1 0 3544 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3731_
timestamp 1597059762
transform -1 0 3608 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4227_
timestamp 1597059762
transform -1 0 3800 0 -1 4610
box -4 -6 196 206
use FILL  SFILL38000x44100
timestamp 1597059762
transform -1 0 3816 0 -1 4610
box -4 -6 20 206
use FILL  SFILL38160x44100
timestamp 1597059762
transform -1 0 3832 0 -1 4610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert32
timestamp 1597059762
transform 1 0 3864 0 -1 4610
box -4 -6 148 206
use AOI21X1  _3859_
timestamp 1597059762
transform 1 0 4008 0 -1 4610
box -4 -6 68 206
use FILL  SFILL38320x44100
timestamp 1597059762
transform -1 0 3848 0 -1 4610
box -4 -6 20 206
use FILL  SFILL38480x44100
timestamp 1597059762
transform -1 0 3864 0 -1 4610
box -4 -6 20 206
use AOI21X1  _3848_
timestamp 1597059762
transform 1 0 4072 0 -1 4610
box -4 -6 68 206
use AOI21X1  _3892_
timestamp 1597059762
transform 1 0 4136 0 -1 4610
box -4 -6 68 206
use AOI21X1  _3925_
timestamp 1597059762
transform 1 0 4200 0 -1 4610
box -4 -6 68 206
use OAI21X1  _3924_
timestamp 1597059762
transform -1 0 4328 0 -1 4610
box -4 -6 68 206
use DFFPOSX1  _4330_
timestamp 1597059762
transform 1 0 4328 0 -1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert98
timestamp 1597059762
transform 1 0 4520 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert160
timestamp 1597059762
transform 1 0 4568 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert1
timestamp 1597059762
transform 1 0 4616 0 -1 4610
box -4 -6 52 206
use XNOR2X1  _2507_
timestamp 1597059762
transform -1 0 4776 0 -1 4610
box -4 -6 116 206
use INVX1  _2516_
timestamp 1597059762
transform 1 0 4776 0 -1 4610
box -4 -6 36 206
use OAI21X1  _2517_
timestamp 1597059762
transform 1 0 4808 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2509_
timestamp 1597059762
transform 1 0 4872 0 -1 4610
box -4 -6 52 206
use INVX1  _2508_
timestamp 1597059762
transform -1 0 4952 0 -1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert215
timestamp 1597059762
transform -1 0 5000 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2340_
timestamp 1597059762
transform -1 0 5048 0 -1 4610
box -4 -6 52 206
use OR2X2  _2609_
timestamp 1597059762
transform 1 0 5048 0 -1 4610
box -4 -6 68 206
use OAI22X1  _2344_
timestamp 1597059762
transform 1 0 5112 0 -1 4610
box -4 -6 84 206
use AND2X2  _2343_
timestamp 1597059762
transform -1 0 5256 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2342_
timestamp 1597059762
transform 1 0 5320 0 -1 4610
box -4 -6 52 206
use AOI21X1  _2672_
timestamp 1597059762
transform -1 0 5432 0 -1 4610
box -4 -6 68 206
use FILL  SFILL52560x44100
timestamp 1597059762
transform -1 0 5272 0 -1 4610
box -4 -6 20 206
use FILL  SFILL52720x44100
timestamp 1597059762
transform -1 0 5288 0 -1 4610
box -4 -6 20 206
use FILL  SFILL52880x44100
timestamp 1597059762
transform -1 0 5304 0 -1 4610
box -4 -6 20 206
use FILL  SFILL53040x44100
timestamp 1597059762
transform -1 0 5320 0 -1 4610
box -4 -6 20 206
use BUFX2  BUFX2_insert3
timestamp 1597059762
transform 1 0 5432 0 -1 4610
box -4 -6 52 206
use INVX1  _2791_
timestamp 1597059762
transform 1 0 5480 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2610_
timestamp 1597059762
transform 1 0 5512 0 -1 4610
box -4 -6 52 206
use AOI21X1  _2673_
timestamp 1597059762
transform -1 0 5624 0 -1 4610
box -4 -6 68 206
use INVX1  _2669_
timestamp 1597059762
transform -1 0 5656 0 -1 4610
box -4 -6 36 206
use AOI22X1  _2613_
timestamp 1597059762
transform 1 0 5656 0 -1 4610
box -4 -6 84 206
use OR2X2  _2611_
timestamp 1597059762
transform -1 0 5800 0 -1 4610
box -4 -6 68 206
use INVX1  _2758_
timestamp 1597059762
transform 1 0 5800 0 -1 4610
box -4 -6 36 206
use NOR2X1  _2759_
timestamp 1597059762
transform -1 0 5880 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2854_
timestamp 1597059762
transform -1 0 5944 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2796_
timestamp 1597059762
transform 1 0 5944 0 -1 4610
box -4 -6 52 206
use INVX1  _2698_
timestamp 1597059762
transform 1 0 5992 0 -1 4610
box -4 -6 36 206
use AOI21X1  _2761_
timestamp 1597059762
transform -1 0 6088 0 -1 4610
box -4 -6 68 206
use INVX1  _2760_
timestamp 1597059762
transform -1 0 6120 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2699_
timestamp 1597059762
transform -1 0 6168 0 -1 4610
box -4 -6 52 206
use NAND3X1  _2701_
timestamp 1597059762
transform 1 0 6168 0 -1 4610
box -4 -6 68 206
use AOI21X1  _2862_
timestamp 1597059762
transform -1 0 6296 0 -1 4610
box -4 -6 68 206
use INVX1  _2802_
timestamp 1597059762
transform 1 0 6296 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2810_
timestamp 1597059762
transform -1 0 6376 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2860_
timestamp 1597059762
transform 1 0 6376 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2803_
timestamp 1597059762
transform 1 0 6440 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2859_
timestamp 1597059762
transform -1 0 6552 0 -1 4610
box -4 -6 68 206
use NAND3X1  _2808_
timestamp 1597059762
transform 1 0 6552 0 -1 4610
box -4 -6 68 206
use OR2X2  _2805_
timestamp 1597059762
transform 1 0 6616 0 -1 4610
box -4 -6 68 206
use AND2X2  _2777_
timestamp 1597059762
transform 1 0 6680 0 -1 4610
box -4 -6 68 206
use NAND3X1  _2713_
timestamp 1597059762
transform 1 0 6808 0 -1 4610
box -4 -6 68 206
use FILL  SFILL67440x44100
timestamp 1597059762
transform -1 0 6760 0 -1 4610
box -4 -6 20 206
use FILL  SFILL67600x44100
timestamp 1597059762
transform -1 0 6776 0 -1 4610
box -4 -6 20 206
use FILL  SFILL67760x44100
timestamp 1597059762
transform -1 0 6792 0 -1 4610
box -4 -6 20 206
use FILL  SFILL67920x44100
timestamp 1597059762
transform -1 0 6808 0 -1 4610
box -4 -6 20 206
use NAND2X1  _2768_
timestamp 1597059762
transform 1 0 6872 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2778_
timestamp 1597059762
transform -1 0 6984 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert244
timestamp 1597059762
transform -1 0 7032 0 -1 4610
box -4 -6 52 206
use NAND3X1  _2625_
timestamp 1597059762
transform 1 0 7032 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert214
timestamp 1597059762
transform 1 0 7096 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2164_
timestamp 1597059762
transform -1 0 7208 0 -1 4610
box -4 -6 68 206
use INVX1  _2160_
timestamp 1597059762
transform 1 0 7208 0 -1 4610
box -4 -6 36 206
use OR2X2  _2162_
timestamp 1597059762
transform 1 0 7240 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2161_
timestamp 1597059762
transform -1 0 7352 0 -1 4610
box -4 -6 52 206
use NOR3X1  _2556_
timestamp 1597059762
transform 1 0 7352 0 -1 4610
box -4 -6 132 206
use OAI21X1  _2578_
timestamp 1597059762
transform 1 0 7480 0 -1 4610
box -4 -6 68 206
use FILL  FILL72240x44100
timestamp 1597059762
transform -1 0 7560 0 -1 4610
box -4 -6 20 206
use DFFPOSX1  _4229_
timestamp 1597059762
transform 1 0 8 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4228_
timestamp 1597059762
transform 1 0 200 0 1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert38
timestamp 1597059762
transform -1 0 440 0 1 4610
box -4 -6 52 206
use OAI22X1  _3867_
timestamp 1597059762
transform -1 0 520 0 1 4610
box -4 -6 84 206
use OAI21X1  _3866_
timestamp 1597059762
transform -1 0 584 0 1 4610
box -4 -6 68 206
use OAI21X1  _4078_
timestamp 1597059762
transform 1 0 584 0 1 4610
box -4 -6 68 206
use OAI22X1  _4079_
timestamp 1597059762
transform 1 0 648 0 1 4610
box -4 -6 84 206
use OAI21X1  _3601_
timestamp 1597059762
transform 1 0 792 0 1 4610
box -4 -6 68 206
use FILL  SFILL7280x46100
timestamp 1597059762
transform 1 0 728 0 1 4610
box -4 -6 20 206
use FILL  SFILL7440x46100
timestamp 1597059762
transform 1 0 744 0 1 4610
box -4 -6 20 206
use FILL  SFILL7600x46100
timestamp 1597059762
transform 1 0 760 0 1 4610
box -4 -6 20 206
use FILL  SFILL7760x46100
timestamp 1597059762
transform 1 0 776 0 1 4610
box -4 -6 20 206
use NAND2X1  _3600_
timestamp 1597059762
transform -1 0 904 0 1 4610
box -4 -6 52 206
use MUX2X1  _4080_
timestamp 1597059762
transform 1 0 904 0 1 4610
box -4 -6 100 206
use OAI21X1  _3862_
timestamp 1597059762
transform 1 0 1000 0 1 4610
box -4 -6 68 206
use OAI22X1  _3863_
timestamp 1597059762
transform 1 0 1064 0 1 4610
box -4 -6 84 206
use MUX2X1  _3868_
timestamp 1597059762
transform 1 0 1144 0 1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert37
timestamp 1597059762
transform 1 0 1240 0 1 4610
box -4 -6 52 206
use OAI21X1  _3605_
timestamp 1597059762
transform 1 0 1288 0 1 4610
box -4 -6 68 206
use NAND2X1  _3604_
timestamp 1597059762
transform -1 0 1400 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4215_
timestamp 1597059762
transform 1 0 1400 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4231_
timestamp 1597059762
transform 1 0 1592 0 1 4610
box -4 -6 196 206
use OAI21X1  _4096_
timestamp 1597059762
transform 1 0 1784 0 1 4610
box -4 -6 68 206
use OAI22X1  _4097_
timestamp 1597059762
transform -1 0 1928 0 1 4610
box -4 -6 84 206
use OAI21X1  _4100_
timestamp 1597059762
transform 1 0 1928 0 1 4610
box -4 -6 68 206
use NOR2X1  _4095_
timestamp 1597059762
transform 1 0 1992 0 1 4610
box -4 -6 52 206
use OAI22X1  _4101_
timestamp 1597059762
transform 1 0 2040 0 1 4610
box -4 -6 84 206
use NOR2X1  _4099_
timestamp 1597059762
transform 1 0 2120 0 1 4610
box -4 -6 52 206
use MUX2X1  _4102_
timestamp 1597059762
transform 1 0 2168 0 1 4610
box -4 -6 100 206
use DFFPOSX1  _4201_
timestamp 1597059762
transform 1 0 2328 0 1 4610
box -4 -6 196 206
use FILL  SFILL22640x46100
timestamp 1597059762
transform 1 0 2264 0 1 4610
box -4 -6 20 206
use FILL  SFILL22800x46100
timestamp 1597059762
transform 1 0 2280 0 1 4610
box -4 -6 20 206
use FILL  SFILL22960x46100
timestamp 1597059762
transform 1 0 2296 0 1 4610
box -4 -6 20 206
use FILL  SFILL23120x46100
timestamp 1597059762
transform 1 0 2312 0 1 4610
box -4 -6 20 206
use NOR2X1  _4121_
timestamp 1597059762
transform -1 0 2568 0 1 4610
box -4 -6 52 206
use OAI22X1  _4123_
timestamp 1597059762
transform 1 0 2568 0 1 4610
box -4 -6 84 206
use OAI21X1  _4122_
timestamp 1597059762
transform -1 0 2712 0 1 4610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert35
timestamp 1597059762
transform 1 0 2712 0 1 4610
box -4 -6 148 206
use NOR2X1  _3742_
timestamp 1597059762
transform 1 0 2856 0 1 4610
box -4 -6 52 206
use AOI21X1  _3743_
timestamp 1597059762
transform -1 0 2968 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4195_
timestamp 1597059762
transform 1 0 2968 0 1 4610
box -4 -6 196 206
use NOR2X1  _4055_
timestamp 1597059762
transform -1 0 3208 0 1 4610
box -4 -6 52 206
use OAI21X1  _4056_
timestamp 1597059762
transform 1 0 3208 0 1 4610
box -4 -6 68 206
use OAI22X1  _4057_
timestamp 1597059762
transform 1 0 3272 0 1 4610
box -4 -6 84 206
use MUX2X1  _4058_
timestamp 1597059762
transform -1 0 3448 0 1 4610
box -4 -6 100 206
use AOI21X1  _4060_
timestamp 1597059762
transform 1 0 3448 0 1 4610
box -4 -6 68 206
use OAI21X1  _4059_
timestamp 1597059762
transform -1 0 3576 0 1 4610
box -4 -6 68 206
use AOI21X1  _4071_
timestamp 1597059762
transform 1 0 3576 0 1 4610
box -4 -6 68 206
use OAI21X1  _4070_
timestamp 1597059762
transform -1 0 3704 0 1 4610
box -4 -6 68 206
use AOI21X1  _4082_
timestamp 1597059762
transform 1 0 3704 0 1 4610
box -4 -6 68 206
use FILL  SFILL37680x46100
timestamp 1597059762
transform 1 0 3768 0 1 4610
box -4 -6 20 206
use FILL  SFILL37840x46100
timestamp 1597059762
transform 1 0 3784 0 1 4610
box -4 -6 20 206
use FILL  SFILL38000x46100
timestamp 1597059762
transform 1 0 3800 0 1 4610
box -4 -6 20 206
use FILL  SFILL38160x46100
timestamp 1597059762
transform 1 0 3816 0 1 4610
box -4 -6 20 206
use OAI21X1  _4081_
timestamp 1597059762
transform -1 0 3896 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4307_
timestamp 1597059762
transform 1 0 3896 0 1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert64
timestamp 1597059762
transform -1 0 4136 0 1 4610
box -4 -6 52 206
use OAI21X1  _3847_
timestamp 1597059762
transform -1 0 4200 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4327_
timestamp 1597059762
transform 1 0 4200 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4309_
timestamp 1597059762
transform 1 0 4392 0 1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert56
timestamp 1597059762
transform 1 0 4584 0 1 4610
box -4 -6 52 206
use XNOR2X1  _2506_
timestamp 1597059762
transform 1 0 4632 0 1 4610
box -4 -6 116 206
use BUFX2  _2046_
timestamp 1597059762
transform -1 0 4792 0 1 4610
box -4 -6 52 206
use AND2X2  _2341_
timestamp 1597059762
transform 1 0 4792 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert116
timestamp 1597059762
transform 1 0 4856 0 1 4610
box -4 -6 52 206
use INVX1  _2670_
timestamp 1597059762
transform 1 0 4904 0 1 4610
box -4 -6 36 206
use NAND2X1  _2671_
timestamp 1597059762
transform -1 0 4984 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert57
timestamp 1597059762
transform 1 0 4984 0 1 4610
box -4 -6 52 206
use INVX1  _2465_
timestamp 1597059762
transform 1 0 5032 0 1 4610
box -4 -6 36 206
use OR2X2  _2475_
timestamp 1597059762
transform -1 0 5128 0 1 4610
box -4 -6 68 206
use AND2X2  _2473_
timestamp 1597059762
transform -1 0 5192 0 1 4610
box -4 -6 68 206
use NOR2X1  _2474_
timestamp 1597059762
transform -1 0 5240 0 1 4610
box -4 -6 52 206
use INVX1  _2479_
timestamp 1597059762
transform 1 0 5240 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert117
timestamp 1597059762
transform 1 0 5336 0 1 4610
box -4 -6 52 206
use NAND2X1  _2612_
timestamp 1597059762
transform 1 0 5384 0 1 4610
box -4 -6 52 206
use FILL  SFILL52720x46100
timestamp 1597059762
transform 1 0 5272 0 1 4610
box -4 -6 20 206
use FILL  SFILL52880x46100
timestamp 1597059762
transform 1 0 5288 0 1 4610
box -4 -6 20 206
use FILL  SFILL53040x46100
timestamp 1597059762
transform 1 0 5304 0 1 4610
box -4 -6 20 206
use FILL  SFILL53200x46100
timestamp 1597059762
transform 1 0 5320 0 1 4610
box -4 -6 20 206
use OR2X2  _2792_
timestamp 1597059762
transform -1 0 5496 0 1 4610
box -4 -6 68 206
use NAND2X1  _2793_
timestamp 1597059762
transform 1 0 5496 0 1 4610
box -4 -6 52 206
use NOR2X1  _2846_
timestamp 1597059762
transform -1 0 5592 0 1 4610
box -4 -6 52 206
use AOI21X1  _2849_
timestamp 1597059762
transform -1 0 5656 0 1 4610
box -4 -6 68 206
use INVX1  _2847_
timestamp 1597059762
transform 1 0 5656 0 1 4610
box -4 -6 36 206
use NOR2X1  _2848_
timestamp 1597059762
transform -1 0 5736 0 1 4610
box -4 -6 52 206
use NAND3X1  _2795_
timestamp 1597059762
transform 1 0 5736 0 1 4610
box -4 -6 68 206
use XNOR2X1  _2794_
timestamp 1597059762
transform -1 0 5912 0 1 4610
box -4 -6 116 206
use INVX1  _2696_
timestamp 1597059762
transform 1 0 5912 0 1 4610
box -4 -6 36 206
use NAND2X1  _2697_
timestamp 1597059762
transform -1 0 5992 0 1 4610
box -4 -6 52 206
use INVX1  _2472_
timestamp 1597059762
transform -1 0 6024 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert159
timestamp 1597059762
transform 1 0 6024 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert216
timestamp 1597059762
transform 1 0 6072 0 1 4610
box -4 -6 52 206
use XNOR2X1  _2356_
timestamp 1597059762
transform -1 0 6232 0 1 4610
box -4 -6 116 206
use NAND2X1  _2358_
timestamp 1597059762
transform 1 0 6232 0 1 4610
box -4 -6 52 206
use XNOR2X1  _2357_
timestamp 1597059762
transform -1 0 6392 0 1 4610
box -4 -6 116 206
use OAI21X1  _2861_
timestamp 1597059762
transform -1 0 6456 0 1 4610
box -4 -6 68 206
use NOR2X1  _2809_
timestamp 1597059762
transform 1 0 6456 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert158
timestamp 1597059762
transform 1 0 6504 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert161
timestamp 1597059762
transform 1 0 6552 0 1 4610
box -4 -6 52 206
use OR2X2  _2704_
timestamp 1597059762
transform 1 0 6600 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert63
timestamp 1597059762
transform 1 0 6664 0 1 4610
box -4 -6 52 206
use AOI22X1  _2706_
timestamp 1597059762
transform -1 0 6792 0 1 4610
box -4 -6 84 206
use FILL  SFILL67920x46100
timestamp 1597059762
transform 1 0 6792 0 1 4610
box -4 -6 20 206
use FILL  SFILL68080x46100
timestamp 1597059762
transform 1 0 6808 0 1 4610
box -4 -6 20 206
use FILL  SFILL68240x46100
timestamp 1597059762
transform 1 0 6824 0 1 4610
box -4 -6 20 206
use OR2X2  _2702_
timestamp 1597059762
transform -1 0 6920 0 1 4610
box -4 -6 68 206
use NAND2X1  _2703_
timestamp 1597059762
transform -1 0 6968 0 1 4610
box -4 -6 52 206
use NOR2X1  _2154_
timestamp 1597059762
transform -1 0 7016 0 1 4610
box -4 -6 52 206
use NAND2X1  _2152_
timestamp 1597059762
transform 1 0 7016 0 1 4610
box -4 -6 52 206
use FILL  SFILL68400x46100
timestamp 1597059762
transform 1 0 6840 0 1 4610
box -4 -6 20 206
use NAND2X1  _2159_
timestamp 1597059762
transform 1 0 7064 0 1 4610
box -4 -6 52 206
use INVX1  _2551_
timestamp 1597059762
transform 1 0 7112 0 1 4610
box -4 -6 36 206
use NOR2X1  _2569_
timestamp 1597059762
transform -1 0 7192 0 1 4610
box -4 -6 52 206
use OAI21X1  _2555_
timestamp 1597059762
transform 1 0 7192 0 1 4610
box -4 -6 68 206
use OAI21X1  _2553_
timestamp 1597059762
transform 1 0 7256 0 1 4610
box -4 -6 68 206
use NAND2X1  _2552_
timestamp 1597059762
transform 1 0 7320 0 1 4610
box -4 -6 52 206
use NOR2X1  _2570_
timestamp 1597059762
transform -1 0 7416 0 1 4610
box -4 -6 52 206
use AOI21X1  _2571_
timestamp 1597059762
transform 1 0 7416 0 1 4610
box -4 -6 68 206
use NOR2X1  _2545_
timestamp 1597059762
transform 1 0 7480 0 1 4610
box -4 -6 52 206
use INVX1  _2102_
timestamp 1597059762
transform 1 0 7528 0 1 4610
box -4 -6 36 206
use DFFPOSX1  _4293_
timestamp 1597059762
transform 1 0 8 0 -1 5010
box -4 -6 196 206
use AOI21X1  _4160_
timestamp 1597059762
transform 1 0 200 0 -1 5010
box -4 -6 68 206
use NOR2X1  _4159_
timestamp 1597059762
transform 1 0 264 0 -1 5010
box -4 -6 52 206
use MUX2X1  _3864_
timestamp 1597059762
transform -1 0 408 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4076_
timestamp 1597059762
transform -1 0 504 0 -1 5010
box -4 -6 100 206
use DFFPOSX1  _4213_
timestamp 1597059762
transform 1 0 504 0 -1 5010
box -4 -6 196 206
use MUX2X1  _4072_
timestamp 1597059762
transform 1 0 696 0 -1 5010
box -4 -6 100 206
use FILL  SFILL7920x48100
timestamp 1597059762
transform -1 0 808 0 -1 5010
box -4 -6 20 206
use FILL  SFILL8080x48100
timestamp 1597059762
transform -1 0 824 0 -1 5010
box -4 -6 20 206
use MUX2X1  _3860_
timestamp 1597059762
transform 1 0 856 0 -1 5010
box -4 -6 100 206
use NAND2X1  _3634_
timestamp 1597059762
transform 1 0 952 0 -1 5010
box -4 -6 52 206
use OAI21X1  _3645_
timestamp 1597059762
transform 1 0 1000 0 -1 5010
box -4 -6 68 206
use FILL  SFILL8240x48100
timestamp 1597059762
transform -1 0 840 0 -1 5010
box -4 -6 20 206
use FILL  SFILL8400x48100
timestamp 1597059762
transform -1 0 856 0 -1 5010
box -4 -6 20 206
use NAND2X1  _3644_
timestamp 1597059762
transform -1 0 1112 0 -1 5010
box -4 -6 52 206
use OAI21X1  _3639_
timestamp 1597059762
transform -1 0 1176 0 -1 5010
box -4 -6 68 206
use NAND2X1  _3638_
timestamp 1597059762
transform -1 0 1224 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4247_
timestamp 1597059762
transform 1 0 1224 0 -1 5010
box -4 -6 196 206
use MUX2X1  _3882_
timestamp 1597059762
transform -1 0 1512 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4094_
timestamp 1597059762
transform -1 0 1608 0 -1 5010
box -4 -6 100 206
use AOI21X1  _4164_
timestamp 1597059762
transform 1 0 1608 0 -1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert72
timestamp 1597059762
transform 1 0 1672 0 -1 5010
box -4 -6 52 206
use NOR2X1  _4163_
timestamp 1597059762
transform -1 0 1768 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4295_
timestamp 1597059762
transform 1 0 1768 0 -1 5010
box -4 -6 196 206
use MUX2X1  _3886_
timestamp 1597059762
transform 1 0 1960 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4098_
timestamp 1597059762
transform 1 0 2056 0 -1 5010
box -4 -6 100 206
use CLKBUF1  CLKBUF1_insert22
timestamp 1597059762
transform -1 0 2296 0 -1 5010
box -4 -6 148 206
use MUX2X1  _3908_
timestamp 1597059762
transform 1 0 2360 0 -1 5010
box -4 -6 100 206
use FILL  SFILL22960x48100
timestamp 1597059762
transform -1 0 2312 0 -1 5010
box -4 -6 20 206
use FILL  SFILL23120x48100
timestamp 1597059762
transform -1 0 2328 0 -1 5010
box -4 -6 20 206
use FILL  SFILL23280x48100
timestamp 1597059762
transform -1 0 2344 0 -1 5010
box -4 -6 20 206
use FILL  SFILL23440x48100
timestamp 1597059762
transform -1 0 2360 0 -1 5010
box -4 -6 20 206
use NOR2X1  _4167_
timestamp 1597059762
transform 1 0 2456 0 -1 5010
box -4 -6 52 206
use MUX2X1  _4120_
timestamp 1597059762
transform -1 0 2600 0 -1 5010
box -4 -6 100 206
use AOI21X1  _3676_
timestamp 1597059762
transform 1 0 2600 0 -1 5010
box -4 -6 68 206
use NOR2X1  _3675_
timestamp 1597059762
transform -1 0 2712 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4224_
timestamp 1597059762
transform 1 0 2712 0 -1 5010
box -4 -6 196 206
use AOI21X1  _3725_
timestamp 1597059762
transform 1 0 2904 0 -1 5010
box -4 -6 68 206
use NOR2X1  _3724_
timestamp 1597059762
transform -1 0 3016 0 -1 5010
box -4 -6 52 206
use AOI21X1  _4150_
timestamp 1597059762
transform 1 0 3016 0 -1 5010
box -4 -6 68 206
use NOR2X1  _4149_
timestamp 1597059762
transform -1 0 3128 0 -1 5010
box -4 -6 52 206
use MUX2X1  _4021_
timestamp 1597059762
transform 1 0 3128 0 -1 5010
box -4 -6 100 206
use MUX2X1  _3809_
timestamp 1597059762
transform 1 0 3224 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4054_
timestamp 1597059762
transform -1 0 3416 0 -1 5010
box -4 -6 100 206
use MUX2X1  _3842_
timestamp 1597059762
transform -1 0 3512 0 -1 5010
box -4 -6 100 206
use NOR2X1  _3938_
timestamp 1597059762
transform 1 0 3512 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3939_
timestamp 1597059762
transform -1 0 3624 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4272_
timestamp 1597059762
transform -1 0 3816 0 -1 5010
box -4 -6 196 206
use FILL  SFILL38160x48100
timestamp 1597059762
transform -1 0 3832 0 -1 5010
box -4 -6 20 206
use BUFX2  BUFX2_insert271
timestamp 1597059762
transform 1 0 3880 0 -1 5010
box -4 -6 52 206
use AOI21X1  _4104_
timestamp 1597059762
transform 1 0 3928 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4103_
timestamp 1597059762
transform -1 0 4056 0 -1 5010
box -4 -6 68 206
use FILL  SFILL38320x48100
timestamp 1597059762
transform -1 0 3848 0 -1 5010
box -4 -6 20 206
use FILL  SFILL38480x48100
timestamp 1597059762
transform -1 0 3864 0 -1 5010
box -4 -6 20 206
use FILL  SFILL38640x48100
timestamp 1597059762
transform -1 0 3880 0 -1 5010
box -4 -6 20 206
use AOI21X1  _3870_
timestamp 1597059762
transform 1 0 4056 0 -1 5010
box -4 -6 68 206
use OAI21X1  _3869_
timestamp 1597059762
transform -1 0 4184 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4311_
timestamp 1597059762
transform 1 0 4184 0 -1 5010
box -4 -6 196 206
use DFFPOSX1  _4323_
timestamp 1597059762
transform 1 0 4376 0 -1 5010
box -4 -6 196 206
use DFFPOSX1  _4324_
timestamp 1597059762
transform 1 0 4568 0 -1 5010
box -4 -6 196 206
use OAI21X1  _2512_
timestamp 1597059762
transform -1 0 4824 0 -1 5010
box -4 -6 68 206
use AOI21X1  _2505_
timestamp 1597059762
transform -1 0 4888 0 -1 5010
box -4 -6 68 206
use XNOR2X1  _2502_
timestamp 1597059762
transform 1 0 4888 0 -1 5010
box -4 -6 116 206
use NOR2X1  _2503_
timestamp 1597059762
transform -1 0 5048 0 -1 5010
box -4 -6 52 206
use XNOR2X1  _2487_
timestamp 1597059762
transform -1 0 5160 0 -1 5010
box -4 -6 116 206
use INVX1  _2510_
timestamp 1597059762
transform 1 0 5160 0 -1 5010
box -4 -6 36 206
use AOI21X1  _2511_
timestamp 1597059762
transform -1 0 5256 0 -1 5010
box -4 -6 68 206
use AND2X2  _2495_
timestamp 1597059762
transform 1 0 5320 0 -1 5010
box -4 -6 68 206
use XNOR2X1  _2476_
timestamp 1597059762
transform 1 0 5384 0 -1 5010
box -4 -6 116 206
use FILL  SFILL52560x48100
timestamp 1597059762
transform -1 0 5272 0 -1 5010
box -4 -6 20 206
use FILL  SFILL52720x48100
timestamp 1597059762
transform -1 0 5288 0 -1 5010
box -4 -6 20 206
use FILL  SFILL52880x48100
timestamp 1597059762
transform -1 0 5304 0 -1 5010
box -4 -6 20 206
use FILL  SFILL53040x48100
timestamp 1597059762
transform -1 0 5320 0 -1 5010
box -4 -6 20 206
use OAI21X1  _2480_
timestamp 1597059762
transform 1 0 5496 0 -1 5010
box -4 -6 68 206
use NOR2X1  _2477_
timestamp 1597059762
transform -1 0 5608 0 -1 5010
box -4 -6 52 206
use AOI21X1  _2481_
timestamp 1597059762
transform -1 0 5672 0 -1 5010
box -4 -6 68 206
use AND2X2  _2493_
timestamp 1597059762
transform -1 0 5736 0 -1 5010
box -4 -6 68 206
use OAI21X1  _2482_
timestamp 1597059762
transform -1 0 5800 0 -1 5010
box -4 -6 68 206
use NAND2X1  _2478_
timestamp 1597059762
transform -1 0 5848 0 -1 5010
box -4 -6 52 206
use XNOR2X1  _2452_
timestamp 1597059762
transform 1 0 5848 0 -1 5010
box -4 -6 116 206
use XNOR2X1  _2458_
timestamp 1597059762
transform 1 0 5960 0 -1 5010
box -4 -6 116 206
use INVX1  _2451_
timestamp 1597059762
transform -1 0 6104 0 -1 5010
box -4 -6 36 206
use NOR2X1  _2456_
timestamp 1597059762
transform 1 0 6104 0 -1 5010
box -4 -6 52 206
use AND2X2  _2455_
timestamp 1597059762
transform -1 0 6216 0 -1 5010
box -4 -6 68 206
use INVX1  _2454_
timestamp 1597059762
transform -1 0 6248 0 -1 5010
box -4 -6 36 206
use NOR2X1  _2324_
timestamp 1597059762
transform 1 0 6248 0 -1 5010
box -4 -6 52 206
use OAI22X1  _2326_
timestamp 1597059762
transform -1 0 6376 0 -1 5010
box -4 -6 84 206
use AND2X2  _2325_
timestamp 1597059762
transform -1 0 6440 0 -1 5010
box -4 -6 68 206
use INVX1  _2797_
timestamp 1597059762
transform 1 0 6440 0 -1 5010
box -4 -6 36 206
use OR2X2  _2798_
timestamp 1597059762
transform 1 0 6472 0 -1 5010
box -4 -6 68 206
use NAND3X1  _2801_
timestamp 1597059762
transform 1 0 6536 0 -1 5010
box -4 -6 68 206
use NAND2X1  _2799_
timestamp 1597059762
transform -1 0 6648 0 -1 5010
box -4 -6 52 206
use NOR2X1  _2855_
timestamp 1597059762
transform -1 0 6696 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert65
timestamp 1597059762
transform -1 0 6744 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert62
timestamp 1597059762
transform 1 0 6808 0 -1 5010
box -4 -6 52 206
use FILL  SFILL67440x48100
timestamp 1597059762
transform -1 0 6760 0 -1 5010
box -4 -6 20 206
use FILL  SFILL67600x48100
timestamp 1597059762
transform -1 0 6776 0 -1 5010
box -4 -6 20 206
use FILL  SFILL67760x48100
timestamp 1597059762
transform -1 0 6792 0 -1 5010
box -4 -6 20 206
use FILL  SFILL67920x48100
timestamp 1597059762
transform -1 0 6808 0 -1 5010
box -4 -6 20 206
use NAND2X1  _2705_
timestamp 1597059762
transform -1 0 6904 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert44
timestamp 1597059762
transform 1 0 6904 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert43
timestamp 1597059762
transform 1 0 6952 0 -1 5010
box -4 -6 52 206
use OR2X2  _2616_
timestamp 1597059762
transform 1 0 7000 0 -1 5010
box -4 -6 68 206
use NAND2X1  _2617_
timestamp 1597059762
transform -1 0 7112 0 -1 5010
box -4 -6 52 206
use INVX1  _2550_
timestamp 1597059762
transform 1 0 7112 0 -1 5010
box -4 -6 36 206
use AOI21X1  _2618_
timestamp 1597059762
transform 1 0 7144 0 -1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert217
timestamp 1597059762
transform 1 0 7208 0 -1 5010
box -4 -6 52 206
use NAND2X1  _2554_
timestamp 1597059762
transform -1 0 7304 0 -1 5010
box -4 -6 52 206
use XOR2X1  _2615_
timestamp 1597059762
transform -1 0 7416 0 -1 5010
box -4 -6 116 206
use BUFX2  _2033_
timestamp 1597059762
transform -1 0 7464 0 -1 5010
box -4 -6 52 206
use INVX1  _2575_
timestamp 1597059762
transform -1 0 7496 0 -1 5010
box -4 -6 36 206
use OAI21X1  _2866_
timestamp 1597059762
transform 1 0 7496 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4277_
timestamp 1597059762
transform 1 0 8 0 1 5010
box -4 -6 196 206
use AOI21X1  _3949_
timestamp 1597059762
transform 1 0 200 0 1 5010
box -4 -6 68 206
use NOR2X1  _3948_
timestamp 1597059762
transform -1 0 312 0 1 5010
box -4 -6 52 206
use NOR2X1  _3958_
timestamp 1597059762
transform -1 0 360 0 1 5010
box -4 -6 52 206
use AOI21X1  _3959_
timestamp 1597059762
transform -1 0 424 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4282_
timestamp 1597059762
transform 1 0 424 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4261_
timestamp 1597059762
transform -1 0 808 0 1 5010
box -4 -6 196 206
use FILL  SFILL8080x50100
timestamp 1597059762
transform 1 0 808 0 1 5010
box -4 -6 20 206
use AOI21X1  _3668_
timestamp 1597059762
transform 1 0 872 0 1 5010
box -4 -6 68 206
use NOR2X1  _3667_
timestamp 1597059762
transform 1 0 936 0 1 5010
box -4 -6 52 206
use OAI21X1  _3635_
timestamp 1597059762
transform -1 0 1048 0 1 5010
box -4 -6 68 206
use FILL  SFILL8240x50100
timestamp 1597059762
transform 1 0 824 0 1 5010
box -4 -6 20 206
use FILL  SFILL8400x50100
timestamp 1597059762
transform 1 0 840 0 1 5010
box -4 -6 20 206
use FILL  SFILL8560x50100
timestamp 1597059762
transform 1 0 856 0 1 5010
box -4 -6 20 206
use DFFPOSX1  _4245_
timestamp 1597059762
transform 1 0 1048 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4250_
timestamp 1597059762
transform 1 0 1240 0 1 5010
box -4 -6 196 206
use NOR2X1  _3677_
timestamp 1597059762
transform 1 0 1432 0 1 5010
box -4 -6 52 206
use AOI21X1  _3678_
timestamp 1597059762
transform -1 0 1544 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4266_
timestamp 1597059762
transform -1 0 1736 0 1 5010
box -4 -6 196 206
use NOR2X1  _3671_
timestamp 1597059762
transform -1 0 1784 0 1 5010
box -4 -6 52 206
use AOI21X1  _3672_
timestamp 1597059762
transform 1 0 1784 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4263_
timestamp 1597059762
transform -1 0 2040 0 1 5010
box -4 -6 196 206
use AOI21X1  _3953_
timestamp 1597059762
transform 1 0 2040 0 1 5010
box -4 -6 68 206
use NOR2X1  _3952_
timestamp 1597059762
transform 1 0 2104 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4279_
timestamp 1597059762
transform -1 0 2344 0 1 5010
box -4 -6 196 206
use NOR2X1  _3956_
timestamp 1597059762
transform -1 0 2456 0 1 5010
box -4 -6 52 206
use FILL  SFILL23440x50100
timestamp 1597059762
transform 1 0 2344 0 1 5010
box -4 -6 20 206
use FILL  SFILL23600x50100
timestamp 1597059762
transform 1 0 2360 0 1 5010
box -4 -6 20 206
use FILL  SFILL23760x50100
timestamp 1597059762
transform 1 0 2376 0 1 5010
box -4 -6 20 206
use FILL  SFILL23920x50100
timestamp 1597059762
transform 1 0 2392 0 1 5010
box -4 -6 20 206
use AOI21X1  _3957_
timestamp 1597059762
transform -1 0 2520 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4281_
timestamp 1597059762
transform 1 0 2520 0 1 5010
box -4 -6 196 206
use AOI21X1  _4168_
timestamp 1597059762
transform -1 0 2776 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4297_
timestamp 1597059762
transform -1 0 2968 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4265_
timestamp 1597059762
transform -1 0 3160 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4288_
timestamp 1597059762
transform 1 0 3160 0 1 5010
box -4 -6 196 206
use NOR2X1  _4155_
timestamp 1597059762
transform -1 0 3400 0 1 5010
box -4 -6 52 206
use AOI21X1  _4156_
timestamp 1597059762
transform -1 0 3464 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4291_
timestamp 1597059762
transform -1 0 3656 0 1 5010
box -4 -6 196 206
use AOI21X1  _3945_
timestamp 1597059762
transform 1 0 3656 0 1 5010
box -4 -6 68 206
use NOR2X1  _3944_
timestamp 1597059762
transform -1 0 3768 0 1 5010
box -4 -6 52 206
use FILL  SFILL37680x50100
timestamp 1597059762
transform 1 0 3768 0 1 5010
box -4 -6 20 206
use FILL  SFILL37840x50100
timestamp 1597059762
transform 1 0 3784 0 1 5010
box -4 -6 20 206
use FILL  SFILL38000x50100
timestamp 1597059762
transform 1 0 3800 0 1 5010
box -4 -6 20 206
use FILL  SFILL38160x50100
timestamp 1597059762
transform 1 0 3816 0 1 5010
box -4 -6 20 206
use DFFPOSX1  _4275_
timestamp 1597059762
transform -1 0 4024 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4308_
timestamp 1597059762
transform 1 0 4024 0 1 5010
box -4 -6 196 206
use BUFX2  _2040_
timestamp 1597059762
transform -1 0 4264 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4325_
timestamp 1597059762
transform 1 0 4264 0 1 5010
box -4 -6 196 206
use BUFX2  _2042_
timestamp 1597059762
transform -1 0 4504 0 1 5010
box -4 -6 52 206
use BUFX2  _2047_
timestamp 1597059762
transform -1 0 4552 0 1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert42
timestamp 1597059762
transform -1 0 4600 0 1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert12
timestamp 1597059762
transform -1 0 4648 0 1 5010
box -4 -6 52 206
use BUFX2  _2045_
timestamp 1597059762
transform 1 0 4648 0 1 5010
box -4 -6 52 206
use INVX1  _2497_
timestamp 1597059762
transform 1 0 4696 0 1 5010
box -4 -6 36 206
use NAND2X1  _2500_
timestamp 1597059762
transform -1 0 4776 0 1 5010
box -4 -6 52 206
use NOR2X1  _2498_
timestamp 1597059762
transform -1 0 4824 0 1 5010
box -4 -6 52 206
use OAI21X1  _2504_
timestamp 1597059762
transform -1 0 4888 0 1 5010
box -4 -6 68 206
use INVX1  _2499_
timestamp 1597059762
transform 1 0 4888 0 1 5010
box -4 -6 36 206
use NAND2X1  _2501_
timestamp 1597059762
transform 1 0 4920 0 1 5010
box -4 -6 52 206
use OAI21X1  _2496_
timestamp 1597059762
transform -1 0 5032 0 1 5010
box -4 -6 68 206
use NAND2X1  _2486_
timestamp 1597059762
transform -1 0 5080 0 1 5010
box -4 -6 52 206
use OR2X2  _2485_
timestamp 1597059762
transform -1 0 5144 0 1 5010
box -4 -6 68 206
use NAND2X1  _2484_
timestamp 1597059762
transform -1 0 5192 0 1 5010
box -4 -6 52 206
use INVX1  _2483_
timestamp 1597059762
transform -1 0 5224 0 1 5010
box -4 -6 36 206
use BUFX2  _2044_
timestamp 1597059762
transform 1 0 5224 0 1 5010
box -4 -6 52 206
use NAND2X1  _2467_
timestamp 1597059762
transform 1 0 5336 0 1 5010
box -4 -6 52 206
use OAI21X1  _2471_
timestamp 1597059762
transform 1 0 5384 0 1 5010
box -4 -6 68 206
use FILL  SFILL52720x50100
timestamp 1597059762
transform 1 0 5272 0 1 5010
box -4 -6 20 206
use FILL  SFILL52880x50100
timestamp 1597059762
transform 1 0 5288 0 1 5010
box -4 -6 20 206
use FILL  SFILL53040x50100
timestamp 1597059762
transform 1 0 5304 0 1 5010
box -4 -6 20 206
use FILL  SFILL53200x50100
timestamp 1597059762
transform 1 0 5320 0 1 5010
box -4 -6 20 206
use OR2X2  _2466_
timestamp 1597059762
transform 1 0 5448 0 1 5010
box -4 -6 68 206
use NAND3X1  _2470_
timestamp 1597059762
transform 1 0 5512 0 1 5010
box -4 -6 68 206
use NAND2X1  _2468_
timestamp 1597059762
transform 1 0 5576 0 1 5010
box -4 -6 52 206
use XNOR2X1  _2469_
timestamp 1597059762
transform -1 0 5736 0 1 5010
box -4 -6 116 206
use INVX1  _2461_
timestamp 1597059762
transform 1 0 5736 0 1 5010
box -4 -6 36 206
use OAI21X1  _2464_
timestamp 1597059762
transform -1 0 5832 0 1 5010
box -4 -6 68 206
use INVX1  _2463_
timestamp 1597059762
transform -1 0 5864 0 1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert66
timestamp 1597059762
transform -1 0 5912 0 1 5010
box -4 -6 52 206
use NOR2X1  _2462_
timestamp 1597059762
transform -1 0 5960 0 1 5010
box -4 -6 52 206
use OAI21X1  _2453_
timestamp 1597059762
transform 1 0 5960 0 1 5010
box -4 -6 68 206
use OAI21X1  _2460_
timestamp 1597059762
transform -1 0 6088 0 1 5010
box -4 -6 68 206
use OR2X2  _2457_
timestamp 1597059762
transform -1 0 6152 0 1 5010
box -4 -6 68 206
use INVX1  _2459_
timestamp 1597059762
transform -1 0 6184 0 1 5010
box -4 -6 36 206
use NAND2X1  _2450_
timestamp 1597059762
transform -1 0 6232 0 1 5010
box -4 -6 52 206
use OR2X2  _2448_
timestamp 1597059762
transform -1 0 6296 0 1 5010
box -4 -6 68 206
use NAND2X1  _2449_
timestamp 1597059762
transform -1 0 6344 0 1 5010
box -4 -6 52 206
use INVX1  _2447_
timestamp 1597059762
transform -1 0 6376 0 1 5010
box -4 -6 36 206
use NOR2X1  _2322_
timestamp 1597059762
transform 1 0 6376 0 1 5010
box -4 -6 52 206
use AND2X2  _2323_
timestamp 1597059762
transform -1 0 6488 0 1 5010
box -4 -6 68 206
use XNOR2X1  _2800_
timestamp 1597059762
transform -1 0 6600 0 1 5010
box -4 -6 116 206
use AOI21X1  _2858_
timestamp 1597059762
transform 1 0 6600 0 1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert41
timestamp 1597059762
transform -1 0 6712 0 1 5010
box -4 -6 52 206
use INVX1  _2856_
timestamp 1597059762
transform 1 0 6712 0 1 5010
box -4 -6 36 206
use NOR2X1  _2857_
timestamp 1597059762
transform -1 0 6856 0 1 5010
box -4 -6 52 206
use FILL  SFILL67440x50100
timestamp 1597059762
transform 1 0 6744 0 1 5010
box -4 -6 20 206
use FILL  SFILL67600x50100
timestamp 1597059762
transform 1 0 6760 0 1 5010
box -4 -6 20 206
use FILL  SFILL67760x50100
timestamp 1597059762
transform 1 0 6776 0 1 5010
box -4 -6 20 206
use FILL  SFILL67920x50100
timestamp 1597059762
transform 1 0 6792 0 1 5010
box -4 -6 20 206
use NOR2X1  _2772_
timestamp 1597059762
transform 1 0 6856 0 1 5010
box -4 -6 52 206
use INVX1  _2771_
timestamp 1597059762
transform -1 0 6936 0 1 5010
box -4 -6 36 206
use AOI21X1  _2774_
timestamp 1597059762
transform 1 0 6936 0 1 5010
box -4 -6 68 206
use NOR2X1  _2773_
timestamp 1597059762
transform 1 0 7000 0 1 5010
box -4 -6 52 206
use NAND2X1  _2770_
timestamp 1597059762
transform -1 0 7096 0 1 5010
box -4 -6 52 206
use INVX1  _2681_
timestamp 1597059762
transform 1 0 7096 0 1 5010
box -4 -6 36 206
use NOR2X1  _2682_
timestamp 1597059762
transform 1 0 7128 0 1 5010
box -4 -6 52 206
use INVX1  _2769_
timestamp 1597059762
transform -1 0 7208 0 1 5010
box -4 -6 36 206
use AOI21X1  _2684_
timestamp 1597059762
transform 1 0 7208 0 1 5010
box -4 -6 68 206
use NOR2X1  _2683_
timestamp 1597059762
transform 1 0 7272 0 1 5010
box -4 -6 52 206
use NAND2X1  _2680_
timestamp 1597059762
transform 1 0 7320 0 1 5010
box -4 -6 52 206
use INVX1  _2679_
timestamp 1597059762
transform -1 0 7400 0 1 5010
box -4 -6 36 206
use AOI21X1  _2590_
timestamp 1597059762
transform -1 0 7464 0 1 5010
box -4 -6 68 206
use BUFX2  _2041_
timestamp 1597059762
transform -1 0 7512 0 1 5010
box -4 -6 52 206
use NOR2X1  _2103_
timestamp 1597059762
transform 1 0 7512 0 1 5010
box -4 -6 52 206
<< labels >>
flabel metal4 s 2240 -10 2304 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 736 -10 800 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 3245 -23 3251 -17 7 FreeSans 24 270 0 0 adrs_bus[15]
port 2 nsew
flabel metal2 s 3629 -23 3635 -17 7 FreeSans 24 270 0 0 adrs_bus[14]
port 3 nsew
flabel metal2 s 3293 -23 3299 -17 7 FreeSans 24 270 0 0 adrs_bus[13]
port 4 nsew
flabel metal2 s 5709 -23 5715 -17 7 FreeSans 24 270 0 0 adrs_bus[12]
port 5 nsew
flabel metal2 s 3581 -23 3587 -17 7 FreeSans 24 270 0 0 adrs_bus[11]
port 6 nsew
flabel metal2 s 4029 -23 4035 -17 7 FreeSans 24 270 0 0 adrs_bus[10]
port 7 nsew
flabel metal2 s 4077 -23 4083 -17 7 FreeSans 24 270 0 0 adrs_bus[9]
port 8 nsew
flabel metal2 s 4909 -23 4915 -17 7 FreeSans 24 270 0 0 adrs_bus[8]
port 9 nsew
flabel metal2 s 6349 -23 6355 -17 7 FreeSans 24 270 0 0 adrs_bus[7]
port 10 nsew
flabel metal2 s 5997 -23 6003 -17 7 FreeSans 24 270 0 0 adrs_bus[6]
port 11 nsew
flabel metal2 s 6397 -23 6403 -17 7 FreeSans 24 270 0 0 adrs_bus[5]
port 12 nsew
flabel metal2 s 6077 -23 6083 -17 7 FreeSans 24 270 0 0 adrs_bus[4]
port 13 nsew
flabel metal2 s 5741 -23 5747 -17 7 FreeSans 24 270 0 0 adrs_bus[3]
port 14 nsew
flabel metal2 s 5677 -23 5683 -17 7 FreeSans 24 270 0 0 adrs_bus[2]
port 15 nsew
flabel metal2 s 5773 -23 5779 -17 7 FreeSans 24 270 0 0 adrs_bus[1]
port 16 nsew
flabel metal2 s 5821 -23 5827 -17 7 FreeSans 24 270 0 0 adrs_bus[0]
port 17 nsew
flabel metal3 s -35 3477 -29 3483 7 FreeSans 24 0 0 0 clock
port 18 nsew
flabel metal2 s 989 -23 995 -17 7 FreeSans 24 270 0 0 data_in[15]
port 19 nsew
flabel metal2 s 1261 -23 1267 -17 7 FreeSans 24 270 0 0 data_in[14]
port 20 nsew
flabel metal2 s 685 -23 691 -17 7 FreeSans 24 270 0 0 data_in[13]
port 21 nsew
flabel metal2 s 1037 -23 1043 -17 7 FreeSans 24 270 0 0 data_in[12]
port 22 nsew
flabel metal3 s -35 957 -29 963 7 FreeSans 24 0 0 0 data_in[11]
port 23 nsew
flabel metal3 s -35 997 -29 1003 7 FreeSans 24 0 0 0 data_in[10]
port 24 nsew
flabel metal2 s 829 -23 835 -17 7 FreeSans 24 270 0 0 data_in[9]
port 25 nsew
flabel metal2 s 1677 -23 1683 -17 7 FreeSans 24 270 0 0 data_in[8]
port 26 nsew
flabel metal2 s 253 -23 259 -17 7 FreeSans 24 270 0 0 data_in[7]
port 27 nsew
flabel metal2 s 1165 -23 1171 -17 7 FreeSans 24 270 0 0 data_in[6]
port 28 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 data_in[5]
port 29 nsew
flabel metal3 s -35 917 -29 923 7 FreeSans 24 0 0 0 data_in[4]
port 30 nsew
flabel metal2 s 1645 -23 1651 -17 7 FreeSans 24 270 0 0 data_in[3]
port 31 nsew
flabel metal2 s 861 -23 867 -17 7 FreeSans 24 270 0 0 data_in[2]
port 32 nsew
flabel metal2 s 1213 -23 1219 -17 7 FreeSans 24 270 0 0 data_in[1]
port 33 nsew
flabel metal2 s 1597 -23 1603 -17 7 FreeSans 24 270 0 0 data_in[0]
port 34 nsew
flabel metal2 s 4525 5257 4531 5263 3 FreeSans 24 90 0 0 data_out[15]
port 35 nsew
flabel metal2 s 4765 5257 4771 5263 3 FreeSans 24 90 0 0 data_out[14]
port 36 nsew
flabel metal2 s 4669 5257 4675 5263 3 FreeSans 24 90 0 0 data_out[13]
port 37 nsew
flabel metal2 s 5341 5257 5347 5263 3 FreeSans 24 90 0 0 data_out[12]
port 38 nsew
flabel metal3 s 7597 3897 7603 3903 3 FreeSans 24 0 0 0 data_out[11]
port 39 nsew
flabel metal2 s 4477 5257 4483 5263 3 FreeSans 24 90 0 0 data_out[10]
port 40 nsew
flabel metal2 s 7485 5257 7491 5263 3 FreeSans 24 90 0 0 data_out[9]
port 41 nsew
flabel metal2 s 4237 5257 4243 5263 3 FreeSans 24 90 0 0 data_out[8]
port 42 nsew
flabel metal2 s 7181 -23 7187 -17 7 FreeSans 24 270 0 0 data_out[7]
port 43 nsew
flabel metal3 s 7597 1297 7603 1303 3 FreeSans 24 0 0 0 data_out[6]
port 44 nsew
flabel metal2 s 6445 -23 6451 -17 7 FreeSans 24 270 0 0 data_out[5]
port 45 nsew
flabel metal2 s 6605 -23 6611 -17 7 FreeSans 24 270 0 0 data_out[4]
port 46 nsew
flabel metal3 s 7597 2297 7603 2303 3 FreeSans 24 0 0 0 data_out[3]
port 47 nsew
flabel metal3 s 7597 1497 7603 1503 3 FreeSans 24 0 0 0 data_out[2]
port 48 nsew
flabel metal3 s 7597 3677 7603 3683 3 FreeSans 24 0 0 0 data_out[1]
port 49 nsew
flabel metal3 s 7597 3717 7603 3723 3 FreeSans 24 0 0 0 data_out[0]
port 50 nsew
flabel metal2 s 1565 -23 1571 -17 7 FreeSans 24 270 0 0 mem_rd
port 51 nsew
flabel metal2 s 2525 -23 2531 -17 7 FreeSans 24 270 0 0 mem_wr
port 52 nsew
flabel metal2 s 3885 5257 3891 5263 3 FreeSans 24 90 0 0 reset
port 53 nsew
<< end >>
