magic
tech scmos
magscale 1 2
timestamp 1591628762
<< metal1 >>
rect 1754 1414 1766 1416
rect 1739 1406 1741 1414
rect 1749 1406 1751 1414
rect 1759 1406 1761 1414
rect 1769 1406 1771 1414
rect 1779 1406 1781 1414
rect 1754 1404 1766 1406
rect 1789 1377 1804 1383
rect 1116 1337 1140 1343
rect 1405 1337 1443 1343
rect 1485 1337 1500 1343
rect 1517 1337 1555 1343
rect 404 1317 419 1323
rect 676 1317 707 1323
rect 1236 1317 1251 1323
rect 1444 1317 1459 1323
rect 1581 1317 1596 1323
rect 1812 1317 1875 1323
rect 2381 1277 2396 1283
rect 618 1214 630 1216
rect 603 1206 605 1214
rect 613 1206 615 1214
rect 623 1206 625 1214
rect 633 1206 635 1214
rect 643 1206 645 1214
rect 618 1204 630 1206
rect 394 1176 396 1184
rect 1188 1176 1190 1184
rect 1418 1176 1420 1184
rect 852 1116 860 1124
rect 916 1116 924 1124
rect 1012 1116 1020 1124
rect 1277 1117 1292 1123
rect 1716 1117 1795 1123
rect 1805 1117 1843 1123
rect 1860 1116 1868 1124
rect 317 1097 332 1103
rect 349 1097 364 1103
rect 413 1097 435 1103
rect 138 1076 140 1084
rect 308 1077 339 1083
rect 413 1077 419 1097
rect 692 1097 771 1103
rect 973 1097 1004 1103
rect 1172 1097 1187 1103
rect 1341 1103 1347 1116
rect 1309 1097 1347 1103
rect 692 1077 755 1083
rect 813 1077 828 1083
rect 1085 1083 1091 1096
rect 2365 1097 2380 1103
rect 1069 1077 1091 1083
rect 1444 1077 1459 1083
rect 1476 1077 1507 1083
rect 1533 1077 1564 1083
rect 2004 1076 2006 1084
rect 2317 1077 2332 1083
rect 1469 1057 1475 1076
rect 1700 1057 1772 1063
rect 1754 1014 1766 1016
rect 1739 1006 1741 1014
rect 1749 1006 1751 1014
rect 1759 1006 1761 1014
rect 1769 1006 1771 1014
rect 1779 1006 1781 1014
rect 1754 1004 1766 1006
rect 605 977 668 983
rect 2365 957 2396 963
rect 628 937 691 943
rect 724 937 739 943
rect 781 937 796 943
rect 1085 937 1100 943
rect 1133 937 1148 943
rect 1485 937 1500 943
rect 1796 937 1811 943
rect 244 917 275 923
rect 285 917 300 923
rect 701 917 739 923
rect 765 917 796 923
rect 221 897 259 903
rect 605 897 684 903
rect 733 897 739 917
rect 861 917 924 923
rect 1085 917 1123 923
rect 1421 917 1436 923
rect 1085 897 1091 917
rect 1485 917 1523 923
rect 1485 897 1491 917
rect 1652 917 1667 923
rect 1796 917 1827 923
rect 1837 917 1852 923
rect 2100 877 2115 883
rect 618 814 630 816
rect 603 806 605 814
rect 613 806 615 814
rect 623 806 625 814
rect 633 806 635 814
rect 643 806 645 814
rect 618 804 630 806
rect 282 776 284 784
rect 2020 736 2022 744
rect 573 717 611 723
rect 676 717 691 723
rect 708 716 716 724
rect 772 716 780 724
rect 388 697 467 703
rect 605 697 636 703
rect 740 697 771 703
rect 941 703 947 723
rect 941 697 979 703
rect 1405 703 1411 723
rect 1405 697 1443 703
rect 1469 684 1475 703
rect 1533 697 1548 703
rect 2093 703 2099 723
rect 2093 697 2108 703
rect 301 677 323 683
rect 404 677 435 683
rect 333 657 355 663
rect 429 657 435 677
rect 861 677 876 683
rect 1341 677 1356 683
rect 1453 677 1468 683
rect 1677 677 1740 683
rect 1932 677 1955 683
rect 1932 672 1940 677
rect 2116 677 2131 683
rect 482 637 524 643
rect 1754 614 1766 616
rect 1739 606 1741 614
rect 1749 606 1751 614
rect 1759 606 1761 614
rect 1769 606 1771 614
rect 1779 606 1781 614
rect 1754 604 1766 606
rect 1741 577 1804 583
rect 1898 576 1900 584
rect 1972 556 1980 564
rect 77 537 108 543
rect 317 537 332 543
rect 125 517 179 523
rect 317 517 323 537
rect 1276 537 1300 543
rect 1844 537 1859 543
rect 349 517 387 523
rect 381 497 387 517
rect 644 517 707 523
rect 813 517 828 523
rect 1357 517 1388 523
rect 1853 517 1859 537
rect 1981 537 1996 543
rect 1924 517 1939 523
rect 404 496 412 504
rect 2084 497 2099 503
rect 2132 456 2134 464
rect 618 414 630 416
rect 603 406 605 414
rect 613 406 615 414
rect 623 406 625 414
rect 633 406 635 414
rect 643 406 645 414
rect 618 404 630 406
rect 1050 376 1052 384
rect 2004 336 2006 344
rect 2196 337 2211 343
rect 253 303 259 323
rect 349 317 371 323
rect 221 297 259 303
rect 285 297 316 303
rect 813 303 819 323
rect 1652 317 1667 323
rect 788 297 819 303
rect 852 297 867 303
rect 1556 297 1571 303
rect 1988 297 2003 303
rect 2036 297 2060 303
rect 2093 303 2099 323
rect 2093 297 2131 303
rect 692 277 755 283
rect 1156 277 1171 283
rect 1181 277 1212 283
rect 1229 277 1283 283
rect 1389 277 1427 283
rect 1725 277 1804 283
rect 2093 277 2108 283
rect 2141 277 2156 283
rect 1741 257 1820 263
rect 1828 257 1843 263
rect 1853 257 1868 263
rect 1876 257 1891 263
rect 340 236 342 244
rect 1754 214 1766 216
rect 1739 206 1741 214
rect 1749 206 1751 214
rect 1759 206 1761 214
rect 1769 206 1771 214
rect 1779 206 1781 214
rect 1754 204 1766 206
rect 276 176 278 184
rect 1812 177 1859 183
rect 333 143 339 163
rect 948 157 963 163
rect 1076 157 1091 163
rect 308 137 339 143
rect 525 137 547 143
rect 612 137 691 143
rect 1396 137 1411 143
rect 1453 137 1475 143
rect 1869 137 1884 143
rect 1981 137 2019 143
rect 573 117 668 123
rect 909 117 940 123
rect 1092 117 1107 123
rect 1373 117 1411 123
rect 1437 117 1452 123
rect 589 97 604 103
rect 1405 97 1411 117
rect 1876 117 1907 123
rect 1933 117 1948 123
rect 1933 97 1939 117
rect 2068 117 2099 123
rect 618 14 630 16
rect 603 6 605 14
rect 613 6 615 14
rect 623 6 625 14
rect 633 6 635 14
rect 643 6 645 14
rect 618 4 630 6
<< m2contact >>
rect 1731 1406 1739 1414
rect 1741 1406 1749 1414
rect 1751 1406 1759 1414
rect 1761 1406 1769 1414
rect 1771 1406 1779 1414
rect 1781 1406 1789 1414
rect 252 1376 260 1384
rect 732 1376 740 1384
rect 892 1376 900 1384
rect 1356 1376 1364 1384
rect 1804 1376 1812 1384
rect 1900 1376 1908 1384
rect 2140 1376 2148 1384
rect 1420 1356 1428 1364
rect 1532 1356 1540 1364
rect 220 1336 228 1344
rect 428 1336 436 1344
rect 460 1336 468 1344
rect 492 1336 500 1344
rect 620 1336 628 1344
rect 748 1336 756 1344
rect 1388 1336 1396 1344
rect 1500 1336 1508 1344
rect 2188 1336 2196 1344
rect 2332 1336 2340 1344
rect 44 1316 52 1324
rect 172 1316 180 1324
rect 284 1316 292 1324
rect 396 1316 404 1324
rect 668 1316 676 1324
rect 876 1316 884 1324
rect 924 1316 932 1324
rect 1004 1316 1012 1324
rect 1068 1318 1076 1326
rect 1180 1318 1188 1326
rect 1228 1316 1236 1324
rect 1324 1316 1332 1324
rect 1372 1316 1380 1324
rect 1436 1316 1444 1324
rect 1500 1316 1508 1324
rect 1564 1316 1572 1324
rect 1596 1316 1604 1324
rect 1660 1318 1668 1326
rect 1724 1316 1732 1324
rect 1804 1316 1812 1324
rect 1964 1318 1972 1326
rect 2028 1316 2036 1324
rect 2108 1316 2116 1324
rect 2204 1316 2212 1324
rect 2348 1316 2356 1324
rect 1484 1296 1492 1304
rect 1596 1296 1604 1304
rect 2156 1296 2164 1304
rect 12 1276 20 1284
rect 60 1276 68 1284
rect 300 1276 308 1284
rect 940 1276 948 1284
rect 1308 1276 1316 1284
rect 2092 1276 2100 1284
rect 2396 1276 2404 1284
rect 2172 1236 2180 1244
rect 595 1206 603 1214
rect 605 1206 613 1214
rect 615 1206 623 1214
rect 625 1206 633 1214
rect 635 1206 643 1214
rect 645 1206 653 1214
rect 396 1176 404 1184
rect 668 1176 676 1184
rect 1180 1176 1188 1184
rect 1356 1176 1364 1184
rect 1420 1176 1428 1184
rect 1532 1176 1540 1184
rect 1260 1156 1268 1164
rect 12 1136 20 1144
rect 60 1136 68 1144
rect 1244 1136 1252 1144
rect 2268 1136 2276 1144
rect 364 1116 372 1124
rect 780 1116 788 1124
rect 844 1116 852 1124
rect 876 1116 884 1124
rect 908 1116 916 1124
rect 940 1116 948 1124
rect 1004 1116 1012 1124
rect 1036 1116 1044 1124
rect 1132 1116 1140 1124
rect 1212 1116 1220 1124
rect 1292 1116 1300 1124
rect 1324 1116 1332 1124
rect 1340 1116 1348 1124
rect 1388 1116 1396 1124
rect 1708 1116 1716 1124
rect 1868 1116 1876 1124
rect 44 1096 52 1104
rect 188 1094 196 1102
rect 252 1096 260 1104
rect 284 1096 292 1104
rect 332 1096 340 1104
rect 364 1096 372 1104
rect 396 1096 404 1104
rect 140 1076 148 1084
rect 220 1076 228 1084
rect 268 1076 276 1084
rect 300 1076 308 1084
rect 556 1096 564 1104
rect 684 1096 692 1104
rect 844 1096 852 1104
rect 908 1096 916 1104
rect 1004 1096 1012 1104
rect 1084 1096 1092 1104
rect 1148 1096 1156 1104
rect 1164 1096 1172 1104
rect 1260 1096 1268 1104
rect 1420 1096 1428 1104
rect 1484 1096 1492 1104
rect 1548 1096 1556 1104
rect 1564 1096 1572 1104
rect 1596 1096 1604 1104
rect 1628 1096 1636 1104
rect 1868 1096 1876 1104
rect 460 1080 468 1088
rect 476 1076 484 1084
rect 572 1076 580 1084
rect 684 1076 692 1084
rect 828 1076 836 1084
rect 892 1076 900 1084
rect 988 1076 996 1084
rect 1948 1094 1956 1102
rect 2012 1096 2020 1104
rect 2156 1096 2164 1104
rect 2204 1096 2212 1104
rect 2284 1096 2292 1104
rect 2380 1096 2388 1104
rect 1100 1076 1108 1084
rect 1132 1076 1140 1084
rect 1164 1076 1172 1084
rect 1292 1076 1300 1084
rect 1372 1076 1380 1084
rect 1436 1076 1444 1084
rect 1468 1076 1476 1084
rect 1564 1076 1572 1084
rect 1580 1076 1588 1084
rect 1612 1076 1620 1084
rect 1676 1076 1684 1084
rect 1820 1076 1828 1084
rect 1884 1076 1892 1084
rect 1996 1076 2004 1084
rect 2332 1076 2340 1084
rect 956 1056 964 1064
rect 1644 1056 1652 1064
rect 1772 1056 1780 1064
rect 2332 1056 2340 1064
rect 796 1036 804 1044
rect 1052 1036 1060 1044
rect 1660 1036 1668 1044
rect 2076 1036 2084 1044
rect 2348 1036 2356 1044
rect 1731 1006 1739 1014
rect 1741 1006 1749 1014
rect 1751 1006 1759 1014
rect 1761 1006 1769 1014
rect 1771 1006 1779 1014
rect 1781 1006 1789 1014
rect 12 976 20 984
rect 316 976 324 984
rect 556 976 564 984
rect 668 976 676 984
rect 844 976 852 984
rect 940 976 948 984
rect 1020 976 1028 984
rect 1180 976 1188 984
rect 1372 976 1380 984
rect 1388 976 1396 984
rect 1548 976 1556 984
rect 1868 976 1876 984
rect 2060 976 2068 984
rect 140 956 148 964
rect 428 956 436 964
rect 892 956 900 964
rect 956 956 964 964
rect 1244 956 1252 964
rect 1676 956 1684 964
rect 1996 956 2004 964
rect 2076 956 2084 964
rect 2396 956 2404 964
rect 172 936 180 944
rect 236 936 244 944
rect 300 936 308 944
rect 364 936 372 944
rect 572 936 580 944
rect 620 936 628 944
rect 716 936 724 944
rect 796 936 804 944
rect 876 936 884 944
rect 972 936 980 944
rect 1036 936 1044 944
rect 1100 936 1108 944
rect 1148 936 1156 944
rect 1436 936 1444 944
rect 1500 936 1508 944
rect 1532 936 1540 944
rect 1788 936 1796 944
rect 2092 936 2100 944
rect 2204 936 2212 944
rect 140 918 148 926
rect 236 916 244 924
rect 300 916 308 924
rect 348 916 356 924
rect 444 916 452 924
rect 204 896 212 904
rect 316 896 324 904
rect 684 896 692 904
rect 716 896 724 904
rect 796 916 804 924
rect 924 916 932 924
rect 988 916 996 924
rect 1052 916 1060 924
rect 1244 918 1252 926
rect 1436 916 1444 924
rect 1452 916 1460 924
rect 1100 896 1108 904
rect 1180 896 1188 904
rect 1644 916 1652 924
rect 1788 916 1796 924
rect 1852 916 1860 924
rect 1980 916 1988 924
rect 2204 916 2212 924
rect 2332 916 2340 924
rect 1500 896 1508 904
rect 1852 896 1860 904
rect 2124 896 2132 904
rect 2092 876 2100 884
rect 2316 876 2324 884
rect 595 806 603 814
rect 605 806 613 814
rect 615 806 623 814
rect 625 806 633 814
rect 635 806 643 814
rect 645 806 653 814
rect 284 776 292 784
rect 1004 776 1012 784
rect 2364 776 2372 784
rect 60 736 68 744
rect 1052 736 1060 744
rect 1276 736 1284 744
rect 1628 736 1636 744
rect 1932 736 1940 744
rect 2012 736 2020 744
rect 252 716 260 724
rect 348 716 356 724
rect 668 716 676 724
rect 716 716 724 724
rect 764 716 772 724
rect 796 716 804 724
rect 44 696 52 704
rect 188 694 196 702
rect 284 696 292 704
rect 380 696 388 704
rect 636 696 644 704
rect 716 696 724 704
rect 732 696 740 704
rect 812 696 820 704
rect 844 696 852 704
rect 876 696 884 704
rect 908 696 916 704
rect 956 716 964 724
rect 1292 716 1300 724
rect 1036 696 1044 704
rect 1164 696 1172 704
rect 1244 696 1252 704
rect 1324 696 1332 704
rect 1372 696 1380 704
rect 1420 716 1428 724
rect 1484 716 1492 724
rect 1644 716 1652 724
rect 1964 716 1972 724
rect 1980 716 1988 724
rect 2044 716 2052 724
rect 2076 716 2084 724
rect 1548 696 1556 704
rect 1580 696 1588 704
rect 1596 696 1604 704
rect 1804 694 1812 702
rect 2012 696 2020 704
rect 2108 696 2116 704
rect 2172 696 2180 704
rect 2252 696 2260 704
rect 12 676 20 684
rect 172 676 180 684
rect 396 676 404 684
rect 444 676 452 684
rect 540 676 548 684
rect 732 676 740 684
rect 748 676 756 684
rect 828 676 836 684
rect 876 676 884 684
rect 892 676 900 684
rect 940 676 948 684
rect 988 676 996 684
rect 1164 676 1172 684
rect 1356 676 1364 684
rect 1388 676 1396 684
rect 1468 676 1476 684
rect 1484 676 1492 684
rect 1516 676 1524 684
rect 1740 676 1748 684
rect 1836 676 1844 684
rect 1996 676 2004 684
rect 2060 676 2068 684
rect 2108 676 2116 684
rect 2156 676 2164 684
rect 2268 676 2276 684
rect 556 656 564 664
rect 588 656 596 664
rect 1548 656 1556 664
rect 1564 656 1572 664
rect 524 636 532 644
rect 1292 636 1300 644
rect 1644 636 1652 644
rect 2140 636 2148 644
rect 1731 606 1739 614
rect 1741 606 1749 614
rect 1751 606 1759 614
rect 1761 606 1769 614
rect 1771 606 1779 614
rect 1781 606 1789 614
rect 204 576 212 584
rect 236 576 244 584
rect 284 576 292 584
rect 620 576 628 584
rect 716 576 724 584
rect 748 576 756 584
rect 860 576 868 584
rect 1084 576 1092 584
rect 1100 576 1108 584
rect 1468 576 1476 584
rect 1484 576 1492 584
rect 1628 576 1636 584
rect 1804 576 1812 584
rect 1900 576 1908 584
rect 60 556 68 564
rect 220 556 228 564
rect 732 556 740 564
rect 764 556 772 564
rect 1068 556 1076 564
rect 1980 556 1988 564
rect 2028 556 2036 564
rect 2172 556 2180 564
rect 2188 556 2196 564
rect 12 536 20 544
rect 108 536 116 544
rect 140 536 148 544
rect 156 536 164 544
rect 268 536 276 544
rect 300 536 308 544
rect 92 516 100 524
rect 252 516 260 524
rect 332 536 340 544
rect 428 536 436 544
rect 460 536 468 544
rect 924 536 932 544
rect 1564 536 1572 544
rect 1612 536 1620 544
rect 1676 536 1684 544
rect 1692 536 1700 544
rect 1836 536 1844 544
rect 44 496 52 504
rect 108 496 116 504
rect 204 496 212 504
rect 364 496 372 504
rect 412 516 420 524
rect 492 518 500 526
rect 636 516 644 524
rect 828 516 836 524
rect 908 516 916 524
rect 1036 516 1044 524
rect 1164 516 1172 524
rect 1228 518 1236 526
rect 1388 516 1396 524
rect 1516 516 1524 524
rect 1532 516 1540 524
rect 1580 516 1588 524
rect 1660 516 1668 524
rect 1708 516 1716 524
rect 1868 536 1876 544
rect 1900 536 1908 544
rect 1948 536 1956 544
rect 1996 536 2004 544
rect 2108 536 2116 544
rect 2204 536 2212 544
rect 2236 536 2244 544
rect 1916 516 1924 524
rect 1996 516 2004 524
rect 2076 516 2084 524
rect 2124 516 2132 524
rect 2220 516 2228 524
rect 412 496 420 504
rect 1628 496 1636 504
rect 2076 496 2084 504
rect 2156 496 2164 504
rect 28 476 36 484
rect 2044 476 2052 484
rect 2060 476 2068 484
rect 2124 456 2132 464
rect 780 436 788 444
rect 876 436 884 444
rect 1820 436 1828 444
rect 2012 436 2020 444
rect 2348 436 2356 444
rect 595 406 603 414
rect 605 406 613 414
rect 615 406 623 414
rect 625 406 633 414
rect 635 406 643 414
rect 645 406 653 414
rect 364 376 372 384
rect 1052 376 1060 384
rect 1900 376 1908 384
rect 2172 376 2180 384
rect 1100 356 1108 364
rect 380 336 388 344
rect 1116 336 1124 344
rect 1996 336 2004 344
rect 2188 336 2196 344
rect 236 316 244 324
rect 412 316 420 324
rect 748 316 756 324
rect 140 294 148 302
rect 316 296 324 304
rect 396 296 404 304
rect 476 296 484 304
rect 620 294 628 302
rect 780 296 788 304
rect 828 316 836 324
rect 908 316 916 324
rect 924 316 932 324
rect 988 316 996 324
rect 1020 316 1028 324
rect 1084 316 1092 324
rect 1244 316 1252 324
rect 1340 316 1348 324
rect 1644 316 1652 324
rect 1964 316 1972 324
rect 2028 316 2036 324
rect 844 296 852 304
rect 940 296 948 304
rect 1004 296 1012 304
rect 1052 296 1060 304
rect 1100 296 1108 304
rect 1196 296 1204 304
rect 1260 296 1268 304
rect 1292 296 1300 304
rect 1324 296 1332 304
rect 1372 296 1380 304
rect 1436 296 1444 304
rect 1548 296 1556 304
rect 1708 296 1716 304
rect 1868 296 1876 304
rect 1932 296 1940 304
rect 1980 296 1988 304
rect 2028 296 2036 304
rect 2060 296 2068 304
rect 2108 316 2116 324
rect 2156 316 2164 324
rect 2316 296 2324 304
rect 172 276 180 284
rect 204 276 212 284
rect 252 276 260 284
rect 300 276 308 284
rect 316 276 324 284
rect 460 276 468 284
rect 652 276 660 284
rect 684 276 692 284
rect 796 276 804 284
rect 844 276 852 284
rect 892 276 900 284
rect 956 276 964 284
rect 988 276 996 284
rect 1068 276 1076 284
rect 1148 276 1156 284
rect 1212 276 1220 284
rect 1308 276 1316 284
rect 1356 276 1364 284
rect 1612 276 1620 284
rect 1804 276 1812 284
rect 1916 276 1924 284
rect 1948 276 1956 284
rect 1980 276 1988 284
rect 2044 276 2052 284
rect 2108 276 2116 284
rect 2156 276 2164 284
rect 2188 276 2196 284
rect 2268 276 2276 284
rect 2332 276 2340 284
rect 428 256 436 264
rect 876 256 884 264
rect 1148 256 1156 264
rect 1404 256 1412 264
rect 1820 256 1828 264
rect 1868 256 1876 264
rect 12 236 20 244
rect 332 236 340 244
rect 444 236 452 244
rect 492 236 500 244
rect 1452 236 1460 244
rect 1731 206 1739 214
rect 1741 206 1749 214
rect 1751 206 1759 214
rect 1761 206 1769 214
rect 1771 206 1779 214
rect 1781 206 1789 214
rect 268 176 276 184
rect 348 176 356 184
rect 460 176 468 184
rect 716 176 724 184
rect 1004 176 1012 184
rect 1052 176 1060 184
rect 1292 176 1300 184
rect 1340 176 1348 184
rect 1804 176 1812 184
rect 2044 176 2052 184
rect 2140 176 2148 184
rect 2332 176 2340 184
rect 172 136 180 144
rect 268 136 276 144
rect 300 136 308 144
rect 508 156 516 164
rect 844 156 852 164
rect 924 156 932 164
rect 940 156 948 164
rect 972 156 980 164
rect 988 156 996 164
rect 1068 156 1076 164
rect 1164 156 1172 164
rect 1484 156 1492 164
rect 2060 156 2068 164
rect 2268 156 2276 164
rect 380 136 388 144
rect 412 136 420 144
rect 444 136 452 144
rect 476 136 484 144
rect 604 136 612 144
rect 700 136 708 144
rect 1308 136 1316 144
rect 1356 136 1364 144
rect 1388 136 1396 144
rect 1756 136 1764 144
rect 1884 136 1892 144
rect 1932 136 1940 144
rect 2028 136 2036 144
rect 2076 136 2084 144
rect 2124 136 2132 144
rect 2380 136 2388 144
rect 44 116 52 124
rect 188 118 196 126
rect 252 116 260 124
rect 316 116 324 124
rect 396 116 404 124
rect 428 116 436 124
rect 492 116 500 124
rect 556 116 564 124
rect 668 116 676 124
rect 828 116 836 124
rect 940 116 948 124
rect 1020 116 1028 124
rect 1036 116 1044 124
rect 1084 116 1092 124
rect 1180 116 1188 124
rect 364 96 372 104
rect 604 96 612 104
rect 668 96 676 104
rect 1340 96 1348 104
rect 1388 96 1396 104
rect 1452 116 1460 124
rect 1500 116 1508 124
rect 1580 116 1588 124
rect 1724 118 1732 126
rect 1868 116 1876 124
rect 1948 116 1956 124
rect 1964 116 1972 124
rect 2060 116 2068 124
rect 2252 116 2260 124
rect 2364 116 2372 124
rect 1948 96 1956 104
rect 1996 96 2004 104
rect 2124 96 2132 104
rect 2332 96 2340 104
rect 12 76 20 84
rect 60 76 68 84
rect 1596 76 1604 84
rect 1532 36 1540 44
rect 1548 36 1556 44
rect 595 6 603 14
rect 605 6 613 14
rect 615 6 623 14
rect 625 6 633 14
rect 635 6 643 14
rect 645 6 653 14
<< metal2 >>
rect 253 1457 275 1463
rect 717 1457 739 1463
rect 253 1384 259 1457
rect 733 1384 739 1457
rect 829 1457 851 1463
rect 893 1457 915 1463
rect 13 1284 19 1296
rect 45 1283 51 1316
rect 45 1277 60 1283
rect 45 1137 60 1143
rect 45 1104 51 1137
rect 189 1084 195 1094
rect 221 1084 227 1336
rect 285 1283 291 1316
rect 285 1277 300 1283
rect 397 1184 403 1316
rect 285 1104 291 1116
rect 141 964 147 1076
rect 253 1043 259 1096
rect 301 1084 307 1096
rect 237 1037 259 1043
rect 237 984 243 1037
rect 237 944 243 976
rect 45 737 60 743
rect 45 704 51 737
rect 13 684 19 696
rect 61 544 67 556
rect 141 544 147 776
rect 173 684 179 936
rect 189 702 195 716
rect 173 564 179 676
rect 205 584 211 616
rect 237 584 243 636
rect 253 624 259 716
rect 269 684 275 1076
rect 285 784 291 1076
rect 317 984 323 1096
rect 317 784 323 896
rect 285 664 291 696
rect 45 444 51 496
rect 61 404 67 536
rect 93 444 99 516
rect 109 484 115 496
rect 141 302 147 316
rect 173 284 179 556
rect 221 544 227 556
rect 221 504 227 536
rect 253 524 259 596
rect 285 584 291 616
rect 301 544 307 676
rect 205 484 211 496
rect 237 304 243 316
rect 253 284 259 316
rect 13 204 19 236
rect 173 144 179 276
rect 205 204 211 276
rect 189 126 195 156
rect 253 124 259 196
rect 269 184 275 476
rect 301 423 307 536
rect 285 417 307 423
rect 285 144 291 417
rect 301 284 307 396
rect 317 323 323 776
rect 333 604 339 1096
rect 349 924 355 1136
rect 365 1084 371 1096
rect 365 944 371 1076
rect 429 964 435 1336
rect 461 1324 467 1336
rect 477 1084 483 1136
rect 573 1084 579 1316
rect 618 1214 630 1216
rect 603 1206 605 1214
rect 613 1206 615 1214
rect 623 1206 625 1214
rect 633 1206 635 1214
rect 643 1206 645 1214
rect 618 1204 630 1206
rect 669 1184 675 1316
rect 669 1077 684 1083
rect 669 984 675 1077
rect 557 943 563 976
rect 557 937 572 943
rect 349 744 355 916
rect 349 704 355 716
rect 349 644 355 696
rect 333 544 339 576
rect 365 524 371 916
rect 381 704 387 736
rect 397 684 403 936
rect 717 924 723 936
rect 618 814 630 816
rect 603 806 605 814
rect 613 806 615 814
rect 623 806 625 814
rect 633 806 635 814
rect 643 806 645 814
rect 618 804 630 806
rect 365 504 371 516
rect 365 384 371 436
rect 381 344 387 636
rect 429 544 435 696
rect 445 684 451 696
rect 541 684 547 776
rect 669 724 675 776
rect 685 684 691 896
rect 749 864 755 1336
rect 829 1084 835 1457
rect 893 1384 899 1457
rect 925 1283 931 1316
rect 925 1277 940 1283
rect 1037 1104 1043 1116
rect 845 1084 851 1096
rect 877 1077 892 1083
rect 797 944 803 1036
rect 845 984 851 1016
rect 877 944 883 1077
rect 893 1064 899 1076
rect 909 1044 915 1096
rect 1005 1084 1011 1096
rect 941 1063 947 1076
rect 989 1064 995 1076
rect 941 1057 956 1063
rect 941 984 947 1057
rect 1021 984 1027 1056
rect 973 924 979 936
rect 989 924 995 956
rect 1053 943 1059 1036
rect 1044 937 1059 943
rect 1037 924 1043 936
rect 797 904 803 916
rect 724 717 739 723
rect 733 704 739 717
rect 845 704 851 716
rect 877 704 883 736
rect 756 677 771 683
rect 733 663 739 676
rect 765 664 771 677
rect 733 657 755 663
rect 589 644 595 656
rect 461 544 467 556
rect 637 524 643 636
rect 717 584 723 656
rect 749 644 755 657
rect 749 584 755 636
rect 797 564 803 696
rect 813 604 819 696
rect 829 684 835 696
rect 493 504 499 518
rect 618 414 630 416
rect 603 406 605 414
rect 613 406 615 414
rect 623 406 625 414
rect 633 406 635 414
rect 643 406 645 414
rect 618 404 630 406
rect 381 324 387 336
rect 317 317 339 323
rect 333 283 339 317
rect 324 277 339 283
rect 301 224 307 276
rect 276 137 284 143
rect 13 84 19 96
rect 45 83 51 116
rect 45 77 60 83
rect 301 -23 307 136
rect 333 104 339 236
rect 349 184 355 216
rect 365 104 371 196
rect 397 164 403 296
rect 413 284 419 316
rect 477 304 483 316
rect 381 144 387 156
rect 413 144 419 176
rect 429 163 435 256
rect 445 184 451 236
rect 461 184 467 196
rect 429 157 444 163
rect 445 144 451 156
rect 397 104 403 116
rect 445 -23 451 136
rect 493 124 499 136
rect 557 124 563 296
rect 685 284 691 296
rect 733 284 739 556
rect 829 524 835 656
rect 861 584 867 696
rect 861 524 867 576
rect 877 524 883 676
rect 893 644 899 676
rect 909 524 915 576
rect 925 544 931 856
rect 941 684 947 716
rect 957 704 963 716
rect 781 304 787 436
rect 877 304 883 436
rect 925 324 931 516
rect 973 364 979 916
rect 1053 904 1059 916
rect 989 684 995 736
rect 1037 704 1043 756
rect 1069 723 1075 1318
rect 1101 1243 1107 1463
rect 1341 1457 1363 1463
rect 1357 1384 1363 1457
rect 1421 1424 1427 1463
rect 1533 1424 1539 1463
rect 1885 1457 1907 1463
rect 2125 1457 2147 1463
rect 1421 1364 1427 1416
rect 1389 1344 1395 1356
rect 1085 1237 1107 1243
rect 1085 1104 1091 1237
rect 1181 1184 1187 1318
rect 1421 1317 1436 1323
rect 1165 1104 1171 1116
rect 1108 1077 1123 1083
rect 1117 1044 1123 1077
rect 1165 1064 1171 1076
rect 1053 717 1075 723
rect 1053 384 1059 717
rect 1085 644 1091 1036
rect 1101 924 1107 936
rect 1069 564 1075 596
rect 1085 584 1091 636
rect 1117 604 1123 1036
rect 1181 984 1187 1116
rect 1229 1003 1235 1316
rect 1325 1283 1331 1316
rect 1316 1277 1331 1283
rect 1357 1184 1363 1256
rect 1373 1164 1379 1316
rect 1421 1184 1427 1317
rect 1261 1144 1267 1156
rect 1245 1024 1251 1136
rect 1325 1124 1331 1156
rect 1373 1117 1388 1123
rect 1261 1084 1267 1096
rect 1293 1084 1299 1116
rect 1293 1064 1299 1076
rect 1325 1024 1331 1116
rect 1373 1104 1379 1117
rect 1373 1084 1379 1096
rect 1229 997 1251 1003
rect 1149 944 1155 976
rect 1245 964 1251 997
rect 1389 984 1395 1116
rect 1421 1104 1427 1116
rect 1469 1084 1475 1416
rect 1533 1364 1539 1416
rect 1533 1184 1539 1296
rect 1565 1264 1571 1316
rect 1437 944 1443 1076
rect 1485 1044 1491 1096
rect 1549 984 1555 1096
rect 1581 1084 1587 1416
rect 1754 1414 1766 1416
rect 1739 1406 1741 1414
rect 1749 1406 1751 1414
rect 1759 1406 1761 1414
rect 1769 1406 1771 1414
rect 1779 1406 1781 1414
rect 1754 1404 1766 1406
rect 1901 1384 1907 1457
rect 2141 1384 2147 1457
rect 1661 1326 1667 1336
rect 1805 1324 1811 1376
rect 2301 1344 2307 1463
rect 2013 1317 2028 1323
rect 1597 1104 1603 1296
rect 1725 1284 1731 1316
rect 2013 1284 2019 1317
rect 2109 1283 2115 1316
rect 2100 1277 2115 1283
rect 1709 1104 1715 1116
rect 1677 1084 1683 1096
rect 1533 977 1548 983
rect 1533 944 1539 977
rect 1501 924 1507 936
rect 1165 704 1171 716
rect 1181 684 1187 896
rect 1277 744 1283 896
rect 1437 764 1443 916
rect 1453 904 1459 916
rect 1277 704 1283 736
rect 1421 704 1427 716
rect 653 184 659 276
rect 701 177 716 183
rect 701 144 707 177
rect 557 104 563 116
rect 605 104 611 136
rect 781 104 787 296
rect 797 284 803 296
rect 925 283 931 316
rect 925 277 947 283
rect 845 244 851 276
rect 877 244 883 256
rect 845 164 851 176
rect 493 -23 499 56
rect 877 44 883 236
rect 941 164 947 277
rect 973 283 979 356
rect 989 304 995 316
rect 1005 304 1011 376
rect 1069 304 1075 556
rect 1165 524 1171 676
rect 1245 664 1251 696
rect 1325 644 1331 696
rect 1229 526 1235 576
rect 1117 304 1123 336
rect 973 277 988 283
rect 1005 184 1011 196
rect 1053 184 1059 276
rect 1069 264 1075 276
rect 1101 244 1107 296
rect 1133 277 1148 283
rect 1133 264 1139 277
rect 1149 244 1155 256
rect 1165 184 1171 516
rect 1261 384 1267 596
rect 1293 584 1299 636
rect 1357 624 1363 676
rect 1389 524 1395 676
rect 1437 524 1443 756
rect 1469 584 1475 676
rect 1517 624 1523 676
rect 1549 664 1555 696
rect 1565 684 1571 1076
rect 1581 1064 1587 1076
rect 1581 704 1587 1036
rect 1661 944 1667 1036
rect 1677 964 1683 1036
rect 1709 904 1715 1096
rect 1725 1044 1731 1276
rect 1949 1102 1955 1116
rect 2013 1104 2019 1276
rect 2157 1084 2163 1096
rect 1821 1044 1827 1076
rect 1754 1014 1766 1016
rect 1739 1006 1741 1014
rect 1749 1006 1751 1014
rect 1759 1006 1761 1014
rect 1769 1006 1771 1014
rect 1779 1006 1781 1014
rect 1754 1004 1766 1006
rect 1789 904 1795 916
rect 1837 903 1843 1056
rect 1869 984 1875 1076
rect 1885 1004 1891 1076
rect 1997 964 2003 1076
rect 2084 1037 2099 1043
rect 2061 984 2067 996
rect 2077 924 2083 956
rect 2093 944 2099 1037
rect 2173 1024 2179 1236
rect 1837 897 1852 903
rect 1629 744 1635 896
rect 1629 723 1635 736
rect 1629 717 1644 723
rect 1485 584 1491 596
rect 1533 524 1539 656
rect 1549 604 1555 656
rect 1581 584 1587 696
rect 1597 664 1603 696
rect 1629 584 1635 696
rect 1741 684 1747 716
rect 1821 663 1827 736
rect 1933 724 1939 736
rect 1805 657 1827 663
rect 1213 284 1219 316
rect 1245 304 1251 316
rect 1261 304 1267 376
rect 1293 304 1299 316
rect 1213 264 1219 276
rect 1325 264 1331 296
rect 1341 184 1347 316
rect 1373 304 1379 316
rect 1549 284 1555 296
rect 1453 224 1459 236
rect 1165 164 1171 176
rect 1293 163 1299 176
rect 1485 164 1491 256
rect 1293 157 1308 163
rect 941 144 947 156
rect 941 104 947 116
rect 618 14 630 16
rect 603 6 605 14
rect 613 6 615 14
rect 623 6 625 14
rect 633 6 635 14
rect 643 6 645 14
rect 618 4 630 6
rect 893 -23 899 16
rect 925 -23 931 36
rect 957 -23 963 156
rect 973 124 979 156
rect 1037 104 1043 116
rect 1069 -17 1075 156
rect 1309 144 1315 156
rect 1357 144 1363 156
rect 1341 104 1347 136
rect 1389 124 1395 136
rect 1453 124 1459 156
rect 1453 104 1459 116
rect 1485 -17 1491 156
rect 1501 124 1507 216
rect 1565 164 1571 536
rect 1613 524 1619 536
rect 1645 503 1651 636
rect 1754 614 1766 616
rect 1739 606 1741 614
rect 1749 606 1751 614
rect 1759 606 1761 614
rect 1769 606 1771 614
rect 1779 606 1781 614
rect 1754 604 1766 606
rect 1805 584 1811 657
rect 1837 644 1843 676
rect 1901 584 1907 696
rect 1981 684 1987 716
rect 1997 684 2003 736
rect 1869 544 1875 576
rect 1661 524 1667 536
rect 1677 504 1683 536
rect 1636 497 1651 503
rect 1693 484 1699 536
rect 1709 504 1715 516
rect 1645 304 1651 316
rect 1709 304 1715 476
rect 1821 444 1827 496
rect 1613 184 1619 276
rect 1754 214 1766 216
rect 1739 206 1741 214
rect 1749 206 1751 214
rect 1759 206 1761 214
rect 1769 206 1771 214
rect 1779 206 1781 214
rect 1754 204 1766 206
rect 1805 184 1811 276
rect 1821 264 1827 436
rect 1757 144 1763 176
rect 1581 83 1587 116
rect 1581 77 1596 83
rect 1533 -17 1539 36
rect 1053 -23 1075 -17
rect 1469 -23 1491 -17
rect 1517 -23 1539 -17
rect 1549 -17 1555 36
rect 1837 -17 1843 536
rect 1869 304 1875 476
rect 1901 384 1907 536
rect 1901 304 1907 376
rect 1933 304 1939 616
rect 1997 584 2003 656
rect 2061 623 2067 676
rect 2045 617 2067 623
rect 1997 544 2003 576
rect 2029 544 2035 556
rect 2013 537 2028 543
rect 1949 484 1955 536
rect 2013 523 2019 537
rect 2004 517 2019 523
rect 1965 324 1971 336
rect 1869 124 1875 256
rect 1885 -17 1891 136
rect 1933 103 1939 136
rect 1949 124 1955 276
rect 1981 204 1987 276
rect 1997 104 2003 316
rect 2013 284 2019 436
rect 2029 324 2035 516
rect 2045 504 2051 617
rect 2061 484 2067 536
rect 2077 524 2083 696
rect 2061 344 2067 456
rect 2061 304 2067 336
rect 2029 164 2035 296
rect 2077 283 2083 496
rect 2061 277 2083 283
rect 2045 184 2051 256
rect 2061 164 2067 277
rect 2036 157 2051 163
rect 2045 123 2051 157
rect 2077 144 2083 196
rect 2045 117 2060 123
rect 2093 104 2099 876
rect 2109 704 2115 916
rect 2125 684 2131 896
rect 2189 764 2195 1336
rect 2205 1104 2211 1316
rect 2276 1137 2291 1143
rect 2285 1104 2291 1137
rect 2205 944 2211 1096
rect 2205 804 2211 916
rect 2301 864 2307 1336
rect 2333 1084 2339 1096
rect 2349 1063 2355 1316
rect 2397 1284 2403 1296
rect 2349 1057 2371 1063
rect 2333 883 2339 916
rect 2324 877 2339 883
rect 2157 684 2163 716
rect 2109 664 2115 676
rect 2173 663 2179 696
rect 2157 657 2179 663
rect 2109 544 2115 556
rect 2125 524 2131 536
rect 2109 324 2115 336
rect 2109 284 2115 296
rect 2141 224 2147 636
rect 2157 524 2163 657
rect 2157 463 2163 496
rect 2173 484 2179 556
rect 2205 544 2211 696
rect 2237 544 2243 856
rect 2253 704 2259 736
rect 2269 644 2275 676
rect 2221 504 2227 516
rect 2157 457 2179 463
rect 2173 384 2179 457
rect 2189 284 2195 336
rect 2269 284 2275 636
rect 2349 463 2355 1036
rect 2365 784 2371 1057
rect 2381 924 2387 1096
rect 2349 457 2371 463
rect 2349 383 2355 436
rect 2333 377 2355 383
rect 2333 284 2339 377
rect 2141 184 2147 196
rect 2269 184 2275 276
rect 2333 184 2339 256
rect 2269 164 2275 176
rect 2253 124 2259 136
rect 2349 123 2355 216
rect 2365 143 2371 457
rect 2365 137 2380 143
rect 2349 117 2364 123
rect 2125 104 2131 116
rect 1933 97 1948 103
rect 1549 -23 1571 -17
rect 1837 -23 1859 -17
rect 1885 -23 1907 -17
<< m3contact >>
rect 220 1336 228 1344
rect 492 1336 500 1344
rect 620 1336 628 1344
rect 748 1336 756 1344
rect 172 1316 180 1324
rect 12 1296 20 1304
rect 12 1136 20 1144
rect 348 1136 356 1144
rect 284 1116 292 1124
rect 300 1096 308 1104
rect 316 1096 324 1104
rect 188 1076 196 1084
rect 12 976 20 984
rect 284 1076 292 1084
rect 236 976 244 984
rect 140 918 148 924
rect 140 916 148 918
rect 140 776 148 784
rect 12 696 20 704
rect 236 916 244 924
rect 204 896 212 904
rect 188 716 196 724
rect 236 636 244 644
rect 204 616 212 624
rect 300 936 308 944
rect 300 916 308 924
rect 316 776 324 784
rect 268 676 276 684
rect 300 676 308 684
rect 284 656 292 664
rect 252 616 260 624
rect 284 616 292 624
rect 252 596 260 604
rect 172 556 180 564
rect 12 536 20 544
rect 60 536 68 544
rect 108 536 116 544
rect 156 536 164 544
rect 28 476 36 484
rect 44 436 52 444
rect 108 476 116 484
rect 92 436 100 444
rect 60 396 68 404
rect 140 316 148 324
rect 220 536 228 544
rect 268 536 276 544
rect 220 496 228 504
rect 204 476 212 484
rect 268 476 276 484
rect 252 316 260 324
rect 236 296 244 304
rect 12 196 20 204
rect 204 196 212 204
rect 252 196 260 204
rect 188 156 196 164
rect 300 396 308 404
rect 364 1116 372 1124
rect 396 1096 404 1104
rect 364 1076 372 1084
rect 460 1316 468 1324
rect 572 1316 580 1324
rect 476 1136 484 1144
rect 556 1096 564 1104
rect 595 1206 603 1214
rect 605 1206 613 1214
rect 615 1206 623 1214
rect 625 1206 633 1214
rect 635 1206 643 1214
rect 645 1206 653 1214
rect 684 1096 692 1104
rect 460 1080 468 1084
rect 460 1076 468 1080
rect 364 936 372 944
rect 396 936 404 944
rect 572 936 580 944
rect 620 936 628 944
rect 364 916 372 924
rect 348 736 356 744
rect 348 696 356 704
rect 348 636 356 644
rect 332 596 340 604
rect 332 576 340 584
rect 380 736 388 744
rect 444 916 452 924
rect 716 916 724 924
rect 716 896 724 904
rect 595 806 603 814
rect 605 806 613 814
rect 615 806 623 814
rect 625 806 633 814
rect 635 806 643 814
rect 645 806 653 814
rect 540 776 548 784
rect 668 776 676 784
rect 428 696 436 704
rect 444 696 452 704
rect 380 636 388 644
rect 364 516 372 524
rect 364 436 372 444
rect 636 696 644 704
rect 780 1116 788 1124
rect 876 1316 884 1324
rect 1004 1316 1012 1324
rect 844 1116 852 1124
rect 876 1116 884 1124
rect 908 1116 916 1124
rect 940 1116 948 1124
rect 1004 1116 1012 1124
rect 1036 1096 1044 1104
rect 844 1076 852 1084
rect 844 1016 852 1024
rect 892 1056 900 1064
rect 940 1076 948 1084
rect 1004 1076 1012 1084
rect 908 1036 916 1044
rect 988 1056 996 1064
rect 1020 1056 1028 1064
rect 892 956 900 964
rect 956 956 964 964
rect 988 956 996 964
rect 796 936 804 944
rect 876 936 884 944
rect 924 916 932 924
rect 972 916 980 924
rect 988 916 996 924
rect 1036 916 1044 924
rect 796 896 804 904
rect 748 856 756 864
rect 924 856 932 864
rect 876 736 884 744
rect 764 716 772 724
rect 796 716 804 724
rect 844 716 852 724
rect 716 696 724 704
rect 796 696 804 704
rect 828 696 836 704
rect 860 696 868 704
rect 908 696 916 704
rect 684 676 692 684
rect 556 656 564 664
rect 716 656 724 664
rect 524 636 532 644
rect 588 636 596 644
rect 636 636 644 644
rect 620 576 628 584
rect 460 556 468 564
rect 412 516 420 524
rect 764 656 772 664
rect 748 636 756 644
rect 828 656 836 664
rect 812 596 820 604
rect 732 556 740 564
rect 764 556 772 564
rect 796 556 804 564
rect 412 496 420 504
rect 492 496 500 504
rect 595 406 603 414
rect 605 406 613 414
rect 615 406 623 414
rect 625 406 633 414
rect 635 406 643 414
rect 645 406 653 414
rect 316 296 324 304
rect 380 316 388 324
rect 476 316 484 324
rect 300 216 308 224
rect 284 136 292 144
rect 12 96 20 104
rect 316 116 324 124
rect 348 216 356 224
rect 364 196 372 204
rect 556 296 564 304
rect 620 302 628 304
rect 620 296 628 302
rect 684 296 692 304
rect 412 276 420 284
rect 460 276 468 284
rect 412 176 420 184
rect 380 156 388 164
rect 396 156 404 164
rect 492 236 500 244
rect 460 196 468 204
rect 444 176 452 184
rect 444 156 452 164
rect 508 156 516 164
rect 476 136 484 144
rect 492 136 500 144
rect 428 116 436 124
rect 332 96 340 104
rect 396 96 404 104
rect 876 676 884 684
rect 892 636 900 644
rect 908 576 916 584
rect 940 716 948 724
rect 956 696 964 704
rect 860 516 868 524
rect 876 516 884 524
rect 924 516 932 524
rect 748 316 756 324
rect 828 316 836 324
rect 1052 896 1060 904
rect 1004 776 1012 784
rect 1036 756 1044 764
rect 988 736 996 744
rect 1052 736 1060 744
rect 1420 1416 1428 1424
rect 1468 1416 1476 1424
rect 1532 1416 1540 1424
rect 1580 1416 1588 1424
rect 1388 1356 1396 1364
rect 1372 1316 1380 1324
rect 1132 1116 1140 1124
rect 1164 1116 1172 1124
rect 1180 1116 1188 1124
rect 1212 1116 1220 1124
rect 1148 1096 1156 1104
rect 1132 1076 1140 1084
rect 1164 1056 1172 1064
rect 1084 1036 1092 1044
rect 1116 1036 1124 1044
rect 1036 516 1044 524
rect 1100 916 1108 924
rect 1100 896 1108 904
rect 1084 636 1092 644
rect 1068 596 1076 604
rect 1356 1256 1364 1264
rect 1324 1156 1332 1164
rect 1372 1156 1380 1164
rect 1260 1136 1268 1144
rect 1340 1116 1348 1124
rect 1260 1076 1268 1084
rect 1292 1056 1300 1064
rect 1420 1116 1428 1124
rect 1372 1096 1380 1104
rect 1244 1016 1252 1024
rect 1324 1016 1332 1024
rect 1148 976 1156 984
rect 1532 1356 1540 1364
rect 1500 1336 1508 1344
rect 1500 1316 1508 1324
rect 1484 1296 1492 1304
rect 1532 1296 1540 1304
rect 1564 1256 1572 1264
rect 1484 1096 1492 1104
rect 1564 1096 1572 1104
rect 1468 1076 1476 1084
rect 1372 976 1380 984
rect 1484 1036 1492 1044
rect 1731 1406 1739 1414
rect 1741 1406 1749 1414
rect 1751 1406 1759 1414
rect 1761 1406 1769 1414
rect 1771 1406 1779 1414
rect 1781 1406 1789 1414
rect 1660 1336 1668 1344
rect 1596 1316 1604 1324
rect 2300 1336 2308 1344
rect 2332 1336 2340 1344
rect 1964 1318 1972 1324
rect 1964 1316 1972 1318
rect 2028 1316 2036 1324
rect 1724 1276 1732 1284
rect 2012 1276 2020 1284
rect 2156 1296 2164 1304
rect 1628 1096 1636 1104
rect 1676 1096 1684 1104
rect 1708 1096 1716 1104
rect 1564 1076 1572 1084
rect 1612 1076 1620 1084
rect 1676 1076 1684 1084
rect 1244 918 1252 924
rect 1244 916 1252 918
rect 1500 916 1508 924
rect 1276 896 1284 904
rect 1164 716 1172 724
rect 1452 896 1460 904
rect 1500 896 1508 904
rect 1436 756 1444 764
rect 1292 716 1300 724
rect 1276 696 1284 704
rect 1372 696 1380 704
rect 1420 696 1428 704
rect 1180 676 1188 684
rect 1116 596 1124 604
rect 1100 576 1108 584
rect 1004 376 1012 384
rect 972 356 980 364
rect 908 316 916 324
rect 796 296 804 304
rect 844 296 852 304
rect 876 296 884 304
rect 732 276 740 284
rect 652 176 660 184
rect 700 136 708 144
rect 668 116 676 124
rect 844 276 852 284
rect 892 276 900 284
rect 940 296 948 304
rect 844 236 852 244
rect 876 236 884 244
rect 844 176 852 184
rect 828 116 836 124
rect 556 96 564 104
rect 668 96 676 104
rect 780 96 788 104
rect 492 56 500 64
rect 956 276 964 284
rect 1020 316 1028 324
rect 1244 656 1252 664
rect 1324 636 1332 644
rect 1260 596 1268 604
rect 1228 576 1236 584
rect 1164 516 1172 524
rect 1100 356 1108 364
rect 1084 316 1092 324
rect 988 296 996 304
rect 1052 296 1060 304
rect 1068 296 1076 304
rect 1116 296 1124 304
rect 1052 276 1060 284
rect 1004 196 1012 204
rect 1068 256 1076 264
rect 1132 256 1140 264
rect 1100 236 1108 244
rect 1148 236 1156 244
rect 1356 616 1364 624
rect 1292 576 1300 584
rect 1484 716 1492 724
rect 1484 676 1492 684
rect 1580 1056 1588 1064
rect 1644 1056 1652 1064
rect 1580 1036 1588 1044
rect 1676 1036 1684 1044
rect 1660 936 1668 944
rect 1644 916 1652 924
rect 1868 1116 1876 1124
rect 1948 1116 1956 1124
rect 1868 1096 1876 1104
rect 1868 1076 1876 1084
rect 2156 1076 2164 1084
rect 1772 1056 1780 1064
rect 1836 1056 1844 1064
rect 1724 1036 1732 1044
rect 1820 1036 1828 1044
rect 1731 1006 1739 1014
rect 1741 1006 1749 1014
rect 1751 1006 1759 1014
rect 1761 1006 1769 1014
rect 1771 1006 1779 1014
rect 1781 1006 1789 1014
rect 1788 936 1796 944
rect 1628 896 1636 904
rect 1708 896 1716 904
rect 1788 896 1796 904
rect 1884 996 1892 1004
rect 2076 1036 2084 1044
rect 2060 996 2068 1004
rect 2172 1016 2180 1024
rect 1852 916 1860 924
rect 1980 916 1988 924
rect 2076 916 2084 924
rect 2108 916 2116 924
rect 1820 736 1828 744
rect 1996 736 2004 744
rect 2012 736 2020 744
rect 1740 716 1748 724
rect 1628 696 1636 704
rect 1564 676 1572 684
rect 1532 656 1540 664
rect 1564 656 1572 664
rect 1516 616 1524 624
rect 1484 596 1492 604
rect 1548 596 1556 604
rect 1596 656 1604 664
rect 1804 702 1812 704
rect 1804 696 1812 702
rect 1932 716 1940 724
rect 1964 716 1972 724
rect 1900 696 1908 704
rect 1580 576 1588 584
rect 1564 536 1572 544
rect 1436 516 1444 524
rect 1516 516 1524 524
rect 1260 376 1268 384
rect 1212 316 1220 324
rect 1196 296 1204 304
rect 1292 316 1300 324
rect 1372 316 1380 324
rect 1244 296 1252 304
rect 1308 276 1316 284
rect 1212 256 1220 264
rect 1324 256 1332 264
rect 1436 296 1444 304
rect 1356 276 1364 284
rect 1548 276 1556 284
rect 1404 256 1412 264
rect 1484 256 1492 264
rect 1452 216 1460 224
rect 1164 176 1172 184
rect 924 156 932 164
rect 956 156 964 164
rect 988 156 996 164
rect 1500 216 1508 224
rect 1308 156 1316 164
rect 1356 156 1364 164
rect 1452 156 1460 164
rect 940 136 948 144
rect 940 96 948 104
rect 876 36 884 44
rect 924 36 932 44
rect 892 16 900 24
rect 595 6 603 14
rect 605 6 613 14
rect 615 6 623 14
rect 625 6 633 14
rect 635 6 643 14
rect 645 6 653 14
rect 972 116 980 124
rect 1020 116 1028 124
rect 1036 96 1044 104
rect 1340 136 1348 144
rect 1084 116 1092 124
rect 1180 116 1188 124
rect 1388 116 1396 124
rect 1388 96 1396 104
rect 1452 96 1460 104
rect 1580 516 1588 524
rect 1612 516 1620 524
rect 1731 606 1739 614
rect 1741 606 1749 614
rect 1751 606 1759 614
rect 1761 606 1769 614
rect 1771 606 1779 614
rect 1781 606 1789 614
rect 1836 636 1844 644
rect 2044 716 2052 724
rect 2076 716 2084 724
rect 2012 696 2020 704
rect 2076 696 2084 704
rect 1980 676 1988 684
rect 1996 656 2004 664
rect 1932 616 1940 624
rect 1868 576 1876 584
rect 1660 536 1668 544
rect 1676 496 1684 504
rect 1708 496 1716 504
rect 1820 496 1828 504
rect 1692 476 1700 484
rect 1708 476 1716 484
rect 1644 296 1652 304
rect 1804 276 1812 284
rect 1731 206 1739 214
rect 1741 206 1749 214
rect 1751 206 1759 214
rect 1761 206 1769 214
rect 1771 206 1779 214
rect 1781 206 1789 214
rect 1612 176 1620 184
rect 1756 176 1764 184
rect 1564 156 1572 164
rect 1724 118 1732 124
rect 1724 116 1732 118
rect 1868 476 1876 484
rect 1916 516 1924 524
rect 1996 576 2004 584
rect 1980 556 1988 564
rect 2028 536 2036 544
rect 2028 516 2036 524
rect 1948 476 1956 484
rect 1964 336 1972 344
rect 1996 336 2004 344
rect 1996 316 2004 324
rect 1900 296 1908 304
rect 1980 296 1988 304
rect 1916 276 1924 284
rect 1980 276 1988 284
rect 1980 196 1988 204
rect 1964 116 1972 124
rect 2060 536 2068 544
rect 2044 496 2052 504
rect 2076 496 2084 504
rect 2044 476 2052 484
rect 2060 476 2068 484
rect 2060 456 2068 464
rect 2060 336 2068 344
rect 2012 276 2020 284
rect 2044 276 2052 284
rect 2044 256 2052 264
rect 2076 196 2084 204
rect 2028 156 2036 164
rect 2028 136 2036 144
rect 2108 696 2116 704
rect 2204 1316 2212 1324
rect 2332 1096 2340 1104
rect 2332 1056 2340 1064
rect 2396 1296 2404 1304
rect 2236 856 2244 864
rect 2300 856 2308 864
rect 2204 796 2212 804
rect 2188 756 2196 764
rect 2156 716 2164 724
rect 2204 696 2212 704
rect 2124 676 2132 684
rect 2108 656 2116 664
rect 2108 556 2116 564
rect 2124 536 2132 544
rect 2124 456 2132 464
rect 2108 336 2116 344
rect 2108 296 2116 304
rect 2188 556 2196 564
rect 2156 516 2164 524
rect 2252 736 2260 744
rect 2268 636 2276 644
rect 2220 496 2228 504
rect 2172 476 2180 484
rect 2156 316 2164 324
rect 2396 956 2404 964
rect 2380 916 2388 924
rect 2316 296 2324 304
rect 2156 276 2164 284
rect 2188 276 2196 284
rect 2140 216 2148 224
rect 2140 196 2148 204
rect 2332 256 2340 264
rect 2348 216 2356 224
rect 2268 176 2276 184
rect 2124 136 2132 144
rect 2252 136 2260 144
rect 2124 116 2132 124
rect 2092 96 2100 104
rect 2332 96 2340 104
<< metal3 >>
rect 1428 1417 1468 1423
rect 1540 1417 1580 1423
rect 1730 1414 1790 1416
rect 1730 1406 1731 1414
rect 1740 1406 1741 1414
rect 1779 1406 1780 1414
rect 1789 1406 1790 1414
rect 1730 1404 1790 1406
rect 1396 1357 1532 1363
rect 228 1337 492 1343
rect 628 1337 748 1343
rect 1508 1337 1660 1343
rect 2308 1337 2332 1343
rect 468 1317 572 1323
rect 580 1317 876 1323
rect 884 1317 1004 1323
rect 1380 1317 1500 1323
rect 1604 1317 1964 1323
rect 2036 1317 2204 1323
rect -35 1297 12 1303
rect 1492 1297 1532 1303
rect 2004 1297 2156 1303
rect 2404 1297 2435 1303
rect 1732 1277 2012 1283
rect 1364 1257 1564 1263
rect 594 1214 654 1216
rect 594 1206 595 1214
rect 604 1206 605 1214
rect 643 1206 644 1214
rect 653 1206 654 1214
rect 594 1204 654 1206
rect 1332 1157 1372 1163
rect -35 1137 12 1143
rect 356 1137 476 1143
rect 484 1137 1260 1143
rect 292 1117 364 1123
rect 788 1117 844 1123
rect 884 1117 908 1123
rect 948 1117 1004 1123
rect 1140 1117 1164 1123
rect 1188 1117 1212 1123
rect 1348 1117 1420 1123
rect 1876 1117 1948 1123
rect -35 1097 300 1103
rect 324 1097 396 1103
rect 564 1097 684 1103
rect 1044 1097 1148 1103
rect 1156 1097 1372 1103
rect 1492 1097 1564 1103
rect 1636 1097 1676 1103
rect 1716 1097 1868 1103
rect 2340 1097 2435 1103
rect 196 1077 284 1083
rect 372 1077 460 1083
rect 852 1077 940 1083
rect 1012 1077 1132 1083
rect 1268 1077 1468 1083
rect 1572 1077 1612 1083
rect 1684 1077 1868 1083
rect 2164 1077 2284 1083
rect 900 1057 988 1063
rect 1028 1057 1164 1063
rect 1300 1057 1580 1063
rect 1588 1057 1644 1063
rect 1780 1057 1836 1063
rect 2340 1057 2380 1063
rect 2388 1057 2435 1063
rect 916 1037 1084 1043
rect 1124 1037 1484 1043
rect 1492 1037 1580 1043
rect 1684 1037 1724 1043
rect 1828 1037 2076 1043
rect 852 1017 1244 1023
rect 1252 1017 1324 1023
rect 2068 1017 2172 1023
rect 1730 1014 1790 1016
rect 1730 1006 1731 1014
rect 1740 1006 1741 1014
rect 1779 1006 1780 1014
rect 1789 1006 1790 1014
rect 1730 1004 1790 1006
rect 1892 997 2060 1003
rect 20 977 236 983
rect 1156 977 1372 983
rect 900 957 956 963
rect 964 957 988 963
rect 2404 957 2435 963
rect 308 937 364 943
rect 372 937 396 943
rect 580 937 620 943
rect 804 937 876 943
rect 1668 937 1788 943
rect 148 917 236 923
rect 308 917 364 923
rect 452 917 716 923
rect 932 917 972 923
rect 996 917 1036 923
rect 1108 917 1244 923
rect 1508 917 1644 923
rect 1860 917 1980 923
rect 2084 917 2108 923
rect 2116 917 2380 923
rect 2388 917 2435 923
rect 301 903 307 916
rect 212 897 307 903
rect 724 897 796 903
rect 804 897 1052 903
rect 1060 897 1100 903
rect 1108 897 1276 903
rect 1460 897 1500 903
rect 1508 897 1628 903
rect 1636 897 1708 903
rect 1716 897 1788 903
rect 756 857 924 863
rect 932 857 2236 863
rect 2244 857 2300 863
rect 594 814 654 816
rect 594 806 595 814
rect 604 806 605 814
rect 643 806 644 814
rect 653 806 654 814
rect 594 804 654 806
rect 2212 797 2220 803
rect 148 777 316 783
rect 324 777 540 783
rect 548 777 668 783
rect 676 777 1004 783
rect 1012 757 1036 763
rect 1044 757 1436 763
rect 2100 757 2188 763
rect 356 737 380 743
rect 884 737 988 743
rect 996 737 1052 743
rect 1828 737 1996 743
rect 2020 737 2252 743
rect 196 717 764 723
rect 804 717 844 723
rect 948 717 1164 723
rect 1300 717 1484 723
rect 1748 717 1932 723
rect 1972 717 2044 723
rect 2084 717 2156 723
rect -35 697 12 703
rect 356 697 428 703
rect 436 697 444 703
rect 644 697 716 703
rect 804 697 828 703
rect 868 697 908 703
rect 916 697 956 703
rect 1284 697 1372 703
rect 1380 697 1420 703
rect 1636 697 1804 703
rect 1908 697 2012 703
rect 2084 697 2108 703
rect 2116 697 2204 703
rect 276 677 300 683
rect 308 677 684 683
rect 692 677 876 683
rect 884 677 1180 683
rect 1188 677 1484 683
rect 1492 677 1564 683
rect 1572 677 1980 683
rect 1988 677 2124 683
rect 2132 677 2156 683
rect 292 657 556 663
rect 724 657 764 663
rect 836 657 1244 663
rect 1252 657 1532 663
rect 1540 657 1564 663
rect 1572 657 1596 663
rect 2004 657 2108 663
rect 244 637 348 643
rect 388 637 524 643
rect 532 637 588 643
rect 596 637 636 643
rect 756 637 892 643
rect 1092 637 1324 643
rect 1332 637 1827 643
rect 180 617 204 623
rect 260 617 284 623
rect 1364 617 1516 623
rect 1821 623 1827 637
rect 1844 637 2268 643
rect 1821 617 1932 623
rect 1730 614 1790 616
rect 1730 606 1731 614
rect 1740 606 1741 614
rect 1779 606 1780 614
rect 1789 606 1790 614
rect 1730 604 1790 606
rect 260 597 332 603
rect 340 597 428 603
rect 436 597 812 603
rect 820 597 1068 603
rect 1076 597 1116 603
rect 1268 597 1484 603
rect 1492 597 1548 603
rect 340 577 620 583
rect 916 577 1100 583
rect 1236 577 1292 583
rect 1588 577 1868 583
rect 1876 577 1996 583
rect 180 557 460 563
rect 740 557 764 563
rect 772 557 796 563
rect 1988 557 2099 563
rect 20 537 60 543
rect 116 537 156 543
rect 228 537 268 543
rect 1572 537 1660 543
rect 2036 537 2060 543
rect 2093 543 2099 557
rect 2116 557 2188 563
rect 2093 537 2124 543
rect 372 517 412 523
rect 420 517 860 523
rect 884 517 924 523
rect 1044 517 1164 523
rect 1444 517 1516 523
rect 1524 517 1580 523
rect 1620 517 1916 523
rect 1924 517 2028 523
rect 2036 517 2156 523
rect -35 497 220 503
rect 420 497 492 503
rect 1684 497 1708 503
rect 1716 497 1820 503
rect 2052 497 2076 503
rect 2084 497 2220 503
rect 2228 497 2380 503
rect 36 477 108 483
rect 212 477 268 483
rect 1700 477 1708 483
rect 1716 477 1868 483
rect 1876 477 1948 483
rect 1956 477 2044 483
rect 2068 477 2172 483
rect 2429 483 2435 503
rect 2180 477 2435 483
rect 2004 457 2060 463
rect 2132 457 2220 463
rect 52 437 92 443
rect 100 437 364 443
rect 594 414 654 416
rect 594 406 595 414
rect 604 406 605 414
rect 643 406 644 414
rect 653 406 654 414
rect 594 404 654 406
rect 68 397 300 403
rect 1012 377 1260 383
rect 980 357 1100 363
rect 1972 337 1996 343
rect 2068 337 2108 343
rect 148 317 252 323
rect 388 317 476 323
rect 756 317 828 323
rect 916 317 1020 323
rect 1092 317 1212 323
rect 1300 317 1372 323
rect 2004 317 2156 323
rect 244 297 316 303
rect 324 297 556 303
rect 628 297 684 303
rect 804 297 844 303
rect 996 297 1052 303
rect 1124 297 1196 303
rect 1204 297 1244 303
rect 1252 297 1436 303
rect 1444 297 1644 303
rect 1908 297 1980 303
rect 2116 297 2316 303
rect 420 277 460 283
rect 468 277 492 283
rect 500 277 732 283
rect 852 277 892 283
rect 964 277 1052 283
rect 1069 283 1075 296
rect 1060 277 1308 283
rect 1364 277 1548 283
rect 1812 277 1916 283
rect 1924 277 1980 283
rect 2020 277 2044 283
rect 2164 277 2188 283
rect 1076 257 1132 263
rect 1220 257 1324 263
rect 1332 257 1404 263
rect 1412 257 1484 263
rect 1524 257 2044 263
rect 2292 257 2332 263
rect 500 237 844 243
rect 884 237 940 243
rect 948 237 1100 243
rect 1108 237 1148 243
rect 308 217 348 223
rect 1460 217 1500 223
rect 2148 217 2348 223
rect 1730 214 1790 216
rect 1730 206 1731 214
rect 1740 206 1741 214
rect 1779 206 1780 214
rect 1789 206 1790 214
rect 1730 204 1790 206
rect 20 197 204 203
rect 212 197 252 203
rect 372 197 460 203
rect 1988 197 2076 203
rect 2100 197 2140 203
rect 420 177 444 183
rect 660 177 844 183
rect 852 177 1164 183
rect 1620 177 1756 183
rect 1764 177 2268 183
rect 196 157 380 163
rect 404 157 444 163
rect 452 157 508 163
rect 932 157 956 163
rect 964 157 988 163
rect 1316 157 1356 163
rect 1460 157 1564 163
rect 1572 157 2028 163
rect 292 137 476 143
rect 500 137 700 143
rect 948 137 1340 143
rect 2036 137 2092 143
rect 2132 137 2252 143
rect 324 117 428 123
rect 676 117 828 123
rect 980 117 1020 123
rect 1028 117 1084 123
rect 1188 117 1388 123
rect 1732 117 1964 123
rect 2068 117 2124 123
rect -35 97 12 103
rect 340 97 396 103
rect 564 97 668 103
rect 676 97 780 103
rect 948 97 1036 103
rect 1396 97 1452 103
rect 2100 97 2332 103
rect 884 37 924 43
rect 884 17 892 23
rect 594 14 654 16
rect 594 6 595 14
rect 604 6 605 14
rect 643 6 644 14
rect 653 6 654 14
rect 594 4 654 6
<< m4contact >>
rect 1732 1406 1739 1414
rect 1739 1406 1740 1414
rect 1744 1406 1749 1414
rect 1749 1406 1751 1414
rect 1751 1406 1752 1414
rect 1756 1406 1759 1414
rect 1759 1406 1761 1414
rect 1761 1406 1764 1414
rect 1768 1406 1769 1414
rect 1769 1406 1771 1414
rect 1771 1406 1776 1414
rect 1780 1406 1781 1414
rect 1781 1406 1788 1414
rect 172 1316 180 1324
rect 1996 1296 2004 1304
rect 596 1206 603 1214
rect 603 1206 604 1214
rect 608 1206 613 1214
rect 613 1206 615 1214
rect 615 1206 616 1214
rect 620 1206 623 1214
rect 623 1206 625 1214
rect 625 1206 628 1214
rect 632 1206 633 1214
rect 633 1206 635 1214
rect 635 1206 640 1214
rect 644 1206 645 1214
rect 645 1206 652 1214
rect 2284 1076 2292 1084
rect 2380 1056 2388 1064
rect 2060 1016 2068 1024
rect 1732 1006 1739 1014
rect 1739 1006 1740 1014
rect 1744 1006 1749 1014
rect 1749 1006 1751 1014
rect 1751 1006 1752 1014
rect 1756 1006 1759 1014
rect 1759 1006 1761 1014
rect 1761 1006 1764 1014
rect 1768 1006 1769 1014
rect 1769 1006 1771 1014
rect 1771 1006 1776 1014
rect 1780 1006 1781 1014
rect 1781 1006 1788 1014
rect 596 806 603 814
rect 603 806 604 814
rect 608 806 613 814
rect 613 806 615 814
rect 615 806 616 814
rect 620 806 623 814
rect 623 806 625 814
rect 625 806 628 814
rect 632 806 633 814
rect 633 806 635 814
rect 635 806 640 814
rect 644 806 645 814
rect 645 806 652 814
rect 2220 796 2228 804
rect 1004 756 1012 764
rect 2092 756 2100 764
rect 2156 676 2164 684
rect 172 616 180 624
rect 1516 616 1524 624
rect 1732 606 1739 614
rect 1739 606 1740 614
rect 1744 606 1749 614
rect 1749 606 1751 614
rect 1751 606 1752 614
rect 1756 606 1759 614
rect 1759 606 1761 614
rect 1761 606 1764 614
rect 1768 606 1769 614
rect 1769 606 1771 614
rect 1771 606 1776 614
rect 1780 606 1781 614
rect 1781 606 1788 614
rect 428 596 436 604
rect 2380 496 2388 504
rect 1996 456 2004 464
rect 2220 456 2228 464
rect 596 406 603 414
rect 603 406 604 414
rect 608 406 613 414
rect 613 406 615 414
rect 615 406 616 414
rect 620 406 623 414
rect 623 406 625 414
rect 625 406 628 414
rect 632 406 633 414
rect 633 406 635 414
rect 635 406 640 414
rect 644 406 645 414
rect 645 406 652 414
rect 2156 316 2164 324
rect 876 296 884 304
rect 940 296 948 304
rect 492 276 500 284
rect 1516 256 1524 264
rect 2284 256 2292 264
rect 940 236 948 244
rect 1732 206 1739 214
rect 1739 206 1740 214
rect 1744 206 1749 214
rect 1749 206 1751 214
rect 1751 206 1752 214
rect 1756 206 1759 214
rect 1759 206 1761 214
rect 1761 206 1764 214
rect 1768 206 1769 214
rect 1769 206 1771 214
rect 1771 206 1776 214
rect 1780 206 1781 214
rect 1781 206 1788 214
rect 1004 196 1012 204
rect 2092 196 2100 204
rect 2092 136 2100 144
rect 428 116 436 124
rect 2060 116 2068 124
rect 492 56 500 64
rect 876 16 884 24
rect 596 6 603 14
rect 603 6 604 14
rect 608 6 613 14
rect 613 6 615 14
rect 615 6 616 14
rect 620 6 623 14
rect 623 6 625 14
rect 625 6 628 14
rect 632 6 633 14
rect 633 6 635 14
rect 635 6 640 14
rect 644 6 645 14
rect 645 6 652 14
<< metal4 >>
rect 170 1324 182 1326
rect 170 1316 172 1324
rect 180 1316 182 1324
rect 170 624 182 1316
rect 170 616 172 624
rect 180 616 182 624
rect 170 614 182 616
rect 592 1214 656 1416
rect 592 1206 596 1214
rect 604 1206 608 1214
rect 616 1206 620 1214
rect 628 1206 632 1214
rect 640 1206 644 1214
rect 652 1206 656 1214
rect 592 814 656 1206
rect 592 806 596 814
rect 604 806 608 814
rect 616 806 620 814
rect 628 806 632 814
rect 640 806 644 814
rect 652 806 656 814
rect 426 604 438 606
rect 426 596 428 604
rect 436 596 438 604
rect 426 124 438 596
rect 592 414 656 806
rect 1728 1414 1792 1416
rect 1728 1406 1732 1414
rect 1740 1406 1744 1414
rect 1752 1406 1756 1414
rect 1764 1406 1768 1414
rect 1776 1406 1780 1414
rect 1788 1406 1792 1414
rect 1728 1014 1792 1406
rect 1728 1006 1732 1014
rect 1740 1006 1744 1014
rect 1752 1006 1756 1014
rect 1764 1006 1768 1014
rect 1776 1006 1780 1014
rect 1788 1006 1792 1014
rect 592 406 596 414
rect 604 406 608 414
rect 616 406 620 414
rect 628 406 632 414
rect 640 406 644 414
rect 652 406 656 414
rect 426 116 428 124
rect 436 116 438 124
rect 426 114 438 116
rect 490 284 502 286
rect 490 276 492 284
rect 500 276 502 284
rect 490 64 502 276
rect 490 56 492 64
rect 500 56 502 64
rect 490 54 502 56
rect 592 14 656 406
rect 1002 764 1014 766
rect 1002 756 1004 764
rect 1012 756 1014 764
rect 874 304 886 306
rect 874 296 876 304
rect 884 296 886 304
rect 874 24 886 296
rect 938 304 950 306
rect 938 296 940 304
rect 948 296 950 304
rect 938 244 950 296
rect 938 236 940 244
rect 948 236 950 244
rect 938 234 950 236
rect 1002 204 1014 756
rect 1514 624 1526 626
rect 1514 616 1516 624
rect 1524 616 1526 624
rect 1514 264 1526 616
rect 1514 256 1516 264
rect 1524 256 1526 264
rect 1514 254 1526 256
rect 1728 614 1792 1006
rect 1728 606 1732 614
rect 1740 606 1744 614
rect 1752 606 1756 614
rect 1764 606 1768 614
rect 1776 606 1780 614
rect 1788 606 1792 614
rect 1002 196 1004 204
rect 1012 196 1014 204
rect 1002 194 1014 196
rect 1728 214 1792 606
rect 1994 1304 2006 1306
rect 1994 1296 1996 1304
rect 2004 1296 2006 1304
rect 1994 464 2006 1296
rect 2282 1084 2294 1086
rect 2282 1076 2284 1084
rect 2292 1076 2294 1084
rect 1994 456 1996 464
rect 2004 456 2006 464
rect 1994 454 2006 456
rect 2058 1024 2070 1026
rect 2058 1016 2060 1024
rect 2068 1016 2070 1024
rect 1728 206 1732 214
rect 1740 206 1744 214
rect 1752 206 1756 214
rect 1764 206 1768 214
rect 1776 206 1780 214
rect 1788 206 1792 214
rect 874 16 876 24
rect 884 16 886 24
rect 874 14 886 16
rect 592 6 596 14
rect 604 6 608 14
rect 616 6 620 14
rect 628 6 632 14
rect 640 6 644 14
rect 652 6 656 14
rect 592 -10 656 6
rect 1728 -10 1792 206
rect 2058 124 2070 1016
rect 2218 804 2230 806
rect 2218 796 2220 804
rect 2228 796 2230 804
rect 2090 764 2102 766
rect 2090 756 2092 764
rect 2100 756 2102 764
rect 2090 204 2102 756
rect 2154 684 2166 686
rect 2154 676 2156 684
rect 2164 676 2166 684
rect 2154 324 2166 676
rect 2218 464 2230 796
rect 2218 456 2220 464
rect 2228 456 2230 464
rect 2218 454 2230 456
rect 2154 316 2156 324
rect 2164 316 2166 324
rect 2154 314 2166 316
rect 2282 264 2294 1076
rect 2378 1064 2390 1066
rect 2378 1056 2380 1064
rect 2388 1056 2390 1064
rect 2378 504 2390 1056
rect 2378 496 2380 504
rect 2388 496 2390 504
rect 2378 494 2390 496
rect 2282 256 2284 264
rect 2292 256 2294 264
rect 2282 254 2294 256
rect 2090 196 2092 204
rect 2100 196 2102 204
rect 2090 144 2102 196
rect 2090 136 2092 144
rect 2100 136 2102 144
rect 2090 134 2102 136
rect 2058 116 2060 124
rect 2068 116 2070 124
rect 2058 114 2070 116
use BUFX2  _257_
timestamp 1591628762
transform -1 0 56 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _273_
timestamp 1591628762
transform -1 0 248 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _290_
timestamp 1591628762
transform -1 0 200 0 1 210
box -4 -6 196 206
use NAND2X1  _158_
timestamp 1591628762
transform 1 0 200 0 1 210
box -4 -6 52 206
use AOI22X1  _241_
timestamp 1591628762
transform -1 0 328 0 -1 210
box -4 -6 84 206
use INVX1  _157_
timestamp 1591628762
transform 1 0 328 0 -1 210
box -4 -6 36 206
use OAI21X1  _237_
timestamp 1591628762
transform -1 0 424 0 -1 210
box -4 -6 68 206
use OAI21X1  _159_
timestamp 1591628762
transform -1 0 312 0 1 210
box -4 -6 68 206
use NAND2X1  _235_
timestamp 1591628762
transform 1 0 312 0 1 210
box -4 -6 52 206
use NAND3X1  _234_
timestamp 1591628762
transform -1 0 424 0 1 210
box -4 -6 68 206
use AOI22X1  _236_
timestamp 1591628762
transform 1 0 424 0 -1 210
box -4 -6 84 206
use INVX1  _154_
timestamp 1591628762
transform 1 0 504 0 -1 210
box -4 -6 36 206
use OAI21X1  _156_
timestamp 1591628762
transform 1 0 536 0 -1 210
box -4 -6 68 206
use AOI21X1  _233_
timestamp 1591628762
transform -1 0 488 0 1 210
box -4 -6 68 206
use DFFPOSX1  _281_
timestamp 1591628762
transform -1 0 680 0 1 210
box -4 -6 196 206
use FILL  SFILL6000x100
timestamp 1591628762
transform -1 0 616 0 -1 210
box -4 -6 20 206
use FILL  SFILL6960x2100
timestamp 1591628762
transform 1 0 696 0 1 210
box -4 -6 20 206
use FILL  SFILL6800x2100
timestamp 1591628762
transform 1 0 680 0 1 210
box -4 -6 20 206
use FILL  SFILL6480x100
timestamp 1591628762
transform -1 0 664 0 -1 210
box -4 -6 20 206
use FILL  SFILL6320x100
timestamp 1591628762
transform -1 0 648 0 -1 210
box -4 -6 20 206
use FILL  SFILL6160x100
timestamp 1591628762
transform -1 0 632 0 -1 210
box -4 -6 20 206
use NAND2X1  _155_
timestamp 1591628762
transform -1 0 712 0 -1 210
box -4 -6 52 206
use FILL  SFILL7280x2100
timestamp 1591628762
transform 1 0 728 0 1 210
box -4 -6 20 206
use FILL  SFILL7120x2100
timestamp 1591628762
transform 1 0 712 0 1 210
box -4 -6 20 206
use NAND2X1  _131_
timestamp 1591628762
transform -1 0 856 0 1 210
box -4 -6 52 206
use OAI21X1  _132_
timestamp 1591628762
transform -1 0 808 0 1 210
box -4 -6 68 206
use DFFPOSX1  _289_
timestamp 1591628762
transform -1 0 904 0 -1 210
box -4 -6 196 206
use INVX1  _110_
timestamp 1591628762
transform -1 0 936 0 -1 210
box -4 -6 36 206
use NOR2X1  _161_
timestamp 1591628762
transform -1 0 984 0 -1 210
box -4 -6 52 206
use NOR2X1  _109_
timestamp 1591628762
transform 1 0 984 0 -1 210
box -4 -6 52 206
use INVX1  _130_
timestamp 1591628762
transform -1 0 888 0 1 210
box -4 -6 36 206
use NAND2X1  _191_
timestamp 1591628762
transform 1 0 888 0 1 210
box -4 -6 52 206
use AOI22X1  _194_
timestamp 1591628762
transform 1 0 936 0 1 210
box -4 -6 84 206
use NOR2X1  _111_
timestamp 1591628762
transform -1 0 1080 0 -1 210
box -4 -6 52 206
use INVX1  _108_
timestamp 1591628762
transform 1 0 1080 0 -1 210
box -4 -6 36 206
use DFFPOSX1  _280_
timestamp 1591628762
transform 1 0 1112 0 -1 210
box -4 -6 196 206
use OAI21X1  _195_
timestamp 1591628762
transform -1 0 1080 0 1 210
box -4 -6 68 206
use NAND3X1  _193_
timestamp 1591628762
transform 1 0 1080 0 1 210
box -4 -6 68 206
use AOI21X1  _192_
timestamp 1591628762
transform -1 0 1208 0 1 210
box -4 -6 68 206
use NAND2X1  _188_
timestamp 1591628762
transform 1 0 1208 0 1 210
box -4 -6 52 206
use NAND2X1  _185_
timestamp 1591628762
transform 1 0 1304 0 -1 210
box -4 -6 52 206
use NAND2X1  _128_
timestamp 1591628762
transform 1 0 1352 0 -1 210
box -4 -6 52 206
use OAI21X1  _129_
timestamp 1591628762
transform -1 0 1464 0 -1 210
box -4 -6 68 206
use AOI22X1  _189_
timestamp 1591628762
transform -1 0 1336 0 1 210
box -4 -6 84 206
use OAI21X1  _190_
timestamp 1591628762
transform -1 0 1400 0 1 210
box -4 -6 68 206
use NOR2X1  _187_
timestamp 1591628762
transform 1 0 1400 0 1 210
box -4 -6 52 206
use INVX1  _127_
timestamp 1591628762
transform -1 0 1496 0 -1 210
box -4 -6 36 206
use BUFX2  _248_
timestamp 1591628762
transform 1 0 1496 0 -1 210
box -4 -6 52 206
use BUFX2  _247_
timestamp 1591628762
transform -1 0 1592 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _263_
timestamp 1591628762
transform -1 0 1784 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _264_
timestamp 1591628762
transform -1 0 1640 0 1 210
box -4 -6 196 206
use NOR3X1  _186_
timestamp 1591628762
transform -1 0 1768 0 1 210
box -4 -6 132 206
use FILL  SFILL17840x100
timestamp 1591628762
transform -1 0 1800 0 -1 210
box -4 -6 20 206
use FILL  SFILL18000x100
timestamp 1591628762
transform -1 0 1816 0 -1 210
box -4 -6 20 206
use FILL  SFILL17680x2100
timestamp 1591628762
transform 1 0 1768 0 1 210
box -4 -6 20 206
use FILL  SFILL17840x2100
timestamp 1591628762
transform 1 0 1784 0 1 210
box -4 -6 20 206
use FILL  SFILL18000x2100
timestamp 1591628762
transform 1 0 1800 0 1 210
box -4 -6 20 206
use FILL  SFILL18160x2100
timestamp 1591628762
transform 1 0 1816 0 1 210
box -4 -6 20 206
use FILL  SFILL18320x100
timestamp 1591628762
transform -1 0 1848 0 -1 210
box -4 -6 20 206
use FILL  SFILL18160x100
timestamp 1591628762
transform -1 0 1832 0 -1 210
box -4 -6 20 206
use INVX1  _177_
timestamp 1591628762
transform 1 0 1880 0 1 210
box -4 -6 36 206
use NOR2X1  _176_
timestamp 1591628762
transform 1 0 1832 0 1 210
box -4 -6 52 206
use OAI21X1  _183_
timestamp 1591628762
transform 1 0 1880 0 -1 210
box -4 -6 68 206
use INVX2  _124_
timestamp 1591628762
transform -1 0 1880 0 -1 210
box -4 -6 36 206
use OAI21X1  _182_
timestamp 1591628762
transform 1 0 1912 0 1 210
box -4 -6 68 206
use NAND2X1  _184_
timestamp 1591628762
transform -1 0 1992 0 -1 210
box -4 -6 52 206
use OAI21X1  _181_
timestamp 1591628762
transform 1 0 1976 0 1 210
box -4 -6 68 206
use NAND2X1  _180_
timestamp 1591628762
transform -1 0 2040 0 -1 210
box -4 -6 52 206
use INVX1  _107_
timestamp 1591628762
transform -1 0 2072 0 -1 210
box -4 -6 36 206
use OAI21X1  _126_
timestamp 1591628762
transform 1 0 2072 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _279_
timestamp 1591628762
transform -1 0 2328 0 -1 210
box -4 -6 196 206
use OAI21X1  _120_
timestamp 1591628762
transform 1 0 2040 0 1 210
box -4 -6 68 206
use NAND2X1  _119_
timestamp 1591628762
transform -1 0 2152 0 1 210
box -4 -6 52 206
use NAND2X1  _169_
timestamp 1591628762
transform -1 0 2200 0 1 210
box -4 -6 52 206
use DFFPOSX1  _277_
timestamp 1591628762
transform -1 0 2392 0 1 210
box -4 -6 196 206
use OAI21X1  _168_
timestamp 1591628762
transform -1 0 2392 0 -1 210
box -4 -6 68 206
use NAND2X1  _239_
timestamp 1591628762
transform 1 0 8 0 -1 610
box -4 -6 52 206
use NOR2X1  _238_
timestamp 1591628762
transform 1 0 56 0 -1 610
box -4 -6 52 206
use NAND2X1  _240_
timestamp 1591628762
transform -1 0 152 0 -1 610
box -4 -6 52 206
use OAI21X1  _242_
timestamp 1591628762
transform 1 0 152 0 -1 610
box -4 -6 68 206
use INVX1  _148_
timestamp 1591628762
transform 1 0 216 0 -1 610
box -4 -6 36 206
use AOI22X1  _227_
timestamp 1591628762
transform 1 0 248 0 -1 610
box -4 -6 84 206
use NAND2X1  _149_
timestamp 1591628762
transform 1 0 328 0 -1 610
box -4 -6 52 206
use OAI21X1  _150_
timestamp 1591628762
transform -1 0 440 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _287_
timestamp 1591628762
transform 1 0 440 0 -1 610
box -4 -6 196 206
use NOR2X1  _229_
timestamp 1591628762
transform -1 0 744 0 -1 610
box -4 -6 52 206
use INVX1  _151_
timestamp 1591628762
transform -1 0 776 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert8
timestamp 1591628762
transform -1 0 824 0 -1 610
box -4 -6 52 206
use FILL  SFILL6320x4100
timestamp 1591628762
transform -1 0 648 0 -1 610
box -4 -6 20 206
use FILL  SFILL6480x4100
timestamp 1591628762
transform -1 0 664 0 -1 610
box -4 -6 20 206
use FILL  SFILL6640x4100
timestamp 1591628762
transform -1 0 680 0 -1 610
box -4 -6 20 206
use FILL  SFILL6800x4100
timestamp 1591628762
transform -1 0 696 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert7
timestamp 1591628762
transform 1 0 824 0 -1 610
box -4 -6 52 206
use BUFX2  _243_
timestamp 1591628762
transform -1 0 920 0 -1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert4
timestamp 1591628762
transform 1 0 920 0 -1 610
box -4 -6 148 206
use INVX1  _160_
timestamp 1591628762
transform 1 0 1064 0 -1 610
box -4 -6 36 206
use DFFPOSX1  _259_
timestamp 1591628762
transform -1 0 1288 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _275_
timestamp 1591628762
transform 1 0 1288 0 -1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert12
timestamp 1591628762
transform -1 0 1528 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert5
timestamp 1591628762
transform 1 0 1528 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert11
timestamp 1591628762
transform 1 0 1576 0 -1 610
box -4 -6 52 206
use OAI21X1  _123_
timestamp 1591628762
transform -1 0 1688 0 -1 610
box -4 -6 68 206
use AND2X2  _175_
timestamp 1591628762
transform 1 0 1688 0 -1 610
box -4 -6 68 206
use FILL  SFILL17520x4100
timestamp 1591628762
transform -1 0 1768 0 -1 610
box -4 -6 20 206
use FILL  SFILL17680x4100
timestamp 1591628762
transform -1 0 1784 0 -1 610
box -4 -6 20 206
use FILL  SFILL17840x4100
timestamp 1591628762
transform -1 0 1800 0 -1 610
box -4 -6 20 206
use FILL  SFILL18000x4100
timestamp 1591628762
transform -1 0 1816 0 -1 610
box -4 -6 20 206
use INVX2  _121_
timestamp 1591628762
transform -1 0 1848 0 -1 610
box -4 -6 36 206
use AOI22X1  _178_
timestamp 1591628762
transform 1 0 1848 0 -1 610
box -4 -6 84 206
use AOI22X1  _172_
timestamp 1591628762
transform 1 0 1928 0 -1 610
box -4 -6 84 206
use INVX1  _118_
timestamp 1591628762
transform -1 0 2040 0 -1 610
box -4 -6 36 206
use NAND3X1  _171_
timestamp 1591628762
transform -1 0 2104 0 -1 610
box -4 -6 68 206
use OAI21X1  _173_
timestamp 1591628762
transform 1 0 2104 0 -1 610
box -4 -6 68 206
use AOI21X1  _170_
timestamp 1591628762
transform -1 0 2232 0 -1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert3
timestamp 1591628762
transform 1 0 2232 0 -1 610
box -4 -6 148 206
use FILL  FILL22480x4100
timestamp 1591628762
transform -1 0 2392 0 -1 610
box -4 -6 20 206
use BUFX2  _256_
timestamp 1591628762
transform -1 0 56 0 1 610
box -4 -6 52 206
use DFFPOSX1  _272_
timestamp 1591628762
transform -1 0 248 0 1 610
box -4 -6 196 206
use OAI21X1  _228_
timestamp 1591628762
transform -1 0 312 0 1 610
box -4 -6 68 206
use INVX1  _223_
timestamp 1591628762
transform -1 0 344 0 1 610
box -4 -6 36 206
use OAI21X1  _222_
timestamp 1591628762
transform -1 0 408 0 1 610
box -4 -6 68 206
use NOR3X1  _224_
timestamp 1591628762
transform 1 0 408 0 1 610
box -4 -6 132 206
use NAND2X1  _226_
timestamp 1591628762
transform 1 0 536 0 1 610
box -4 -6 52 206
use INVX1  _225_
timestamp 1591628762
transform 1 0 584 0 1 610
box -4 -6 36 206
use OAI21X1  _230_
timestamp 1591628762
transform -1 0 744 0 1 610
box -4 -6 68 206
use OAI21X1  _232_
timestamp 1591628762
transform 1 0 744 0 1 610
box -4 -6 68 206
use AOI22X1  _231_
timestamp 1591628762
transform 1 0 808 0 1 610
box -4 -6 84 206
use FILL  SFILL6160x6100
timestamp 1591628762
transform 1 0 616 0 1 610
box -4 -6 20 206
use FILL  SFILL6320x6100
timestamp 1591628762
transform 1 0 632 0 1 610
box -4 -6 20 206
use FILL  SFILL6480x6100
timestamp 1591628762
transform 1 0 648 0 1 610
box -4 -6 20 206
use FILL  SFILL6640x6100
timestamp 1591628762
transform 1 0 664 0 1 610
box -4 -6 20 206
use OAI21X1  _153_
timestamp 1591628762
transform 1 0 888 0 1 610
box -4 -6 68 206
use NAND2X1  _152_
timestamp 1591628762
transform -1 0 1000 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert10
timestamp 1591628762
transform -1 0 1048 0 1 610
box -4 -6 52 206
use DFFPOSX1  _288_
timestamp 1591628762
transform -1 0 1240 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert9
timestamp 1591628762
transform 1 0 1240 0 1 610
box -4 -6 52 206
use OAI21X1  _163_
timestamp 1591628762
transform -1 0 1352 0 1 610
box -4 -6 68 206
use OAI21X1  _114_
timestamp 1591628762
transform 1 0 1352 0 1 610
box -4 -6 68 206
use NAND2X1  _113_
timestamp 1591628762
transform -1 0 1464 0 1 610
box -4 -6 52 206
use AOI22X1  _162_
timestamp 1591628762
transform -1 0 1544 0 1 610
box -4 -6 84 206
use NOR2X1  _112_
timestamp 1591628762
transform 1 0 1544 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert6
timestamp 1591628762
transform 1 0 1592 0 1 610
box -4 -6 52 206
use NAND2X1  _122_
timestamp 1591628762
transform -1 0 1688 0 1 610
box -4 -6 52 206
use DFFPOSX1  _278_
timestamp 1591628762
transform 1 0 1752 0 1 610
box -4 -6 196 206
use FILL  SFILL16880x6100
timestamp 1591628762
transform 1 0 1688 0 1 610
box -4 -6 20 206
use FILL  SFILL17040x6100
timestamp 1591628762
transform 1 0 1704 0 1 610
box -4 -6 20 206
use FILL  SFILL17200x6100
timestamp 1591628762
transform 1 0 1720 0 1 610
box -4 -6 20 206
use FILL  SFILL17360x6100
timestamp 1591628762
transform 1 0 1736 0 1 610
box -4 -6 20 206
use NAND2X1  _174_
timestamp 1591628762
transform 1 0 1944 0 1 610
box -4 -6 52 206
use OAI21X1  _179_
timestamp 1591628762
transform 1 0 1992 0 1 610
box -4 -6 68 206
use NAND2X1  _166_
timestamp 1591628762
transform 1 0 2056 0 1 610
box -4 -6 52 206
use AOI22X1  _167_
timestamp 1591628762
transform -1 0 2184 0 1 610
box -4 -6 84 206
use DFFPOSX1  _262_
timestamp 1591628762
transform 1 0 2184 0 1 610
box -4 -6 196 206
use FILL  FILL22480x6100
timestamp 1591628762
transform 1 0 2376 0 1 610
box -4 -6 20 206
use DFFPOSX1  _286_
timestamp 1591628762
transform -1 0 200 0 -1 1010
box -4 -6 196 206
use NAND2X1  _146_
timestamp 1591628762
transform -1 0 248 0 -1 1010
box -4 -6 52 206
use OAI21X1  _147_
timestamp 1591628762
transform -1 0 312 0 -1 1010
box -4 -6 68 206
use OAI21X1  _219_
timestamp 1591628762
transform -1 0 376 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _283_
timestamp 1591628762
transform 1 0 376 0 -1 1010
box -4 -6 196 206
use NAND2X1  _202_
timestamp 1591628762
transform 1 0 568 0 -1 1010
box -4 -6 52 206
use NAND2X1  _137_
timestamp 1591628762
transform 1 0 680 0 -1 1010
box -4 -6 52 206
use OAI21X1  _138_
timestamp 1591628762
transform -1 0 792 0 -1 1010
box -4 -6 68 206
use NOR3X1  _207_
timestamp 1591628762
transform -1 0 920 0 -1 1010
box -4 -6 132 206
use FILL  SFILL6160x8100
timestamp 1591628762
transform -1 0 632 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6320x8100
timestamp 1591628762
transform -1 0 648 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6480x8100
timestamp 1591628762
transform -1 0 664 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6640x8100
timestamp 1591628762
transform -1 0 680 0 -1 1010
box -4 -6 20 206
use NOR2X1  _198_
timestamp 1591628762
transform -1 0 968 0 -1 1010
box -4 -6 52 206
use AND2X2  _197_
timestamp 1591628762
transform 1 0 968 0 -1 1010
box -4 -6 68 206
use OAI21X1  _135_
timestamp 1591628762
transform 1 0 1032 0 -1 1010
box -4 -6 68 206
use NAND2X1  _134_
timestamp 1591628762
transform -1 0 1144 0 -1 1010
box -4 -6 52 206
use NAND2X1  _196_
timestamp 1591628762
transform 1 0 1144 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _282_
timestamp 1591628762
transform 1 0 1192 0 -1 1010
box -4 -6 196 206
use BUFX2  BUFX2_insert13
timestamp 1591628762
transform -1 0 1432 0 -1 1010
box -4 -6 52 206
use OAI21X1  _144_
timestamp 1591628762
transform 1 0 1432 0 -1 1010
box -4 -6 68 206
use NAND2X1  _143_
timestamp 1591628762
transform -1 0 1544 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _285_
timestamp 1591628762
transform -1 0 1736 0 -1 1010
box -4 -6 196 206
use OAI21X1  _141_
timestamp 1591628762
transform 1 0 1800 0 -1 1010
box -4 -6 68 206
use FILL  SFILL17360x8100
timestamp 1591628762
transform -1 0 1752 0 -1 1010
box -4 -6 20 206
use FILL  SFILL17520x8100
timestamp 1591628762
transform -1 0 1768 0 -1 1010
box -4 -6 20 206
use FILL  SFILL17680x8100
timestamp 1591628762
transform -1 0 1784 0 -1 1010
box -4 -6 20 206
use FILL  SFILL17840x8100
timestamp 1591628762
transform -1 0 1800 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  _284_
timestamp 1591628762
transform -1 0 2056 0 -1 1010
box -4 -6 196 206
use INVX1  _115_
timestamp 1591628762
transform -1 0 2088 0 -1 1010
box -4 -6 36 206
use NAND2X1  _164_
timestamp 1591628762
transform 1 0 2088 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _261_
timestamp 1591628762
transform 1 0 2136 0 -1 1010
box -4 -6 196 206
use BUFX2  _245_
timestamp 1591628762
transform 1 0 2328 0 -1 1010
box -4 -6 52 206
use FILL  FILL22480x8100
timestamp 1591628762
transform -1 0 2392 0 -1 1010
box -4 -6 20 206
use BUFX2  _255_
timestamp 1591628762
transform -1 0 56 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _271_
timestamp 1591628762
transform -1 0 248 0 1 1010
box -4 -6 196 206
use AOI22X1  _220_
timestamp 1591628762
transform -1 0 328 0 1 1010
box -4 -6 84 206
use INVX2  _145_
timestamp 1591628762
transform 1 0 328 0 1 1010
box -4 -6 36 206
use OAI21X1  _221_
timestamp 1591628762
transform -1 0 424 0 1 1010
box -4 -6 68 206
use AND2X2  _218_
timestamp 1591628762
transform -1 0 488 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _267_
timestamp 1591628762
transform 1 0 488 0 1 1010
box -4 -6 196 206
use NAND2X1  _206_
timestamp 1591628762
transform 1 0 744 0 1 1010
box -4 -6 52 206
use INVX2  _136_
timestamp 1591628762
transform -1 0 824 0 1 1010
box -4 -6 36 206
use FILL  SFILL6800x10100
timestamp 1591628762
transform 1 0 680 0 1 1010
box -4 -6 20 206
use FILL  SFILL6960x10100
timestamp 1591628762
transform 1 0 696 0 1 1010
box -4 -6 20 206
use FILL  SFILL7120x10100
timestamp 1591628762
transform 1 0 712 0 1 1010
box -4 -6 20 206
use FILL  SFILL7280x10100
timestamp 1591628762
transform 1 0 728 0 1 1010
box -4 -6 20 206
use OAI21X1  _205_
timestamp 1591628762
transform 1 0 824 0 1 1010
box -4 -6 68 206
use OAI21X1  _204_
timestamp 1591628762
transform 1 0 888 0 1 1010
box -4 -6 68 206
use INVX1  _199_
timestamp 1591628762
transform 1 0 952 0 1 1010
box -4 -6 36 206
use OAI21X1  _203_
timestamp 1591628762
transform 1 0 984 0 1 1010
box -4 -6 68 206
use INVX2  _133_
timestamp 1591628762
transform -1 0 1080 0 1 1010
box -4 -6 36 206
use AOI22X1  _200_
timestamp 1591628762
transform 1 0 1080 0 1 1010
box -4 -6 84 206
use OAI21X1  _201_
timestamp 1591628762
transform 1 0 1160 0 1 1010
box -4 -6 68 206
use NAND3X1  _217_
timestamp 1591628762
transform -1 0 1288 0 1 1010
box -4 -6 68 206
use NAND2X1  _209_
timestamp 1591628762
transform 1 0 1288 0 1 1010
box -4 -6 52 206
use NAND2X1  _210_
timestamp 1591628762
transform -1 0 1384 0 1 1010
box -4 -6 52 206
use OAI21X1  _214_
timestamp 1591628762
transform -1 0 1448 0 1 1010
box -4 -6 68 206
use INVX1  _142_
timestamp 1591628762
transform -1 0 1480 0 1 1010
box -4 -6 36 206
use AOI22X1  _215_
timestamp 1591628762
transform 1 0 1480 0 1 1010
box -4 -6 84 206
use AOI22X1  _211_
timestamp 1591628762
transform 1 0 1560 0 1 1010
box -4 -6 84 206
use INVX1  _139_
timestamp 1591628762
transform 1 0 1640 0 1 1010
box -4 -6 36 206
use NAND2X1  _140_
timestamp 1591628762
transform 1 0 1672 0 1 1010
box -4 -6 52 206
use NAND2X1  _116_
timestamp 1591628762
transform -1 0 1832 0 1 1010
box -4 -6 52 206
use FILL  SFILL17200x10100
timestamp 1591628762
transform 1 0 1720 0 1 1010
box -4 -6 20 206
use FILL  SFILL17360x10100
timestamp 1591628762
transform 1 0 1736 0 1 1010
box -4 -6 20 206
use FILL  SFILL17520x10100
timestamp 1591628762
transform 1 0 1752 0 1 1010
box -4 -6 20 206
use FILL  SFILL17680x10100
timestamp 1591628762
transform 1 0 1768 0 1 1010
box -4 -6 20 206
use OAI21X1  _117_
timestamp 1591628762
transform -1 0 1896 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _276_
timestamp 1591628762
transform 1 0 1896 0 1 1010
box -4 -6 196 206
use DFFPOSX1  _260_
timestamp 1591628762
transform 1 0 2088 0 1 1010
box -4 -6 196 206
use BUFX2  _244_
timestamp 1591628762
transform 1 0 2280 0 1 1010
box -4 -6 52 206
use NOR2X1  _165_
timestamp 1591628762
transform 1 0 2328 0 1 1010
box -4 -6 52 206
use FILL  FILL22480x10100
timestamp 1591628762
transform 1 0 2376 0 1 1010
box -4 -6 20 206
use BUFX2  _258_
timestamp 1591628762
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _274_
timestamp 1591628762
transform -1 0 248 0 -1 1410
box -4 -6 196 206
use BUFX2  _254_
timestamp 1591628762
transform -1 0 296 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _270_
timestamp 1591628762
transform -1 0 488 0 -1 1410
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert1
timestamp 1591628762
transform -1 0 632 0 -1 1410
box -4 -6 148 206
use BUFX2  _251_
timestamp 1591628762
transform 1 0 696 0 -1 1410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert2
timestamp 1591628762
transform 1 0 744 0 -1 1410
box -4 -6 148 206
use FILL  SFILL6320x12100
timestamp 1591628762
transform -1 0 648 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6480x12100
timestamp 1591628762
transform -1 0 664 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6640x12100
timestamp 1591628762
transform -1 0 680 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6800x12100
timestamp 1591628762
transform -1 0 696 0 -1 1410
box -4 -6 20 206
use BUFX2  _249_
timestamp 1591628762
transform -1 0 936 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _265_
timestamp 1591628762
transform -1 0 1128 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _266_
timestamp 1591628762
transform 1 0 1128 0 -1 1410
box -4 -6 196 206
use BUFX2  _250_
timestamp 1591628762
transform 1 0 1320 0 -1 1410
box -4 -6 52 206
use AOI21X1  _213_
timestamp 1591628762
transform 1 0 1368 0 -1 1410
box -4 -6 68 206
use OAI21X1  _216_
timestamp 1591628762
transform 1 0 1432 0 -1 1410
box -4 -6 68 206
use NOR2X1  _208_
timestamp 1591628762
transform -1 0 1544 0 -1 1410
box -4 -6 52 206
use OAI21X1  _212_
timestamp 1591628762
transform 1 0 1544 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _269_
timestamp 1591628762
transform 1 0 1608 0 -1 1410
box -4 -6 196 206
use FILL  SFILL18000x12100
timestamp 1591628762
transform -1 0 1816 0 -1 1410
box -4 -6 20 206
use BUFX2  _253_
timestamp 1591628762
transform 1 0 1864 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _268_
timestamp 1591628762
transform 1 0 1912 0 -1 1410
box -4 -6 196 206
use FILL  SFILL18160x12100
timestamp 1591628762
transform -1 0 1832 0 -1 1410
box -4 -6 20 206
use FILL  SFILL18320x12100
timestamp 1591628762
transform -1 0 1848 0 -1 1410
box -4 -6 20 206
use FILL  SFILL18480x12100
timestamp 1591628762
transform -1 0 1864 0 -1 1410
box -4 -6 20 206
use BUFX2  _252_
timestamp 1591628762
transform 1 0 2104 0 -1 1410
box -4 -6 52 206
use NAND2X1  _125_
timestamp 1591628762
transform -1 0 2200 0 -1 1410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert0
timestamp 1591628762
transform -1 0 2344 0 -1 1410
box -4 -6 148 206
use BUFX2  _246_
timestamp 1591628762
transform 1 0 2344 0 -1 1410
box -4 -6 52 206
<< labels >>
flabel metal4 s 1728 -10 1792 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 592 -10 656 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 2301 1457 2307 1463 3 FreeSans 24 90 0 0 clock
port 2 nsew
flabel metal2 s 1053 -23 1059 -17 7 FreeSans 24 270 0 0 opcode[1]
port 3 nsew
flabel metal2 s 957 -23 963 -17 7 FreeSans 24 270 0 0 opcode[0]
port 4 nsew
flabel metal2 s 301 -23 307 -17 7 FreeSans 24 270 0 0 pc_in[15]
port 5 nsew
flabel metal2 s 445 -23 451 -17 7 FreeSans 24 270 0 0 pc_in[14]
port 6 nsew
flabel metal2 s 493 -23 499 -17 7 FreeSans 24 270 0 0 pc_in[13]
port 7 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 pc_in[12]
port 8 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 pc_in[11]
port 9 nsew
flabel metal2 s 1421 1457 1427 1463 3 FreeSans 24 90 0 0 pc_in[10]
port 10 nsew
flabel metal2 s 1533 1457 1539 1463 3 FreeSans 24 90 0 0 pc_in[9]
port 11 nsew
flabel metal2 s 845 1457 851 1463 3 FreeSans 24 90 0 0 pc_in[8]
port 12 nsew
flabel metal2 s 1101 1457 1107 1463 3 FreeSans 24 90 0 0 pc_in[7]
port 13 nsew
flabel metal2 s 925 -23 931 -17 7 FreeSans 24 270 0 0 pc_in[6]
port 14 nsew
flabel metal2 s 1469 -23 1475 -17 7 FreeSans 24 270 0 0 pc_in[5]
port 15 nsew
flabel metal2 s 1901 -23 1907 -17 7 FreeSans 24 270 0 0 pc_in[4]
port 16 nsew
flabel metal2 s 1853 -23 1859 -17 7 FreeSans 24 270 0 0 pc_in[3]
port 17 nsew
flabel metal3 s 2429 497 2435 503 3 FreeSans 24 0 0 0 pc_in[2]
port 18 nsew
flabel metal3 s 2429 917 2435 923 3 FreeSans 24 0 0 0 pc_in[1]
port 19 nsew
flabel metal3 s 2429 1057 2435 1063 3 FreeSans 24 0 0 0 pc_in[0]
port 20 nsew
flabel metal3 s -35 1297 -29 1303 7 FreeSans 24 0 0 0 pc_out[15]
port 21 nsew
flabel metal3 s -35 97 -29 103 7 FreeSans 24 0 0 0 pc_out[14]
port 22 nsew
flabel metal3 s -35 697 -29 703 7 FreeSans 24 0 0 0 pc_out[13]
port 23 nsew
flabel metal3 s -35 1137 -29 1143 7 FreeSans 24 0 0 0 pc_out[12]
port 24 nsew
flabel metal2 s 269 1457 275 1463 3 FreeSans 24 90 0 0 pc_out[11]
port 25 nsew
flabel metal2 s 1885 1457 1891 1463 3 FreeSans 24 90 0 0 pc_out[10]
port 26 nsew
flabel metal2 s 2125 1457 2131 1463 3 FreeSans 24 90 0 0 pc_out[9]
port 27 nsew
flabel metal2 s 717 1457 723 1463 3 FreeSans 24 90 0 0 pc_out[8]
port 28 nsew
flabel metal2 s 1341 1457 1347 1463 3 FreeSans 24 90 0 0 pc_out[7]
port 29 nsew
flabel metal2 s 909 1457 915 1463 3 FreeSans 24 90 0 0 pc_out[6]
port 30 nsew
flabel metal2 s 1517 -23 1523 -17 7 FreeSans 24 270 0 0 pc_out[5]
port 31 nsew
flabel metal2 s 1565 -23 1571 -17 7 FreeSans 24 270 0 0 pc_out[4]
port 32 nsew
flabel metal3 s 2429 1297 2435 1303 3 FreeSans 24 0 0 0 pc_out[3]
port 33 nsew
flabel metal3 s 2429 957 2435 963 3 FreeSans 24 0 0 0 pc_out[2]
port 34 nsew
flabel metal3 s 2429 1097 2435 1103 3 FreeSans 24 0 0 0 pc_out[1]
port 35 nsew
flabel metal2 s 893 -23 899 -17 7 FreeSans 24 270 0 0 pc_out[0]
port 36 nsew
<< end >>
