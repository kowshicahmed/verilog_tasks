magic
tech scmos
magscale 1 2
timestamp 1591630448
<< metal1 >>
rect 442 1214 454 1216
rect 427 1206 429 1214
rect 437 1206 439 1214
rect 447 1206 449 1214
rect 457 1206 459 1214
rect 467 1206 469 1214
rect 442 1204 454 1206
rect 60 1132 68 1136
rect 140 1132 148 1136
rect 844 1132 852 1136
rect 1036 1132 1044 1136
rect 1084 1132 1092 1136
rect 1276 1132 1284 1136
rect 77 1117 108 1123
rect 996 1116 1004 1124
rect 189 1097 204 1103
rect 221 1097 259 1103
rect 388 1097 419 1103
rect 1021 1103 1027 1123
rect 957 1097 995 1103
rect 1021 1097 1059 1103
rect 1284 1097 1299 1103
rect 1564 1103 1572 1106
rect 1564 1097 1587 1103
rect 93 1077 108 1083
rect 858 1036 860 1044
rect 1098 1036 1100 1044
rect 1268 1036 1270 1044
rect 1210 1014 1222 1016
rect 1195 1006 1197 1014
rect 1205 1006 1207 1014
rect 1215 1006 1217 1014
rect 1225 1006 1227 1014
rect 1235 1006 1237 1014
rect 1210 1004 1222 1006
rect 436 937 468 943
rect 1197 937 1283 943
rect 221 917 259 923
rect 333 917 371 923
rect 1005 917 1036 923
rect 1197 923 1203 937
rect 1165 917 1203 923
rect 1325 917 1363 923
rect 292 897 307 903
rect 442 814 454 816
rect 427 806 429 814
rect 437 806 439 814
rect 447 806 449 814
rect 457 806 459 814
rect 467 806 469 814
rect 442 804 454 806
rect 1517 737 1532 743
rect 1005 697 1043 703
rect 1149 697 1164 703
rect 1405 697 1420 703
rect 1549 697 1587 703
rect 333 677 355 683
rect 1261 637 1324 643
rect 1210 614 1222 616
rect 1195 606 1197 614
rect 1205 606 1207 614
rect 1215 606 1217 614
rect 1225 606 1227 614
rect 1235 606 1237 614
rect 1210 604 1222 606
rect 1188 577 1251 583
rect 1556 576 1558 584
rect 1469 537 1491 543
rect 45 517 60 523
rect 244 517 275 523
rect 909 517 940 523
rect 1053 517 1091 523
rect 1277 517 1315 523
rect 1380 517 1395 523
rect 1372 484 1380 488
rect 1021 477 1036 483
rect 1564 484 1572 488
rect 548 437 563 443
rect 442 414 454 416
rect 427 406 429 414
rect 437 406 439 414
rect 447 406 449 414
rect 457 406 459 414
rect 467 406 469 414
rect 442 404 454 406
rect 29 317 60 323
rect 1645 317 1660 323
rect 77 297 92 303
rect 221 297 252 303
rect 733 297 787 303
rect 1053 297 1084 303
rect 1453 297 1491 303
rect 749 277 764 283
rect 340 237 396 243
rect 1546 236 1548 244
rect 1210 214 1222 216
rect 1195 206 1197 214
rect 1205 206 1207 214
rect 1215 206 1217 214
rect 1225 206 1227 214
rect 1235 206 1237 214
rect 1210 204 1222 206
rect 164 117 179 123
rect 308 117 323 123
rect 452 117 515 123
rect 813 117 851 123
rect 877 117 915 123
rect 877 97 883 117
rect 932 117 947 123
rect 1053 117 1091 123
rect 1117 117 1155 123
rect 1085 97 1091 117
rect 1172 117 1251 123
rect 1453 117 1484 123
rect 348 84 356 88
rect 588 84 596 88
rect 892 84 900 88
rect 781 77 796 83
rect 1068 84 1076 88
rect 429 37 492 43
rect 442 14 454 16
rect 427 6 429 14
rect 437 6 439 14
rect 447 6 449 14
rect 457 6 459 14
rect 467 6 469 14
rect 442 4 454 6
<< m2contact >>
rect 419 1206 427 1214
rect 429 1206 437 1214
rect 439 1206 447 1214
rect 449 1206 457 1214
rect 459 1206 467 1214
rect 469 1206 477 1214
rect 156 1176 164 1184
rect 588 1176 596 1184
rect 636 1176 644 1184
rect 924 1176 932 1184
rect 1164 1176 1172 1184
rect 1324 1176 1332 1184
rect 1372 1176 1380 1184
rect 1612 1176 1620 1184
rect 60 1136 68 1144
rect 140 1136 148 1144
rect 300 1136 308 1144
rect 828 1136 836 1144
rect 844 1136 852 1144
rect 1036 1136 1044 1144
rect 1084 1136 1092 1144
rect 1276 1136 1284 1144
rect 108 1116 116 1124
rect 284 1116 292 1124
rect 988 1116 996 1124
rect 44 1096 52 1104
rect 204 1096 212 1104
rect 380 1096 388 1104
rect 556 1096 564 1104
rect 604 1096 612 1104
rect 716 1096 724 1104
rect 892 1096 900 1104
rect 1132 1096 1140 1104
rect 1276 1096 1284 1104
rect 1340 1096 1348 1104
rect 1452 1096 1460 1104
rect 12 1076 20 1084
rect 108 1076 116 1084
rect 236 1076 244 1084
rect 284 1076 292 1084
rect 668 1076 676 1084
rect 876 1076 884 1084
rect 972 1076 980 1084
rect 1068 1076 1076 1084
rect 1116 1076 1124 1084
rect 1244 1076 1252 1084
rect 1404 1076 1412 1084
rect 204 1056 212 1064
rect 428 1056 436 1064
rect 940 1056 948 1064
rect 140 1036 148 1044
rect 860 1036 868 1044
rect 1100 1036 1108 1044
rect 1260 1036 1268 1044
rect 1564 1036 1572 1044
rect 1187 1006 1195 1014
rect 1197 1006 1205 1014
rect 1207 1006 1215 1014
rect 1217 1006 1225 1014
rect 1227 1006 1235 1014
rect 1237 1006 1245 1014
rect 12 976 20 984
rect 636 976 644 984
rect 652 976 660 984
rect 1116 976 1124 984
rect 1628 976 1636 984
rect 204 956 212 964
rect 380 956 388 964
rect 844 956 852 964
rect 1260 956 1268 964
rect 1372 956 1380 964
rect 172 936 180 944
rect 236 936 244 944
rect 348 936 356 944
rect 428 936 436 944
rect 924 936 932 944
rect 956 936 964 944
rect 1180 936 1188 944
rect 140 918 148 926
rect 268 916 276 924
rect 316 916 324 924
rect 508 918 516 926
rect 572 916 580 924
rect 716 916 724 924
rect 780 918 788 926
rect 892 916 900 924
rect 908 916 916 924
rect 1036 916 1044 924
rect 1148 916 1156 924
rect 1340 936 1348 944
rect 1404 936 1412 944
rect 1580 936 1588 944
rect 1308 916 1316 924
rect 1436 918 1444 926
rect 1596 916 1604 924
rect 284 896 292 904
rect 860 896 868 904
rect 876 896 884 904
rect 1132 896 1140 904
rect 1292 896 1300 904
rect 1628 896 1636 904
rect 1564 836 1572 844
rect 419 806 427 814
rect 429 806 437 814
rect 439 806 447 814
rect 449 806 457 814
rect 459 806 467 814
rect 469 806 477 814
rect 348 776 356 784
rect 572 776 580 784
rect 716 776 724 784
rect 780 776 788 784
rect 12 736 20 744
rect 60 736 68 744
rect 1532 736 1540 744
rect 284 716 292 724
rect 1068 716 1076 724
rect 1612 716 1620 724
rect 44 696 52 704
rect 188 694 196 702
rect 300 696 308 704
rect 316 696 324 704
rect 380 696 388 704
rect 748 696 756 704
rect 860 696 868 704
rect 924 694 932 702
rect 1052 696 1060 704
rect 1164 696 1172 704
rect 1420 696 1428 704
rect 1596 696 1604 704
rect 172 676 180 684
rect 268 676 276 684
rect 460 676 468 684
rect 604 676 612 684
rect 956 676 964 684
rect 1020 676 1028 684
rect 1100 676 1108 684
rect 1356 676 1364 684
rect 1404 676 1412 684
rect 1564 676 1572 684
rect 252 656 260 664
rect 988 656 996 664
rect 1532 656 1540 664
rect 796 636 804 644
rect 1324 636 1332 644
rect 1187 606 1195 614
rect 1197 606 1205 614
rect 1207 606 1215 614
rect 1217 606 1225 614
rect 1227 606 1235 614
rect 1237 606 1245 614
rect 156 576 164 584
rect 1180 576 1188 584
rect 1420 576 1428 584
rect 1548 576 1556 584
rect 1612 576 1620 584
rect 60 556 68 564
rect 1036 556 1044 564
rect 1116 556 1124 564
rect 1324 556 1332 564
rect 1356 556 1364 564
rect 1596 556 1604 564
rect 76 536 84 544
rect 140 536 148 544
rect 268 536 276 544
rect 316 536 324 544
rect 348 536 356 544
rect 476 536 484 544
rect 604 536 612 544
rect 732 536 740 544
rect 860 536 868 544
rect 1068 536 1076 544
rect 1164 536 1172 544
rect 1292 536 1300 544
rect 1340 536 1348 544
rect 1532 536 1540 544
rect 60 516 68 524
rect 108 516 116 524
rect 124 516 132 524
rect 236 516 244 524
rect 588 516 596 524
rect 748 516 756 524
rect 828 516 836 524
rect 940 516 948 524
rect 1132 516 1140 524
rect 1372 516 1380 524
rect 1436 516 1444 524
rect 1644 516 1652 524
rect 92 496 100 504
rect 1116 496 1124 504
rect 1244 496 1252 504
rect 1516 496 1524 504
rect 12 476 20 484
rect 1036 476 1044 484
rect 1372 476 1380 484
rect 1564 476 1572 484
rect 540 436 548 444
rect 780 436 788 444
rect 796 436 804 444
rect 1468 436 1476 444
rect 1500 436 1508 444
rect 1580 436 1588 444
rect 419 406 427 414
rect 429 406 437 414
rect 439 406 447 414
rect 449 406 457 414
rect 459 406 467 414
rect 469 406 477 414
rect 1580 376 1588 384
rect 1628 376 1636 384
rect 12 316 20 324
rect 60 316 68 324
rect 92 316 100 324
rect 636 316 644 324
rect 700 316 708 324
rect 1516 316 1524 324
rect 1532 316 1540 324
rect 1660 316 1668 324
rect 92 296 100 304
rect 124 296 132 304
rect 252 296 260 304
rect 268 296 276 304
rect 476 296 484 304
rect 524 296 532 304
rect 668 296 676 304
rect 716 296 724 304
rect 844 294 852 302
rect 1084 296 1092 304
rect 1100 296 1108 304
rect 1308 296 1316 304
rect 1372 294 1380 302
rect 1500 296 1508 304
rect 44 276 52 284
rect 140 276 148 284
rect 172 276 180 284
rect 572 276 580 284
rect 620 276 628 284
rect 636 276 644 284
rect 684 276 692 284
rect 764 276 772 284
rect 860 276 868 284
rect 1004 276 1012 284
rect 1404 276 1412 284
rect 1468 276 1476 284
rect 1564 276 1572 284
rect 1612 276 1620 284
rect 60 256 68 264
rect 604 256 612 264
rect 764 256 772 264
rect 1436 256 1444 264
rect 1596 256 1604 264
rect 92 236 100 244
rect 332 236 340 244
rect 396 236 404 244
rect 412 236 420 244
rect 972 236 980 244
rect 1164 236 1172 244
rect 1244 236 1252 244
rect 1548 236 1556 244
rect 1187 206 1195 214
rect 1197 206 1205 214
rect 1207 206 1215 214
rect 1217 206 1225 214
rect 1227 206 1235 214
rect 1237 206 1245 214
rect 300 176 308 184
rect 588 176 596 184
rect 1084 176 1092 184
rect 332 156 340 164
rect 796 156 804 164
rect 1164 156 1172 164
rect 1436 156 1444 164
rect 172 136 180 144
rect 252 136 260 144
rect 380 136 388 144
rect 556 136 564 144
rect 620 136 628 144
rect 828 136 836 144
rect 860 136 868 144
rect 924 136 932 144
rect 1036 136 1044 144
rect 1132 136 1140 144
rect 1580 136 1588 144
rect 44 116 52 124
rect 156 116 164 124
rect 268 116 276 124
rect 300 116 308 124
rect 396 116 404 124
rect 444 116 452 124
rect 668 116 676 124
rect 300 96 308 104
rect 364 96 372 104
rect 924 116 932 124
rect 988 116 996 124
rect 1164 116 1172 124
rect 1292 116 1300 124
rect 1372 116 1380 124
rect 1484 116 1492 124
rect 1596 116 1604 124
rect 1612 116 1620 124
rect 1628 96 1636 104
rect 12 76 20 84
rect 60 76 68 84
rect 348 76 356 84
rect 588 76 596 84
rect 796 76 804 84
rect 892 76 900 84
rect 1068 76 1076 84
rect 1564 76 1572 84
rect 492 36 500 44
rect 540 36 548 44
rect 972 36 980 44
rect 1020 36 1028 44
rect 1276 36 1284 44
rect 1324 36 1332 44
rect 1340 36 1348 44
rect 419 6 427 14
rect 429 6 437 14
rect 439 6 447 14
rect 449 6 457 14
rect 459 6 467 14
rect 469 6 477 14
<< metal2 >>
rect 125 1257 147 1263
rect 141 1144 147 1257
rect 157 1257 179 1263
rect 573 1257 595 1263
rect 621 1257 643 1263
rect 157 1184 163 1257
rect 442 1214 454 1216
rect 427 1206 429 1214
rect 437 1206 439 1214
rect 447 1206 449 1214
rect 457 1206 459 1214
rect 467 1206 469 1214
rect 442 1204 454 1206
rect 589 1184 595 1257
rect 637 1184 643 1257
rect 845 1257 867 1263
rect 909 1257 931 1263
rect 845 1144 851 1257
rect 925 1184 931 1257
rect 1037 1257 1059 1263
rect 1085 1257 1107 1263
rect 1149 1257 1171 1263
rect 1037 1144 1043 1257
rect 1085 1144 1091 1257
rect 1165 1184 1171 1257
rect 1277 1144 1283 1263
rect 1309 1257 1331 1263
rect 1357 1257 1379 1263
rect 1597 1257 1619 1263
rect 1325 1184 1331 1257
rect 1373 1184 1379 1257
rect 1613 1184 1619 1257
rect 205 1104 211 1136
rect 717 1104 723 1116
rect 829 1104 835 1136
rect 13 1084 19 1096
rect 45 984 51 1096
rect 205 1064 211 1096
rect 381 1084 387 1096
rect 141 964 147 1036
rect 205 964 211 976
rect 237 944 243 1076
rect 381 964 387 976
rect 173 924 179 936
rect 141 904 147 918
rect 45 737 60 743
rect 13 724 19 736
rect 45 704 51 737
rect 45 684 51 696
rect 173 684 179 916
rect 269 904 275 916
rect 285 904 291 956
rect 429 944 435 1056
rect 557 984 563 1096
rect 317 904 323 916
rect 349 784 355 936
rect 429 924 435 936
rect 573 924 579 1076
rect 605 1004 611 1096
rect 653 984 659 996
rect 845 964 851 996
rect 509 904 515 918
rect 861 923 867 1036
rect 925 944 931 1076
rect 941 1064 947 1096
rect 861 917 883 923
rect 442 814 454 816
rect 427 806 429 814
rect 437 806 439 814
rect 447 806 449 814
rect 457 806 459 814
rect 467 806 469 814
rect 442 804 454 806
rect 573 784 579 916
rect 717 784 723 916
rect 877 904 883 917
rect 909 904 915 916
rect 925 884 931 936
rect 781 784 787 876
rect 717 704 723 776
rect 317 684 323 696
rect 253 664 259 676
rect 61 564 67 576
rect 61 524 67 556
rect 125 524 131 536
rect 13 484 19 496
rect 93 324 99 496
rect 13 304 19 316
rect 141 284 147 536
rect 269 304 275 536
rect 381 524 387 696
rect 461 664 467 676
rect 461 543 467 656
rect 605 544 611 676
rect 461 537 476 543
rect 749 524 755 696
rect 957 684 963 936
rect 1085 743 1091 976
rect 1101 904 1107 1036
rect 1133 983 1139 1096
rect 1124 977 1139 983
rect 1133 964 1139 977
rect 1165 943 1171 1076
rect 1210 1014 1222 1016
rect 1195 1006 1197 1014
rect 1205 1006 1207 1014
rect 1215 1006 1217 1014
rect 1225 1006 1227 1014
rect 1235 1006 1237 1014
rect 1210 1004 1222 1006
rect 1261 984 1267 1036
rect 1165 937 1180 943
rect 1069 737 1091 743
rect 1069 724 1075 737
rect 989 644 995 656
rect 829 524 835 636
rect 442 414 454 416
rect 427 406 429 414
rect 437 406 439 414
rect 447 406 449 414
rect 457 406 459 414
rect 467 406 469 414
rect 442 404 454 406
rect 13 84 19 96
rect 45 83 51 116
rect 61 84 67 256
rect 141 144 147 276
rect 157 124 163 236
rect 173 144 179 276
rect 253 184 259 296
rect 333 164 339 236
rect 397 124 403 236
rect 445 124 451 236
rect 541 144 547 436
rect 637 284 643 296
rect 669 284 675 296
rect 573 144 579 276
rect 605 244 611 256
rect 701 224 707 316
rect 781 283 787 436
rect 797 343 803 436
rect 797 337 819 343
rect 772 277 787 283
rect 589 184 595 216
rect 548 137 556 143
rect 669 124 675 156
rect 781 144 787 277
rect 797 124 803 156
rect 797 84 803 116
rect 45 77 60 83
rect 349 -17 355 76
rect 442 14 454 16
rect 427 6 429 14
rect 437 6 439 14
rect 447 6 449 14
rect 457 6 459 14
rect 467 6 469 14
rect 442 4 454 6
rect 493 -17 499 36
rect 349 -23 371 -17
rect 493 -23 515 -17
rect 541 -23 547 36
rect 589 -17 595 76
rect 573 -23 595 -17
rect 813 -23 819 337
rect 861 284 867 536
rect 941 524 947 556
rect 1021 544 1027 676
rect 1037 564 1043 576
rect 1037 484 1043 556
rect 1101 304 1107 676
rect 1165 583 1171 696
rect 1210 614 1222 616
rect 1195 606 1197 614
rect 1205 606 1207 614
rect 1215 606 1217 614
rect 1225 606 1227 614
rect 1235 606 1237 614
rect 1210 604 1222 606
rect 1277 584 1283 1096
rect 1293 904 1299 976
rect 1341 964 1347 1096
rect 1341 884 1347 936
rect 1165 577 1180 583
rect 1245 504 1251 556
rect 1293 544 1299 876
rect 1373 844 1379 956
rect 1405 944 1411 1076
rect 1453 1064 1459 1096
rect 1405 684 1411 936
rect 1565 863 1571 1036
rect 1629 984 1635 1056
rect 1581 884 1587 936
rect 1565 857 1587 863
rect 1533 664 1539 736
rect 1325 564 1331 636
rect 1421 584 1427 656
rect 1325 504 1331 556
rect 1373 504 1379 516
rect 1117 484 1123 496
rect 1373 464 1379 476
rect 973 244 979 256
rect 980 237 995 243
rect 861 144 867 156
rect 989 124 995 237
rect 1085 184 1091 296
rect 1252 237 1267 243
rect 1165 164 1171 236
rect 1261 224 1267 237
rect 1210 214 1222 216
rect 1195 206 1197 214
rect 1205 206 1207 214
rect 1215 206 1217 214
rect 1225 206 1227 214
rect 1235 206 1237 214
rect 1210 204 1222 206
rect 1165 124 1171 156
rect 1293 124 1299 216
rect 1405 164 1411 276
rect 1437 224 1443 256
rect 1373 84 1379 116
rect 1453 84 1459 576
rect 1517 504 1523 596
rect 1533 564 1539 656
rect 1549 584 1555 716
rect 1533 504 1539 536
rect 1565 504 1571 676
rect 1581 543 1587 857
rect 1613 584 1619 616
rect 1597 564 1603 576
rect 1581 537 1603 543
rect 1501 444 1507 476
rect 1469 324 1475 436
rect 1501 323 1507 436
rect 1533 324 1539 496
rect 1565 437 1580 443
rect 1501 317 1516 323
rect 1469 284 1475 316
rect 1533 144 1539 316
rect 1565 303 1571 437
rect 1581 384 1587 416
rect 1565 297 1587 303
rect 1549 104 1555 236
rect 1581 163 1587 297
rect 1597 264 1603 537
rect 1613 284 1619 536
rect 1629 384 1635 896
rect 1645 524 1651 556
rect 1661 524 1667 696
rect 1581 157 1603 163
rect 1597 124 1603 157
rect 893 -17 899 76
rect 973 -17 979 36
rect 1021 -17 1027 36
rect 1069 -17 1075 76
rect 893 -23 915 -17
rect 957 -23 979 -17
rect 1005 -23 1027 -17
rect 1053 -23 1075 -17
rect 1277 -23 1283 36
rect 1325 -17 1331 36
rect 1309 -23 1331 -17
rect 1341 -17 1347 36
rect 1341 -23 1363 -17
<< m3contact >>
rect 419 1206 427 1214
rect 429 1206 437 1214
rect 439 1206 447 1214
rect 449 1206 457 1214
rect 459 1206 467 1214
rect 469 1206 477 1214
rect 60 1136 68 1144
rect 204 1136 212 1144
rect 300 1136 308 1144
rect 108 1116 116 1124
rect 284 1116 292 1124
rect 716 1116 724 1124
rect 988 1116 996 1124
rect 12 1096 20 1104
rect 828 1096 836 1104
rect 892 1096 900 1104
rect 940 1096 948 1104
rect 108 1076 116 1084
rect 236 1076 244 1084
rect 284 1076 292 1084
rect 380 1076 388 1084
rect 12 976 20 984
rect 44 976 52 984
rect 204 976 212 984
rect 140 956 148 964
rect 380 976 388 984
rect 284 956 292 964
rect 236 936 244 944
rect 172 916 180 924
rect 140 896 148 904
rect 12 716 20 724
rect 572 1076 580 1084
rect 556 976 564 984
rect 348 936 356 944
rect 268 896 276 904
rect 316 896 324 904
rect 428 916 436 924
rect 668 1076 676 1084
rect 876 1076 884 1084
rect 924 1076 932 1084
rect 604 996 612 1004
rect 652 996 660 1004
rect 844 996 852 1004
rect 636 976 644 984
rect 780 918 788 924
rect 780 916 788 918
rect 972 1076 980 1084
rect 1068 1076 1076 1084
rect 1116 1076 1124 1084
rect 1084 976 1092 984
rect 508 896 516 904
rect 419 806 427 814
rect 429 806 437 814
rect 439 806 447 814
rect 449 806 457 814
rect 459 806 467 814
rect 469 806 477 814
rect 892 916 900 924
rect 860 896 868 904
rect 908 896 916 904
rect 780 876 788 884
rect 924 876 932 884
rect 284 716 292 724
rect 188 702 196 704
rect 188 696 196 702
rect 300 696 308 704
rect 716 696 724 704
rect 860 696 868 704
rect 924 702 932 704
rect 924 696 932 702
rect 44 676 52 684
rect 252 676 260 684
rect 268 676 276 684
rect 316 676 324 684
rect 60 576 68 584
rect 156 576 164 584
rect 76 536 84 544
rect 124 536 132 544
rect 316 536 324 544
rect 348 536 356 544
rect 108 516 116 524
rect 12 496 20 504
rect 60 316 68 324
rect 92 316 100 324
rect 12 296 20 304
rect 92 296 100 304
rect 124 296 132 304
rect 236 516 244 524
rect 460 656 468 664
rect 476 536 484 544
rect 604 536 612 544
rect 732 536 740 544
rect 1036 916 1044 924
rect 1164 1076 1172 1084
rect 1244 1076 1252 1084
rect 1132 956 1140 964
rect 1187 1006 1195 1014
rect 1197 1006 1205 1014
rect 1207 1006 1215 1014
rect 1217 1006 1225 1014
rect 1227 1006 1235 1014
rect 1237 1006 1245 1014
rect 1260 976 1268 984
rect 1260 956 1268 964
rect 1148 916 1156 924
rect 1100 896 1108 904
rect 1132 896 1140 904
rect 1052 696 1060 704
rect 956 676 964 684
rect 796 636 804 644
rect 828 636 836 644
rect 988 636 996 644
rect 940 556 948 564
rect 860 536 868 544
rect 380 516 388 524
rect 588 516 596 524
rect 748 516 756 524
rect 419 406 427 414
rect 429 406 437 414
rect 439 406 447 414
rect 449 406 457 414
rect 459 406 467 414
rect 469 406 477 414
rect 268 296 276 304
rect 476 296 484 304
rect 524 296 532 304
rect 44 276 52 284
rect 140 276 148 284
rect 12 96 20 104
rect 92 236 100 244
rect 156 236 164 244
rect 140 136 148 144
rect 412 236 420 244
rect 444 236 452 244
rect 252 176 260 184
rect 300 176 308 184
rect 252 136 260 144
rect 380 136 388 144
rect 636 316 644 324
rect 700 316 708 324
rect 636 296 644 304
rect 620 276 628 284
rect 668 276 676 284
rect 684 276 692 284
rect 604 236 612 244
rect 716 296 724 304
rect 764 276 772 284
rect 764 256 772 264
rect 588 216 596 224
rect 700 216 708 224
rect 668 156 676 164
rect 540 136 548 144
rect 572 136 580 144
rect 620 136 628 144
rect 780 136 788 144
rect 268 116 276 124
rect 300 116 308 124
rect 796 116 804 124
rect 300 96 308 104
rect 364 96 372 104
rect 419 6 427 14
rect 429 6 437 14
rect 439 6 447 14
rect 449 6 457 14
rect 459 6 467 14
rect 469 6 477 14
rect 844 302 852 304
rect 844 296 852 302
rect 1036 576 1044 584
rect 1020 536 1028 544
rect 1068 536 1076 544
rect 1187 606 1195 614
rect 1197 606 1205 614
rect 1207 606 1215 614
rect 1217 606 1225 614
rect 1227 606 1235 614
rect 1237 606 1245 614
rect 1292 976 1300 984
rect 1340 956 1348 964
rect 1372 956 1380 964
rect 1308 916 1316 924
rect 1292 876 1300 884
rect 1340 876 1348 884
rect 1276 576 1284 584
rect 1116 556 1124 564
rect 1244 556 1252 564
rect 1164 536 1172 544
rect 1132 516 1140 524
rect 1452 1056 1460 1064
rect 1628 1056 1636 1064
rect 1372 836 1380 844
rect 1436 918 1444 924
rect 1436 916 1444 918
rect 1596 916 1604 924
rect 1580 876 1588 884
rect 1564 836 1572 844
rect 1420 696 1428 704
rect 1356 676 1364 684
rect 1548 716 1556 724
rect 1420 656 1428 664
rect 1516 596 1524 604
rect 1452 576 1460 584
rect 1356 556 1364 564
rect 1292 536 1300 544
rect 1340 536 1348 544
rect 1436 516 1444 524
rect 1324 496 1332 504
rect 1372 496 1380 504
rect 1116 476 1124 484
rect 1372 456 1380 464
rect 1100 296 1108 304
rect 1308 296 1316 304
rect 1372 302 1380 304
rect 1372 296 1380 302
rect 860 276 868 284
rect 1004 276 1012 284
rect 972 256 980 264
rect 860 156 868 164
rect 828 136 836 144
rect 924 136 932 144
rect 1260 216 1268 224
rect 1292 216 1300 224
rect 1187 206 1195 214
rect 1197 206 1205 214
rect 1207 206 1215 214
rect 1217 206 1225 214
rect 1227 206 1235 214
rect 1237 206 1245 214
rect 1036 136 1044 144
rect 1132 136 1140 144
rect 1436 216 1444 224
rect 1404 156 1412 164
rect 1436 156 1444 164
rect 924 116 932 124
rect 1532 556 1540 564
rect 1612 716 1620 724
rect 1596 696 1604 704
rect 1612 616 1620 624
rect 1596 576 1604 584
rect 1532 496 1540 504
rect 1564 496 1572 504
rect 1500 476 1508 484
rect 1468 316 1476 324
rect 1564 476 1572 484
rect 1532 316 1540 324
rect 1500 296 1508 304
rect 1580 416 1588 424
rect 1564 276 1572 284
rect 1532 136 1540 144
rect 1484 116 1492 124
rect 1612 536 1620 544
rect 1660 696 1668 704
rect 1644 556 1652 564
rect 1660 516 1668 524
rect 1660 316 1668 324
rect 1580 136 1588 144
rect 1612 116 1620 124
rect 1548 96 1556 104
rect 1628 96 1636 104
rect 1372 76 1380 84
rect 1452 76 1460 84
rect 1564 76 1572 84
<< metal3 >>
rect 418 1214 478 1216
rect 418 1206 419 1214
rect 428 1206 429 1214
rect 467 1206 468 1214
rect 477 1206 478 1214
rect 418 1204 478 1206
rect -35 1137 60 1143
rect 212 1137 300 1143
rect 116 1117 268 1123
rect 276 1117 284 1123
rect 724 1117 988 1123
rect -35 1097 12 1103
rect 836 1097 892 1103
rect 900 1097 940 1103
rect 116 1077 236 1083
rect 292 1077 380 1083
rect 580 1077 668 1083
rect 884 1077 924 1083
rect 932 1077 972 1083
rect 980 1077 1068 1083
rect 1076 1077 1116 1083
rect 1124 1077 1164 1083
rect 1172 1077 1244 1083
rect 1460 1057 1628 1063
rect 1186 1014 1246 1016
rect 1186 1006 1187 1014
rect 1196 1006 1197 1014
rect 1235 1006 1236 1014
rect 1245 1006 1246 1014
rect 1186 1004 1246 1006
rect 612 997 652 1003
rect 660 997 844 1003
rect 20 977 44 983
rect 52 977 204 983
rect 388 977 556 983
rect 564 977 636 983
rect 1092 977 1260 983
rect 1268 977 1292 983
rect 148 957 284 963
rect 1140 957 1260 963
rect 1348 957 1372 963
rect 244 937 348 943
rect 180 917 428 923
rect 788 917 892 923
rect 1044 917 1148 923
rect 1316 917 1436 923
rect 1604 917 1612 923
rect 148 897 268 903
rect 324 897 508 903
rect 868 897 908 903
rect 1108 897 1132 903
rect 788 877 924 883
rect 1300 877 1340 883
rect 1348 877 1580 883
rect 1380 837 1564 843
rect 418 814 478 816
rect 418 806 419 814
rect 428 806 429 814
rect 467 806 468 814
rect 477 806 478 814
rect 418 804 478 806
rect -35 717 12 723
rect 276 717 284 723
rect 1556 717 1612 723
rect 196 697 300 703
rect 724 697 860 703
rect 932 697 1052 703
rect 1428 697 1596 703
rect 1668 697 1699 703
rect -35 663 -29 683
rect 52 677 252 683
rect 276 677 316 683
rect 964 677 1356 683
rect -35 657 460 663
rect 1428 657 1699 663
rect 804 637 828 643
rect 836 637 988 643
rect 1620 617 1699 623
rect 1186 614 1246 616
rect 1186 606 1187 614
rect 1196 606 1197 614
rect 1235 606 1236 614
rect 1245 606 1246 614
rect 1186 604 1246 606
rect 1524 597 1644 603
rect 68 577 156 583
rect 1044 577 1276 583
rect 1460 577 1596 583
rect 948 557 1116 563
rect 1252 557 1356 563
rect 1540 557 1644 563
rect 1693 563 1699 583
rect 1693 557 1715 563
rect 84 537 124 543
rect 324 537 348 543
rect 484 537 604 543
rect 740 537 860 543
rect 1028 537 1068 543
rect 1076 537 1164 543
rect 1172 537 1292 543
rect 1300 537 1340 543
rect 1348 537 1612 543
rect 1652 537 1699 543
rect 116 517 236 523
rect 388 517 588 523
rect 596 517 748 523
rect 756 517 1132 523
rect 1140 517 1436 523
rect 1444 517 1660 523
rect -35 497 12 503
rect 1332 497 1372 503
rect 1540 497 1564 503
rect 1645 497 1699 503
rect 1124 477 1500 483
rect 1645 483 1651 497
rect 1572 477 1651 483
rect 1709 463 1715 557
rect 1380 457 1715 463
rect 1588 417 1612 423
rect 418 414 478 416
rect 418 406 419 414
rect 428 406 429 414
rect 467 406 468 414
rect 477 406 478 414
rect 418 404 478 406
rect 68 317 92 323
rect 644 317 700 323
rect 1476 317 1532 323
rect 1668 317 1699 323
rect -35 297 12 303
rect 100 297 124 303
rect 276 297 476 303
rect 532 297 636 303
rect 724 297 844 303
rect 1108 297 1308 303
rect 1380 297 1500 303
rect 52 277 140 283
rect 628 277 668 283
rect 692 277 764 283
rect 868 277 1004 283
rect 1572 277 1699 283
rect 772 257 972 263
rect 100 237 156 243
rect 420 237 444 243
rect 452 237 604 243
rect 596 217 700 223
rect 1268 217 1292 223
rect 1300 217 1436 223
rect 1186 214 1246 216
rect 1186 206 1187 214
rect 1196 206 1197 214
rect 1235 206 1236 214
rect 1245 206 1246 214
rect 1186 204 1246 206
rect 260 177 300 183
rect 676 157 860 163
rect 1412 157 1436 163
rect 148 137 252 143
rect 260 137 380 143
rect 388 137 540 143
rect 580 137 620 143
rect 788 137 828 143
rect 836 137 924 143
rect 932 137 1036 143
rect 1044 137 1132 143
rect 1540 137 1580 143
rect 276 117 300 123
rect 804 117 924 123
rect 1492 117 1612 123
rect -35 97 12 103
rect 308 97 364 103
rect 1556 97 1628 103
rect 1380 77 1452 83
rect 1460 77 1564 83
rect 418 14 478 16
rect 418 6 419 14
rect 428 6 429 14
rect 467 6 468 14
rect 477 6 478 14
rect 418 4 478 6
<< m4contact >>
rect 420 1206 427 1214
rect 427 1206 428 1214
rect 432 1206 437 1214
rect 437 1206 439 1214
rect 439 1206 440 1214
rect 444 1206 447 1214
rect 447 1206 449 1214
rect 449 1206 452 1214
rect 456 1206 457 1214
rect 457 1206 459 1214
rect 459 1206 464 1214
rect 468 1206 469 1214
rect 469 1206 476 1214
rect 268 1116 276 1124
rect 1188 1006 1195 1014
rect 1195 1006 1196 1014
rect 1200 1006 1205 1014
rect 1205 1006 1207 1014
rect 1207 1006 1208 1014
rect 1212 1006 1215 1014
rect 1215 1006 1217 1014
rect 1217 1006 1220 1014
rect 1224 1006 1225 1014
rect 1225 1006 1227 1014
rect 1227 1006 1232 1014
rect 1236 1006 1237 1014
rect 1237 1006 1244 1014
rect 1612 916 1620 924
rect 420 806 427 814
rect 427 806 428 814
rect 432 806 437 814
rect 437 806 439 814
rect 439 806 440 814
rect 444 806 447 814
rect 447 806 449 814
rect 449 806 452 814
rect 456 806 457 814
rect 457 806 459 814
rect 459 806 464 814
rect 468 806 469 814
rect 469 806 476 814
rect 268 716 276 724
rect 1188 606 1195 614
rect 1195 606 1196 614
rect 1200 606 1205 614
rect 1205 606 1207 614
rect 1207 606 1208 614
rect 1212 606 1215 614
rect 1215 606 1217 614
rect 1217 606 1220 614
rect 1224 606 1225 614
rect 1225 606 1227 614
rect 1227 606 1232 614
rect 1236 606 1237 614
rect 1237 606 1244 614
rect 1644 596 1652 604
rect 1644 536 1652 544
rect 1612 416 1620 424
rect 420 406 427 414
rect 427 406 428 414
rect 432 406 437 414
rect 437 406 439 414
rect 439 406 440 414
rect 444 406 447 414
rect 447 406 449 414
rect 449 406 452 414
rect 456 406 457 414
rect 457 406 459 414
rect 459 406 464 414
rect 468 406 469 414
rect 469 406 476 414
rect 1188 206 1195 214
rect 1195 206 1196 214
rect 1200 206 1205 214
rect 1205 206 1207 214
rect 1207 206 1208 214
rect 1212 206 1215 214
rect 1215 206 1217 214
rect 1217 206 1220 214
rect 1224 206 1225 214
rect 1225 206 1227 214
rect 1227 206 1232 214
rect 1236 206 1237 214
rect 1237 206 1244 214
rect 420 6 427 14
rect 427 6 428 14
rect 432 6 437 14
rect 437 6 439 14
rect 439 6 440 14
rect 444 6 447 14
rect 447 6 449 14
rect 449 6 452 14
rect 456 6 457 14
rect 457 6 459 14
rect 459 6 464 14
rect 468 6 469 14
rect 469 6 476 14
<< metal4 >>
rect 416 1214 480 1216
rect 416 1206 420 1214
rect 428 1206 432 1214
rect 440 1206 444 1214
rect 452 1206 456 1214
rect 464 1206 468 1214
rect 476 1206 480 1214
rect 266 1124 278 1126
rect 266 1116 268 1124
rect 276 1116 278 1124
rect 266 724 278 1116
rect 266 716 268 724
rect 276 716 278 724
rect 266 714 278 716
rect 416 814 480 1206
rect 416 806 420 814
rect 428 806 432 814
rect 440 806 444 814
rect 452 806 456 814
rect 464 806 468 814
rect 476 806 480 814
rect 416 414 480 806
rect 416 406 420 414
rect 428 406 432 414
rect 440 406 444 414
rect 452 406 456 414
rect 464 406 468 414
rect 476 406 480 414
rect 416 14 480 406
rect 416 6 420 14
rect 428 6 432 14
rect 440 6 444 14
rect 452 6 456 14
rect 464 6 468 14
rect 476 6 480 14
rect 416 -10 480 6
rect 1184 1014 1248 1216
rect 1184 1006 1188 1014
rect 1196 1006 1200 1014
rect 1208 1006 1212 1014
rect 1220 1006 1224 1014
rect 1232 1006 1236 1014
rect 1244 1006 1248 1014
rect 1184 614 1248 1006
rect 1184 606 1188 614
rect 1196 606 1200 614
rect 1208 606 1212 614
rect 1220 606 1224 614
rect 1232 606 1236 614
rect 1244 606 1248 614
rect 1184 214 1248 606
rect 1610 924 1622 926
rect 1610 916 1612 924
rect 1620 916 1622 924
rect 1610 424 1622 916
rect 1642 604 1654 606
rect 1642 596 1644 604
rect 1652 596 1654 604
rect 1642 544 1654 596
rect 1642 536 1644 544
rect 1652 536 1654 544
rect 1642 534 1654 536
rect 1610 416 1612 424
rect 1620 416 1622 424
rect 1610 414 1622 416
rect 1184 206 1188 214
rect 1196 206 1200 214
rect 1208 206 1212 214
rect 1220 206 1224 214
rect 1232 206 1236 214
rect 1244 206 1248 214
rect 1184 -10 1248 206
use BUFX2  _125_
timestamp 1591630448
transform -1 0 56 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _133_
timestamp 1591630448
transform -1 0 248 0 -1 210
box -4 -6 196 206
use NAND2X1  _75_
timestamp 1591630448
transform -1 0 56 0 1 210
box -4 -6 52 206
use INVX1  _87_
timestamp 1591630448
transform 1 0 56 0 1 210
box -4 -6 36 206
use OAI21X1  _88_
timestamp 1591630448
transform -1 0 152 0 1 210
box -4 -6 68 206
use DFFPOSX1  _150_
timestamp 1591630448
transform 1 0 152 0 1 210
box -4 -6 196 206
use OAI21X1  _91_
timestamp 1591630448
transform 1 0 248 0 -1 210
box -4 -6 68 206
use INVX1  _89_
timestamp 1591630448
transform -1 0 344 0 -1 210
box -4 -6 36 206
use NAND2X1  _90_
timestamp 1591630448
transform -1 0 392 0 -1 210
box -4 -6 52 206
use BUFX2  _129_
timestamp 1591630448
transform 1 0 392 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _153_
timestamp 1591630448
transform -1 0 600 0 1 210
box -4 -6 196 206
use FILL  SFILL3440x2100
timestamp 1591630448
transform 1 0 344 0 1 210
box -4 -6 20 206
use FILL  SFILL3600x2100
timestamp 1591630448
transform 1 0 360 0 1 210
box -4 -6 20 206
use FILL  SFILL3760x2100
timestamp 1591630448
transform 1 0 376 0 1 210
box -4 -6 20 206
use FILL  SFILL3920x2100
timestamp 1591630448
transform 1 0 392 0 1 210
box -4 -6 20 206
use BUFX2  _123_
timestamp 1591630448
transform 1 0 504 0 -1 210
box -4 -6 52 206
use NAND2X1  _69_
timestamp 1591630448
transform 1 0 552 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _146_
timestamp 1591630448
transform 1 0 600 0 -1 210
box -4 -6 196 206
use INVX1  _83_
timestamp 1591630448
transform 1 0 600 0 1 210
box -4 -6 36 206
use FILL  SFILL4400x100
timestamp 1591630448
transform -1 0 456 0 -1 210
box -4 -6 20 206
use FILL  SFILL4560x100
timestamp 1591630448
transform -1 0 472 0 -1 210
box -4 -6 20 206
use FILL  SFILL4720x100
timestamp 1591630448
transform -1 0 488 0 -1 210
box -4 -6 20 206
use FILL  SFILL4880x100
timestamp 1591630448
transform -1 0 504 0 -1 210
box -4 -6 20 206
use INVX1  _98_
timestamp 1591630448
transform 1 0 792 0 -1 210
box -4 -6 36 206
use OAI21X1  _84_
timestamp 1591630448
transform -1 0 696 0 1 210
box -4 -6 68 206
use OAI21X1  _70_
timestamp 1591630448
transform -1 0 760 0 1 210
box -4 -6 68 206
use INVX1  _68_
timestamp 1591630448
transform 1 0 760 0 1 210
box -4 -6 36 206
use DFFPOSX1  _142_
timestamp 1591630448
transform 1 0 792 0 1 210
box -4 -6 196 206
use OAI21X1  _100_
timestamp 1591630448
transform 1 0 824 0 -1 210
box -4 -6 68 206
use NAND2X1  _99_
timestamp 1591630448
transform -1 0 936 0 -1 210
box -4 -6 52 206
use BUFX2  _119_
timestamp 1591630448
transform 1 0 936 0 -1 210
box -4 -6 52 206
use BUFX2  _116_
timestamp 1591630448
transform 1 0 984 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _138_
timestamp 1591630448
transform 1 0 984 0 1 210
box -4 -6 196 206
use NAND2X1  _57_
timestamp 1591630448
transform 1 0 1032 0 -1 210
box -4 -6 52 206
use OAI21X1  _58_
timestamp 1591630448
transform -1 0 1144 0 -1 210
box -4 -6 68 206
use INVX1  _56_
timestamp 1591630448
transform -1 0 1176 0 -1 210
box -4 -6 36 206
use FILL  SFILL11760x100
timestamp 1591630448
transform -1 0 1192 0 -1 210
box -4 -6 20 206
use FILL  SFILL11920x100
timestamp 1591630448
transform -1 0 1208 0 -1 210
box -4 -6 20 206
use FILL  SFILL12080x100
timestamp 1591630448
transform -1 0 1224 0 -1 210
box -4 -6 20 206
use FILL  SFILL11760x2100
timestamp 1591630448
transform 1 0 1176 0 1 210
box -4 -6 20 206
use FILL  SFILL11920x2100
timestamp 1591630448
transform 1 0 1192 0 1 210
box -4 -6 20 206
use FILL  SFILL12080x2100
timestamp 1591630448
transform 1 0 1208 0 1 210
box -4 -6 20 206
use BUFX2  _112_
timestamp 1591630448
transform 1 0 1240 0 -1 210
box -4 -6 52 206
use BUFX2  _126_
timestamp 1591630448
transform 1 0 1288 0 -1 210
box -4 -6 52 206
use BUFX2  _110_
timestamp 1591630448
transform -1 0 1384 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _145_
timestamp 1591630448
transform 1 0 1384 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _134_
timestamp 1591630448
transform -1 0 1432 0 1 210
box -4 -6 196 206
use FILL  SFILL12240x100
timestamp 1591630448
transform -1 0 1240 0 -1 210
box -4 -6 20 206
use FILL  SFILL12240x2100
timestamp 1591630448
transform 1 0 1224 0 1 210
box -4 -6 20 206
use OAI21X1  _52_
timestamp 1591630448
transform 1 0 1576 0 -1 210
box -4 -6 68 206
use INVX1  _77_
timestamp 1591630448
transform 1 0 1432 0 1 210
box -4 -6 36 206
use OAI21X1  _78_
timestamp 1591630448
transform 1 0 1464 0 1 210
box -4 -6 68 206
use NAND2X1  _51_
timestamp 1591630448
transform -1 0 1576 0 1 210
box -4 -6 52 206
use INVX1  _107_
timestamp 1591630448
transform -1 0 1608 0 1 210
box -4 -6 36 206
use NAND2X1  _108_
timestamp 1591630448
transform 1 0 1608 0 1 210
box -4 -6 52 206
use FILL  FILL15120x100
timestamp 1591630448
transform -1 0 1656 0 -1 210
box -4 -6 20 206
use BUFX2  _118_
timestamp 1591630448
transform -1 0 56 0 -1 610
box -4 -6 52 206
use INVX1  _74_
timestamp 1591630448
transform 1 0 56 0 -1 610
box -4 -6 36 206
use OAI21X1  _76_
timestamp 1591630448
transform -1 0 152 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _144_
timestamp 1591630448
transform -1 0 344 0 -1 610
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert2
timestamp 1591630448
transform -1 0 488 0 -1 610
box -4 -6 148 206
use BUFX2  BUFX2_insert6
timestamp 1591630448
transform -1 0 600 0 -1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert0
timestamp 1591630448
transform 1 0 600 0 -1 610
box -4 -6 148 206
use FILL  SFILL4880x4100
timestamp 1591630448
transform -1 0 504 0 -1 610
box -4 -6 20 206
use FILL  SFILL5040x4100
timestamp 1591630448
transform -1 0 520 0 -1 610
box -4 -6 20 206
use FILL  SFILL5200x4100
timestamp 1591630448
transform -1 0 536 0 -1 610
box -4 -6 20 206
use FILL  SFILL5360x4100
timestamp 1591630448
transform -1 0 552 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert9
timestamp 1591630448
transform 1 0 744 0 -1 610
box -4 -6 52 206
use BUFX2  _124_
timestamp 1591630448
transform -1 0 840 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _139_
timestamp 1591630448
transform 1 0 840 0 -1 610
box -4 -6 196 206
use INVX1  _59_
timestamp 1591630448
transform 1 0 1032 0 -1 610
box -4 -6 36 206
use OAI21X1  _61_
timestamp 1591630448
transform 1 0 1064 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert4
timestamp 1591630448
transform 1 0 1128 0 -1 610
box -4 -6 52 206
use FILL  SFILL11760x4100
timestamp 1591630448
transform -1 0 1192 0 -1 610
box -4 -6 20 206
use FILL  SFILL11920x4100
timestamp 1591630448
transform -1 0 1208 0 -1 610
box -4 -6 20 206
use FILL  SFILL12080x4100
timestamp 1591630448
transform -1 0 1224 0 -1 610
box -4 -6 20 206
use OAI21X1  _94_
timestamp 1591630448
transform -1 0 1304 0 -1 610
box -4 -6 68 206
use INVX1  _92_
timestamp 1591630448
transform -1 0 1336 0 -1 610
box -4 -6 36 206
use NAND2X1  _93_
timestamp 1591630448
transform 1 0 1336 0 -1 610
box -4 -6 52 206
use BUFX2  _130_
timestamp 1591630448
transform 1 0 1384 0 -1 610
box -4 -6 52 206
use FILL  SFILL12240x4100
timestamp 1591630448
transform -1 0 1240 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert7
timestamp 1591630448
transform 1 0 1432 0 -1 610
box -4 -6 52 206
use NAND2X1  _60_
timestamp 1591630448
transform 1 0 1480 0 -1 610
box -4 -6 52 206
use NAND2X1  _102_
timestamp 1591630448
transform 1 0 1528 0 -1 610
box -4 -6 52 206
use INVX1  _50_
timestamp 1591630448
transform -1 0 1608 0 -1 610
box -4 -6 36 206
use BUFX2  _120_
timestamp 1591630448
transform -1 0 1656 0 -1 610
box -4 -6 52 206
use BUFX2  _115_
timestamp 1591630448
transform -1 0 56 0 1 610
box -4 -6 52 206
use DFFPOSX1  _141_
timestamp 1591630448
transform -1 0 248 0 1 610
box -4 -6 196 206
use INVX1  _65_
timestamp 1591630448
transform 1 0 248 0 1 610
box -4 -6 36 206
use OAI21X1  _67_
timestamp 1591630448
transform -1 0 344 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert8
timestamp 1591630448
transform -1 0 392 0 1 610
box -4 -6 52 206
use FILL  SFILL3920x6100
timestamp 1591630448
transform 1 0 392 0 1 610
box -4 -6 20 206
use FILL  SFILL4080x6100
timestamp 1591630448
transform 1 0 408 0 1 610
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert3
timestamp 1591630448
transform 1 0 456 0 1 610
box -4 -6 148 206
use CLKBUF1  CLKBUF1_insert1
timestamp 1591630448
transform 1 0 600 0 1 610
box -4 -6 148 206
use FILL  SFILL4240x6100
timestamp 1591630448
transform 1 0 424 0 1 610
box -4 -6 20 206
use FILL  SFILL4400x6100
timestamp 1591630448
transform 1 0 440 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert5
timestamp 1591630448
transform 1 0 744 0 1 610
box -4 -6 52 206
use DFFPOSX1  _132_
timestamp 1591630448
transform -1 0 984 0 1 610
box -4 -6 196 206
use INVX1  _85_
timestamp 1591630448
transform 1 0 984 0 1 610
box -4 -6 36 206
use OAI21X1  _86_
timestamp 1591630448
transform 1 0 1016 0 1 610
box -4 -6 68 206
use DFFPOSX1  _151_
timestamp 1591630448
transform 1 0 1080 0 1 610
box -4 -6 196 206
use DFFPOSX1  _147_
timestamp 1591630448
transform 1 0 1336 0 1 610
box -4 -6 196 206
use FILL  SFILL12720x6100
timestamp 1591630448
transform 1 0 1272 0 1 610
box -4 -6 20 206
use FILL  SFILL12880x6100
timestamp 1591630448
transform 1 0 1288 0 1 610
box -4 -6 20 206
use FILL  SFILL13040x6100
timestamp 1591630448
transform 1 0 1304 0 1 610
box -4 -6 20 206
use FILL  SFILL13200x6100
timestamp 1591630448
transform 1 0 1320 0 1 610
box -4 -6 20 206
use INVX1  _101_
timestamp 1591630448
transform 1 0 1528 0 1 610
box -4 -6 36 206
use OAI21X1  _103_
timestamp 1591630448
transform 1 0 1560 0 1 610
box -4 -6 68 206
use FILL  FILL14960x6100
timestamp 1591630448
transform 1 0 1624 0 1 610
box -4 -6 20 206
use FILL  FILL15120x6100
timestamp 1591630448
transform 1 0 1640 0 1 610
box -4 -6 20 206
use DFFPOSX1  _140_
timestamp 1591630448
transform -1 0 200 0 -1 1010
box -4 -6 196 206
use INVX1  _62_
timestamp 1591630448
transform 1 0 200 0 -1 1010
box -4 -6 36 206
use OAI21X1  _64_
timestamp 1591630448
transform 1 0 232 0 -1 1010
box -4 -6 68 206
use OAI21X1  _80_
timestamp 1591630448
transform -1 0 360 0 -1 1010
box -4 -6 68 206
use INVX1  _79_
timestamp 1591630448
transform -1 0 392 0 -1 1010
box -4 -6 36 206
use FILL  SFILL3920x8100
timestamp 1591630448
transform -1 0 408 0 -1 1010
box -4 -6 20 206
use FILL  SFILL4080x8100
timestamp 1591630448
transform -1 0 424 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  _135_
timestamp 1591630448
transform 1 0 456 0 -1 1010
box -4 -6 196 206
use FILL  SFILL4240x8100
timestamp 1591630448
transform -1 0 440 0 -1 1010
box -4 -6 20 206
use FILL  SFILL4400x8100
timestamp 1591630448
transform -1 0 456 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  _152_
timestamp 1591630448
transform -1 0 840 0 -1 1010
box -4 -6 196 206
use INVX1  _95_
timestamp 1591630448
transform 1 0 840 0 -1 1010
box -4 -6 36 206
use OAI21X1  _97_
timestamp 1591630448
transform -1 0 936 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _137_
timestamp 1591630448
transform 1 0 936 0 -1 1010
box -4 -6 196 206
use OAI21X1  _55_
timestamp 1591630448
transform -1 0 1192 0 -1 1010
box -4 -6 68 206
use FILL  SFILL11920x8100
timestamp 1591630448
transform -1 0 1208 0 -1 1010
box -4 -6 20 206
use FILL  SFILL12080x8100
timestamp 1591630448
transform -1 0 1224 0 -1 1010
box -4 -6 20 206
use INVX1  _53_
timestamp 1591630448
transform 1 0 1256 0 -1 1010
box -4 -6 36 206
use OAI21X1  _73_
timestamp 1591630448
transform -1 0 1352 0 -1 1010
box -4 -6 68 206
use INVX1  _71_
timestamp 1591630448
transform -1 0 1384 0 -1 1010
box -4 -6 36 206
use DFFPOSX1  _143_
timestamp 1591630448
transform 1 0 1384 0 -1 1010
box -4 -6 196 206
use FILL  SFILL12240x8100
timestamp 1591630448
transform -1 0 1240 0 -1 1010
box -4 -6 20 206
use FILL  SFILL12400x8100
timestamp 1591630448
transform -1 0 1256 0 -1 1010
box -4 -6 20 206
use OAI21X1  _109_
timestamp 1591630448
transform 1 0 1576 0 -1 1010
box -4 -6 68 206
use FILL  FILL15120x8100
timestamp 1591630448
transform -1 0 1656 0 -1 1010
box -4 -6 20 206
use BUFX2  _114_
timestamp 1591630448
transform -1 0 56 0 1 1010
box -4 -6 52 206
use NAND2X1  _66_
timestamp 1591630448
transform -1 0 104 0 1 1010
box -4 -6 52 206
use NAND2X1  _63_
timestamp 1591630448
transform 1 0 104 0 1 1010
box -4 -6 52 206
use BUFX2  _128_
timestamp 1591630448
transform -1 0 200 0 1 1010
box -4 -6 52 206
use INVX1  _81_
timestamp 1591630448
transform 1 0 200 0 1 1010
box -4 -6 36 206
use OAI21X1  _82_
timestamp 1591630448
transform 1 0 232 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _136_
timestamp 1591630448
transform -1 0 488 0 1 1010
box -4 -6 196 206
use BUFX2  _127_
timestamp 1591630448
transform 1 0 552 0 1 1010
box -4 -6 52 206
use BUFX2  _131_
timestamp 1591630448
transform 1 0 600 0 1 1010
box -4 -6 52 206
use FILL  SFILL4880x10100
timestamp 1591630448
transform 1 0 488 0 1 1010
box -4 -6 20 206
use FILL  SFILL5040x10100
timestamp 1591630448
transform 1 0 504 0 1 1010
box -4 -6 20 206
use FILL  SFILL5200x10100
timestamp 1591630448
transform 1 0 520 0 1 1010
box -4 -6 20 206
use FILL  SFILL5360x10100
timestamp 1591630448
transform 1 0 536 0 1 1010
box -4 -6 20 206
use DFFPOSX1  _148_
timestamp 1591630448
transform 1 0 648 0 1 1010
box -4 -6 196 206
use NAND2X1  _96_
timestamp 1591630448
transform -1 0 888 0 1 1010
box -4 -6 52 206
use BUFX2  _121_
timestamp 1591630448
transform 1 0 888 0 1 1010
box -4 -6 52 206
use INVX1  _104_
timestamp 1591630448
transform 1 0 936 0 1 1010
box -4 -6 36 206
use OAI21X1  _106_
timestamp 1591630448
transform 1 0 968 0 1 1010
box -4 -6 68 206
use NAND2X1  _105_
timestamp 1591630448
transform -1 0 1080 0 1 1010
box -4 -6 52 206
use NAND2X1  _54_
timestamp 1591630448
transform -1 0 1128 0 1 1010
box -4 -6 52 206
use BUFX2  _111_
timestamp 1591630448
transform 1 0 1128 0 1 1010
box -4 -6 52 206
use FILL  SFILL11760x10100
timestamp 1591630448
transform 1 0 1176 0 1 1010
box -4 -6 20 206
use FILL  SFILL11920x10100
timestamp 1591630448
transform 1 0 1192 0 1 1010
box -4 -6 20 206
use FILL  SFILL12080x10100
timestamp 1591630448
transform 1 0 1208 0 1 1010
box -4 -6 20 206
use NAND2X1  _72_
timestamp 1591630448
transform 1 0 1240 0 1 1010
box -4 -6 52 206
use BUFX2  _113_
timestamp 1591630448
transform 1 0 1288 0 1 1010
box -4 -6 52 206
use BUFX2  _117_
timestamp 1591630448
transform 1 0 1336 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _149_
timestamp 1591630448
transform 1 0 1384 0 1 1010
box -4 -6 196 206
use FILL  SFILL12240x10100
timestamp 1591630448
transform 1 0 1224 0 1 1010
box -4 -6 20 206
use BUFX2  _122_
timestamp 1591630448
transform 1 0 1576 0 1 1010
box -4 -6 52 206
use FILL  FILL14960x10100
timestamp 1591630448
transform 1 0 1624 0 1 1010
box -4 -6 20 206
use FILL  FILL15120x10100
timestamp 1591630448
transform 1 0 1640 0 1 1010
box -4 -6 20 206
<< labels >>
flabel metal4 s 1184 -10 1248 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 416 -10 480 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal3 s -35 677 -29 683 7 FreeSans 24 0 0 0 clock
port 2 nsew
flabel metal3 s 1693 697 1699 703 3 FreeSans 24 0 0 0 enable
port 3 nsew
flabel metal2 s 1357 -23 1363 -17 7 FreeSans 24 270 0 0 flag
port 4 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 imm[7]
port 5 nsew
flabel metal2 s 1357 1257 1363 1263 3 FreeSans 24 90 0 0 imm[6]
port 6 nsew
flabel metal2 s 1005 -23 1011 -17 7 FreeSans 24 270 0 0 imm[5]
port 7 nsew
flabel metal3 s -35 717 -29 723 7 FreeSans 24 0 0 0 imm[4]
port 8 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 imm[3]
port 9 nsew
flabel metal2 s 1309 1257 1315 1263 3 FreeSans 24 90 0 0 imm[2]
port 10 nsew
flabel metal2 s 1277 -23 1283 -17 7 FreeSans 24 270 0 0 imm[1]
port 11 nsew
flabel metal2 s 1149 1257 1155 1263 3 FreeSans 24 90 0 0 imm[0]
port 12 nsew
flabel metal3 s 1693 317 1699 323 3 FreeSans 24 0 0 0 instruct[15]
port 13 nsew
flabel metal2 s 1053 1257 1059 1263 3 FreeSans 24 90 0 0 instruct[14]
port 14 nsew
flabel metal3 s 1693 497 1699 503 3 FreeSans 24 0 0 0 instruct[13]
port 15 nsew
flabel metal2 s 909 -23 915 -17 7 FreeSans 24 270 0 0 instruct[12]
port 16 nsew
flabel metal2 s 861 1257 867 1263 3 FreeSans 24 90 0 0 instruct[11]
port 17 nsew
flabel metal3 s 1693 577 1699 583 3 FreeSans 24 0 0 0 instruct[10]
port 18 nsew
flabel metal2 s 365 -23 371 -17 7 FreeSans 24 270 0 0 instruct[9]
port 19 nsew
flabel metal3 s 1693 277 1699 283 3 FreeSans 24 0 0 0 instruct[8]
port 20 nsew
flabel metal3 s -35 297 -29 303 7 FreeSans 24 0 0 0 instruct[7]
port 21 nsew
flabel metal2 s 1277 1257 1283 1263 3 FreeSans 24 90 0 0 instruct[6]
port 22 nsew
flabel metal2 s 573 -23 579 -17 7 FreeSans 24 270 0 0 instruct[5]
port 23 nsew
flabel metal3 s -35 1137 -29 1143 7 FreeSans 24 0 0 0 instruct[4]
port 24 nsew
flabel metal2 s 125 1257 131 1263 3 FreeSans 24 90 0 0 instruct[3]
port 25 nsew
flabel metal3 s 1693 537 1699 543 3 FreeSans 24 0 0 0 instruct[2]
port 26 nsew
flabel metal2 s 1053 -23 1059 -17 7 FreeSans 24 270 0 0 instruct[1]
port 27 nsew
flabel metal2 s 1101 1257 1107 1263 3 FreeSans 24 90 0 0 instruct[0]
port 28 nsew
flabel metal2 s 1597 1257 1603 1263 3 FreeSans 24 90 0 0 opcode[3]
port 29 nsew
flabel metal2 s 909 1257 915 1263 3 FreeSans 24 90 0 0 opcode[2]
port 30 nsew
flabel metal3 s 1693 617 1699 623 3 FreeSans 24 0 0 0 opcode[1]
port 31 nsew
flabel metal2 s 957 -23 963 -17 7 FreeSans 24 270 0 0 opcode[0]
port 32 nsew
flabel metal3 s -35 97 -29 103 7 FreeSans 24 0 0 0 rAadrs[2]
port 33 nsew
flabel metal2 s 813 -23 819 -17 7 FreeSans 24 270 0 0 rAadrs[1]
port 34 nsew
flabel metal2 s 541 -23 547 -17 7 FreeSans 24 270 0 0 rAadrs[0]
port 35 nsew
flabel metal2 s 173 1257 179 1263 3 FreeSans 24 90 0 0 rBadrs[2]
port 36 nsew
flabel metal2 s 573 1257 579 1263 3 FreeSans 24 90 0 0 rBadrs[1]
port 37 nsew
flabel metal2 s 1309 -23 1315 -17 7 FreeSans 24 270 0 0 rBadrs[0]
port 38 nsew
flabel metal2 s 621 1257 627 1263 3 FreeSans 24 90 0 0 rDadrs[2]
port 39 nsew
flabel metal3 s 1693 657 1699 663 3 FreeSans 24 0 0 0 rDadrs[1]
port 40 nsew
flabel metal2 s 509 -23 515 -17 7 FreeSans 24 270 0 0 rDadrs[0]
port 41 nsew
<< end >>
