magic
tech scmos
magscale 1 2
timestamp 1591632351
<< metal1 >>
rect 2570 3414 2582 3416
rect 2555 3406 2557 3414
rect 2565 3406 2567 3414
rect 2575 3406 2577 3414
rect 2585 3406 2587 3414
rect 2595 3406 2597 3414
rect 2570 3404 2582 3406
rect 2628 3357 2691 3363
rect 1172 3337 1203 3343
rect 1236 3337 1251 3343
rect 1540 3337 1555 3343
rect 1917 3337 1939 3343
rect 2701 3337 2723 3343
rect 3901 3337 3923 3343
rect 4317 3337 4339 3343
rect 4765 3337 4787 3343
rect 333 3317 348 3323
rect 509 3317 524 3323
rect 1213 3317 1251 3323
rect 324 3296 332 3304
rect 1245 3297 1251 3317
rect 1517 3317 1555 3323
rect 1340 3304 1348 3314
rect 1549 3297 1555 3317
rect 2189 3317 2227 3323
rect 1828 3296 1836 3304
rect 2221 3297 2227 3317
rect 2788 3317 2803 3323
rect 3060 3317 3075 3323
rect 3373 3317 3411 3323
rect 3405 3297 3411 3317
rect 4916 3317 4931 3323
rect 4172 3312 4180 3316
rect 4236 3312 4244 3316
rect 4652 3312 4660 3316
rect 3940 3296 3948 3304
rect 4285 3297 4300 3303
rect 4637 3297 4659 3303
rect 524 3277 547 3283
rect 3434 3276 3436 3284
rect 4180 3277 4211 3283
rect 4221 3277 4252 3283
rect 4605 3277 4684 3283
rect 4804 3277 4819 3283
rect 3012 3236 3014 3244
rect 1066 3214 1078 3216
rect 4074 3214 4086 3216
rect 1051 3206 1053 3214
rect 1061 3206 1063 3214
rect 1071 3206 1073 3214
rect 1081 3206 1083 3214
rect 1091 3206 1093 3214
rect 4059 3206 4061 3214
rect 4069 3206 4071 3214
rect 4079 3206 4081 3214
rect 4089 3206 4091 3214
rect 4099 3206 4101 3214
rect 1066 3204 1078 3206
rect 4074 3204 4086 3206
rect 596 3176 598 3184
rect 650 3176 652 3184
rect 756 3176 758 3184
rect 1236 3176 1238 3184
rect 2682 3176 2684 3184
rect 538 3156 540 3164
rect 820 3136 822 3144
rect 2244 3136 2246 3144
rect 3796 3136 3802 3144
rect 4356 3137 4371 3143
rect 468 3116 476 3124
rect 653 3097 668 3103
rect 717 3097 732 3103
rect 1149 3103 1155 3123
rect 1117 3097 1155 3103
rect 1332 3097 1363 3103
rect 1444 3097 1459 3103
rect 1965 3103 1971 3123
rect 1988 3116 1996 3124
rect 2932 3116 2940 3124
rect 1933 3097 1971 3103
rect 2276 3097 2291 3103
rect 2388 3097 2403 3103
rect 2509 3097 2547 3103
rect 669 3077 691 3083
rect 1044 3077 1107 3083
rect 1277 3077 1299 3083
rect 2445 3077 2460 3083
rect 2541 3083 2547 3097
rect 2724 3097 2739 3103
rect 2877 3097 2892 3103
rect 3277 3103 3283 3123
rect 3245 3097 3283 3103
rect 3389 3103 3395 3123
rect 3357 3097 3395 3103
rect 3517 3097 3532 3103
rect 3693 3103 3699 3123
rect 4292 3116 4300 3124
rect 3661 3097 3699 3103
rect 4301 3097 4316 3103
rect 4468 3097 4483 3103
rect 4788 3097 4803 3103
rect 4813 3097 4828 3103
rect 2541 3077 2627 3083
rect 2996 3077 3011 3083
rect 3684 3077 3699 3083
rect 4317 3077 4339 3083
rect 4829 3077 4851 3083
rect 1021 3037 1036 3043
rect 1396 3036 1398 3044
rect 2570 3014 2582 3016
rect 2555 3006 2557 3014
rect 2565 3006 2567 3014
rect 2575 3006 2577 3014
rect 2585 3006 2587 3014
rect 2595 3006 2597 3014
rect 2570 3004 2582 3006
rect 1044 2956 1046 2964
rect 1293 2957 1308 2963
rect 596 2937 611 2943
rect 909 2937 931 2943
rect 1268 2937 1283 2943
rect 2532 2937 2611 2943
rect 2653 2937 2668 2943
rect 2925 2937 2940 2943
rect 3092 2937 3107 2943
rect 3165 2937 3187 2943
rect 3914 2936 3916 2944
rect 4301 2937 4316 2943
rect 4637 2937 4659 2943
rect 669 2917 700 2923
rect 765 2917 803 2923
rect 428 2904 436 2914
rect 797 2897 803 2917
rect 868 2917 883 2923
rect 1069 2917 1180 2923
rect 1652 2917 1667 2923
rect 1693 2917 1731 2923
rect 1693 2897 1699 2917
rect 2061 2917 2099 2923
rect 2061 2897 2067 2917
rect 2157 2917 2195 2923
rect 2189 2897 2195 2917
rect 2340 2917 2371 2923
rect 2724 2917 2739 2923
rect 2909 2917 2963 2923
rect 3284 2917 3292 2923
rect 3300 2917 3315 2923
rect 3709 2917 3747 2923
rect 3741 2897 3747 2917
rect 3773 2917 3788 2923
rect 4068 2917 4179 2923
rect 4301 2917 4339 2923
rect 4301 2897 4307 2917
rect 4452 2917 4483 2923
rect 4781 2917 4796 2923
rect 4556 2912 4564 2916
rect 4909 2897 4924 2903
rect 2884 2876 2886 2884
rect 4605 2877 4620 2883
rect 4756 2876 4762 2884
rect 4980 2877 5011 2883
rect 3274 2856 3276 2864
rect 1476 2836 1478 2844
rect 2484 2836 2486 2844
rect 2740 2836 2742 2844
rect 3444 2836 3446 2844
rect 1066 2814 1078 2816
rect 4074 2814 4086 2816
rect 1051 2806 1053 2814
rect 1061 2806 1063 2814
rect 1071 2806 1073 2814
rect 1081 2806 1083 2814
rect 1091 2806 1093 2814
rect 4059 2806 4061 2814
rect 4069 2806 4071 2814
rect 4079 2806 4081 2814
rect 4089 2806 4091 2814
rect 4099 2806 4101 2814
rect 1066 2804 1078 2806
rect 4074 2804 4086 2806
rect 1300 2776 1302 2784
rect 2068 2776 2070 2784
rect 2276 2776 2278 2784
rect 2468 2776 2470 2784
rect 2557 2777 2572 2783
rect 2964 2776 2966 2784
rect 3098 2776 3100 2784
rect 3962 2776 3964 2784
rect 5085 2777 5100 2783
rect 474 2756 476 2764
rect 172 2737 195 2743
rect 794 2736 796 2744
rect 1962 2736 1964 2744
rect 2906 2736 2908 2744
rect 3204 2736 3206 2744
rect 1812 2716 1820 2724
rect 93 2697 140 2703
rect 157 2697 172 2703
rect 253 2697 268 2703
rect 484 2697 531 2703
rect 797 2697 828 2703
rect 884 2697 915 2703
rect 1132 2703 1140 2706
rect 1132 2697 1235 2703
rect 1325 2697 1340 2703
rect 1757 2697 1811 2703
rect 1869 2703 1875 2723
rect 1852 2697 1875 2703
rect 1852 2692 1860 2697
rect 2148 2697 2179 2703
rect 2420 2697 2435 2703
rect 2877 2703 2883 2723
rect 3044 2716 3052 2724
rect 2845 2697 2883 2703
rect 3005 2697 3020 2703
rect 116 2677 131 2683
rect 500 2677 515 2683
rect 1981 2677 1996 2683
rect 2013 2677 2044 2683
rect 3005 2677 3011 2697
rect 3149 2697 3203 2703
rect 3261 2703 3267 2723
rect 3244 2697 3267 2703
rect 3244 2692 3252 2697
rect 3549 2697 3564 2703
rect 3693 2703 3699 2723
rect 3661 2697 3699 2703
rect 3933 2703 3939 2723
rect 3901 2697 3939 2703
rect 3981 2697 3996 2703
rect 3844 2677 3875 2683
rect 3981 2677 3987 2697
rect 4109 2703 4115 2723
rect 4013 2697 4115 2703
rect 4228 2697 4243 2703
rect 4660 2697 4675 2703
rect 4781 2697 4796 2703
rect 5044 2697 5059 2703
rect 4925 2677 4947 2683
rect 4052 2637 4115 2643
rect 4196 2636 4198 2644
rect 2570 2614 2582 2616
rect 2555 2606 2557 2614
rect 2565 2606 2567 2614
rect 2575 2606 2577 2614
rect 2585 2606 2587 2614
rect 2595 2606 2597 2614
rect 2570 2604 2582 2606
rect 2557 2557 2636 2563
rect 621 2537 636 2543
rect 916 2537 931 2543
rect 1053 2537 1132 2543
rect 2301 2537 2323 2543
rect 93 2517 116 2523
rect 108 2514 116 2517
rect 308 2517 323 2523
rect 628 2517 659 2523
rect 749 2517 764 2523
rect 788 2517 803 2523
rect 893 2517 931 2523
rect 925 2497 931 2517
rect 1053 2517 1132 2523
rect 1661 2517 1699 2523
rect 1661 2497 1667 2517
rect 2365 2523 2371 2543
rect 2964 2537 2979 2543
rect 4717 2537 4739 2543
rect 5101 2537 5123 2543
rect 2365 2517 2396 2523
rect 2444 2523 2452 2528
rect 2429 2517 2452 2523
rect 1956 2496 1964 2504
rect 2429 2497 2435 2517
rect 2493 2517 2508 2523
rect 2564 2517 2604 2523
rect 2628 2517 2643 2523
rect 2941 2517 2979 2523
rect 2973 2497 2979 2517
rect 3341 2517 3379 2523
rect 3373 2497 3379 2517
rect 5085 2517 5100 2523
rect 4180 2497 4195 2503
rect 4756 2496 4764 2504
rect 1172 2476 1174 2484
rect 2260 2476 2262 2484
rect 2404 2476 2406 2484
rect 1066 2414 1078 2416
rect 4074 2414 4086 2416
rect 1051 2406 1053 2414
rect 1061 2406 1063 2414
rect 1071 2406 1073 2414
rect 1081 2406 1083 2414
rect 1091 2406 1093 2414
rect 4059 2406 4061 2414
rect 4069 2406 4071 2414
rect 4079 2406 4081 2414
rect 4089 2406 4091 2414
rect 4099 2406 4101 2414
rect 1066 2404 1078 2406
rect 4074 2404 4086 2406
rect 132 2376 134 2384
rect 1428 2376 1430 2384
rect 1540 2376 1542 2384
rect 1930 2356 1932 2364
rect 196 2336 198 2344
rect 220 2337 243 2343
rect 3060 2336 3062 2344
rect 4349 2337 4364 2343
rect 4420 2337 4467 2343
rect 4596 2337 4611 2343
rect 93 2297 108 2303
rect 301 2297 316 2303
rect 484 2297 515 2303
rect 525 2297 579 2303
rect 589 2297 604 2303
rect 845 2297 899 2303
rect 1380 2297 1411 2303
rect 1325 2277 1347 2283
rect 1405 2277 1411 2297
rect 1709 2297 1763 2303
rect 1901 2303 1907 2323
rect 1869 2297 1907 2303
rect 1933 2297 1948 2303
rect 2317 2297 2332 2303
rect 2845 2303 2851 2323
rect 2845 2297 2868 2303
rect 1501 2277 1516 2283
rect 1501 2264 1507 2277
rect 1725 2277 1740 2283
rect 1844 2277 1859 2283
rect 2125 2277 2147 2283
rect 2189 2277 2195 2296
rect 2860 2292 2868 2297
rect 2909 2297 2963 2303
rect 3501 2303 3507 2323
rect 3876 2316 3884 2324
rect 3501 2297 3539 2303
rect 3693 2297 3708 2303
rect 4013 2303 4019 2323
rect 3981 2297 4019 2303
rect 4868 2297 4883 2303
rect 2269 2277 2291 2283
rect 2669 2277 2691 2283
rect 3837 2277 3859 2283
rect 4061 2277 4124 2283
rect 4557 2277 4579 2283
rect 4909 2277 4931 2283
rect 1476 2257 1491 2263
rect 2365 2257 2380 2263
rect 2756 2257 2771 2263
rect 3156 2236 3158 2244
rect 2570 2214 2582 2216
rect 2555 2206 2557 2214
rect 2565 2206 2567 2214
rect 2575 2206 2577 2214
rect 2585 2206 2587 2214
rect 2595 2206 2597 2214
rect 2570 2204 2582 2206
rect 948 2176 950 2184
rect 548 2157 563 2163
rect 573 2157 588 2163
rect 628 2157 643 2163
rect 580 2137 611 2143
rect 1012 2137 1027 2143
rect 1213 2137 1235 2143
rect 2004 2137 2019 2143
rect 4829 2137 4867 2143
rect 372 2117 387 2123
rect 420 2117 435 2123
rect 797 2117 812 2123
rect 989 2117 1027 2123
rect 1021 2097 1027 2117
rect 1981 2117 2019 2123
rect 2013 2097 2019 2117
rect 2141 2117 2179 2123
rect 2173 2097 2179 2117
rect 2509 2117 2588 2123
rect 2797 2117 2835 2123
rect 2861 2117 2876 2123
rect 2532 2097 2572 2103
rect 2829 2097 2835 2117
rect 3149 2117 3164 2123
rect 3517 2117 3555 2123
rect 2852 2096 2860 2104
rect 3492 2096 3500 2104
rect 3517 2097 3523 2117
rect 3853 2117 3891 2123
rect 3885 2097 3891 2117
rect 4013 2117 4115 2123
rect 4141 2117 4156 2123
rect 4109 2097 4115 2117
rect 4909 2117 4924 2123
rect 4132 2096 4140 2104
rect 4436 2097 4451 2103
rect 156 2077 179 2083
rect 461 2077 484 2083
rect 3220 2076 3222 2084
rect 4468 2077 4483 2083
rect 3124 2056 3126 2064
rect 2634 2036 2636 2044
rect 1066 2014 1078 2016
rect 4074 2014 4086 2016
rect 1051 2006 1053 2014
rect 1061 2006 1063 2014
rect 1071 2006 1073 2014
rect 1081 2006 1083 2014
rect 1091 2006 1093 2014
rect 4059 2006 4061 2014
rect 4069 2006 4071 2014
rect 4079 2006 4081 2014
rect 4089 2006 4091 2014
rect 4099 2006 4101 2014
rect 1066 2004 1078 2006
rect 4074 2004 4086 2006
rect 1924 1976 1926 1984
rect 1802 1956 1804 1964
rect 2196 1956 2198 1964
rect 204 1937 227 1943
rect 2676 1937 2691 1943
rect 4269 1937 4300 1943
rect 4396 1932 4404 1936
rect 493 1897 547 1903
rect 644 1897 675 1903
rect 765 1897 780 1903
rect 804 1897 819 1903
rect 989 1903 995 1923
rect 1428 1916 1436 1924
rect 989 1897 1027 1903
rect 1060 1897 1155 1903
rect 1396 1897 1411 1903
rect 141 1877 163 1883
rect 1293 1877 1308 1883
rect 1405 1877 1411 1897
rect 2461 1903 2467 1923
rect 2452 1897 2467 1903
rect 3133 1903 3139 1923
rect 3156 1916 3164 1924
rect 3101 1897 3139 1903
rect 3581 1903 3587 1923
rect 4284 1904 4292 1908
rect 5084 1904 5092 1908
rect 3549 1897 3587 1903
rect 3613 1897 3628 1903
rect 4388 1897 4419 1903
rect 4813 1897 4828 1903
rect 4932 1897 4963 1903
rect 1533 1877 1555 1883
rect 1885 1877 1907 1883
rect 2077 1877 2099 1883
rect 2157 1877 2172 1883
rect 2381 1877 2403 1883
rect 4116 1877 4131 1883
rect 4765 1877 4787 1883
rect 5053 1837 5068 1843
rect 2570 1814 2582 1816
rect 2555 1806 2557 1814
rect 2565 1806 2567 1814
rect 2575 1806 2577 1814
rect 2585 1806 2587 1814
rect 2595 1806 2597 1814
rect 2570 1804 2582 1806
rect 3466 1776 3468 1784
rect 237 1744 243 1763
rect 2557 1757 2636 1763
rect 3180 1757 3203 1763
rect 3180 1754 3188 1757
rect 4477 1757 4492 1763
rect 77 1737 92 1743
rect 125 1737 140 1743
rect 244 1737 259 1743
rect 1117 1724 1123 1743
rect 2532 1737 2547 1743
rect 2564 1737 2659 1743
rect 3885 1737 3900 1743
rect 4026 1736 4028 1744
rect 4148 1737 4211 1743
rect 4461 1737 4476 1743
rect 5069 1737 5091 1743
rect 109 1717 124 1723
rect 765 1717 803 1723
rect 797 1697 803 1717
rect 925 1717 940 1723
rect 1165 1717 1203 1723
rect 1437 1717 1475 1723
rect 1165 1697 1171 1717
rect 1469 1697 1475 1717
rect 2157 1717 2195 1723
rect 2189 1697 2195 1717
rect 2356 1717 2371 1723
rect 2564 1717 2636 1723
rect 2909 1717 2947 1723
rect 2941 1697 2947 1717
rect 3501 1717 3516 1723
rect 3620 1717 3635 1723
rect 4413 1717 4451 1723
rect 4484 1717 4499 1723
rect 4396 1712 4404 1716
rect 4588 1712 4596 1716
rect 4796 1712 4804 1716
rect 4308 1697 4323 1703
rect 4397 1697 4419 1703
rect 3940 1677 3955 1683
rect 4573 1677 4620 1683
rect 2218 1636 2220 1644
rect 3220 1636 3222 1644
rect 1066 1614 1078 1616
rect 4074 1614 4086 1616
rect 1051 1606 1053 1614
rect 1061 1606 1063 1614
rect 1071 1606 1073 1614
rect 1081 1606 1083 1614
rect 1091 1606 1093 1614
rect 4059 1606 4061 1614
rect 4069 1606 4071 1614
rect 4079 1606 4081 1614
rect 4089 1606 4091 1614
rect 4099 1606 4101 1614
rect 1066 1604 1078 1606
rect 4074 1604 4086 1606
rect 180 1576 182 1584
rect 1540 1576 1542 1584
rect 1978 1576 1980 1584
rect 2548 1577 2611 1583
rect 2794 1576 2796 1584
rect 1364 1556 1366 1564
rect 1860 1556 1862 1564
rect 2948 1556 2950 1564
rect 3284 1556 3286 1564
rect 204 1537 227 1543
rect 2596 1537 2611 1543
rect 3098 1536 3100 1544
rect 3644 1537 3660 1543
rect 4132 1536 4138 1544
rect 4980 1536 4986 1544
rect 324 1497 339 1503
rect 669 1497 700 1503
rect 893 1503 899 1523
rect 861 1497 899 1503
rect 1005 1503 1011 1523
rect 1005 1497 1043 1503
rect 1389 1503 1395 1523
rect 1348 1497 1363 1503
rect 1389 1497 1427 1503
rect 1444 1497 1475 1503
rect 1764 1497 1779 1503
rect 1869 1497 1884 1503
rect 2413 1497 2428 1503
rect 2637 1497 2652 1503
rect 2685 1497 2700 1503
rect 2893 1497 2947 1503
rect 3005 1503 3011 1523
rect 2988 1497 3011 1503
rect 3037 1497 3052 1503
rect 141 1477 163 1483
rect 396 1477 420 1483
rect 948 1477 963 1483
rect 1437 1477 1443 1496
rect 2988 1492 2996 1497
rect 3229 1497 3283 1503
rect 3341 1503 3347 1523
rect 3476 1516 3484 1524
rect 3324 1497 3347 1503
rect 3324 1492 3332 1497
rect 3460 1497 3475 1503
rect 3533 1503 3539 1523
rect 3516 1497 3539 1503
rect 3516 1492 3524 1497
rect 3709 1503 3715 1523
rect 3677 1497 3715 1503
rect 3741 1497 3756 1503
rect 3997 1497 4028 1503
rect 4525 1503 4531 1523
rect 4493 1497 4531 1503
rect 4788 1497 4803 1503
rect 1501 1477 1523 1483
rect 1741 1477 1763 1483
rect 2861 1477 2876 1483
rect 4516 1477 4531 1483
rect 4829 1477 4851 1483
rect 1636 1457 1667 1463
rect 1194 1436 1196 1444
rect 2570 1414 2582 1416
rect 2555 1406 2557 1414
rect 2565 1406 2567 1414
rect 2575 1406 2577 1414
rect 2585 1406 2587 1414
rect 2595 1406 2597 1414
rect 2570 1404 2582 1406
rect 836 1357 851 1363
rect 1645 1357 1660 1363
rect 186 1336 188 1344
rect 356 1337 371 1343
rect 1188 1337 1203 1343
rect 1261 1337 1283 1343
rect 1620 1337 1635 1343
rect 1748 1337 1779 1343
rect 2596 1337 2611 1343
rect 3060 1337 3075 1343
rect 3924 1337 3939 1343
rect 4413 1337 4428 1343
rect 4477 1337 4492 1343
rect 4941 1337 4963 1343
rect 340 1317 387 1323
rect 397 1317 412 1323
rect 676 1317 707 1323
rect 724 1317 755 1323
rect 765 1317 796 1323
rect 1245 1317 1276 1323
rect 1469 1317 1500 1323
rect 1981 1317 1996 1323
rect 2093 1317 2131 1323
rect 2125 1297 2131 1317
rect 2292 1317 2307 1323
rect 2509 1317 2611 1323
rect 2605 1297 2611 1317
rect 2989 1317 3004 1323
rect 3421 1317 3436 1323
rect 3533 1317 3564 1323
rect 3693 1317 3708 1323
rect 3901 1317 3916 1323
rect 3924 1317 3955 1323
rect 3965 1317 4003 1323
rect 3997 1297 4003 1317
rect 4356 1317 4387 1323
rect 4477 1317 4515 1323
rect 4333 1297 4371 1303
rect 4477 1297 4483 1317
rect 4644 1317 4659 1323
rect 4964 1317 4979 1323
rect 330 1276 332 1284
rect 412 1277 435 1283
rect 938 1276 940 1284
rect 1220 1276 1222 1284
rect 1524 1276 1526 1284
rect 4532 1277 4547 1283
rect 2154 1256 2156 1264
rect 820 1236 822 1244
rect 2020 1236 2022 1244
rect 3204 1236 3206 1244
rect 3668 1236 3670 1244
rect 3898 1236 3900 1244
rect 1066 1214 1078 1216
rect 4074 1214 4086 1216
rect 1051 1206 1053 1214
rect 1061 1206 1063 1214
rect 1071 1206 1073 1214
rect 1081 1206 1083 1214
rect 1091 1206 1093 1214
rect 4059 1206 4061 1214
rect 4069 1206 4071 1214
rect 4079 1206 4081 1214
rect 4089 1206 4091 1214
rect 4099 1206 4101 1214
rect 1066 1204 1078 1206
rect 4074 1204 4086 1206
rect 330 1176 332 1184
rect 1348 1176 1350 1184
rect 4052 1177 4115 1183
rect 3012 1156 3014 1164
rect 276 1136 278 1144
rect 685 1097 716 1103
rect 861 1103 867 1123
rect 829 1097 867 1103
rect 1133 1097 1148 1103
rect 1629 1103 1635 1123
rect 3556 1116 3564 1124
rect 1597 1097 1635 1103
rect 2132 1097 2147 1103
rect 2157 1097 2172 1103
rect 2269 1097 2284 1103
rect 2372 1097 2403 1103
rect 2436 1097 2451 1103
rect 3076 1097 3091 1103
rect 4589 1103 4595 1123
rect 4964 1116 4972 1124
rect 4557 1097 4595 1103
rect 4948 1097 4963 1103
rect 796 1077 819 1083
rect 796 1072 804 1077
rect 1149 1077 1171 1083
rect 1620 1077 1635 1083
rect 1677 1077 1692 1083
rect 1821 1077 1836 1083
rect 1796 1057 1811 1063
rect 1821 1057 1827 1077
rect 2980 1077 2995 1083
rect 4029 1077 4076 1083
rect 4580 1077 4595 1083
rect 4925 1077 4947 1083
rect 2700 1064 2708 1072
rect 2301 1057 2316 1063
rect 2340 1057 2355 1063
rect 2372 1057 2387 1063
rect 3140 1057 3155 1063
rect 3732 1056 3734 1064
rect 3636 1036 3638 1044
rect 2570 1014 2582 1016
rect 2555 1006 2557 1014
rect 2565 1006 2567 1014
rect 2575 1006 2577 1014
rect 2585 1006 2587 1014
rect 2595 1006 2597 1014
rect 2570 1004 2582 1006
rect 2644 977 2675 983
rect 2100 956 2102 964
rect 3364 956 3366 964
rect 541 937 579 943
rect 644 937 675 943
rect 740 937 755 943
rect 1309 937 1324 943
rect 1437 937 1459 943
rect 1581 937 1603 943
rect 1917 937 1939 943
rect 2612 937 2668 943
rect 2925 937 2947 943
rect 3069 937 3091 943
rect 4474 936 4476 944
rect 4605 937 4627 943
rect 4925 937 4963 943
rect 205 917 220 923
rect 269 917 284 923
rect 877 917 892 923
rect 1053 917 1155 923
rect 1053 897 1059 917
rect 1229 917 1283 923
rect 1565 917 1580 923
rect 1693 917 1708 923
rect 2125 917 2156 923
rect 2164 917 2179 923
rect 2317 917 2355 923
rect 1124 897 1139 903
rect 1796 896 1804 904
rect 1876 896 1886 904
rect 2349 897 2355 917
rect 2884 917 2899 923
rect 3053 917 3084 923
rect 3165 917 3219 923
rect 3389 917 3436 923
rect 3533 917 3587 923
rect 3628 923 3636 928
rect 3628 917 3651 923
rect 2372 896 2380 904
rect 2964 896 2972 904
rect 3645 897 3651 917
rect 3789 917 3827 923
rect 3821 897 3827 917
rect 3972 917 4003 923
rect 4365 917 4380 923
rect 4909 917 4924 923
rect 5085 897 5148 903
rect 138 876 140 884
rect 284 877 307 883
rect 2276 856 2278 864
rect 628 836 630 844
rect 724 836 726 844
rect 1348 836 1350 844
rect 1684 836 1686 844
rect 1738 836 1740 844
rect 2026 836 2028 844
rect 3028 836 3030 844
rect 3588 836 3590 844
rect 1066 814 1078 816
rect 4074 814 4086 816
rect 1051 806 1053 814
rect 1061 806 1063 814
rect 1071 806 1073 814
rect 1081 806 1083 814
rect 1091 806 1093 814
rect 4059 806 4061 814
rect 4069 806 4071 814
rect 4079 806 4081 814
rect 4089 806 4091 814
rect 4099 806 4101 814
rect 1066 804 1078 806
rect 4074 804 4086 806
rect 746 776 748 784
rect 1748 756 1750 764
rect 2372 756 2374 764
rect 426 736 428 744
rect 3581 737 3596 743
rect 541 697 572 703
rect 772 697 787 703
rect 893 697 924 703
rect 1069 703 1075 723
rect 1140 717 1155 723
rect 1069 697 1171 703
rect 1485 703 1491 723
rect 1780 717 1795 723
rect 2756 716 2766 724
rect 1453 697 1491 703
rect 1796 697 1811 703
rect 2205 697 2236 703
rect 2292 697 2323 703
rect 2525 697 2572 703
rect 2781 697 2835 703
rect 2156 692 2164 696
rect 3156 697 3171 703
rect 3293 703 3299 723
rect 3293 697 3331 703
rect 3444 697 3475 703
rect 3869 697 3884 703
rect 4253 703 4259 723
rect 4804 716 4812 724
rect 4221 697 4259 703
rect 4788 697 4803 703
rect 1428 677 1443 683
rect 2141 677 2163 683
rect 2221 677 2243 683
rect 2285 677 2300 683
rect 2541 677 2556 683
rect 2596 677 2643 683
rect 3060 677 3075 683
rect 3341 677 3364 683
rect 3356 672 3364 677
rect 3613 677 3628 683
rect 4148 677 4211 683
rect 4477 677 4499 683
rect 4765 677 4787 683
rect 4925 677 4947 683
rect 2570 614 2582 616
rect 2555 606 2557 614
rect 2565 606 2567 614
rect 2575 606 2577 614
rect 2585 606 2587 614
rect 2595 606 2597 614
rect 2570 604 2582 606
rect 2506 576 2508 584
rect 3380 576 3382 584
rect 684 557 716 563
rect 684 548 692 557
rect 1181 537 1203 543
rect 1434 536 1436 544
rect 2317 537 2339 543
rect 2525 537 2540 543
rect 2717 537 2739 543
rect 2845 537 2860 543
rect 2973 537 2995 543
rect 3037 537 3052 543
rect 3149 537 3171 543
rect 3229 537 3244 543
rect 3428 537 3459 543
rect 3581 537 3596 543
rect 468 517 483 523
rect 493 517 508 523
rect 925 517 940 523
rect 1076 517 1155 523
rect 1236 517 1244 523
rect 1325 517 1340 523
rect 1581 517 1596 523
rect 1645 517 1699 523
rect 1732 517 1763 523
rect 1773 517 1827 523
rect 1837 517 1852 523
rect 1876 517 1891 523
rect 2052 517 2083 523
rect 2093 517 2108 523
rect 2301 517 2332 523
rect 2404 517 2419 523
rect 3044 517 3059 523
rect 3284 517 3299 523
rect 3405 517 3452 523
rect 3565 517 3612 523
rect 3956 517 3987 523
rect 4301 517 4339 523
rect 420 496 428 504
rect 3188 496 3196 504
rect 4333 497 4339 517
rect 4548 517 4563 523
rect 4749 523 4755 543
rect 4749 517 4764 523
rect 4716 512 4724 516
rect 5012 517 5043 523
rect 4764 512 4772 516
rect 4908 512 4916 516
rect 1578 476 1580 484
rect 2026 476 2028 484
rect 3620 476 3622 484
rect 3644 477 3667 483
rect 1322 436 1324 444
rect 2932 436 2934 444
rect 3562 436 3564 444
rect 3988 436 3990 444
rect 1066 414 1078 416
rect 4074 414 4086 416
rect 1051 406 1053 414
rect 1061 406 1063 414
rect 1071 406 1073 414
rect 1081 406 1083 414
rect 1091 406 1093 414
rect 4059 406 4061 414
rect 4069 406 4071 414
rect 4079 406 4081 414
rect 4089 406 4091 414
rect 4099 406 4101 414
rect 1066 404 1078 406
rect 4074 404 4086 406
rect 426 376 428 384
rect 922 376 924 384
rect 1348 376 1350 384
rect 1610 376 1612 384
rect 1668 376 1670 384
rect 3380 376 3382 384
rect 2612 356 2614 364
rect 381 337 404 343
rect 986 336 988 344
rect 1124 337 1139 343
rect 3476 336 3482 344
rect 3860 336 3866 344
rect 269 297 284 303
rect 589 303 595 323
rect 557 297 595 303
rect 925 297 940 303
rect 1053 297 1116 303
rect 1620 297 1667 303
rect 2413 297 2428 303
rect 2708 297 2739 303
rect 3021 303 3027 323
rect 3284 316 3292 324
rect 3021 297 3059 303
rect 3268 297 3283 303
rect 3405 297 3420 303
rect 2140 292 2148 296
rect 3757 303 3763 323
rect 3700 297 3715 303
rect 3725 297 3763 303
rect 4125 303 4131 323
rect 4676 316 4684 324
rect 4029 297 4131 303
rect 4276 297 4307 303
rect 4877 297 4892 303
rect 5012 297 5027 303
rect 516 277 531 283
rect 1636 277 1651 283
rect 2125 277 2147 283
rect 2205 277 2227 283
rect 2580 277 2595 283
rect 3108 277 3123 283
rect 3245 277 3267 283
rect 4637 277 4659 283
rect 4733 277 4755 283
rect 4829 277 4851 283
rect 44 264 52 272
rect 1852 264 1860 272
rect 1946 256 1948 264
rect 3468 263 3476 272
rect 3468 257 3500 263
rect 4586 236 4588 244
rect 2570 214 2582 216
rect 2555 206 2557 214
rect 2565 206 2567 214
rect 2575 206 2577 214
rect 2585 206 2587 214
rect 2595 206 2597 214
rect 2570 204 2582 206
rect 2573 177 2620 183
rect 2644 177 2659 183
rect 3460 157 3475 163
rect 556 148 564 156
rect 2269 137 2291 143
rect 2333 137 2348 143
rect 3437 137 3452 143
rect 420 117 435 123
rect 612 117 643 123
rect 749 117 764 123
rect 893 117 924 123
rect 1165 117 1219 123
rect 1229 117 1244 123
rect 1645 117 1668 123
rect 1660 114 1668 117
rect 2109 117 2147 123
rect 324 96 332 104
rect 2141 97 2147 117
rect 2340 117 2355 123
rect 2461 117 2476 123
rect 2765 117 2780 123
rect 2909 117 2947 123
rect 2941 97 2947 117
rect 3213 117 3251 123
rect 3245 97 3251 117
rect 3372 123 3380 128
rect 3357 117 3380 123
rect 3357 97 3363 117
rect 3444 117 3459 123
rect 3508 117 3523 123
rect 3588 117 3603 123
rect 3780 117 3811 123
rect 4157 117 4195 123
rect 4189 97 4195 117
rect 4493 117 4531 123
rect 4493 97 4499 117
rect 4708 117 4739 123
rect 3636 56 3638 64
rect 1053 37 1116 43
rect 3396 36 3398 44
rect 1066 14 1078 16
rect 4074 14 4086 16
rect 1051 6 1053 14
rect 1061 6 1063 14
rect 1071 6 1073 14
rect 1081 6 1083 14
rect 1091 6 1093 14
rect 4059 6 4061 14
rect 4069 6 4071 14
rect 4079 6 4081 14
rect 4089 6 4091 14
rect 4099 6 4101 14
rect 1066 4 1078 6
rect 4074 4 4086 6
<< m2contact >>
rect 2547 3406 2555 3414
rect 2557 3406 2565 3414
rect 2567 3406 2575 3414
rect 2577 3406 2585 3414
rect 2587 3406 2595 3414
rect 2597 3406 2605 3414
rect 204 3376 212 3384
rect 284 3376 292 3384
rect 428 3376 436 3384
rect 1308 3376 1316 3384
rect 2428 3376 2436 3384
rect 3468 3376 3476 3384
rect 4396 3376 4404 3384
rect 364 3356 372 3364
rect 1932 3356 1940 3364
rect 2620 3356 2628 3364
rect 3884 3356 3892 3364
rect 4300 3356 4308 3364
rect 4796 3356 4804 3364
rect 5004 3356 5012 3364
rect 124 3336 132 3344
rect 348 3336 356 3344
rect 412 3336 420 3344
rect 476 3336 484 3344
rect 732 3336 740 3344
rect 780 3336 788 3344
rect 924 3336 932 3344
rect 1164 3336 1172 3344
rect 1228 3336 1236 3344
rect 1292 3336 1300 3344
rect 1500 3336 1508 3344
rect 1532 3336 1540 3344
rect 1596 3336 1604 3344
rect 1708 3336 1716 3344
rect 1852 3336 1860 3344
rect 1868 3336 1876 3344
rect 1948 3336 1956 3344
rect 2156 3336 2164 3344
rect 2220 3336 2228 3344
rect 2268 3336 2276 3344
rect 2284 3336 2292 3344
rect 2748 3336 2756 3344
rect 2796 3336 2804 3344
rect 3324 3336 3332 3344
rect 3356 3336 3364 3344
rect 3452 3336 3460 3344
rect 3628 3336 3636 3344
rect 3676 3336 3684 3344
rect 3788 3336 3796 3344
rect 4380 3336 4388 3344
rect 4524 3336 4532 3344
rect 4924 3336 4932 3344
rect 5036 3336 5044 3344
rect 5084 3336 5092 3344
rect 140 3318 148 3326
rect 236 3316 244 3324
rect 252 3316 260 3324
rect 348 3316 356 3324
rect 396 3316 404 3324
rect 460 3316 468 3324
rect 492 3316 500 3324
rect 524 3316 532 3324
rect 604 3316 612 3324
rect 668 3318 676 3326
rect 764 3316 772 3324
rect 1004 3316 1012 3324
rect 1068 3318 1076 3326
rect 300 3296 308 3304
rect 332 3296 340 3304
rect 364 3296 372 3304
rect 524 3296 532 3304
rect 732 3296 740 3304
rect 1228 3296 1236 3304
rect 1276 3316 1284 3324
rect 1372 3316 1380 3324
rect 1436 3318 1444 3326
rect 1340 3296 1348 3304
rect 1532 3296 1540 3304
rect 1580 3316 1588 3324
rect 1740 3318 1748 3326
rect 1836 3316 1844 3324
rect 1900 3316 1908 3324
rect 2028 3316 2036 3324
rect 2076 3316 2084 3324
rect 2172 3316 2180 3324
rect 1836 3296 1844 3304
rect 1868 3296 1876 3304
rect 2252 3316 2260 3324
rect 2412 3316 2420 3324
rect 2492 3316 2500 3324
rect 2556 3318 2564 3326
rect 2732 3316 2740 3324
rect 2780 3316 2788 3324
rect 2844 3316 2852 3324
rect 2860 3316 2868 3324
rect 2892 3316 2900 3324
rect 2940 3316 2948 3324
rect 2956 3316 2964 3324
rect 2972 3316 2980 3324
rect 2988 3316 2996 3324
rect 3036 3316 3044 3324
rect 3052 3316 3060 3324
rect 3084 3316 3092 3324
rect 3132 3316 3140 3324
rect 3292 3318 3300 3326
rect 2764 3296 2772 3304
rect 3388 3296 3396 3304
rect 3436 3316 3444 3324
rect 3532 3316 3540 3324
rect 3580 3316 3588 3324
rect 3660 3316 3668 3324
rect 3820 3318 3828 3326
rect 3932 3316 3940 3324
rect 3996 3316 4004 3324
rect 4124 3316 4132 3324
rect 4172 3316 4180 3324
rect 4188 3316 4196 3324
rect 4236 3316 4244 3324
rect 4252 3316 4260 3324
rect 4348 3316 4356 3324
rect 4508 3316 4516 3324
rect 4620 3316 4628 3324
rect 4652 3316 4660 3324
rect 4668 3316 4676 3324
rect 4732 3316 4740 3324
rect 4748 3316 4756 3324
rect 4908 3316 4916 3324
rect 5068 3316 5076 3324
rect 5100 3316 5108 3324
rect 3932 3296 3940 3304
rect 3964 3296 3972 3304
rect 3980 3296 3988 3304
rect 4108 3296 4116 3304
rect 4156 3296 4164 3304
rect 4300 3296 4308 3304
rect 4380 3296 4388 3304
rect 4588 3296 4596 3304
rect 4716 3296 4724 3304
rect 12 3276 20 3284
rect 1612 3276 1620 3284
rect 1804 3276 1812 3284
rect 2140 3276 2148 3284
rect 2204 3276 2212 3284
rect 3164 3276 3172 3284
rect 3436 3276 3444 3284
rect 3692 3276 3700 3284
rect 4012 3276 4020 3284
rect 4140 3276 4148 3284
rect 4172 3276 4180 3284
rect 4252 3276 4260 3284
rect 4268 3276 4276 3284
rect 4684 3276 4692 3284
rect 4796 3276 4804 3284
rect 812 3236 820 3244
rect 940 3236 948 3244
rect 2908 3236 2916 3244
rect 3004 3236 3012 3244
rect 3116 3236 3124 3244
rect 3996 3236 4004 3244
rect 4700 3236 4708 3244
rect 5020 3236 5028 3244
rect 5132 3236 5140 3244
rect 1043 3206 1051 3214
rect 1053 3206 1061 3214
rect 1063 3206 1071 3214
rect 1073 3206 1081 3214
rect 1083 3206 1091 3214
rect 1093 3206 1101 3214
rect 4051 3206 4059 3214
rect 4061 3206 4069 3214
rect 4071 3206 4079 3214
rect 4081 3206 4089 3214
rect 4091 3206 4099 3214
rect 4101 3206 4109 3214
rect 124 3176 132 3184
rect 588 3176 596 3184
rect 652 3176 660 3184
rect 748 3176 756 3184
rect 1228 3176 1236 3184
rect 2204 3176 2212 3184
rect 2684 3176 2692 3184
rect 3996 3176 4004 3184
rect 4924 3176 4932 3184
rect 540 3156 548 3164
rect 60 3136 68 3144
rect 252 3136 260 3144
rect 444 3136 452 3144
rect 812 3136 820 3144
rect 2236 3136 2244 3144
rect 2364 3136 2372 3144
rect 3036 3136 3044 3144
rect 3788 3136 3796 3144
rect 3980 3136 3988 3144
rect 4076 3136 4084 3144
rect 4348 3136 4356 3144
rect 476 3116 484 3124
rect 508 3116 516 3124
rect 620 3116 628 3124
rect 780 3116 788 3124
rect 1132 3116 1140 3124
rect 44 3096 52 3104
rect 92 3096 100 3104
rect 380 3094 388 3102
rect 476 3096 484 3104
rect 540 3096 548 3104
rect 604 3096 612 3104
rect 668 3096 676 3104
rect 732 3096 740 3104
rect 748 3096 756 3104
rect 828 3096 836 3104
rect 908 3096 916 3104
rect 1292 3116 1300 3124
rect 1948 3116 1956 3124
rect 1180 3096 1188 3104
rect 1228 3096 1236 3104
rect 1260 3096 1268 3104
rect 1324 3096 1332 3104
rect 1372 3096 1380 3104
rect 1420 3096 1428 3104
rect 1436 3096 1444 3104
rect 1468 3096 1476 3104
rect 1564 3096 1572 3104
rect 1628 3094 1636 3102
rect 1756 3096 1764 3104
rect 1996 3116 2004 3124
rect 2268 3116 2276 3124
rect 2652 3116 2660 3124
rect 2924 3116 2932 3124
rect 3260 3116 3268 3124
rect 1820 3094 1828 3102
rect 1996 3096 2004 3104
rect 2076 3094 2084 3102
rect 2140 3096 2148 3104
rect 2236 3096 2244 3104
rect 2268 3096 2276 3104
rect 2364 3096 2372 3104
rect 2380 3096 2388 3104
rect 2428 3096 2436 3104
rect 2476 3096 2484 3104
rect 12 3076 20 3084
rect 236 3076 244 3084
rect 364 3076 372 3084
rect 492 3076 500 3084
rect 556 3076 564 3084
rect 732 3076 740 3084
rect 860 3076 868 3084
rect 1036 3076 1044 3084
rect 1148 3076 1156 3084
rect 1196 3076 1204 3084
rect 1212 3076 1220 3084
rect 1340 3076 1348 3084
rect 1916 3076 1924 3084
rect 2012 3076 2020 3084
rect 2044 3076 2052 3084
rect 2220 3076 2228 3084
rect 2380 3076 2388 3084
rect 2460 3076 2468 3084
rect 2524 3076 2532 3084
rect 2604 3096 2612 3104
rect 2684 3096 2692 3104
rect 2716 3096 2724 3104
rect 2780 3096 2788 3104
rect 2796 3096 2804 3104
rect 2812 3096 2820 3104
rect 2828 3096 2836 3104
rect 2892 3096 2900 3104
rect 2924 3096 2932 3104
rect 2956 3096 2964 3104
rect 2988 3096 2996 3104
rect 3372 3116 3380 3124
rect 3164 3094 3172 3102
rect 3308 3096 3316 3104
rect 3676 3116 3684 3124
rect 3404 3096 3412 3104
rect 3420 3096 3428 3104
rect 3532 3096 3540 3104
rect 3948 3116 3956 3124
rect 4268 3116 4276 3124
rect 4300 3116 4308 3124
rect 4780 3116 4788 3124
rect 3580 3094 3588 3102
rect 3724 3096 3732 3104
rect 3884 3094 3892 3102
rect 3964 3096 3972 3104
rect 4204 3094 4212 3102
rect 4316 3096 4324 3104
rect 4460 3096 4468 3104
rect 4716 3094 4724 3102
rect 4780 3096 4788 3104
rect 4828 3096 4836 3104
rect 5052 3096 5060 3104
rect 2700 3076 2708 3084
rect 2732 3076 2740 3084
rect 2876 3076 2884 3084
rect 2908 3076 2916 3084
rect 2972 3076 2980 3084
rect 2988 3076 2996 3084
rect 3228 3076 3236 3084
rect 3276 3076 3284 3084
rect 3324 3076 3332 3084
rect 3340 3076 3348 3084
rect 3436 3076 3444 3084
rect 3612 3076 3620 3084
rect 3644 3076 3652 3084
rect 3676 3076 3684 3084
rect 3740 3076 3748 3084
rect 3916 3076 3924 3084
rect 4188 3076 4196 3084
rect 4524 3076 4532 3084
rect 4572 3076 4580 3084
rect 4652 3076 4660 3084
rect 4748 3076 4756 3084
rect 5036 3076 5044 3084
rect 572 3056 580 3064
rect 796 3056 804 3064
rect 892 3056 900 3064
rect 1484 3056 1492 3064
rect 1884 3056 1892 3064
rect 1900 3056 1908 3064
rect 2332 3056 2340 3064
rect 2636 3056 2644 3064
rect 3020 3056 3028 3064
rect 3164 3056 3172 3064
rect 4348 3056 4356 3064
rect 4860 3056 4868 3064
rect 4876 3056 4884 3064
rect 124 3036 132 3044
rect 684 3036 692 3044
rect 1036 3036 1044 3044
rect 1388 3036 1396 3044
rect 1500 3036 1508 3044
rect 1692 3036 1700 3044
rect 2316 3036 2324 3044
rect 2428 3036 2436 3044
rect 2476 3036 2484 3044
rect 3452 3036 3460 3044
rect 3756 3036 3764 3044
rect 4556 3036 4564 3044
rect 4588 3036 4596 3044
rect 4892 3036 4900 3044
rect 4924 3036 4932 3044
rect 5084 3036 5092 3044
rect 2547 3006 2555 3014
rect 2557 3006 2565 3014
rect 2567 3006 2575 3014
rect 2577 3006 2585 3014
rect 2587 3006 2595 3014
rect 2597 3006 2605 3014
rect 12 2976 20 2984
rect 396 2976 404 2984
rect 716 2976 724 2984
rect 1404 2976 1412 2984
rect 1580 2976 1588 2984
rect 1692 2976 1700 2984
rect 1820 2976 1828 2984
rect 2060 2976 2068 2984
rect 2252 2976 2260 2984
rect 3068 2976 3076 2984
rect 3500 2976 3508 2984
rect 4028 2976 4036 2984
rect 4204 2976 4212 2984
rect 4364 2976 4372 2984
rect 4716 2976 4724 2984
rect 700 2956 708 2964
rect 1036 2956 1044 2964
rect 1308 2956 1316 2964
rect 1596 2956 1604 2964
rect 1772 2956 1780 2964
rect 2668 2956 2676 2964
rect 2940 2956 2948 2964
rect 3084 2956 3092 2964
rect 4620 2956 4628 2964
rect 124 2936 132 2944
rect 364 2936 372 2944
rect 588 2936 596 2944
rect 620 2936 628 2944
rect 652 2936 660 2944
rect 684 2936 692 2944
rect 748 2936 756 2944
rect 844 2936 852 2944
rect 860 2936 868 2944
rect 956 2936 964 2944
rect 988 2936 996 2944
rect 1260 2936 1268 2944
rect 1452 2936 1460 2944
rect 1516 2936 1524 2944
rect 1532 2936 1540 2944
rect 1644 2936 1652 2944
rect 1756 2936 1764 2944
rect 1980 2936 1988 2944
rect 2012 2936 2020 2944
rect 2108 2936 2116 2944
rect 2124 2936 2132 2944
rect 2236 2936 2244 2944
rect 2348 2936 2356 2944
rect 2524 2936 2532 2944
rect 2668 2936 2676 2944
rect 2716 2936 2724 2944
rect 2780 2936 2788 2944
rect 2796 2936 2804 2944
rect 2828 2936 2836 2944
rect 2860 2936 2868 2944
rect 2940 2936 2948 2944
rect 3036 2936 3044 2944
rect 3084 2936 3092 2944
rect 3132 2936 3140 2944
rect 3228 2936 3236 2944
rect 3292 2936 3300 2944
rect 3612 2936 3620 2944
rect 3660 2936 3668 2944
rect 3692 2936 3700 2944
rect 3788 2936 3796 2944
rect 3820 2936 3828 2944
rect 3916 2936 3924 2944
rect 3948 2936 3956 2944
rect 4076 2936 4084 2944
rect 4156 2936 4164 2944
rect 4236 2936 4244 2944
rect 4252 2936 4260 2944
rect 4316 2936 4324 2944
rect 4348 2936 4356 2944
rect 4524 2936 4532 2944
rect 4700 2936 4708 2944
rect 4876 2936 4884 2944
rect 140 2918 148 2926
rect 268 2916 276 2924
rect 332 2918 340 2926
rect 460 2916 468 2924
rect 524 2918 532 2926
rect 700 2916 708 2924
rect 732 2916 740 2924
rect 428 2896 436 2904
rect 636 2896 644 2904
rect 780 2896 788 2904
rect 812 2916 820 2924
rect 828 2916 836 2924
rect 860 2916 868 2924
rect 940 2916 948 2924
rect 972 2916 980 2924
rect 1004 2916 1012 2924
rect 1020 2916 1028 2924
rect 1180 2916 1188 2924
rect 1228 2916 1236 2924
rect 1244 2916 1252 2924
rect 1260 2916 1268 2924
rect 1340 2916 1348 2924
rect 1356 2916 1364 2924
rect 1372 2916 1380 2924
rect 1420 2916 1428 2924
rect 1468 2916 1476 2924
rect 1500 2916 1508 2924
rect 1548 2916 1556 2924
rect 1628 2916 1636 2924
rect 1644 2916 1652 2924
rect 908 2896 916 2904
rect 1580 2896 1588 2904
rect 1612 2896 1620 2904
rect 1740 2916 1748 2924
rect 1804 2916 1812 2924
rect 1948 2918 1956 2926
rect 2028 2916 2036 2924
rect 1708 2896 1716 2904
rect 2140 2916 2148 2924
rect 2076 2896 2084 2904
rect 2172 2896 2180 2904
rect 2204 2916 2212 2924
rect 2220 2916 2228 2924
rect 2332 2916 2340 2924
rect 2444 2916 2452 2924
rect 2460 2916 2468 2924
rect 2508 2916 2516 2924
rect 2636 2916 2644 2924
rect 2700 2916 2708 2924
rect 2716 2916 2724 2924
rect 2764 2916 2772 2924
rect 2812 2916 2820 2924
rect 2876 2916 2884 2924
rect 2972 2916 2980 2924
rect 3004 2916 3012 2924
rect 3020 2916 3028 2924
rect 3052 2916 3060 2924
rect 3116 2916 3124 2924
rect 3148 2916 3156 2924
rect 3212 2916 3220 2924
rect 3276 2916 3284 2924
rect 3292 2916 3300 2924
rect 3324 2916 3332 2924
rect 3372 2916 3380 2924
rect 3404 2916 3412 2924
rect 3420 2916 3428 2924
rect 3468 2916 3476 2924
rect 3612 2916 3620 2924
rect 2604 2896 2612 2904
rect 2844 2896 2852 2904
rect 2988 2896 2996 2904
rect 3180 2896 3188 2904
rect 3244 2896 3252 2904
rect 3356 2896 3364 2904
rect 3724 2896 3732 2904
rect 3756 2916 3764 2924
rect 3788 2916 3796 2924
rect 3964 2918 3972 2926
rect 4060 2916 4068 2924
rect 4268 2916 4276 2924
rect 4028 2896 4036 2904
rect 4204 2896 4212 2904
rect 4444 2916 4452 2924
rect 4556 2916 4564 2924
rect 4572 2916 4580 2924
rect 4668 2916 4676 2924
rect 4796 2916 4804 2924
rect 4828 2916 4836 2924
rect 4924 2916 4932 2924
rect 4988 2916 4996 2924
rect 5052 2916 5060 2924
rect 4316 2896 4324 2904
rect 4700 2896 4708 2904
rect 4924 2896 4932 2904
rect 4972 2896 4980 2904
rect 5036 2896 5044 2904
rect 2700 2876 2708 2884
rect 2876 2876 2884 2884
rect 4588 2876 4596 2884
rect 4620 2876 4628 2884
rect 4748 2876 4756 2884
rect 4940 2876 4948 2884
rect 4972 2876 4980 2884
rect 5068 2876 5076 2884
rect 3276 2856 3284 2864
rect 3804 2856 3812 2864
rect 204 2836 212 2844
rect 1196 2836 1204 2844
rect 1340 2836 1348 2844
rect 1468 2836 1476 2844
rect 2476 2836 2484 2844
rect 2732 2836 2740 2844
rect 3436 2836 3444 2844
rect 3836 2836 3844 2844
rect 4220 2836 4228 2844
rect 4924 2836 4932 2844
rect 4988 2836 4996 2844
rect 5084 2836 5092 2844
rect 1043 2806 1051 2814
rect 1053 2806 1061 2814
rect 1063 2806 1071 2814
rect 1073 2806 1081 2814
rect 1083 2806 1091 2814
rect 1093 2806 1101 2814
rect 4051 2806 4059 2814
rect 4061 2806 4069 2814
rect 4071 2806 4079 2814
rect 4081 2806 4089 2814
rect 4091 2806 4099 2814
rect 4101 2806 4109 2814
rect 1132 2776 1140 2784
rect 1292 2776 1300 2784
rect 1500 2776 1508 2784
rect 2060 2776 2068 2784
rect 2268 2776 2276 2784
rect 2460 2776 2468 2784
rect 2572 2776 2580 2784
rect 2636 2776 2644 2784
rect 2956 2776 2964 2784
rect 3100 2776 3108 2784
rect 3324 2776 3332 2784
rect 3964 2776 3972 2784
rect 4700 2776 4708 2784
rect 5004 2776 5012 2784
rect 5100 2776 5108 2784
rect 476 2756 484 2764
rect 4572 2756 4580 2764
rect 796 2736 804 2744
rect 1964 2736 1972 2744
rect 2908 2736 2916 2744
rect 3196 2736 3204 2744
rect 3756 2736 3764 2744
rect 3916 2736 3924 2744
rect 4588 2736 4596 2744
rect 4620 2736 4628 2744
rect 4716 2736 4724 2744
rect 60 2716 68 2724
rect 172 2716 180 2724
rect 380 2716 388 2724
rect 444 2716 452 2724
rect 556 2716 564 2724
rect 572 2716 580 2724
rect 636 2716 644 2724
rect 700 2716 708 2724
rect 764 2716 772 2724
rect 828 2716 836 2724
rect 892 2716 900 2724
rect 1260 2716 1268 2724
rect 1420 2716 1428 2724
rect 1804 2716 1812 2724
rect 44 2696 52 2704
rect 140 2696 148 2704
rect 172 2696 180 2704
rect 268 2696 276 2704
rect 316 2694 324 2702
rect 412 2696 420 2704
rect 476 2696 484 2704
rect 540 2696 548 2704
rect 588 2696 596 2704
rect 604 2696 612 2704
rect 652 2696 660 2704
rect 668 2696 676 2704
rect 716 2696 724 2704
rect 732 2696 740 2704
rect 828 2696 836 2704
rect 860 2696 868 2704
rect 876 2696 884 2704
rect 924 2696 932 2704
rect 1004 2694 1012 2702
rect 1292 2696 1300 2704
rect 1340 2696 1348 2704
rect 1388 2696 1396 2704
rect 1436 2696 1444 2704
rect 1468 2696 1476 2704
rect 1484 2696 1492 2704
rect 1532 2696 1540 2704
rect 1612 2696 1620 2704
rect 1740 2696 1748 2704
rect 1836 2696 1844 2704
rect 1932 2716 1940 2724
rect 2092 2716 2100 2724
rect 2380 2716 2388 2724
rect 2860 2716 2868 2724
rect 1900 2696 1908 2704
rect 1964 2696 1972 2704
rect 2028 2696 2036 2704
rect 2076 2696 2084 2704
rect 2124 2696 2132 2704
rect 2140 2696 2148 2704
rect 2204 2696 2212 2704
rect 2236 2696 2244 2704
rect 2252 2696 2260 2704
rect 2300 2696 2308 2704
rect 2332 2696 2340 2704
rect 2348 2696 2356 2704
rect 2396 2696 2404 2704
rect 2412 2696 2420 2704
rect 2444 2696 2452 2704
rect 2492 2696 2500 2704
rect 2524 2696 2532 2704
rect 2700 2696 2708 2704
rect 3036 2716 3044 2724
rect 3068 2716 3076 2724
rect 2764 2694 2772 2702
rect 2908 2696 2916 2704
rect 2956 2696 2964 2704
rect 2988 2696 2996 2704
rect 12 2676 20 2684
rect 108 2676 116 2684
rect 380 2676 388 2684
rect 428 2676 436 2684
rect 492 2676 500 2684
rect 620 2676 628 2684
rect 684 2676 692 2684
rect 748 2676 756 2684
rect 812 2676 820 2684
rect 876 2676 884 2684
rect 940 2676 948 2684
rect 1020 2676 1028 2684
rect 1212 2676 1220 2684
rect 1276 2676 1284 2684
rect 1340 2676 1348 2684
rect 1564 2676 1572 2684
rect 1788 2676 1796 2684
rect 1852 2676 1860 2684
rect 1916 2676 1924 2684
rect 1996 2676 2004 2684
rect 2044 2676 2052 2684
rect 2108 2676 2116 2684
rect 2140 2676 2148 2684
rect 2156 2676 2164 2684
rect 2188 2676 2196 2684
rect 2220 2676 2228 2684
rect 2828 2676 2836 2684
rect 2924 2676 2932 2684
rect 2940 2676 2948 2684
rect 3020 2696 3028 2704
rect 3036 2696 3044 2704
rect 3084 2696 3092 2704
rect 3132 2696 3140 2704
rect 3228 2696 3236 2704
rect 3516 2716 3524 2724
rect 3580 2716 3588 2724
rect 3676 2716 3684 2724
rect 3292 2696 3300 2704
rect 3388 2696 3396 2704
rect 3452 2694 3460 2702
rect 3532 2696 3540 2704
rect 3564 2696 3572 2704
rect 3596 2696 3604 2704
rect 3612 2696 3620 2704
rect 3724 2696 3732 2704
rect 3788 2696 3796 2704
rect 3804 2696 3812 2704
rect 3884 2696 3892 2704
rect 4028 2716 4036 2724
rect 3964 2696 3972 2704
rect 3020 2676 3028 2684
rect 3180 2676 3188 2684
rect 3244 2676 3252 2684
rect 3260 2676 3268 2684
rect 3308 2676 3316 2684
rect 3564 2676 3572 2684
rect 3628 2676 3636 2684
rect 3644 2676 3652 2684
rect 3740 2676 3748 2684
rect 3836 2676 3844 2684
rect 3996 2696 4004 2704
rect 4204 2716 4212 2724
rect 4220 2716 4228 2724
rect 4284 2716 4292 2724
rect 4540 2716 4548 2724
rect 4556 2716 4564 2724
rect 4988 2716 4996 2724
rect 4140 2696 4148 2704
rect 4220 2696 4228 2704
rect 4252 2696 4260 2704
rect 4300 2696 4308 2704
rect 4316 2696 4324 2704
rect 4508 2696 4516 2704
rect 4572 2696 4580 2704
rect 4652 2696 4660 2704
rect 4796 2696 4804 2704
rect 4844 2694 4852 2702
rect 4956 2696 4964 2704
rect 5036 2696 5044 2704
rect 3996 2676 4004 2684
rect 4156 2676 4164 2684
rect 4172 2676 4180 2684
rect 4268 2676 4276 2684
rect 4332 2676 4340 2684
rect 4348 2676 4356 2684
rect 4476 2676 4484 2684
rect 4492 2676 4500 2684
rect 4972 2676 4980 2684
rect 828 2656 836 2664
rect 1356 2656 1364 2664
rect 1404 2656 1412 2664
rect 1452 2656 1460 2664
rect 1772 2656 1780 2664
rect 1996 2656 2004 2664
rect 2044 2656 2052 2664
rect 3116 2656 3124 2664
rect 3164 2656 3172 2664
rect 3852 2656 3860 2664
rect 4908 2656 4916 2664
rect 60 2636 68 2644
rect 1260 2636 1268 2644
rect 1372 2636 1380 2644
rect 1500 2636 1508 2644
rect 1724 2636 1732 2644
rect 1868 2636 1876 2644
rect 3692 2636 3700 2644
rect 4044 2636 4052 2644
rect 4188 2636 4196 2644
rect 4540 2636 4548 2644
rect 2547 2606 2555 2614
rect 2557 2606 2565 2614
rect 2567 2606 2575 2614
rect 2577 2606 2585 2614
rect 2587 2606 2595 2614
rect 2597 2606 2605 2614
rect 572 2576 580 2584
rect 860 2576 868 2584
rect 1820 2576 1828 2584
rect 1884 2576 1892 2584
rect 2028 2576 2036 2584
rect 2652 2576 2660 2584
rect 3068 2576 3076 2584
rect 3084 2576 3092 2584
rect 3132 2576 3140 2584
rect 3548 2576 3556 2584
rect 3740 2576 3748 2584
rect 3932 2576 3940 2584
rect 4284 2576 4292 2584
rect 4492 2576 4500 2584
rect 4508 2576 4516 2584
rect 4796 2576 4804 2584
rect 5052 2576 5060 2584
rect 636 2556 644 2564
rect 732 2556 740 2564
rect 1324 2556 1332 2564
rect 1404 2556 1412 2564
rect 1836 2556 1844 2564
rect 2636 2556 2644 2564
rect 2668 2556 2676 2564
rect 2860 2556 2868 2564
rect 3532 2556 3540 2564
rect 4476 2556 4484 2564
rect 4636 2556 4644 2564
rect 4700 2556 4708 2564
rect 5132 2556 5140 2564
rect 60 2536 68 2544
rect 268 2536 276 2544
rect 348 2536 356 2544
rect 364 2536 372 2544
rect 492 2536 500 2544
rect 508 2536 516 2544
rect 556 2536 564 2544
rect 636 2536 644 2544
rect 876 2536 884 2544
rect 908 2536 916 2544
rect 972 2536 980 2544
rect 1132 2536 1140 2544
rect 1148 2536 1156 2544
rect 1212 2536 1220 2544
rect 1580 2536 1588 2544
rect 1612 2536 1620 2544
rect 1660 2536 1668 2544
rect 1724 2536 1732 2544
rect 1980 2536 1988 2544
rect 2236 2536 2244 2544
rect 44 2516 52 2524
rect 236 2518 244 2526
rect 300 2516 308 2524
rect 332 2516 340 2524
rect 540 2516 548 2524
rect 604 2516 612 2524
rect 620 2516 628 2524
rect 668 2516 676 2524
rect 764 2516 772 2524
rect 780 2516 788 2524
rect 300 2496 308 2504
rect 508 2496 516 2504
rect 572 2496 580 2504
rect 908 2496 916 2504
rect 956 2516 964 2524
rect 988 2516 996 2524
rect 1004 2516 1012 2524
rect 1132 2516 1140 2524
rect 1164 2516 1172 2524
rect 1196 2516 1204 2524
rect 1228 2516 1236 2524
rect 1244 2516 1252 2524
rect 1292 2516 1300 2524
rect 1356 2516 1364 2524
rect 1372 2516 1380 2524
rect 1548 2518 1556 2526
rect 1628 2516 1636 2524
rect 1340 2496 1348 2504
rect 1708 2516 1716 2524
rect 1740 2516 1748 2524
rect 1788 2516 1796 2524
rect 1868 2516 1876 2524
rect 1916 2516 1924 2524
rect 1964 2516 1972 2524
rect 1996 2516 2004 2524
rect 2060 2516 2068 2524
rect 2108 2516 2116 2524
rect 2124 2516 2132 2524
rect 2140 2516 2148 2524
rect 2156 2516 2164 2524
rect 2204 2516 2212 2524
rect 2252 2516 2260 2524
rect 2284 2516 2292 2524
rect 2348 2516 2356 2524
rect 2380 2536 2388 2544
rect 2444 2536 2452 2544
rect 2508 2536 2516 2544
rect 2924 2536 2932 2544
rect 2956 2536 2964 2544
rect 3020 2536 3028 2544
rect 3324 2536 3332 2544
rect 3372 2536 3380 2544
rect 3420 2536 3428 2544
rect 3484 2536 3492 2544
rect 3516 2536 3524 2544
rect 3660 2536 3668 2544
rect 3708 2536 3716 2544
rect 3836 2536 3844 2544
rect 4092 2536 4100 2544
rect 4188 2536 4196 2544
rect 4236 2536 4244 2544
rect 4268 2536 4276 2544
rect 4412 2536 4420 2544
rect 2396 2516 2404 2524
rect 1676 2496 1684 2504
rect 1932 2496 1940 2504
rect 1964 2496 1972 2504
rect 2460 2516 2468 2524
rect 2508 2516 2516 2524
rect 2524 2516 2532 2524
rect 2556 2516 2564 2524
rect 2604 2516 2612 2524
rect 2620 2516 2628 2524
rect 2684 2516 2692 2524
rect 2860 2518 2868 2526
rect 2956 2496 2964 2504
rect 3004 2516 3012 2524
rect 3036 2516 3044 2524
rect 3116 2516 3124 2524
rect 3196 2516 3204 2524
rect 3260 2518 3268 2526
rect 3356 2496 3364 2504
rect 3404 2516 3412 2524
rect 3436 2516 3444 2524
rect 3676 2518 3684 2526
rect 3868 2518 3876 2526
rect 4060 2518 4068 2526
rect 4220 2516 4228 2524
rect 4396 2516 4404 2524
rect 4572 2516 4580 2524
rect 4636 2518 4644 2526
rect 4748 2516 4756 2524
rect 4860 2516 4868 2524
rect 4908 2516 4916 2524
rect 5020 2516 5028 2524
rect 5100 2516 5108 2524
rect 4172 2496 4180 2504
rect 4748 2496 4756 2504
rect 4780 2496 4788 2504
rect 5036 2496 5044 2504
rect 5052 2496 5060 2504
rect 12 2476 20 2484
rect 1164 2476 1172 2484
rect 1420 2476 1428 2484
rect 2252 2476 2260 2484
rect 2316 2476 2324 2484
rect 2396 2476 2404 2484
rect 2524 2476 2532 2484
rect 2732 2476 2740 2484
rect 3468 2476 3476 2484
rect 5004 2476 5012 2484
rect 5020 2456 5028 2464
rect 108 2436 116 2444
rect 1276 2436 1284 2444
rect 1372 2436 1380 2444
rect 1772 2436 1780 2444
rect 2076 2436 2084 2444
rect 2188 2436 2196 2444
rect 2476 2436 2484 2444
rect 2716 2436 2724 2444
rect 4252 2436 4260 2444
rect 1043 2406 1051 2414
rect 1053 2406 1061 2414
rect 1063 2406 1071 2414
rect 1073 2406 1081 2414
rect 1083 2406 1091 2414
rect 1093 2406 1101 2414
rect 4051 2406 4059 2414
rect 4061 2406 4069 2414
rect 4071 2406 4079 2414
rect 4081 2406 4089 2414
rect 4091 2406 4099 2414
rect 4101 2406 4109 2414
rect 124 2376 132 2384
rect 1420 2376 1428 2384
rect 1532 2376 1540 2384
rect 1964 2376 1972 2384
rect 2444 2376 2452 2384
rect 3212 2376 3220 2384
rect 3612 2376 3620 2384
rect 3916 2376 3924 2384
rect 4332 2376 4340 2384
rect 620 2356 628 2364
rect 1932 2356 1940 2364
rect 2492 2356 2500 2364
rect 4828 2356 4836 2364
rect 12 2336 20 2344
rect 60 2336 68 2344
rect 156 2336 164 2344
rect 188 2336 196 2344
rect 1244 2336 1252 2344
rect 3052 2336 3060 2344
rect 4364 2336 4372 2344
rect 4412 2336 4420 2344
rect 4588 2336 4596 2344
rect 4812 2336 4820 2344
rect 5132 2336 5140 2344
rect 220 2316 228 2324
rect 476 2316 484 2324
rect 492 2316 500 2324
rect 556 2316 564 2324
rect 812 2316 820 2324
rect 876 2316 884 2324
rect 940 2316 948 2324
rect 1340 2316 1348 2324
rect 1452 2316 1460 2324
rect 1788 2316 1796 2324
rect 1884 2316 1892 2324
rect 44 2296 52 2304
rect 108 2296 116 2304
rect 124 2296 132 2304
rect 188 2296 196 2304
rect 316 2296 324 2304
rect 364 2294 372 2302
rect 444 2296 452 2304
rect 476 2296 484 2304
rect 604 2296 612 2304
rect 684 2296 692 2304
rect 748 2294 756 2302
rect 828 2296 836 2304
rect 908 2296 916 2304
rect 956 2296 964 2304
rect 972 2296 980 2304
rect 1116 2294 1124 2302
rect 1276 2296 1284 2304
rect 1308 2296 1316 2304
rect 1372 2296 1380 2304
rect 108 2276 116 2284
rect 172 2276 180 2284
rect 300 2276 308 2284
rect 428 2276 436 2284
rect 476 2276 484 2284
rect 540 2276 548 2284
rect 604 2276 612 2284
rect 860 2276 868 2284
rect 924 2276 932 2284
rect 988 2276 996 2284
rect 1260 2276 1268 2284
rect 1388 2276 1396 2284
rect 1420 2296 1428 2304
rect 1468 2296 1476 2304
rect 1548 2296 1556 2304
rect 1580 2296 1588 2304
rect 1596 2296 1604 2304
rect 1628 2296 1636 2304
rect 1644 2296 1652 2304
rect 1676 2296 1684 2304
rect 1772 2296 1780 2304
rect 1804 2296 1812 2304
rect 1820 2296 1828 2304
rect 2140 2316 2148 2324
rect 2284 2316 2292 2324
rect 2684 2316 2692 2324
rect 1948 2296 1956 2304
rect 1996 2296 2004 2304
rect 2012 2296 2020 2304
rect 2028 2296 2036 2304
rect 2076 2296 2084 2304
rect 2108 2296 2116 2304
rect 2172 2296 2180 2304
rect 2188 2296 2196 2304
rect 2220 2296 2228 2304
rect 2252 2296 2260 2304
rect 2332 2296 2340 2304
rect 2380 2296 2388 2304
rect 2428 2296 2436 2304
rect 2476 2296 2484 2304
rect 2524 2296 2532 2304
rect 2620 2296 2628 2304
rect 2652 2296 2660 2304
rect 2716 2296 2724 2304
rect 2748 2296 2756 2304
rect 2812 2296 2820 2304
rect 1516 2276 1524 2284
rect 1660 2276 1668 2284
rect 1740 2276 1748 2284
rect 1836 2276 1844 2284
rect 1948 2276 1956 2284
rect 2060 2276 2068 2284
rect 2876 2296 2884 2304
rect 2972 2296 2980 2304
rect 3020 2296 3028 2304
rect 3036 2296 3044 2304
rect 3084 2296 3092 2304
rect 3116 2296 3124 2304
rect 3132 2296 3140 2304
rect 3180 2296 3188 2304
rect 3244 2296 3252 2304
rect 3372 2296 3380 2304
rect 3468 2296 3476 2304
rect 3484 2296 3492 2304
rect 3516 2316 3524 2324
rect 3868 2316 3876 2324
rect 3900 2316 3908 2324
rect 3996 2316 4004 2324
rect 3548 2296 3556 2304
rect 3580 2296 3588 2304
rect 3708 2296 3716 2304
rect 3756 2294 3764 2302
rect 3868 2296 3876 2304
rect 3948 2296 3956 2304
rect 4380 2316 4388 2324
rect 4444 2316 4452 2324
rect 4508 2316 4516 2324
rect 4844 2316 4852 2324
rect 4860 2316 4868 2324
rect 4028 2296 4036 2304
rect 4044 2296 4052 2304
rect 4252 2296 4260 2304
rect 4364 2296 4372 2304
rect 4428 2296 4436 2304
rect 4492 2296 4500 2304
rect 4540 2296 4548 2304
rect 4716 2296 4724 2304
rect 4828 2296 4836 2304
rect 4860 2296 4868 2304
rect 4892 2296 4900 2304
rect 5004 2294 5012 2302
rect 2204 2276 2212 2284
rect 2332 2276 2340 2284
rect 2604 2276 2612 2284
rect 2636 2276 2644 2284
rect 2732 2276 2740 2284
rect 2796 2276 2804 2284
rect 2844 2276 2852 2284
rect 2860 2276 2868 2284
rect 2892 2276 2900 2284
rect 2924 2276 2932 2284
rect 3004 2276 3012 2284
rect 3388 2276 3396 2284
rect 3452 2276 3460 2284
rect 3564 2276 3572 2284
rect 3964 2276 3972 2284
rect 4124 2276 4132 2284
rect 4300 2276 4308 2284
rect 4412 2276 4420 2284
rect 4764 2276 4772 2284
rect 4972 2276 4980 2284
rect 1116 2256 1124 2264
rect 1468 2256 1476 2264
rect 1500 2256 1508 2264
rect 1516 2256 1524 2264
rect 1740 2256 1748 2264
rect 2044 2256 2052 2264
rect 2348 2256 2356 2264
rect 2380 2256 2388 2264
rect 2748 2256 2756 2264
rect 2780 2256 2788 2264
rect 2940 2256 2948 2264
rect 3820 2256 3828 2264
rect 4508 2256 4516 2264
rect 4588 2256 4596 2264
rect 4940 2256 4948 2264
rect 1276 2236 1284 2244
rect 1676 2236 1684 2244
rect 2076 2236 2084 2244
rect 2220 2236 2228 2244
rect 2396 2236 2404 2244
rect 2988 2236 2996 2244
rect 3148 2236 3156 2244
rect 3260 2236 3268 2244
rect 3628 2236 3636 2244
rect 4140 2236 4148 2244
rect 4460 2236 4468 2244
rect 2547 2206 2555 2214
rect 2557 2206 2565 2214
rect 2567 2206 2575 2214
rect 2577 2206 2585 2214
rect 2587 2206 2595 2214
rect 2597 2206 2605 2214
rect 92 2176 100 2184
rect 636 2176 644 2184
rect 684 2176 692 2184
rect 908 2176 916 2184
rect 940 2176 948 2184
rect 1868 2176 1876 2184
rect 2092 2176 2100 2184
rect 2412 2176 2420 2184
rect 2892 2176 2900 2184
rect 3596 2176 3604 2184
rect 3644 2176 3652 2184
rect 3980 2176 3988 2184
rect 4172 2176 4180 2184
rect 4396 2176 4404 2184
rect 4524 2176 4532 2184
rect 4588 2176 4596 2184
rect 4940 2176 4948 2184
rect 300 2156 308 2164
rect 476 2156 484 2164
rect 540 2156 548 2164
rect 588 2156 596 2164
rect 620 2156 628 2164
rect 780 2156 788 2164
rect 1516 2156 1524 2164
rect 2076 2156 2084 2164
rect 2284 2156 2292 2164
rect 4364 2156 4372 2164
rect 4844 2156 4852 2164
rect 108 2136 116 2144
rect 332 2136 340 2144
rect 412 2136 420 2144
rect 524 2136 532 2144
rect 572 2136 580 2144
rect 796 2136 804 2144
rect 924 2136 932 2144
rect 972 2136 980 2144
rect 1004 2136 1012 2144
rect 1068 2136 1076 2144
rect 1148 2136 1156 2144
rect 1276 2136 1284 2144
rect 1308 2136 1316 2144
rect 1692 2136 1700 2144
rect 1964 2136 1972 2144
rect 1996 2136 2004 2144
rect 2060 2136 2068 2144
rect 2124 2136 2132 2144
rect 2220 2136 2228 2144
rect 2780 2136 2788 2144
rect 2876 2136 2884 2144
rect 3052 2136 3060 2144
rect 3388 2136 3396 2144
rect 3468 2136 3476 2144
rect 3580 2136 3588 2144
rect 3836 2136 3844 2144
rect 3884 2136 3892 2144
rect 3932 2136 3940 2144
rect 3996 2136 4004 2144
rect 4156 2136 4164 2144
rect 4332 2136 4340 2144
rect 4380 2136 4388 2144
rect 4428 2136 4436 2144
rect 4508 2136 4516 2144
rect 4748 2136 4756 2144
rect 4876 2136 4884 2144
rect 44 2116 52 2124
rect 60 2116 68 2124
rect 124 2116 132 2124
rect 140 2116 148 2124
rect 300 2118 308 2126
rect 364 2116 372 2124
rect 396 2116 404 2124
rect 412 2116 420 2124
rect 508 2116 516 2124
rect 540 2116 548 2124
rect 620 2116 628 2124
rect 668 2116 676 2124
rect 716 2116 724 2124
rect 812 2116 820 2124
rect 156 2096 164 2104
rect 364 2096 372 2104
rect 956 2096 964 2104
rect 1004 2096 1012 2104
rect 1052 2116 1060 2124
rect 1164 2116 1172 2124
rect 1196 2116 1204 2124
rect 1260 2116 1268 2124
rect 1356 2116 1364 2124
rect 1484 2116 1492 2124
rect 1548 2116 1556 2124
rect 1596 2116 1604 2124
rect 1612 2116 1620 2124
rect 1660 2116 1668 2124
rect 1740 2116 1748 2124
rect 1900 2116 1908 2124
rect 1916 2116 1924 2124
rect 1228 2096 1236 2104
rect 1996 2096 2004 2104
rect 2044 2116 2052 2124
rect 2108 2116 2116 2124
rect 2156 2096 2164 2104
rect 2188 2116 2196 2124
rect 2204 2116 2212 2124
rect 2284 2118 2292 2126
rect 2444 2116 2452 2124
rect 2492 2116 2500 2124
rect 2588 2116 2596 2124
rect 2604 2116 2612 2124
rect 2652 2116 2660 2124
rect 2668 2116 2676 2124
rect 2716 2116 2724 2124
rect 2764 2116 2772 2124
rect 2524 2096 2532 2104
rect 2572 2096 2580 2104
rect 2812 2096 2820 2104
rect 2876 2116 2884 2124
rect 3004 2116 3012 2124
rect 3084 2116 3092 2124
rect 3100 2116 3108 2124
rect 3164 2116 3172 2124
rect 3180 2116 3188 2124
rect 3196 2116 3204 2124
rect 3244 2116 3252 2124
rect 3404 2118 3412 2126
rect 3484 2116 3492 2124
rect 2860 2096 2868 2104
rect 3484 2096 3492 2104
rect 3564 2116 3572 2124
rect 3628 2116 3636 2124
rect 3708 2116 3716 2124
rect 3772 2118 3780 2126
rect 3868 2096 3876 2104
rect 3916 2116 3924 2124
rect 3948 2116 3956 2124
rect 4028 2096 4036 2104
rect 4156 2116 4164 2124
rect 4284 2116 4292 2124
rect 4476 2116 4484 2124
rect 4716 2118 4724 2126
rect 4796 2116 4804 2124
rect 4812 2116 4820 2124
rect 4892 2116 4900 2124
rect 4924 2116 4932 2124
rect 5004 2116 5012 2124
rect 5052 2116 5060 2124
rect 4140 2096 4148 2104
rect 4396 2096 4404 2104
rect 4428 2096 4436 2104
rect 4780 2096 4788 2104
rect 4924 2096 4932 2104
rect 12 2076 20 2084
rect 1180 2076 1188 2084
rect 1468 2076 1476 2084
rect 1484 2076 1492 2084
rect 1628 2076 1636 2084
rect 3212 2076 3220 2084
rect 3532 2076 3540 2084
rect 4460 2076 4468 2084
rect 3116 2056 3124 2064
rect 3276 2056 3284 2064
rect 460 2036 468 2044
rect 1564 2036 1572 2044
rect 1852 2036 1860 2044
rect 1948 2036 1956 2044
rect 2460 2036 2468 2044
rect 2636 2036 2644 2044
rect 2684 2036 2692 2044
rect 2732 2036 2740 2044
rect 4460 2036 4468 2044
rect 4556 2036 4564 2044
rect 1043 2006 1051 2014
rect 1053 2006 1061 2014
rect 1063 2006 1071 2014
rect 1073 2006 1081 2014
rect 1083 2006 1091 2014
rect 1093 2006 1101 2014
rect 4051 2006 4059 2014
rect 4061 2006 4069 2014
rect 4071 2006 4079 2014
rect 4081 2006 4089 2014
rect 4091 2006 4099 2014
rect 4101 2006 4109 2014
rect 140 1976 148 1984
rect 444 1976 452 1984
rect 924 1976 932 1984
rect 1164 1976 1172 1984
rect 1916 1976 1924 1984
rect 2684 1976 2692 1984
rect 2988 1976 2996 1984
rect 3036 1976 3044 1984
rect 3196 1976 3204 1984
rect 3516 1976 3524 1984
rect 4300 1976 4308 1984
rect 4652 1976 4660 1984
rect 4716 1976 4724 1984
rect 1500 1956 1508 1964
rect 1804 1956 1812 1964
rect 1980 1956 1988 1964
rect 2188 1956 2196 1964
rect 2252 1956 2260 1964
rect 2524 1956 2532 1964
rect 4588 1956 4596 1964
rect 5100 1956 5108 1964
rect 876 1936 884 1944
rect 2668 1936 2676 1944
rect 3468 1936 3476 1944
rect 3644 1936 3652 1944
rect 4300 1936 4308 1944
rect 4316 1936 4324 1944
rect 4396 1936 4404 1944
rect 4508 1936 4516 1944
rect 4572 1936 4580 1944
rect 4636 1936 4644 1944
rect 4700 1936 4708 1944
rect 4844 1936 4852 1944
rect 5052 1936 5060 1944
rect 204 1916 212 1924
rect 460 1916 468 1924
rect 524 1916 532 1924
rect 588 1916 596 1924
rect 44 1896 52 1904
rect 60 1896 68 1904
rect 108 1896 116 1904
rect 172 1896 180 1904
rect 348 1894 356 1902
rect 412 1896 420 1904
rect 476 1896 484 1904
rect 556 1896 564 1904
rect 620 1896 628 1904
rect 636 1896 644 1904
rect 684 1896 692 1904
rect 780 1896 788 1904
rect 796 1896 804 1904
rect 892 1896 900 1904
rect 956 1896 964 1904
rect 972 1896 980 1904
rect 1004 1916 1012 1924
rect 1420 1916 1428 1924
rect 1452 1916 1460 1924
rect 1548 1916 1556 1924
rect 1708 1916 1716 1924
rect 1772 1916 1780 1924
rect 1884 1916 1892 1924
rect 2076 1916 2084 1924
rect 2396 1916 2404 1924
rect 1036 1896 1044 1904
rect 1052 1896 1060 1904
rect 1196 1896 1204 1904
rect 1212 1896 1220 1904
rect 1228 1896 1236 1904
rect 1244 1896 1252 1904
rect 1292 1896 1300 1904
rect 1340 1896 1348 1904
rect 1372 1896 1380 1904
rect 1388 1896 1396 1904
rect 12 1876 20 1884
rect 92 1876 100 1884
rect 204 1876 212 1884
rect 332 1876 340 1884
rect 380 1876 388 1884
rect 508 1876 516 1884
rect 572 1876 580 1884
rect 636 1876 644 1884
rect 716 1876 724 1884
rect 940 1876 948 1884
rect 1052 1876 1060 1884
rect 1308 1876 1316 1884
rect 1324 1876 1332 1884
rect 1388 1876 1396 1884
rect 1420 1896 1428 1904
rect 1484 1896 1492 1904
rect 1516 1896 1524 1904
rect 1580 1896 1588 1904
rect 1612 1896 1620 1904
rect 1692 1896 1700 1904
rect 1740 1896 1748 1904
rect 1804 1896 1812 1904
rect 1852 1896 1860 1904
rect 1916 1896 1924 1904
rect 1948 1896 1956 1904
rect 1980 1896 1988 1904
rect 2044 1896 2052 1904
rect 2108 1896 2116 1904
rect 2140 1896 2148 1904
rect 2204 1896 2212 1904
rect 2220 1896 2228 1904
rect 2300 1896 2308 1904
rect 2332 1896 2340 1904
rect 2364 1896 2372 1904
rect 2428 1896 2436 1904
rect 2444 1896 2452 1904
rect 2636 1916 2644 1924
rect 2924 1916 2932 1924
rect 3116 1916 3124 1924
rect 2492 1896 2500 1904
rect 2556 1896 2564 1904
rect 2796 1896 2804 1904
rect 2908 1896 2916 1904
rect 2956 1896 2964 1904
rect 3020 1896 3028 1904
rect 3068 1896 3076 1904
rect 3164 1916 3172 1924
rect 3564 1916 3572 1924
rect 3164 1896 3172 1904
rect 3308 1896 3316 1904
rect 3388 1896 3396 1904
rect 3436 1896 3444 1904
rect 3484 1896 3492 1904
rect 4172 1916 4180 1924
rect 4348 1916 4356 1924
rect 4604 1916 4612 1924
rect 4668 1916 4676 1924
rect 4732 1916 4740 1924
rect 4828 1916 4836 1924
rect 3628 1896 3636 1904
rect 3756 1896 3764 1904
rect 3852 1896 3860 1904
rect 3996 1894 4004 1902
rect 4140 1896 4148 1904
rect 4188 1896 4196 1904
rect 4236 1896 4244 1904
rect 4284 1896 4292 1904
rect 4300 1896 4308 1904
rect 4380 1896 4388 1904
rect 4476 1896 4484 1904
rect 4588 1896 4596 1904
rect 4652 1896 4660 1904
rect 4716 1896 4724 1904
rect 4796 1896 4804 1904
rect 4828 1896 4836 1904
rect 4924 1896 4932 1904
rect 5068 1896 5076 1904
rect 5084 1896 5092 1904
rect 5132 1896 5140 1904
rect 1468 1876 1476 1884
rect 1596 1876 1604 1884
rect 1756 1876 1764 1884
rect 1820 1876 1828 1884
rect 1836 1876 1844 1884
rect 1964 1876 1972 1884
rect 2028 1876 2036 1884
rect 2124 1876 2132 1884
rect 2172 1876 2180 1884
rect 2316 1876 2324 1884
rect 2444 1876 2452 1884
rect 2476 1876 2484 1884
rect 2508 1876 2516 1884
rect 2668 1876 2676 1884
rect 2972 1876 2980 1884
rect 3084 1876 3092 1884
rect 3180 1876 3188 1884
rect 3532 1876 3540 1884
rect 3596 1876 3604 1884
rect 3628 1876 3636 1884
rect 4028 1876 4036 1884
rect 4108 1876 4116 1884
rect 4380 1876 4388 1884
rect 4428 1876 4436 1884
rect 4460 1876 4468 1884
rect 4540 1876 4548 1884
rect 5004 1876 5012 1884
rect 652 1856 660 1864
rect 1644 1856 1652 1864
rect 1660 1856 1668 1864
rect 2012 1856 2020 1864
rect 2172 1856 2180 1864
rect 2812 1856 2820 1864
rect 3324 1856 3332 1864
rect 3772 1856 3780 1864
rect 3836 1856 3844 1864
rect 4748 1856 4756 1864
rect 4972 1856 4980 1864
rect 140 1836 148 1844
rect 588 1836 596 1844
rect 1340 1836 1348 1844
rect 1628 1836 1636 1844
rect 1676 1836 1684 1844
rect 1708 1836 1716 1844
rect 2268 1836 2276 1844
rect 2332 1836 2340 1844
rect 2636 1836 2644 1844
rect 2876 1836 2884 1844
rect 2924 1836 2932 1844
rect 3420 1836 3428 1844
rect 3868 1836 3876 1844
rect 4172 1836 4180 1844
rect 4220 1836 4228 1844
rect 4348 1836 4356 1844
rect 4444 1836 4452 1844
rect 4524 1836 4532 1844
rect 5068 1836 5076 1844
rect 2547 1806 2555 1814
rect 2557 1806 2565 1814
rect 2567 1806 2575 1814
rect 2577 1806 2585 1814
rect 2587 1806 2595 1814
rect 2597 1806 2605 1814
rect 60 1776 68 1784
rect 220 1776 228 1784
rect 284 1776 292 1784
rect 556 1776 564 1784
rect 1036 1776 1044 1784
rect 1228 1776 1236 1784
rect 1532 1776 1540 1784
rect 1580 1776 1588 1784
rect 1772 1776 1780 1784
rect 2076 1776 2084 1784
rect 2252 1776 2260 1784
rect 2460 1776 2468 1784
rect 2684 1776 2692 1784
rect 2940 1776 2948 1784
rect 3356 1776 3364 1784
rect 3468 1776 3476 1784
rect 3772 1776 3780 1784
rect 4268 1776 4276 1784
rect 4364 1776 4372 1784
rect 2636 1756 2644 1764
rect 4332 1756 4340 1764
rect 4428 1756 4436 1764
rect 4492 1756 4500 1764
rect 4508 1756 4516 1764
rect 4524 1756 4532 1764
rect 5052 1756 5060 1764
rect 92 1736 100 1744
rect 140 1736 148 1744
rect 236 1736 244 1744
rect 348 1736 356 1744
rect 380 1736 388 1744
rect 716 1736 724 1744
rect 748 1736 756 1744
rect 796 1736 804 1744
rect 844 1736 852 1744
rect 876 1736 884 1744
rect 1212 1736 1220 1744
rect 1324 1736 1332 1744
rect 1420 1736 1428 1744
rect 1468 1736 1476 1744
rect 1516 1736 1524 1744
rect 2060 1736 2068 1744
rect 2140 1736 2148 1744
rect 2236 1736 2244 1744
rect 2412 1736 2420 1744
rect 2444 1736 2452 1744
rect 2508 1736 2516 1744
rect 2524 1736 2532 1744
rect 2556 1736 2564 1744
rect 2812 1736 2820 1744
rect 2876 1736 2884 1744
rect 2988 1736 2996 1744
rect 3308 1736 3316 1744
rect 3900 1736 3908 1744
rect 3932 1736 3940 1744
rect 4028 1736 4036 1744
rect 4108 1736 4116 1744
rect 4140 1736 4148 1744
rect 4252 1736 4260 1744
rect 4300 1736 4308 1744
rect 4476 1736 4484 1744
rect 4972 1736 4980 1744
rect 5116 1736 5124 1744
rect 124 1716 132 1724
rect 156 1716 164 1724
rect 204 1716 212 1724
rect 316 1716 324 1724
rect 332 1716 340 1724
rect 428 1716 436 1724
rect 668 1716 676 1724
rect 92 1696 100 1704
rect 284 1696 292 1704
rect 300 1696 308 1704
rect 780 1696 788 1704
rect 828 1716 836 1724
rect 940 1716 948 1724
rect 1116 1716 1124 1724
rect 1132 1716 1140 1724
rect 1148 1716 1156 1724
rect 1356 1718 1364 1726
rect 1180 1696 1188 1704
rect 1452 1696 1460 1704
rect 1500 1716 1508 1724
rect 1564 1716 1572 1724
rect 1644 1716 1652 1724
rect 1708 1718 1716 1726
rect 1804 1716 1812 1724
rect 1836 1716 1844 1724
rect 1884 1716 1892 1724
rect 1900 1716 1908 1724
rect 1932 1716 1940 1724
rect 1980 1716 1988 1724
rect 1996 1716 2004 1724
rect 2044 1716 2052 1724
rect 2172 1696 2180 1704
rect 2220 1716 2228 1724
rect 2348 1716 2356 1724
rect 2460 1716 2468 1724
rect 2492 1716 2500 1724
rect 2524 1716 2532 1724
rect 2556 1716 2564 1724
rect 2636 1716 2644 1724
rect 2668 1716 2676 1724
rect 2796 1716 2804 1724
rect 2892 1716 2900 1724
rect 2972 1716 2980 1724
rect 3052 1718 3060 1726
rect 3116 1716 3124 1724
rect 3228 1716 3236 1724
rect 3276 1716 3284 1724
rect 3340 1716 3348 1724
rect 3388 1716 3396 1724
rect 3404 1716 3412 1724
rect 3436 1716 3444 1724
rect 3484 1716 3492 1724
rect 3516 1716 3524 1724
rect 3532 1716 3540 1724
rect 3580 1716 3588 1724
rect 3596 1716 3604 1724
rect 3612 1716 3620 1724
rect 3676 1716 3684 1724
rect 3692 1716 3700 1724
rect 3708 1716 3716 1724
rect 4076 1718 4084 1726
rect 4236 1716 4244 1724
rect 4380 1716 4388 1724
rect 4396 1716 4404 1724
rect 4476 1716 4484 1724
rect 4540 1716 4548 1724
rect 4588 1716 4596 1724
rect 4604 1716 4612 1724
rect 4652 1716 4660 1724
rect 4700 1716 4708 1724
rect 4780 1716 4788 1724
rect 4796 1716 4804 1724
rect 4812 1716 4820 1724
rect 4988 1718 4996 1726
rect 5100 1716 5108 1724
rect 3548 1696 3556 1704
rect 3900 1696 3908 1704
rect 3916 1696 3924 1704
rect 4204 1696 4212 1704
rect 4268 1696 4276 1704
rect 4300 1696 4308 1704
rect 5132 1696 5140 1704
rect 188 1676 196 1684
rect 2924 1676 2932 1684
rect 3932 1676 3940 1684
rect 4364 1676 4372 1684
rect 4620 1676 4628 1684
rect 4684 1676 4692 1684
rect 4732 1676 4740 1684
rect 4764 1676 4772 1684
rect 4860 1676 4868 1684
rect 3740 1656 3748 1664
rect 60 1636 68 1644
rect 540 1636 548 1644
rect 1772 1636 1780 1644
rect 1852 1636 1860 1644
rect 1948 1636 1956 1644
rect 2012 1636 2020 1644
rect 2108 1636 2116 1644
rect 2220 1636 2228 1644
rect 2684 1636 2692 1644
rect 3180 1636 3188 1644
rect 3212 1636 3220 1644
rect 3244 1636 3252 1644
rect 3292 1636 3300 1644
rect 3644 1636 3652 1644
rect 3772 1636 3780 1644
rect 4604 1636 4612 1644
rect 4780 1636 4788 1644
rect 4844 1636 4852 1644
rect 1043 1606 1051 1614
rect 1053 1606 1061 1614
rect 1063 1606 1071 1614
rect 1073 1606 1081 1614
rect 1083 1606 1091 1614
rect 1093 1606 1101 1614
rect 4051 1606 4059 1614
rect 4061 1606 4069 1614
rect 4071 1606 4079 1614
rect 4081 1606 4089 1614
rect 4091 1606 4099 1614
rect 4101 1606 4109 1614
rect 172 1576 180 1584
rect 588 1576 596 1584
rect 1532 1576 1540 1584
rect 1628 1576 1636 1584
rect 1980 1576 1988 1584
rect 2236 1576 2244 1584
rect 2540 1576 2548 1584
rect 2796 1576 2804 1584
rect 4940 1576 4948 1584
rect 1356 1556 1364 1564
rect 1852 1556 1860 1564
rect 2940 1556 2948 1564
rect 3276 1556 3284 1564
rect 4092 1556 4100 1564
rect 2012 1536 2020 1544
rect 2332 1536 2340 1544
rect 2588 1536 2596 1544
rect 2700 1536 2708 1544
rect 3100 1536 3108 1544
rect 3436 1536 3444 1544
rect 3660 1536 3668 1544
rect 3772 1536 3780 1544
rect 4124 1536 4132 1544
rect 4972 1536 4980 1544
rect 204 1516 212 1524
rect 876 1516 884 1524
rect 44 1496 52 1504
rect 60 1496 68 1504
rect 108 1496 116 1504
rect 172 1496 180 1504
rect 316 1496 324 1504
rect 476 1496 484 1504
rect 700 1496 708 1504
rect 828 1496 836 1504
rect 908 1496 916 1504
rect 924 1496 932 1504
rect 972 1496 980 1504
rect 988 1496 996 1504
rect 1020 1516 1028 1524
rect 1308 1516 1316 1524
rect 1052 1496 1060 1504
rect 1164 1496 1172 1504
rect 1212 1496 1220 1504
rect 1228 1496 1236 1504
rect 1276 1496 1284 1504
rect 1324 1496 1332 1504
rect 1340 1496 1348 1504
rect 1404 1516 1412 1524
rect 1500 1516 1508 1524
rect 1740 1516 1748 1524
rect 1884 1516 1892 1524
rect 1948 1516 1956 1524
rect 2764 1516 2772 1524
rect 1436 1496 1444 1504
rect 1532 1496 1540 1504
rect 1564 1496 1572 1504
rect 1628 1496 1636 1504
rect 1644 1496 1652 1504
rect 1708 1496 1716 1504
rect 1756 1496 1764 1504
rect 1804 1496 1812 1504
rect 1884 1496 1892 1504
rect 1900 1496 1908 1504
rect 1916 1496 1924 1504
rect 1980 1496 1988 1504
rect 2124 1496 2132 1504
rect 2204 1496 2212 1504
rect 2284 1496 2292 1504
rect 2300 1496 2308 1504
rect 2428 1496 2436 1504
rect 2460 1496 2468 1504
rect 2652 1496 2660 1504
rect 2668 1496 2676 1504
rect 2700 1496 2708 1504
rect 2748 1496 2756 1504
rect 2796 1496 2804 1504
rect 2828 1496 2836 1504
rect 2876 1496 2884 1504
rect 2972 1496 2980 1504
rect 3068 1516 3076 1524
rect 12 1476 20 1484
rect 92 1476 100 1484
rect 284 1476 292 1484
rect 380 1476 388 1484
rect 524 1476 532 1484
rect 620 1476 628 1484
rect 844 1476 852 1484
rect 940 1476 948 1484
rect 1068 1476 1076 1484
rect 1340 1476 1348 1484
rect 3052 1496 3060 1504
rect 3100 1496 3108 1504
rect 3148 1496 3156 1504
rect 3180 1496 3188 1504
rect 3212 1496 3220 1504
rect 3308 1496 3316 1504
rect 3468 1516 3476 1524
rect 3372 1496 3380 1504
rect 3436 1496 3444 1504
rect 3452 1496 3460 1504
rect 3500 1496 3508 1504
rect 3644 1516 3652 1524
rect 3692 1516 3700 1524
rect 3564 1496 3572 1504
rect 3612 1496 3620 1504
rect 3628 1496 3636 1504
rect 3964 1516 3972 1524
rect 4508 1516 4516 1524
rect 3724 1496 3732 1504
rect 3756 1496 3764 1504
rect 3836 1496 3844 1504
rect 3884 1496 3892 1504
rect 3980 1496 3988 1504
rect 4028 1496 4036 1504
rect 4204 1496 4212 1504
rect 4780 1516 4788 1524
rect 4412 1494 4420 1502
rect 4556 1496 4564 1504
rect 4716 1494 4724 1502
rect 4780 1496 4788 1504
rect 4812 1496 4820 1504
rect 4892 1496 4900 1504
rect 4924 1496 4932 1504
rect 5068 1494 5076 1502
rect 1452 1476 1460 1484
rect 1580 1476 1588 1484
rect 1692 1476 1700 1484
rect 1820 1476 1828 1484
rect 1932 1476 1940 1484
rect 1996 1476 2004 1484
rect 2172 1476 2180 1484
rect 2652 1476 2660 1484
rect 2716 1476 2724 1484
rect 2812 1476 2820 1484
rect 2876 1476 2884 1484
rect 2924 1476 2932 1484
rect 2988 1476 2996 1484
rect 3004 1476 3012 1484
rect 3052 1476 3060 1484
rect 3116 1476 3124 1484
rect 3132 1476 3140 1484
rect 3196 1476 3204 1484
rect 3260 1476 3268 1484
rect 3324 1476 3332 1484
rect 3340 1476 3348 1484
rect 3388 1476 3396 1484
rect 3452 1476 3460 1484
rect 3516 1476 3524 1484
rect 3580 1476 3588 1484
rect 3596 1476 3604 1484
rect 3660 1476 3668 1484
rect 3756 1476 3764 1484
rect 4012 1476 4020 1484
rect 4252 1476 4260 1484
rect 4444 1476 4452 1484
rect 4476 1476 4484 1484
rect 4508 1476 4516 1484
rect 4572 1476 4580 1484
rect 4700 1476 4708 1484
rect 4876 1476 4884 1484
rect 5052 1476 5060 1484
rect 1244 1456 1252 1464
rect 1292 1456 1300 1464
rect 1596 1456 1604 1464
rect 1628 1456 1636 1464
rect 1676 1456 1684 1464
rect 1836 1456 1844 1464
rect 2252 1456 2260 1464
rect 2908 1456 2916 1464
rect 3244 1456 3252 1464
rect 3404 1456 3412 1464
rect 3900 1456 3908 1464
rect 4860 1456 4868 1464
rect 140 1436 148 1444
rect 780 1436 788 1444
rect 796 1436 804 1444
rect 1196 1436 1204 1444
rect 1260 1436 1268 1444
rect 1804 1436 1812 1444
rect 2268 1436 2276 1444
rect 2524 1436 2532 1444
rect 3180 1436 3188 1444
rect 3532 1436 3540 1444
rect 4284 1436 4292 1444
rect 4588 1436 4596 1444
rect 2547 1406 2555 1414
rect 2557 1406 2565 1414
rect 2567 1406 2575 1414
rect 2577 1406 2585 1414
rect 2587 1406 2595 1414
rect 2597 1406 2605 1414
rect 108 1376 116 1384
rect 700 1376 708 1384
rect 1356 1376 1364 1384
rect 1724 1376 1732 1384
rect 1948 1376 1956 1384
rect 2412 1376 2420 1384
rect 3260 1376 3268 1384
rect 3772 1376 3780 1384
rect 4124 1376 4132 1384
rect 4732 1376 4740 1384
rect 5068 1376 5076 1384
rect 620 1356 628 1364
rect 796 1356 804 1364
rect 828 1356 836 1364
rect 1436 1356 1444 1364
rect 1660 1356 1668 1364
rect 1740 1356 1748 1364
rect 1788 1356 1796 1364
rect 1804 1356 1812 1364
rect 2316 1356 2324 1364
rect 2700 1356 2708 1364
rect 2876 1356 2884 1364
rect 2924 1356 2932 1364
rect 3052 1356 3060 1364
rect 3132 1356 3140 1364
rect 3484 1356 3492 1364
rect 3500 1356 3508 1364
rect 4252 1356 4260 1364
rect 4924 1356 4932 1364
rect 12 1336 20 1344
rect 60 1336 68 1344
rect 188 1336 196 1344
rect 268 1336 276 1344
rect 348 1336 356 1344
rect 524 1336 532 1344
rect 668 1336 676 1344
rect 684 1336 692 1344
rect 780 1336 788 1344
rect 892 1336 900 1344
rect 956 1336 964 1344
rect 972 1336 980 1344
rect 1180 1336 1188 1344
rect 1324 1336 1332 1344
rect 1340 1336 1348 1344
rect 1404 1336 1412 1344
rect 1420 1336 1428 1344
rect 1484 1336 1492 1344
rect 1500 1336 1508 1344
rect 1612 1336 1620 1344
rect 1740 1336 1748 1344
rect 1996 1336 2004 1344
rect 2060 1336 2068 1344
rect 2172 1336 2180 1344
rect 2476 1336 2484 1344
rect 2588 1336 2596 1344
rect 2652 1336 2660 1344
rect 2716 1336 2724 1344
rect 2828 1336 2836 1344
rect 2940 1336 2948 1344
rect 3004 1336 3012 1344
rect 3052 1336 3060 1344
rect 3116 1336 3124 1344
rect 3180 1336 3188 1344
rect 3244 1336 3252 1344
rect 3308 1336 3316 1344
rect 3356 1336 3364 1344
rect 3372 1336 3380 1344
rect 3436 1336 3444 1344
rect 3548 1336 3556 1344
rect 3612 1336 3620 1344
rect 3916 1336 3924 1344
rect 4044 1336 4052 1344
rect 4348 1336 4356 1344
rect 4428 1336 4436 1344
rect 4492 1336 4500 1344
rect 4524 1336 4532 1344
rect 4700 1336 4708 1344
rect 4892 1336 4900 1344
rect 4988 1336 4996 1344
rect 5020 1336 5028 1344
rect 44 1316 52 1324
rect 92 1316 100 1324
rect 236 1318 244 1326
rect 332 1316 340 1324
rect 412 1316 420 1324
rect 556 1318 564 1326
rect 652 1316 660 1324
rect 668 1316 676 1324
rect 716 1316 724 1324
rect 796 1316 804 1324
rect 828 1316 836 1324
rect 876 1316 884 1324
rect 940 1316 948 1324
rect 988 1316 996 1324
rect 1004 1316 1012 1324
rect 1100 1316 1108 1324
rect 1116 1316 1124 1324
rect 1148 1316 1156 1324
rect 1164 1316 1172 1324
rect 1212 1316 1220 1324
rect 1276 1316 1284 1324
rect 1308 1316 1316 1324
rect 1356 1316 1364 1324
rect 1388 1316 1396 1324
rect 1436 1316 1444 1324
rect 1500 1316 1508 1324
rect 1516 1316 1524 1324
rect 1596 1316 1604 1324
rect 1612 1316 1620 1324
rect 1692 1316 1700 1324
rect 1708 1316 1716 1324
rect 1756 1316 1764 1324
rect 1836 1316 1844 1324
rect 1884 1316 1892 1324
rect 1932 1316 1940 1324
rect 1996 1316 2004 1324
rect 2012 1316 2020 1324
rect 2076 1316 2084 1324
rect 300 1296 308 1304
rect 412 1296 420 1304
rect 620 1296 628 1304
rect 732 1296 740 1304
rect 844 1296 852 1304
rect 908 1296 916 1304
rect 1020 1296 1028 1304
rect 1276 1296 1284 1304
rect 1548 1296 1556 1304
rect 1676 1296 1684 1304
rect 2156 1316 2164 1324
rect 2284 1316 2292 1324
rect 2380 1316 2388 1324
rect 2460 1316 2468 1324
rect 2492 1316 2500 1324
rect 2524 1296 2532 1304
rect 2636 1316 2644 1324
rect 2668 1316 2676 1324
rect 2796 1316 2804 1324
rect 2844 1316 2852 1324
rect 2892 1316 2900 1324
rect 2956 1316 2964 1324
rect 2972 1316 2980 1324
rect 3004 1316 3012 1324
rect 3020 1316 3028 1324
rect 3100 1316 3108 1324
rect 3164 1316 3172 1324
rect 3196 1316 3204 1324
rect 3228 1316 3236 1324
rect 3292 1316 3300 1324
rect 3324 1316 3332 1324
rect 3388 1316 3396 1324
rect 3436 1316 3444 1324
rect 3452 1316 3460 1324
rect 3564 1316 3572 1324
rect 3580 1316 3588 1324
rect 3596 1316 3604 1324
rect 3628 1316 3636 1324
rect 3644 1316 3652 1324
rect 3708 1316 3716 1324
rect 3724 1316 3732 1324
rect 3740 1316 3748 1324
rect 3788 1316 3796 1324
rect 3852 1316 3860 1324
rect 3916 1316 3924 1324
rect 2908 1296 2916 1304
rect 3068 1296 3076 1304
rect 3260 1296 3268 1304
rect 3500 1296 3508 1304
rect 4012 1316 4020 1324
rect 4028 1316 4036 1324
rect 4252 1318 4260 1326
rect 4348 1316 4356 1324
rect 4396 1316 4404 1324
rect 4444 1316 4452 1324
rect 4316 1296 4324 1304
rect 4636 1316 4644 1324
rect 4860 1318 4868 1326
rect 4956 1316 4964 1324
rect 5036 1316 5044 1324
rect 5100 1316 5108 1324
rect 4492 1296 4500 1304
rect 5004 1296 5012 1304
rect 5068 1296 5076 1304
rect 5084 1296 5092 1304
rect 332 1276 340 1284
rect 940 1276 948 1284
rect 1212 1276 1220 1284
rect 1516 1276 1524 1284
rect 2044 1276 2052 1284
rect 2108 1276 2116 1284
rect 2732 1276 2740 1284
rect 3020 1276 3028 1284
rect 3164 1276 3172 1284
rect 3452 1276 3460 1284
rect 3564 1276 3572 1284
rect 3868 1276 3876 1284
rect 3980 1276 3988 1284
rect 4524 1276 4532 1284
rect 5116 1276 5124 1284
rect 2156 1256 2164 1264
rect 5100 1256 5108 1264
rect 812 1236 820 1244
rect 1564 1236 1572 1244
rect 1852 1236 1860 1244
rect 1900 1236 1908 1244
rect 1948 1236 1956 1244
rect 2012 1236 2020 1244
rect 2188 1236 2196 1244
rect 2412 1236 2420 1244
rect 2428 1236 2436 1244
rect 2844 1236 2852 1244
rect 3196 1236 3204 1244
rect 3404 1236 3412 1244
rect 3660 1236 3668 1244
rect 3820 1236 3828 1244
rect 3900 1236 3908 1244
rect 4124 1236 4132 1244
rect 1043 1206 1051 1214
rect 1053 1206 1061 1214
rect 1063 1206 1071 1214
rect 1073 1206 1081 1214
rect 1083 1206 1091 1214
rect 1093 1206 1101 1214
rect 4051 1206 4059 1214
rect 4061 1206 4069 1214
rect 4071 1206 4079 1214
rect 4081 1206 4089 1214
rect 4091 1206 4099 1214
rect 4101 1206 4109 1214
rect 332 1176 340 1184
rect 1276 1176 1284 1184
rect 1340 1176 1348 1184
rect 2780 1176 2788 1184
rect 3324 1176 3332 1184
rect 3340 1176 3348 1184
rect 3788 1176 3796 1184
rect 4044 1176 4052 1184
rect 4652 1176 4660 1184
rect 5020 1176 5028 1184
rect 5084 1176 5092 1184
rect 3004 1156 3012 1164
rect 268 1136 276 1144
rect 364 1136 372 1144
rect 796 1136 804 1144
rect 1932 1136 1940 1144
rect 2940 1136 2948 1144
rect 3244 1136 3252 1144
rect 4716 1136 4724 1144
rect 5036 1136 5044 1144
rect 5100 1136 5108 1144
rect 300 1116 308 1124
rect 556 1116 564 1124
rect 844 1116 852 1124
rect 44 1096 52 1104
rect 172 1096 180 1104
rect 268 1096 276 1104
rect 316 1096 324 1104
rect 492 1094 500 1102
rect 588 1096 596 1104
rect 716 1096 724 1104
rect 1164 1116 1172 1124
rect 1372 1116 1380 1124
rect 1612 1116 1620 1124
rect 892 1096 900 1104
rect 940 1096 948 1104
rect 956 1096 964 1104
rect 988 1096 996 1104
rect 1004 1096 1012 1104
rect 1100 1096 1108 1104
rect 1148 1096 1156 1104
rect 1196 1096 1204 1104
rect 1228 1096 1236 1104
rect 1244 1096 1252 1104
rect 1292 1096 1300 1104
rect 1340 1096 1348 1104
rect 1452 1096 1460 1104
rect 2124 1116 2132 1124
rect 2476 1116 2484 1124
rect 3116 1116 3124 1124
rect 3228 1116 3236 1124
rect 3548 1116 3556 1124
rect 3580 1116 3588 1124
rect 3980 1116 3988 1124
rect 4332 1116 4340 1124
rect 4572 1116 4580 1124
rect 1516 1094 1524 1102
rect 1660 1096 1668 1104
rect 1692 1096 1700 1104
rect 1740 1096 1748 1104
rect 1788 1096 1796 1104
rect 1868 1096 1876 1104
rect 1916 1096 1924 1104
rect 2060 1094 2068 1102
rect 2124 1096 2132 1104
rect 2172 1096 2180 1104
rect 2220 1096 2228 1104
rect 2284 1096 2292 1104
rect 2316 1096 2324 1104
rect 2332 1096 2340 1104
rect 2364 1096 2372 1104
rect 2412 1096 2420 1104
rect 2428 1096 2436 1104
rect 2460 1096 2468 1104
rect 2604 1094 2612 1102
rect 2748 1096 2756 1104
rect 2812 1096 2820 1104
rect 2860 1096 2868 1104
rect 2876 1096 2884 1104
rect 2892 1096 2900 1104
rect 2908 1096 2916 1104
rect 2956 1096 2964 1104
rect 3004 1096 3012 1104
rect 3036 1096 3044 1104
rect 3068 1096 3076 1104
rect 3132 1096 3140 1104
rect 3196 1096 3204 1104
rect 3276 1096 3284 1104
rect 3292 1096 3300 1104
rect 3468 1094 3476 1102
rect 3548 1096 3556 1104
rect 3596 1096 3604 1104
rect 3612 1096 3620 1104
rect 3660 1096 3668 1104
rect 3692 1096 3700 1104
rect 3708 1096 3716 1104
rect 3756 1096 3764 1104
rect 3900 1096 3908 1104
rect 4012 1096 4020 1104
rect 4220 1096 4228 1104
rect 4956 1116 4964 1124
rect 4988 1116 4996 1124
rect 5004 1116 5012 1124
rect 5068 1116 5076 1124
rect 4476 1094 4484 1102
rect 4620 1096 4628 1104
rect 4844 1094 4852 1102
rect 4940 1096 4948 1104
rect 5020 1096 5028 1104
rect 5084 1096 5092 1104
rect 12 1076 20 1084
rect 188 1076 196 1084
rect 252 1076 260 1084
rect 524 1076 532 1084
rect 556 1076 564 1084
rect 604 1076 612 1084
rect 684 1076 692 1084
rect 860 1076 868 1084
rect 908 1076 916 1084
rect 1084 1076 1092 1084
rect 1212 1076 1220 1084
rect 1324 1076 1332 1084
rect 1580 1076 1588 1084
rect 1612 1076 1620 1084
rect 1692 1076 1700 1084
rect 348 1056 356 1064
rect 1100 1056 1108 1064
rect 1724 1056 1732 1064
rect 1772 1056 1780 1064
rect 1788 1056 1796 1064
rect 1836 1076 1844 1084
rect 2028 1076 2036 1084
rect 2172 1076 2180 1084
rect 2428 1076 2436 1084
rect 2620 1076 2628 1084
rect 2972 1076 2980 1084
rect 3052 1076 3060 1084
rect 3068 1076 3076 1084
rect 3100 1076 3108 1084
rect 3180 1076 3188 1084
rect 3212 1076 3220 1084
rect 3468 1076 3476 1084
rect 3532 1076 3540 1084
rect 3916 1076 3924 1084
rect 3980 1076 3988 1084
rect 4076 1076 4084 1084
rect 4300 1076 4308 1084
rect 4540 1076 4548 1084
rect 4572 1076 4580 1084
rect 4636 1076 4644 1084
rect 4668 1076 4676 1084
rect 4700 1076 4708 1084
rect 1836 1056 1844 1064
rect 1884 1056 1892 1064
rect 2188 1056 2196 1064
rect 2236 1056 2244 1064
rect 2284 1056 2292 1064
rect 2316 1056 2324 1064
rect 2332 1056 2340 1064
rect 2364 1056 2372 1064
rect 2700 1056 2708 1064
rect 3132 1056 3140 1064
rect 3164 1056 3172 1064
rect 3724 1056 3732 1064
rect 4236 1056 4244 1064
rect 4476 1056 4484 1064
rect 4844 1056 4852 1064
rect 4908 1056 4916 1064
rect 60 1036 68 1044
rect 332 1036 340 1044
rect 1388 1036 1396 1044
rect 1708 1036 1716 1044
rect 1756 1036 1764 1044
rect 1852 1036 1860 1044
rect 1900 1036 1908 1044
rect 2204 1036 2212 1044
rect 2252 1036 2260 1044
rect 2732 1036 2740 1044
rect 2828 1036 2836 1044
rect 3628 1036 3636 1044
rect 4332 1036 4340 1044
rect 4348 1036 4356 1044
rect 4684 1036 4692 1044
rect 2547 1006 2555 1014
rect 2557 1006 2565 1014
rect 2567 1006 2575 1014
rect 2577 1006 2585 1014
rect 2587 1006 2595 1014
rect 2597 1006 2605 1014
rect 172 976 180 984
rect 988 976 996 984
rect 1196 976 1204 984
rect 1532 976 1540 984
rect 2412 976 2420 984
rect 2636 976 2644 984
rect 2716 976 2724 984
rect 3452 976 3460 984
rect 4140 976 4148 984
rect 4396 976 4404 984
rect 4684 976 4692 984
rect 556 956 564 964
rect 604 956 612 964
rect 652 956 660 964
rect 700 956 708 964
rect 1324 956 1332 964
rect 1388 956 1396 964
rect 1660 956 1668 964
rect 2092 956 2100 964
rect 2252 956 2260 964
rect 3180 956 3188 964
rect 3356 956 3364 964
rect 3548 956 3556 964
rect 4588 956 4596 964
rect 4876 956 4884 964
rect 4940 956 4948 964
rect 60 936 68 944
rect 156 936 164 944
rect 220 936 228 944
rect 236 936 244 944
rect 492 936 500 944
rect 636 936 644 944
rect 732 936 740 944
rect 796 936 804 944
rect 876 936 884 944
rect 1004 936 1012 944
rect 1036 936 1044 944
rect 1180 936 1188 944
rect 1244 936 1252 944
rect 1324 936 1332 944
rect 1372 936 1380 944
rect 1500 936 1508 944
rect 1516 936 1524 944
rect 1644 936 1652 944
rect 1756 936 1764 944
rect 1772 936 1780 944
rect 1836 936 1844 944
rect 1852 936 1860 944
rect 1980 936 1988 944
rect 2044 936 2052 944
rect 2300 936 2308 944
rect 2396 936 2404 944
rect 2540 936 2548 944
rect 2604 936 2612 944
rect 2668 936 2676 944
rect 2700 936 2708 944
rect 2812 936 2820 944
rect 2844 936 2852 944
rect 2876 936 2884 944
rect 3004 936 3012 944
rect 3132 936 3140 944
rect 3196 936 3204 944
rect 3260 936 3268 944
rect 3308 936 3316 944
rect 3564 936 3572 944
rect 3628 936 3636 944
rect 3644 936 3652 944
rect 3692 936 3700 944
rect 3756 936 3764 944
rect 3868 936 3876 944
rect 4044 936 4052 944
rect 4236 936 4244 944
rect 4300 936 4308 944
rect 4380 936 4388 944
rect 4476 936 4484 944
rect 4556 936 4564 944
rect 4652 936 4660 944
rect 4844 936 4852 944
rect 44 916 52 924
rect 92 916 100 924
rect 140 916 148 924
rect 220 916 228 924
rect 252 916 260 924
rect 284 916 292 924
rect 364 916 372 924
rect 428 918 436 926
rect 524 916 532 924
rect 588 916 596 924
rect 636 916 644 924
rect 684 916 692 924
rect 732 916 740 924
rect 780 916 788 924
rect 892 916 900 924
rect 1020 916 1028 924
rect 108 896 116 904
rect 172 896 180 904
rect 284 896 292 904
rect 492 896 500 904
rect 748 896 756 904
rect 1164 916 1172 924
rect 1292 916 1300 924
rect 1356 916 1364 924
rect 1388 916 1396 924
rect 1420 916 1428 924
rect 1484 916 1492 924
rect 1532 916 1540 924
rect 1580 916 1588 924
rect 1628 916 1636 924
rect 1708 916 1716 924
rect 1740 916 1748 924
rect 1788 916 1796 924
rect 1820 916 1828 924
rect 1868 916 1876 924
rect 1900 916 1908 924
rect 1964 916 1972 924
rect 2028 916 2036 924
rect 2060 916 2068 924
rect 2076 916 2084 924
rect 2156 916 2164 924
rect 2220 916 2228 924
rect 2236 916 2244 924
rect 2284 916 2292 924
rect 1116 896 1124 904
rect 1196 896 1204 904
rect 1260 896 1268 904
rect 1452 896 1460 904
rect 1596 896 1604 904
rect 1708 896 1716 904
rect 1788 896 1796 904
rect 1868 896 1876 904
rect 1932 896 1940 904
rect 1996 896 2004 904
rect 2188 896 2196 904
rect 2332 896 2340 904
rect 2380 916 2388 924
rect 2524 916 2532 924
rect 2748 916 2756 924
rect 2796 916 2804 924
rect 2828 916 2836 924
rect 2860 916 2868 924
rect 2876 916 2884 924
rect 2956 916 2964 924
rect 3020 916 3028 924
rect 3084 916 3092 924
rect 3116 916 3124 924
rect 3148 916 3156 924
rect 3228 916 3236 924
rect 3244 916 3252 924
rect 3276 916 3284 924
rect 3324 916 3332 924
rect 3340 916 3348 924
rect 3436 916 3444 924
rect 3484 916 3492 924
rect 3500 916 3508 924
rect 3516 916 3524 924
rect 3612 916 3620 924
rect 2380 896 2388 904
rect 2668 896 2676 904
rect 2956 896 2964 904
rect 2988 896 2996 904
rect 3084 896 3092 904
rect 3676 916 3684 924
rect 3740 916 3748 924
rect 3772 916 3780 924
rect 3804 896 3812 904
rect 3836 916 3844 924
rect 3852 916 3860 924
rect 3964 916 3972 924
rect 4268 918 4276 926
rect 4348 916 4356 924
rect 4380 916 4388 924
rect 4524 918 4532 926
rect 4636 916 4644 924
rect 4748 916 4756 924
rect 4812 918 4820 926
rect 4924 916 4932 924
rect 4988 916 4996 924
rect 5068 916 5076 924
rect 4332 896 4340 904
rect 4668 896 4676 904
rect 4876 896 4884 904
rect 4972 896 4980 904
rect 5148 896 5156 904
rect 12 876 20 884
rect 140 876 148 884
rect 5004 876 5012 884
rect 5052 876 5060 884
rect 2268 856 2276 864
rect 2924 856 2932 864
rect 4988 856 4996 864
rect 620 836 628 844
rect 716 836 724 844
rect 1340 836 1348 844
rect 1676 836 1684 844
rect 1740 836 1748 844
rect 2028 836 2036 844
rect 2716 836 2724 844
rect 2764 836 2772 844
rect 3020 836 3028 844
rect 3580 836 3588 844
rect 3708 836 3716 844
rect 3884 836 3892 844
rect 5036 836 5044 844
rect 1043 806 1051 814
rect 1053 806 1061 814
rect 1063 806 1071 814
rect 1073 806 1081 814
rect 1083 806 1091 814
rect 1093 806 1101 814
rect 4051 806 4059 814
rect 4061 806 4069 814
rect 4071 806 4079 814
rect 4081 806 4089 814
rect 4091 806 4099 814
rect 4101 806 4109 814
rect 748 776 756 784
rect 812 776 820 784
rect 1004 776 1012 784
rect 1292 776 1300 784
rect 1388 776 1396 784
rect 4876 776 4884 784
rect 5020 776 5028 784
rect 1740 756 1748 764
rect 2364 756 2372 764
rect 3180 756 3188 764
rect 12 736 20 744
rect 156 736 164 744
rect 428 736 436 744
rect 1580 736 1588 744
rect 3356 736 3364 744
rect 3596 736 3604 744
rect 3948 736 3956 744
rect 4556 736 4564 744
rect 4860 736 4868 744
rect 396 716 404 724
rect 508 716 516 724
rect 716 716 724 724
rect 44 696 52 704
rect 60 696 68 704
rect 108 696 116 704
rect 284 694 292 702
rect 348 696 356 704
rect 428 696 436 704
rect 460 696 468 704
rect 524 696 532 704
rect 572 696 580 704
rect 748 696 756 704
rect 764 696 772 704
rect 924 696 932 704
rect 1036 696 1044 704
rect 1052 696 1060 704
rect 1132 716 1140 724
rect 1468 716 1476 724
rect 1196 696 1204 704
rect 1244 696 1252 704
rect 1260 696 1268 704
rect 1308 696 1316 704
rect 1340 696 1348 704
rect 1356 696 1364 704
rect 1404 696 1412 704
rect 1596 716 1604 724
rect 1660 716 1668 724
rect 1772 716 1780 724
rect 2044 716 2052 724
rect 2236 716 2244 724
rect 2476 716 2484 724
rect 2492 716 2500 724
rect 2668 716 2676 724
rect 2748 716 2756 724
rect 1516 696 1524 704
rect 1548 696 1556 704
rect 1628 696 1636 704
rect 1692 696 1700 704
rect 1740 696 1748 704
rect 1788 696 1796 704
rect 1820 696 1828 704
rect 1980 694 1988 702
rect 2060 696 2068 704
rect 2076 696 2084 704
rect 2108 696 2116 704
rect 2156 696 2164 704
rect 2172 696 2180 704
rect 2236 696 2244 704
rect 2268 696 2276 704
rect 2284 696 2292 704
rect 2332 696 2340 704
rect 2364 696 2372 704
rect 2396 696 2404 704
rect 2444 696 2452 704
rect 2572 696 2580 704
rect 2620 696 2628 704
rect 2700 696 2708 704
rect 2748 696 2756 704
rect 2844 696 2852 704
rect 2908 694 2916 702
rect 3068 696 3076 704
rect 3116 696 3124 704
rect 3132 696 3140 704
rect 3148 696 3156 704
rect 3212 696 3220 704
rect 3228 696 3236 704
rect 3260 696 3268 704
rect 3308 716 3316 724
rect 3628 716 3636 724
rect 3836 716 3844 724
rect 4236 716 4244 724
rect 3436 696 3444 704
rect 3548 696 3556 704
rect 3772 694 3780 702
rect 3852 696 3860 704
rect 3884 696 3892 704
rect 3932 696 3940 704
rect 4540 716 4548 724
rect 4796 716 4804 724
rect 4828 716 4836 724
rect 4892 716 4900 724
rect 4988 716 4996 724
rect 4076 694 4084 702
rect 4284 696 4292 704
rect 4508 696 4516 704
rect 4620 696 4628 704
rect 4684 694 4692 702
rect 4780 696 4788 704
rect 4876 696 4884 704
rect 4956 696 4964 704
rect 268 676 276 684
rect 444 676 452 684
rect 556 676 564 684
rect 572 676 580 684
rect 764 676 772 684
rect 844 676 852 684
rect 876 676 884 684
rect 1020 676 1028 684
rect 1180 676 1188 684
rect 1420 676 1428 684
rect 1532 676 1540 684
rect 1644 676 1652 684
rect 1660 676 1668 684
rect 1708 676 1716 684
rect 1724 676 1732 684
rect 1836 676 1844 684
rect 2012 676 2020 684
rect 2092 676 2100 684
rect 2300 676 2308 684
rect 2348 676 2356 684
rect 2412 676 2420 684
rect 2428 676 2436 684
rect 2492 676 2500 684
rect 2556 676 2564 684
rect 2588 676 2596 684
rect 2716 676 2724 684
rect 2732 676 2740 684
rect 2796 676 2804 684
rect 2940 676 2948 684
rect 3052 676 3060 684
rect 3244 676 3252 684
rect 3468 676 3476 684
rect 3596 676 3604 684
rect 3628 676 3636 684
rect 3884 676 3892 684
rect 3900 676 3908 684
rect 4108 676 4116 684
rect 4140 676 4148 684
rect 4252 676 4260 684
rect 4300 676 4308 684
rect 4444 676 4452 684
rect 5132 676 5140 684
rect 380 656 388 664
rect 2172 656 2180 664
rect 2300 656 2308 664
rect 2652 656 2660 664
rect 2812 656 2820 664
rect 3292 656 3300 664
rect 3772 656 3780 664
rect 4460 656 4468 664
rect 4748 656 4756 664
rect 4908 656 4916 664
rect 92 636 100 644
rect 140 636 148 644
rect 492 636 500 644
rect 684 636 692 644
rect 1228 636 1236 644
rect 1484 636 1492 644
rect 1596 636 1604 644
rect 1852 636 1860 644
rect 2476 636 2484 644
rect 2668 636 2676 644
rect 3036 636 3044 644
rect 3580 636 3588 644
rect 3644 636 3652 644
rect 4332 636 4340 644
rect 4540 636 4548 644
rect 4988 636 4996 644
rect 2547 606 2555 614
rect 2557 606 2565 614
rect 2567 606 2575 614
rect 2577 606 2585 614
rect 2587 606 2595 614
rect 2597 606 2605 614
rect 892 576 900 584
rect 1276 576 1284 584
rect 1356 576 1364 584
rect 2476 576 2484 584
rect 2508 576 2516 584
rect 2636 576 2644 584
rect 2796 576 2804 584
rect 3068 576 3076 584
rect 3372 576 3380 584
rect 4092 576 4100 584
rect 4444 576 4452 584
rect 4636 576 4644 584
rect 4828 576 4836 584
rect 4924 576 4932 584
rect 524 556 532 564
rect 716 556 724 564
rect 844 556 852 564
rect 2124 556 2132 564
rect 2268 556 2276 564
rect 2396 556 2404 564
rect 2892 556 2900 564
rect 3084 556 3092 564
rect 3244 556 3252 564
rect 3260 556 3268 564
rect 3324 556 3332 564
rect 4332 556 4340 564
rect 4732 556 4740 564
rect 60 536 68 544
rect 364 536 372 544
rect 444 536 452 544
rect 508 536 516 544
rect 572 536 580 544
rect 588 536 596 544
rect 636 536 644 544
rect 812 536 820 544
rect 940 536 948 544
rect 1004 536 1012 544
rect 1340 536 1348 544
rect 1436 536 1444 544
rect 1452 536 1460 544
rect 1596 536 1604 544
rect 1612 536 1620 544
rect 1660 536 1668 544
rect 1724 536 1732 544
rect 1788 536 1796 544
rect 1852 536 1860 544
rect 1868 536 1876 544
rect 1916 536 1924 544
rect 1980 536 1988 544
rect 2044 536 2052 544
rect 2108 536 2116 544
rect 2172 536 2180 544
rect 2188 536 2196 544
rect 2236 536 2244 544
rect 2252 536 2260 544
rect 2380 536 2388 544
rect 2540 536 2548 544
rect 2604 536 2612 544
rect 2652 536 2660 544
rect 2780 536 2788 544
rect 2860 536 2868 544
rect 2908 536 2916 544
rect 3052 536 3060 544
rect 3100 536 3108 544
rect 3244 536 3252 544
rect 3420 536 3428 544
rect 3596 536 3604 544
rect 3772 536 3780 544
rect 3820 536 3828 544
rect 3852 536 3860 544
rect 3900 536 3908 544
rect 3916 536 3924 544
rect 3964 536 3972 544
rect 4252 536 4260 544
rect 4284 536 4292 544
rect 4380 536 4388 544
rect 4428 536 4436 544
rect 4604 536 4612 544
rect 4652 536 4660 544
rect 44 516 52 524
rect 268 516 276 524
rect 332 518 340 526
rect 428 516 436 524
rect 460 516 468 524
rect 508 516 516 524
rect 556 516 564 524
rect 620 516 628 524
rect 780 518 788 526
rect 876 516 884 524
rect 940 516 948 524
rect 972 516 980 524
rect 988 516 996 524
rect 1052 516 1060 524
rect 1068 516 1076 524
rect 1164 516 1172 524
rect 1228 516 1236 524
rect 1244 516 1252 524
rect 1340 516 1348 524
rect 1420 516 1428 524
rect 1484 518 1492 526
rect 1596 516 1604 524
rect 1708 516 1716 524
rect 1724 516 1732 524
rect 1852 516 1860 524
rect 1868 516 1876 524
rect 1948 516 1956 524
rect 1964 516 1972 524
rect 2028 516 2036 524
rect 2044 516 2052 524
rect 2108 516 2116 524
rect 2156 516 2164 524
rect 2220 516 2228 524
rect 2268 516 2276 524
rect 2332 516 2340 524
rect 2364 516 2372 524
rect 2396 516 2404 524
rect 2428 516 2436 524
rect 2444 516 2452 524
rect 2668 516 2676 524
rect 2700 516 2708 524
rect 2764 516 2772 524
rect 2828 516 2836 524
rect 2860 516 2868 524
rect 2924 516 2932 524
rect 2956 516 2964 524
rect 3020 516 3028 524
rect 3036 516 3044 524
rect 3116 516 3124 524
rect 3180 516 3188 524
rect 3212 516 3220 524
rect 3276 516 3284 524
rect 3340 516 3348 524
rect 3356 516 3364 524
rect 3452 516 3460 524
rect 3500 516 3508 524
rect 3516 516 3524 524
rect 3612 516 3620 524
rect 3788 518 3796 526
rect 3884 516 3892 524
rect 3948 516 3956 524
rect 4220 518 4228 526
rect 428 496 436 504
rect 460 496 468 504
rect 524 496 532 504
rect 588 496 596 504
rect 892 496 900 504
rect 956 496 964 504
rect 1132 496 1140 504
rect 1292 496 1300 504
rect 1548 496 1556 504
rect 1612 496 1620 504
rect 1676 496 1684 504
rect 1740 496 1748 504
rect 1804 496 1812 504
rect 1932 496 1940 504
rect 1996 496 2004 504
rect 2060 496 2068 504
rect 2124 496 2132 504
rect 2188 496 2196 504
rect 2332 496 2340 504
rect 2492 496 2500 504
rect 2636 496 2644 504
rect 2684 496 2692 504
rect 2732 496 2740 504
rect 2796 496 2804 504
rect 2988 496 2996 504
rect 3148 496 3156 504
rect 3180 496 3188 504
rect 3532 496 3540 504
rect 3644 496 3652 504
rect 3852 496 3860 504
rect 3932 496 3940 504
rect 3948 496 3956 504
rect 4012 496 4020 504
rect 4316 496 4324 504
rect 4364 516 4372 524
rect 4396 516 4404 524
rect 4508 516 4516 524
rect 4540 516 4548 524
rect 4700 516 4708 524
rect 4716 516 4724 524
rect 4844 536 4852 544
rect 5020 536 5028 544
rect 4764 516 4772 524
rect 4780 516 4788 524
rect 4892 516 4900 524
rect 4908 516 4916 524
rect 5004 516 5012 524
rect 12 476 20 484
rect 204 476 212 484
rect 396 476 404 484
rect 1580 476 1588 484
rect 1916 476 1924 484
rect 2028 476 2036 484
rect 2860 476 2868 484
rect 3612 476 3620 484
rect 4684 476 4692 484
rect 4796 476 4804 484
rect 4876 476 4884 484
rect 1020 456 1028 464
rect 172 436 180 444
rect 652 436 660 444
rect 1196 436 1204 444
rect 1324 436 1332 444
rect 2924 436 2932 444
rect 3292 436 3300 444
rect 3564 436 3572 444
rect 3980 436 3988 444
rect 4636 436 4644 444
rect 4700 436 4708 444
rect 4780 436 4788 444
rect 4892 436 4900 444
rect 1043 406 1051 414
rect 1053 406 1061 414
rect 1063 406 1071 414
rect 1073 406 1081 414
rect 1083 406 1091 414
rect 1093 406 1101 414
rect 4051 406 4059 414
rect 4061 406 4069 414
rect 4071 406 4079 414
rect 4081 406 4089 414
rect 4091 406 4099 414
rect 4101 406 4109 414
rect 428 376 436 384
rect 924 376 932 384
rect 1340 376 1348 384
rect 1612 376 1620 384
rect 1660 376 1668 384
rect 1884 376 1892 384
rect 2316 376 2324 384
rect 2460 376 2468 384
rect 3372 376 3380 384
rect 3820 376 3828 384
rect 4188 376 4196 384
rect 2604 356 2612 364
rect 3436 356 3444 364
rect 12 336 20 344
rect 460 336 468 344
rect 988 336 996 344
rect 1116 336 1124 344
rect 3468 336 3476 344
rect 3852 336 3860 344
rect 4908 336 4916 344
rect 396 316 404 324
rect 572 316 580 324
rect 140 294 148 302
rect 284 296 292 304
rect 428 296 436 304
rect 476 296 484 304
rect 492 296 500 304
rect 540 296 548 304
rect 892 316 900 324
rect 956 316 964 324
rect 1372 316 1380 324
rect 1580 316 1588 324
rect 1692 316 1700 324
rect 2220 316 2228 324
rect 2716 316 2724 324
rect 620 296 628 304
rect 652 296 660 304
rect 828 294 836 302
rect 940 296 948 304
rect 988 296 996 304
rect 1116 296 1124 304
rect 1244 296 1252 304
rect 1340 296 1348 304
rect 1452 296 1460 304
rect 1516 294 1524 302
rect 1612 296 1620 304
rect 1772 296 1780 304
rect 1916 296 1924 304
rect 1964 296 1972 304
rect 1980 296 1988 304
rect 2012 296 2020 304
rect 2060 296 2068 304
rect 2076 296 2084 304
rect 2092 296 2100 304
rect 2140 296 2148 304
rect 2156 296 2164 304
rect 2188 296 2196 304
rect 2252 296 2260 304
rect 2300 296 2308 304
rect 2348 296 2356 304
rect 2364 296 2372 304
rect 2428 296 2436 304
rect 2444 296 2452 304
rect 2492 296 2500 304
rect 2508 296 2516 304
rect 2604 296 2612 304
rect 2636 296 2644 304
rect 2668 296 2676 304
rect 2684 296 2692 304
rect 2700 296 2708 304
rect 2748 296 2756 304
rect 2892 296 2900 304
rect 2988 296 2996 304
rect 3004 296 3012 304
rect 3036 316 3044 324
rect 3244 316 3252 324
rect 3276 316 3284 324
rect 3628 316 3636 324
rect 3740 316 3748 324
rect 3068 296 3076 304
rect 3116 296 3124 304
rect 3164 296 3172 304
rect 3180 296 3188 304
rect 3212 296 3220 304
rect 3260 296 3268 304
rect 3308 296 3316 304
rect 3340 296 3348 304
rect 3356 296 3364 304
rect 3420 296 3428 304
rect 3564 294 3572 302
rect 3644 296 3652 304
rect 3660 296 3668 304
rect 3692 296 3700 304
rect 4044 316 4052 324
rect 3788 296 3796 304
rect 4572 316 4580 324
rect 4668 316 4676 324
rect 4700 316 4708 324
rect 4796 316 4804 324
rect 4892 316 4900 324
rect 3948 294 3956 302
rect 4140 296 4148 304
rect 4156 296 4164 304
rect 4252 296 4260 304
rect 4268 296 4276 304
rect 4492 296 4500 304
rect 4668 296 4676 304
rect 4764 296 4772 304
rect 4860 296 4868 304
rect 4892 296 4900 304
rect 5004 296 5012 304
rect 172 276 180 284
rect 220 276 228 284
rect 268 276 276 284
rect 444 276 452 284
rect 508 276 516 284
rect 604 276 612 284
rect 636 276 644 284
rect 812 276 820 284
rect 940 276 948 284
rect 1004 276 1012 284
rect 1260 276 1268 284
rect 1324 276 1332 284
rect 1548 276 1556 284
rect 1628 276 1636 284
rect 1724 276 1732 284
rect 2012 276 2020 284
rect 2268 276 2276 284
rect 2572 276 2580 284
rect 2652 276 2660 284
rect 2764 276 2772 284
rect 2908 276 2916 284
rect 2972 276 2980 284
rect 3084 276 3092 284
rect 3100 276 3108 284
rect 3196 276 3204 284
rect 3324 276 3332 284
rect 3596 276 3604 284
rect 3676 276 3684 284
rect 3692 276 3700 284
rect 3772 276 3780 284
rect 3804 276 3812 284
rect 3980 276 3988 284
rect 4012 276 4020 284
rect 4172 276 4180 284
rect 4348 276 4356 284
rect 4508 276 4516 284
rect 4540 276 4548 284
rect 4604 276 4612 284
rect 4972 276 4980 284
rect 5020 276 5028 284
rect 44 256 52 264
rect 1852 256 1860 264
rect 1948 256 1956 264
rect 2380 256 2388 264
rect 2700 256 2708 264
rect 3500 256 3508 264
rect 4620 256 4628 264
rect 4716 256 4724 264
rect 4812 256 4820 264
rect 684 236 692 244
rect 700 236 708 244
rect 1020 236 1028 244
rect 1388 236 1396 244
rect 2156 236 2164 244
rect 2396 236 2404 244
rect 2780 236 2788 244
rect 4380 236 4388 244
rect 4588 236 4596 244
rect 4796 236 4804 244
rect 2547 206 2555 214
rect 2557 206 2565 214
rect 2567 206 2575 214
rect 2577 206 2585 214
rect 2587 206 2595 214
rect 2597 206 2605 214
rect 1260 176 1268 184
rect 1420 176 1428 184
rect 1660 176 1668 184
rect 1900 176 1908 184
rect 2620 176 2628 184
rect 2636 176 2644 184
rect 2700 176 2708 184
rect 3356 176 3364 184
rect 3532 176 3540 184
rect 3692 176 3700 184
rect 4620 176 4628 184
rect 4812 176 4820 184
rect 5020 176 5028 184
rect 556 156 564 164
rect 1548 156 1556 164
rect 2028 156 2036 164
rect 2220 156 2228 164
rect 2380 156 2388 164
rect 3132 156 3140 164
rect 3452 156 3460 164
rect 3484 156 3492 164
rect 4188 156 4196 164
rect 60 136 68 144
rect 220 136 228 144
rect 348 136 356 144
rect 460 136 468 144
rect 716 136 724 144
rect 844 136 852 144
rect 1132 136 1140 144
rect 1180 136 1188 144
rect 1244 136 1252 144
rect 1308 136 1316 144
rect 1820 136 1828 144
rect 2092 136 2100 144
rect 2140 136 2148 144
rect 2188 136 2196 144
rect 2204 136 2212 144
rect 2348 136 2356 144
rect 2412 136 2420 144
rect 2892 136 2900 144
rect 2940 136 2948 144
rect 2988 136 2996 144
rect 3196 136 3204 144
rect 3244 136 3252 144
rect 3292 136 3300 144
rect 3308 136 3316 144
rect 3372 136 3380 144
rect 3452 136 3460 144
rect 3852 136 3860 144
rect 3980 136 3988 144
rect 4140 136 4148 144
rect 4236 136 4244 144
rect 4348 136 4356 144
rect 4444 136 4452 144
rect 4540 136 4548 144
rect 4556 136 4564 144
rect 4604 136 4612 144
rect 4684 136 4692 144
rect 4780 136 4788 144
rect 4876 136 4884 144
rect 4972 136 4980 144
rect 5132 136 5140 144
rect 44 116 52 124
rect 92 116 100 124
rect 172 116 180 124
rect 236 118 244 126
rect 332 116 340 124
rect 396 116 404 124
rect 412 116 420 124
rect 444 116 452 124
rect 508 116 516 124
rect 588 116 596 124
rect 604 116 612 124
rect 732 116 740 124
rect 764 116 772 124
rect 812 116 820 124
rect 924 116 932 124
rect 1020 116 1028 124
rect 1244 116 1252 124
rect 1292 116 1300 124
rect 1356 116 1364 124
rect 1404 116 1412 124
rect 1548 118 1556 126
rect 1724 116 1732 124
rect 1788 118 1796 126
rect 1852 116 1860 124
rect 1964 116 1972 124
rect 2028 118 2036 126
rect 300 96 308 104
rect 332 96 340 104
rect 412 96 420 104
rect 764 96 772 104
rect 1132 96 1140 104
rect 1196 96 1204 104
rect 1260 96 1268 104
rect 2124 96 2132 104
rect 2172 116 2180 124
rect 2220 116 2228 124
rect 2252 116 2260 124
rect 2316 116 2324 124
rect 2332 116 2340 124
rect 2476 116 2484 124
rect 2684 116 2692 124
rect 2780 116 2788 124
rect 2828 118 2836 126
rect 2284 96 2292 104
rect 2924 96 2932 104
rect 2972 116 2980 124
rect 3132 118 3140 126
rect 3228 96 3236 104
rect 3276 116 3284 124
rect 3324 116 3332 124
rect 3388 116 3396 124
rect 3420 116 3428 124
rect 3436 116 3444 124
rect 3500 116 3508 124
rect 3564 116 3572 124
rect 3580 116 3588 124
rect 3612 116 3620 124
rect 3660 116 3668 124
rect 3772 116 3780 124
rect 4012 118 4020 126
rect 4172 96 4180 104
rect 4220 116 4228 124
rect 4380 118 4388 126
rect 4460 116 4468 124
rect 4476 116 4484 124
rect 4572 116 4580 124
rect 4700 116 4708 124
rect 4924 116 4932 124
rect 4508 96 4516 104
rect 4604 96 4612 104
rect 12 76 20 84
rect 108 76 116 84
rect 524 76 532 84
rect 1004 76 1012 84
rect 2348 76 2356 84
rect 3004 76 3012 84
rect 3884 76 3892 84
rect 4252 76 4260 84
rect 3628 56 3636 64
rect 364 36 372 44
rect 476 36 484 44
rect 780 36 788 44
rect 1116 36 1124 44
rect 1324 36 1332 44
rect 1372 36 1380 44
rect 1612 36 1620 44
rect 1884 36 1892 44
rect 3388 36 3396 44
rect 4620 36 4628 44
rect 1043 6 1051 14
rect 1053 6 1061 14
rect 1063 6 1071 14
rect 1073 6 1081 14
rect 1083 6 1091 14
rect 1093 6 1101 14
rect 4051 6 4059 14
rect 4061 6 4069 14
rect 4071 6 4079 14
rect 4081 6 4089 14
rect 4091 6 4099 14
rect 4101 6 4109 14
<< metal2 >>
rect 205 3457 227 3463
rect 269 3457 291 3463
rect 205 3384 211 3457
rect 285 3384 291 3457
rect 429 3457 451 3463
rect 429 3384 435 3457
rect 13 3284 19 3316
rect 125 3184 131 3336
rect 141 3326 147 3356
rect 253 3163 259 3316
rect 301 3304 307 3316
rect 253 3157 275 3163
rect 93 3104 99 3136
rect 13 3084 19 3096
rect 45 3004 51 3096
rect 13 2984 19 2996
rect 45 2743 51 2996
rect 125 2944 131 3036
rect 269 2984 275 3157
rect 349 3104 355 3316
rect 397 3284 403 3316
rect 365 3084 371 3256
rect 413 3244 419 3336
rect 461 3304 467 3316
rect 477 3303 483 3336
rect 669 3326 675 3336
rect 477 3297 499 3303
rect 381 3102 387 3156
rect 365 2944 371 3076
rect 125 2924 131 2936
rect 141 2744 147 2918
rect 205 2784 211 2836
rect 45 2737 67 2743
rect 61 2724 67 2737
rect 45 2704 51 2716
rect 13 2684 19 2696
rect 93 2677 108 2683
rect 45 2524 51 2676
rect 13 2484 19 2496
rect 45 2304 51 2316
rect 61 2304 67 2336
rect 93 2184 99 2677
rect 109 2664 115 2676
rect 125 2384 131 2456
rect 109 2304 115 2356
rect 141 2304 147 2696
rect 205 2684 211 2776
rect 269 2704 275 2916
rect 333 2824 339 2918
rect 429 2723 435 2896
rect 477 2823 483 3096
rect 493 3084 499 3297
rect 605 3264 611 3316
rect 701 3284 707 3463
rect 925 3344 931 3396
rect 1949 3384 1955 3463
rect 1501 3344 1507 3376
rect 1949 3344 1955 3376
rect 2253 3364 2259 3463
rect 2621 3457 2643 3463
rect 2570 3414 2582 3416
rect 2555 3406 2557 3414
rect 2565 3406 2567 3414
rect 2575 3406 2577 3414
rect 2585 3406 2587 3414
rect 2595 3406 2597 3414
rect 2570 3404 2582 3406
rect 2285 3344 2291 3396
rect 2429 3364 2435 3376
rect 749 3317 764 3323
rect 733 3304 739 3316
rect 589 3184 595 3236
rect 653 3184 659 3276
rect 557 3084 563 3136
rect 628 3117 636 3123
rect 461 2817 483 2823
rect 461 2743 467 2817
rect 461 2737 483 2743
rect 429 2717 444 2723
rect 381 2704 387 2716
rect 477 2704 483 2737
rect 317 2684 323 2694
rect 413 2624 419 2696
rect 477 2604 483 2696
rect 493 2684 499 3076
rect 493 2664 499 2676
rect 301 2464 307 2496
rect 157 2344 163 2436
rect 317 2304 323 2536
rect 333 2524 339 2556
rect 349 2524 355 2536
rect 365 2302 371 2316
rect 445 2304 451 2596
rect 509 2563 515 3076
rect 580 3057 595 3063
rect 589 2964 595 3057
rect 605 3024 611 3096
rect 589 2944 595 2956
rect 525 2704 531 2918
rect 637 2904 643 3116
rect 669 3104 675 3156
rect 653 2944 659 3096
rect 685 2944 691 3036
rect 701 2964 707 3036
rect 717 2984 723 3236
rect 733 3104 739 3276
rect 749 3184 755 3317
rect 781 3244 787 3336
rect 813 3184 819 3236
rect 829 3104 835 3176
rect 717 2923 723 2956
rect 733 2944 739 3076
rect 749 3064 755 3096
rect 861 3084 867 3256
rect 909 3104 915 3116
rect 925 3084 931 3336
rect 1069 3326 1075 3336
rect 1069 3317 1075 3318
rect 1005 3304 1011 3316
rect 1005 3264 1011 3296
rect 1165 3244 1171 3336
rect 1229 3304 1235 3316
rect 1293 3284 1299 3336
rect 1533 3324 1539 3336
rect 1373 3304 1379 3316
rect 1066 3214 1078 3216
rect 1051 3206 1053 3214
rect 1061 3206 1063 3214
rect 1071 3206 1073 3214
rect 1081 3206 1083 3214
rect 1091 3206 1093 3214
rect 1066 3204 1078 3206
rect 1133 3104 1139 3116
rect 1149 3084 1155 3116
rect 797 3044 803 3056
rect 845 2944 851 2996
rect 708 2917 723 2923
rect 637 2884 643 2896
rect 733 2844 739 2916
rect 781 2904 787 2916
rect 557 2724 563 2776
rect 541 2704 547 2716
rect 573 2644 579 2716
rect 589 2704 595 2736
rect 653 2704 659 2816
rect 669 2704 675 2736
rect 701 2724 707 2756
rect 733 2704 739 2756
rect 765 2724 771 2876
rect 605 2684 611 2696
rect 749 2684 755 2696
rect 573 2584 579 2616
rect 493 2557 515 2563
rect 493 2544 499 2557
rect 493 2384 499 2536
rect 541 2484 547 2516
rect 564 2497 572 2503
rect 477 2324 483 2356
rect 493 2324 499 2336
rect 557 2324 563 2496
rect 109 2144 115 2276
rect 125 2124 131 2296
rect 461 2303 467 2316
rect 461 2297 476 2303
rect 61 2104 67 2116
rect 13 2084 19 2096
rect 45 1904 51 1916
rect 109 1904 115 2096
rect 125 1904 131 2116
rect 141 2104 147 2116
rect 157 2104 163 2116
rect 173 2044 179 2276
rect 301 2164 307 2276
rect 141 1984 147 2036
rect 13 1884 19 1896
rect 61 1864 67 1896
rect 93 1884 99 1896
rect 61 1784 67 1856
rect 93 1704 99 1736
rect 45 1504 51 1516
rect 61 1504 67 1636
rect 109 1504 115 1896
rect 141 1744 147 1836
rect 221 1784 227 1816
rect 285 1784 291 1936
rect 333 1884 339 2136
rect 397 2124 403 2156
rect 413 1924 419 2116
rect 445 1984 451 2296
rect 541 2164 547 2276
rect 525 2144 531 2156
rect 509 2084 515 2116
rect 461 1964 467 2036
rect 541 1984 547 2116
rect 557 1964 563 2316
rect 589 2164 595 2596
rect 605 2524 611 2616
rect 621 2584 627 2676
rect 685 2644 691 2676
rect 637 2564 643 2596
rect 765 2564 771 2716
rect 813 2704 819 2916
rect 861 2904 867 2916
rect 893 2824 899 3056
rect 941 2924 947 2956
rect 973 2924 979 2936
rect 989 2924 995 2936
rect 1005 2924 1011 3056
rect 1037 3044 1043 3076
rect 1037 2944 1043 2956
rect 1165 2924 1171 3236
rect 1181 3104 1187 3256
rect 1197 3084 1203 3276
rect 1181 2924 1187 2996
rect 1197 2984 1203 3076
rect 909 2904 915 2916
rect 1005 2904 1011 2916
rect 845 2703 851 2756
rect 861 2704 867 2776
rect 909 2744 915 2896
rect 877 2704 883 2736
rect 836 2697 851 2703
rect 781 2643 787 2696
rect 797 2663 803 2676
rect 797 2657 828 2663
rect 909 2643 915 2716
rect 925 2704 931 2796
rect 932 2677 940 2683
rect 781 2637 915 2643
rect 861 2563 867 2576
rect 861 2557 876 2563
rect 877 2544 883 2556
rect 605 2304 611 2336
rect 605 2263 611 2276
rect 605 2257 627 2263
rect 621 2164 627 2257
rect 637 2184 643 2536
rect 765 2524 771 2536
rect 669 2504 675 2516
rect 685 2184 691 2256
rect 781 2164 787 2516
rect 909 2504 915 2516
rect 813 2284 819 2316
rect 861 2284 867 2436
rect 877 2264 883 2316
rect 909 2304 915 2316
rect 925 2284 931 2676
rect 973 2563 979 2896
rect 1021 2684 1027 2816
rect 1066 2814 1078 2816
rect 1051 2806 1053 2814
rect 1061 2806 1063 2814
rect 1071 2806 1073 2814
rect 1081 2806 1083 2814
rect 1091 2806 1093 2814
rect 1066 2804 1078 2806
rect 1037 2664 1043 2696
rect 1117 2684 1123 2796
rect 1133 2784 1139 2856
rect 1149 2784 1155 2856
rect 973 2557 995 2563
rect 973 2383 979 2536
rect 989 2524 995 2557
rect 1005 2524 1011 2556
rect 1149 2544 1155 2736
rect 1197 2664 1203 2836
rect 1213 2744 1219 3076
rect 1229 2984 1235 3096
rect 1293 3084 1299 3116
rect 1309 2964 1315 3156
rect 1325 3064 1331 3096
rect 1341 3084 1347 3296
rect 1533 3224 1539 3296
rect 1565 3104 1571 3296
rect 1581 3224 1587 3316
rect 1597 3277 1612 3283
rect 1245 2924 1251 2956
rect 1245 2684 1251 2916
rect 1325 2804 1331 3056
rect 1373 3044 1379 3096
rect 1421 3064 1427 3096
rect 1341 2924 1347 2936
rect 1357 2924 1363 2956
rect 1373 2924 1379 3036
rect 1389 2984 1395 3036
rect 1421 2924 1427 3056
rect 1437 2924 1443 3096
rect 1485 3064 1491 3076
rect 1501 3004 1507 3036
rect 1293 2784 1299 2796
rect 1261 2724 1267 2776
rect 1277 2684 1283 2776
rect 1341 2704 1347 2836
rect 1389 2704 1395 2836
rect 1453 2784 1459 2936
rect 1469 2924 1475 2976
rect 1517 2944 1523 2976
rect 1533 2944 1539 2956
rect 1501 2904 1507 2916
rect 1437 2704 1443 2716
rect 1229 2544 1235 2676
rect 1293 2664 1299 2696
rect 1453 2683 1459 2736
rect 1469 2724 1475 2836
rect 1501 2784 1507 2796
rect 1485 2704 1491 2716
rect 1501 2684 1507 2756
rect 1533 2684 1539 2696
rect 1565 2684 1571 3096
rect 1597 3084 1603 3277
rect 1709 3104 1715 3336
rect 1837 3324 1843 3336
rect 1853 3244 1859 3336
rect 1869 3324 1875 3336
rect 2029 3284 2035 3316
rect 2077 3304 2083 3316
rect 2157 3244 2163 3336
rect 2173 3324 2179 3336
rect 1629 3102 1635 3103
rect 1597 2964 1603 3076
rect 1629 2984 1635 3094
rect 1693 3044 1699 3056
rect 1725 3004 1731 3136
rect 1629 2924 1635 2936
rect 1629 2904 1635 2916
rect 1581 2784 1587 2896
rect 1645 2883 1651 2916
rect 1629 2877 1651 2883
rect 1437 2677 1459 2683
rect 1341 2664 1347 2676
rect 1309 2643 1315 2656
rect 1268 2637 1315 2643
rect 1261 2584 1267 2616
rect 1165 2524 1171 2536
rect 1197 2504 1203 2516
rect 1066 2414 1078 2416
rect 1051 2406 1053 2414
rect 1061 2406 1063 2414
rect 1071 2406 1073 2414
rect 1081 2406 1083 2414
rect 1091 2406 1093 2414
rect 1066 2404 1078 2406
rect 1117 2404 1123 2496
rect 1213 2484 1219 2536
rect 1229 2524 1235 2536
rect 1245 2524 1251 2576
rect 1325 2564 1331 2596
rect 1357 2524 1363 2616
rect 1405 2564 1411 2596
rect 1373 2484 1379 2516
rect 973 2377 988 2383
rect 589 2004 595 2156
rect 621 2124 627 2136
rect 669 2124 675 2156
rect 925 2144 931 2256
rect 941 2184 947 2316
rect 973 2224 979 2296
rect 989 2284 995 2376
rect 957 2217 972 2223
rect 525 1924 531 1956
rect 589 1924 595 1956
rect 349 1744 355 1776
rect 381 1744 387 1876
rect 413 1864 419 1896
rect 461 1884 467 1916
rect 621 1904 627 2056
rect 509 1884 515 1896
rect 557 1864 563 1896
rect 157 1704 163 1716
rect 173 1584 179 1696
rect 285 1684 291 1696
rect 317 1504 323 1716
rect 13 1484 19 1496
rect 93 1484 99 1496
rect 109 1404 115 1496
rect 45 1324 51 1376
rect 141 1344 147 1436
rect 285 1383 291 1476
rect 269 1377 291 1383
rect 61 1304 67 1336
rect 93 1304 99 1316
rect 45 1104 51 1116
rect 13 1084 19 1096
rect 45 1037 60 1043
rect 45 924 51 1037
rect 173 984 179 1096
rect 189 1084 195 1336
rect 237 1326 243 1356
rect 269 1344 275 1377
rect 301 1304 307 1376
rect 333 1324 339 1496
rect 381 1484 387 1736
rect 429 1524 435 1716
rect 333 1303 339 1316
rect 317 1297 339 1303
rect 221 944 227 1156
rect 317 1104 323 1297
rect 333 1184 339 1256
rect 253 943 259 1076
rect 244 937 259 943
rect 269 923 275 1096
rect 349 1084 355 1336
rect 365 1124 371 1136
rect 349 1064 355 1076
rect 260 917 275 923
rect 93 904 99 916
rect 109 904 115 916
rect 13 884 19 896
rect 173 884 179 896
rect 221 764 227 916
rect 333 844 339 1036
rect 429 926 435 936
rect 45 704 51 736
rect 349 704 355 716
rect 61 544 67 676
rect 141 624 147 636
rect 269 524 275 676
rect 333 526 339 556
rect 365 544 371 916
rect 397 724 403 736
rect 461 724 467 1856
rect 557 1784 563 1836
rect 589 1724 595 1836
rect 653 1644 659 1856
rect 669 1764 675 2116
rect 685 1904 691 1956
rect 797 1904 803 2136
rect 813 2124 819 2136
rect 541 1624 547 1636
rect 477 1504 483 1556
rect 653 1484 659 1636
rect 525 1344 531 1476
rect 525 1084 531 1336
rect 653 1324 659 1396
rect 669 1344 675 1436
rect 685 1424 691 1876
rect 717 1744 723 1876
rect 749 1744 755 1836
rect 701 1504 707 1536
rect 685 1344 691 1416
rect 701 1384 707 1476
rect 557 1284 563 1318
rect 557 1124 563 1136
rect 589 1104 595 1136
rect 557 1084 563 1096
rect 557 964 563 1016
rect 605 964 611 1016
rect 525 924 531 936
rect 589 924 595 956
rect 637 944 643 1076
rect 669 963 675 1316
rect 717 1144 723 1316
rect 717 1104 723 1116
rect 685 984 691 1076
rect 733 1023 739 1296
rect 733 1017 755 1023
rect 701 964 707 1016
rect 660 957 675 963
rect 493 904 499 916
rect 509 724 515 736
rect 461 704 467 716
rect 429 664 435 696
rect 557 684 563 876
rect 580 697 595 703
rect 429 524 435 656
rect 445 644 451 676
rect 445 544 451 636
rect 13 484 19 496
rect 45 484 51 516
rect 141 302 147 356
rect 173 284 179 436
rect 269 284 275 516
rect 285 304 291 516
rect 429 384 435 476
rect 45 124 51 256
rect 173 124 179 276
rect 221 144 227 276
rect 333 124 339 196
rect 349 144 355 276
rect 397 124 403 316
rect 429 204 435 296
rect 445 284 451 536
rect 461 484 467 496
rect 477 304 483 456
rect 493 384 499 636
rect 493 304 499 376
rect 541 304 547 656
rect 589 644 595 697
rect 557 524 563 576
rect 621 544 627 836
rect 637 544 643 736
rect 653 544 659 836
rect 685 804 691 916
rect 749 904 755 1017
rect 749 863 755 896
rect 733 857 755 863
rect 717 744 723 836
rect 589 523 595 536
rect 685 524 691 636
rect 717 564 723 716
rect 733 564 739 857
rect 749 784 755 836
rect 765 704 771 1756
rect 797 1724 803 1736
rect 813 1704 819 1996
rect 925 1984 931 2116
rect 957 2104 963 2217
rect 973 2144 979 2176
rect 1053 2124 1059 2156
rect 1117 2144 1123 2256
rect 1053 2104 1059 2116
rect 1069 2044 1075 2136
rect 877 1924 883 1936
rect 900 1897 915 1903
rect 845 1744 851 1756
rect 781 1684 787 1696
rect 781 1384 787 1436
rect 797 1424 803 1436
rect 813 1403 819 1696
rect 829 1684 835 1716
rect 829 1484 835 1496
rect 797 1397 819 1403
rect 797 1364 803 1397
rect 829 1364 835 1396
rect 845 1384 851 1476
rect 813 1323 819 1356
rect 804 1317 819 1323
rect 829 1264 835 1316
rect 813 1164 819 1236
rect 861 1163 867 1676
rect 909 1643 915 1897
rect 941 1884 947 2036
rect 1066 2014 1078 2016
rect 1051 2006 1053 2014
rect 1061 2006 1063 2014
rect 1071 2006 1073 2014
rect 1081 2006 1083 2014
rect 1091 2006 1093 2014
rect 1066 2004 1078 2006
rect 1053 1904 1059 1916
rect 941 1764 947 1876
rect 893 1637 915 1643
rect 877 1504 883 1516
rect 893 1484 899 1637
rect 909 1504 915 1536
rect 877 1164 883 1316
rect 909 1304 915 1316
rect 925 1184 931 1496
rect 941 1484 947 1536
rect 957 1503 963 1896
rect 1037 1884 1043 1896
rect 989 1504 995 1516
rect 957 1497 972 1503
rect 973 1484 979 1496
rect 1005 1464 1011 1876
rect 1117 1744 1123 2136
rect 1133 1884 1139 2456
rect 1245 2324 1251 2336
rect 1149 2144 1155 2276
rect 1229 2243 1235 2316
rect 1245 2264 1251 2316
rect 1277 2304 1283 2436
rect 1373 2424 1379 2436
rect 1309 2304 1315 2416
rect 1341 2304 1347 2316
rect 1261 2284 1267 2296
rect 1229 2237 1276 2243
rect 1149 2104 1155 2136
rect 1197 2124 1203 2196
rect 1165 1984 1171 2116
rect 1213 1904 1219 2116
rect 1197 1884 1203 1896
rect 1245 1884 1251 1896
rect 1277 1884 1283 2136
rect 1341 2043 1347 2296
rect 1357 2124 1363 2356
rect 1373 2304 1379 2316
rect 1389 2284 1395 2536
rect 1405 2463 1411 2496
rect 1421 2484 1427 2516
rect 1405 2457 1427 2463
rect 1421 2384 1427 2457
rect 1437 2323 1443 2677
rect 1453 2424 1459 2656
rect 1437 2317 1452 2323
rect 1485 2303 1491 2616
rect 1501 2504 1507 2636
rect 1581 2544 1587 2556
rect 1476 2297 1491 2303
rect 1501 2283 1507 2476
rect 1581 2443 1587 2536
rect 1565 2437 1587 2443
rect 1533 2384 1539 2436
rect 1517 2284 1523 2336
rect 1485 2277 1507 2283
rect 1325 2037 1347 2043
rect 1293 1904 1299 1916
rect 1309 1884 1315 1916
rect 1325 1884 1331 2037
rect 1341 1904 1347 1916
rect 1373 1904 1379 2096
rect 1389 1904 1395 2276
rect 1469 2204 1475 2256
rect 1485 2124 1491 2277
rect 1501 2163 1507 2256
rect 1517 2204 1523 2256
rect 1549 2164 1555 2296
rect 1501 2157 1516 2163
rect 1565 2144 1571 2437
rect 1581 2304 1587 2416
rect 1613 2384 1619 2536
rect 1629 2524 1635 2877
rect 1661 2864 1667 2896
rect 1629 2504 1635 2516
rect 1645 2504 1651 2576
rect 1661 2524 1667 2536
rect 1677 2504 1683 2536
rect 1693 2464 1699 2936
rect 1709 2904 1715 2996
rect 1805 2983 1811 3196
rect 1821 3102 1827 3136
rect 1917 3084 1923 3176
rect 1949 3124 1955 3216
rect 1949 3104 1955 3116
rect 1981 3083 1987 3116
rect 2013 3084 2019 3216
rect 2045 3104 2051 3176
rect 2077 3102 2083 3116
rect 1981 3077 2003 3083
rect 1997 3063 2003 3077
rect 1997 3057 2019 3063
rect 2013 3043 2019 3057
rect 2013 3037 2051 3043
rect 2045 3023 2051 3037
rect 2045 3017 2083 3023
rect 2077 2984 2083 3017
rect 1805 2977 1820 2983
rect 1988 2977 2051 2983
rect 1949 2926 1955 2956
rect 2013 2944 2019 2956
rect 2045 2944 2051 2977
rect 2093 2944 2099 3076
rect 2109 2964 2115 3216
rect 2141 3104 2147 3116
rect 2173 3023 2179 3316
rect 2141 3017 2179 3023
rect 1949 2917 1955 2918
rect 1741 2864 1747 2916
rect 1805 2904 1811 2916
rect 1709 2564 1715 2856
rect 1965 2837 2003 2843
rect 1965 2783 1971 2837
rect 1997 2824 2003 2837
rect 1821 2777 1971 2783
rect 1821 2764 1827 2777
rect 1837 2757 1955 2763
rect 1837 2704 1843 2757
rect 1748 2697 1763 2703
rect 1725 2584 1731 2636
rect 1709 2524 1715 2556
rect 1725 2464 1731 2536
rect 1741 2524 1747 2676
rect 1757 2624 1763 2697
rect 1853 2684 1859 2736
rect 1869 2704 1875 2736
rect 1949 2724 1955 2757
rect 1981 2744 1987 2816
rect 2013 2723 2019 2936
rect 2029 2884 2035 2916
rect 2125 2903 2131 2936
rect 2141 2924 2147 3017
rect 2109 2897 2131 2903
rect 2077 2884 2083 2896
rect 2093 2863 2099 2876
rect 2061 2857 2099 2863
rect 2061 2844 2067 2857
rect 2061 2784 2067 2816
rect 1997 2717 2019 2723
rect 1796 2677 1843 2683
rect 1773 2584 1779 2656
rect 1821 2584 1827 2656
rect 1837 2643 1843 2677
rect 1853 2664 1859 2676
rect 1837 2637 1868 2643
rect 1885 2584 1891 2656
rect 1901 2544 1907 2696
rect 1917 2664 1923 2676
rect 1981 2664 1987 2696
rect 1997 2684 2003 2717
rect 2077 2704 2083 2836
rect 2109 2784 2115 2897
rect 2141 2864 2147 2916
rect 2141 2824 2147 2856
rect 2093 2724 2099 2756
rect 2109 2717 2147 2723
rect 2013 2697 2028 2703
rect 1821 2444 1827 2536
rect 1645 2304 1651 2436
rect 1773 2337 1811 2343
rect 1773 2323 1779 2337
rect 1757 2317 1779 2323
rect 1757 2303 1763 2317
rect 1789 2304 1795 2316
rect 1805 2304 1811 2337
rect 1821 2304 1827 2436
rect 1741 2297 1763 2303
rect 1581 2124 1587 2296
rect 1629 2184 1635 2296
rect 1741 2284 1747 2297
rect 1661 2264 1667 2276
rect 1725 2257 1740 2263
rect 1597 2124 1603 2176
rect 1613 2103 1619 2116
rect 1597 2097 1619 2103
rect 1485 2084 1491 2096
rect 1405 1917 1420 1923
rect 1405 1883 1411 1917
rect 1421 1884 1427 1896
rect 1469 1884 1475 1916
rect 1485 1904 1491 2016
rect 1396 1877 1411 1883
rect 1197 1844 1203 1876
rect 1277 1804 1283 1876
rect 1229 1784 1235 1796
rect 1213 1744 1219 1776
rect 1021 1524 1027 1616
rect 1066 1614 1078 1616
rect 1051 1606 1053 1614
rect 1061 1606 1063 1614
rect 1071 1606 1073 1614
rect 1081 1606 1083 1614
rect 1091 1606 1093 1614
rect 1066 1604 1078 1606
rect 1117 1544 1123 1716
rect 1133 1684 1139 1716
rect 1181 1684 1187 1696
rect 1021 1444 1027 1516
rect 957 1344 963 1416
rect 845 1157 867 1163
rect 845 1124 851 1157
rect 845 1104 851 1116
rect 861 1084 867 1116
rect 781 924 787 1076
rect 797 944 803 1056
rect 877 944 883 976
rect 797 883 803 936
rect 829 884 835 916
rect 797 877 819 883
rect 749 664 755 696
rect 765 624 771 676
rect 573 517 595 523
rect 573 364 579 517
rect 589 464 595 496
rect 621 484 627 516
rect 445 124 451 176
rect 461 144 467 156
rect 541 124 547 296
rect 573 283 579 316
rect 621 304 627 336
rect 653 304 659 436
rect 637 284 643 296
rect 765 284 771 616
rect 781 526 787 816
rect 813 784 819 877
rect 813 724 819 776
rect 877 684 883 936
rect 893 924 899 936
rect 909 864 915 1076
rect 941 1024 947 1096
rect 973 1064 979 1336
rect 989 1284 995 1316
rect 1037 1243 1043 1476
rect 1053 1464 1059 1496
rect 1069 1244 1075 1476
rect 1085 1424 1091 1516
rect 1101 1364 1107 1416
rect 1117 1324 1123 1496
rect 1165 1444 1171 1496
rect 1181 1444 1187 1676
rect 1213 1504 1219 1736
rect 1293 1704 1299 1856
rect 1325 1804 1331 1876
rect 1421 1744 1427 1876
rect 1469 1804 1475 1876
rect 1517 1844 1523 1896
rect 1533 1823 1539 2036
rect 1549 1924 1555 2096
rect 1565 2024 1571 2036
rect 1517 1817 1539 1823
rect 1476 1797 1491 1803
rect 1469 1724 1475 1736
rect 1460 1697 1475 1703
rect 1245 1464 1251 1636
rect 1277 1504 1283 1596
rect 1293 1464 1299 1696
rect 1341 1504 1347 1516
rect 1325 1463 1331 1496
rect 1357 1483 1363 1536
rect 1405 1524 1411 1676
rect 1348 1477 1363 1483
rect 1325 1457 1347 1463
rect 1021 1237 1043 1243
rect 989 1104 995 1136
rect 1005 1024 1011 1096
rect 989 984 995 1016
rect 989 924 995 976
rect 1005 864 1011 936
rect 1021 924 1027 1237
rect 1066 1214 1078 1216
rect 1051 1206 1053 1214
rect 1061 1206 1063 1214
rect 1071 1206 1073 1214
rect 1081 1206 1083 1214
rect 1091 1206 1093 1214
rect 1066 1204 1078 1206
rect 1133 1203 1139 1356
rect 1149 1324 1155 1336
rect 1165 1324 1171 1436
rect 1181 1304 1187 1336
rect 1133 1197 1155 1203
rect 1117 1164 1123 1196
rect 1117 924 1123 1056
rect 1117 904 1123 916
rect 1066 814 1078 816
rect 1051 806 1053 814
rect 1061 806 1063 814
rect 1071 806 1073 814
rect 1081 806 1083 814
rect 1091 806 1093 814
rect 1066 804 1078 806
rect 1021 783 1027 796
rect 1021 777 1043 783
rect 1037 763 1043 777
rect 1037 757 1075 763
rect 1069 744 1075 757
rect 925 704 931 736
rect 845 664 851 676
rect 813 544 819 656
rect 781 517 787 518
rect 813 284 819 536
rect 877 524 883 536
rect 893 504 899 556
rect 909 504 915 556
rect 941 544 947 716
rect 1037 704 1043 716
rect 1053 704 1059 736
rect 1133 724 1139 1176
rect 1149 1104 1155 1197
rect 1165 1084 1171 1116
rect 1181 1084 1187 1296
rect 1197 1164 1203 1436
rect 1213 1324 1219 1336
rect 1197 1024 1203 1096
rect 1213 1084 1219 1116
rect 1245 1104 1251 1136
rect 1213 924 1219 1076
rect 1005 544 1011 576
rect 1053 524 1059 536
rect 829 302 835 456
rect 925 384 931 496
rect 941 423 947 516
rect 973 464 979 516
rect 989 504 995 516
rect 1069 504 1075 516
rect 1133 464 1139 496
rect 941 417 963 423
rect 957 384 963 417
rect 941 324 947 376
rect 1021 364 1027 456
rect 1066 414 1078 416
rect 1051 406 1053 414
rect 1061 406 1063 414
rect 1071 406 1073 414
rect 1081 406 1083 414
rect 1091 406 1093 414
rect 1066 404 1078 406
rect 957 324 963 356
rect 1117 344 1123 436
rect 557 277 579 283
rect 557 164 563 277
rect 589 124 595 136
rect 605 124 611 276
rect 13 84 19 96
rect 93 83 99 116
rect 109 84 115 96
rect 93 77 108 83
rect 509 83 515 116
rect 509 77 524 83
rect 365 -17 371 36
rect 477 -17 483 36
rect 685 -17 691 236
rect 717 144 723 276
rect 797 123 803 236
rect 813 144 819 276
rect 893 244 899 316
rect 941 304 947 316
rect 1117 304 1123 336
rect 989 224 995 296
rect 1005 244 1011 276
rect 1021 143 1027 236
rect 1133 204 1139 456
rect 1149 164 1155 796
rect 1181 784 1187 916
rect 1197 844 1203 896
rect 1181 684 1187 776
rect 1165 524 1171 596
rect 1197 244 1203 436
rect 1021 137 1043 143
rect 925 124 931 136
rect 797 117 812 123
rect 1005 84 1011 96
rect 1021 83 1027 116
rect 1012 77 1027 83
rect 1037 44 1043 137
rect 1133 104 1139 116
rect 1197 104 1203 196
rect 1213 144 1219 836
rect 1229 703 1235 1016
rect 1261 943 1267 1436
rect 1341 1424 1347 1457
rect 1421 1424 1427 1516
rect 1437 1504 1443 1556
rect 1453 1484 1459 1496
rect 1325 1403 1331 1416
rect 1325 1397 1363 1403
rect 1357 1384 1363 1397
rect 1325 1344 1331 1376
rect 1453 1364 1459 1476
rect 1389 1357 1436 1363
rect 1389 1343 1395 1357
rect 1373 1337 1395 1343
rect 1284 1317 1299 1323
rect 1293 1304 1299 1317
rect 1277 1184 1283 1276
rect 1293 1064 1299 1096
rect 1309 1024 1315 1316
rect 1357 1284 1363 1316
rect 1341 1184 1347 1216
rect 1373 1163 1379 1337
rect 1405 1224 1411 1336
rect 1357 1157 1379 1163
rect 1341 1104 1347 1116
rect 1325 1084 1331 1096
rect 1252 937 1267 943
rect 1293 924 1299 976
rect 1293 784 1299 896
rect 1309 704 1315 736
rect 1325 704 1331 936
rect 1341 924 1347 1056
rect 1357 984 1363 1157
rect 1421 1144 1427 1336
rect 1437 1284 1443 1316
rect 1469 1263 1475 1697
rect 1485 1523 1491 1797
rect 1517 1744 1523 1817
rect 1549 1803 1555 1856
rect 1533 1797 1555 1803
rect 1533 1784 1539 1797
rect 1565 1724 1571 1936
rect 1581 1904 1587 2076
rect 1597 1884 1603 2097
rect 1629 2084 1635 2096
rect 1597 1724 1603 1876
rect 1629 1863 1635 2016
rect 1709 1924 1715 1956
rect 1725 1924 1731 2257
rect 1741 2124 1747 2136
rect 1757 2103 1763 2276
rect 1741 2097 1763 2103
rect 1645 1864 1651 1916
rect 1741 1904 1747 2097
rect 1613 1857 1635 1863
rect 1533 1584 1539 1596
rect 1485 1517 1500 1523
rect 1501 1504 1507 1516
rect 1565 1504 1571 1576
rect 1540 1497 1555 1503
rect 1549 1483 1555 1497
rect 1581 1484 1587 1496
rect 1549 1477 1571 1483
rect 1565 1463 1571 1477
rect 1597 1464 1603 1636
rect 1613 1483 1619 1857
rect 1645 1784 1651 1856
rect 1645 1724 1651 1736
rect 1645 1643 1651 1656
rect 1661 1644 1667 1856
rect 1677 1764 1683 1836
rect 1693 1764 1699 1896
rect 1709 1726 1715 1836
rect 1741 1804 1747 1896
rect 1757 1884 1763 2036
rect 1773 1944 1779 2276
rect 1789 2264 1795 2296
rect 1869 2284 1875 2516
rect 1901 2323 1907 2496
rect 1892 2317 1907 2323
rect 1773 1784 1779 1896
rect 1789 1823 1795 2196
rect 1805 1864 1811 1896
rect 1821 1884 1827 2096
rect 1837 2084 1843 2276
rect 1901 2264 1907 2317
rect 1853 2164 1859 2196
rect 1869 2184 1875 2196
rect 1853 1924 1859 2036
rect 1869 1964 1875 2116
rect 1885 2024 1891 2196
rect 1901 2124 1907 2156
rect 1917 2124 1923 2516
rect 1933 2504 1939 2576
rect 1949 2483 1955 2616
rect 1997 2584 2003 2656
rect 1965 2524 1971 2556
rect 1981 2544 1987 2556
rect 1981 2524 1987 2536
rect 1997 2503 2003 2516
rect 1981 2497 2003 2503
rect 1949 2477 1971 2483
rect 1965 2384 1971 2477
rect 1949 2324 1955 2356
rect 1956 2297 1971 2303
rect 1933 2277 1948 2283
rect 1901 1964 1907 2076
rect 1933 2044 1939 2277
rect 1965 2264 1971 2297
rect 1981 2264 1987 2497
rect 2013 2444 2019 2697
rect 2109 2703 2115 2717
rect 2141 2704 2147 2717
rect 2157 2704 2163 2936
rect 2173 2904 2179 2976
rect 2173 2864 2179 2896
rect 2189 2843 2195 3236
rect 2269 3184 2275 3336
rect 2349 3304 2355 3316
rect 2525 3304 2531 3396
rect 2621 3383 2627 3457
rect 2589 3377 2627 3383
rect 2557 3326 2563 3336
rect 2285 3123 2291 3236
rect 2333 3144 2339 3276
rect 2276 3117 2291 3123
rect 2221 3064 2227 3076
rect 2253 3044 2259 3076
rect 2205 2903 2211 2916
rect 2253 2903 2259 2936
rect 2269 2924 2275 3096
rect 2333 3064 2339 3136
rect 2349 3124 2355 3296
rect 2372 3137 2387 3143
rect 2205 2897 2259 2903
rect 2173 2837 2195 2843
rect 2093 2697 2115 2703
rect 2093 2683 2099 2697
rect 2052 2677 2099 2683
rect 2125 2677 2140 2683
rect 2109 2664 2115 2676
rect 2029 2584 2035 2656
rect 2045 2644 2051 2656
rect 2013 2304 2019 2436
rect 1997 2163 2003 2296
rect 1981 2157 2003 2163
rect 1949 2004 1955 2036
rect 1917 1984 1923 1996
rect 1837 1884 1843 1916
rect 1789 1817 1811 1823
rect 1805 1724 1811 1817
rect 1805 1704 1811 1716
rect 1629 1637 1651 1643
rect 1629 1584 1635 1637
rect 1645 1523 1651 1596
rect 1629 1517 1651 1523
rect 1629 1504 1635 1517
rect 1677 1483 1683 1616
rect 1693 1484 1699 1556
rect 1709 1524 1715 1556
rect 1757 1504 1763 1556
rect 1613 1477 1651 1483
rect 1565 1457 1587 1463
rect 1581 1443 1587 1457
rect 1629 1443 1635 1456
rect 1581 1437 1635 1443
rect 1501 1344 1507 1356
rect 1485 1284 1491 1336
rect 1517 1324 1523 1376
rect 1581 1337 1612 1343
rect 1581 1323 1587 1337
rect 1533 1317 1587 1323
rect 1501 1303 1507 1316
rect 1533 1303 1539 1317
rect 1501 1297 1539 1303
rect 1469 1257 1491 1263
rect 1373 1124 1379 1136
rect 1373 944 1379 1076
rect 1389 984 1395 1036
rect 1389 944 1395 956
rect 1373 924 1379 936
rect 1421 924 1427 1036
rect 1453 1023 1459 1096
rect 1437 1017 1459 1023
rect 1341 724 1347 836
rect 1357 824 1363 916
rect 1389 904 1395 916
rect 1405 883 1411 896
rect 1389 877 1411 883
rect 1389 784 1395 877
rect 1405 704 1411 736
rect 1229 697 1244 703
rect 1261 684 1267 696
rect 1229 584 1235 636
rect 1245 524 1251 656
rect 1277 584 1283 696
rect 1325 664 1331 696
rect 1357 684 1363 696
rect 1341 544 1347 616
rect 1357 584 1363 676
rect 1437 544 1443 1017
rect 1453 904 1459 916
rect 1469 724 1475 1216
rect 1485 1184 1491 1257
rect 1485 1024 1491 1156
rect 1549 1144 1555 1296
rect 1597 1284 1603 1316
rect 1565 1164 1571 1236
rect 1581 1164 1587 1196
rect 1517 1023 1523 1056
rect 1517 1017 1539 1023
rect 1485 924 1491 1016
rect 1533 984 1539 1017
rect 1581 984 1587 1076
rect 1501 944 1507 976
rect 1517 924 1523 936
rect 1597 924 1603 1136
rect 1613 1084 1619 1096
rect 1645 1003 1651 1477
rect 1661 1477 1683 1483
rect 1661 1364 1667 1477
rect 1677 1424 1683 1456
rect 1725 1424 1731 1496
rect 1741 1364 1747 1376
rect 1773 1324 1779 1636
rect 1805 1504 1811 1596
rect 1821 1524 1827 1836
rect 1853 1824 1859 1896
rect 1837 1724 1843 1736
rect 1853 1584 1859 1636
rect 1821 1484 1827 1516
rect 1837 1504 1843 1516
rect 1837 1464 1843 1496
rect 1805 1424 1811 1436
rect 1869 1403 1875 1956
rect 1885 1904 1891 1916
rect 1917 1904 1923 1956
rect 1965 1924 1971 2136
rect 1981 1983 1987 2157
rect 1997 2004 2003 2096
rect 1981 1977 2003 1983
rect 1997 1964 2003 1977
rect 2013 1943 2019 2276
rect 2045 2264 2051 2596
rect 2061 2504 2067 2516
rect 2077 2483 2083 2576
rect 2061 2477 2083 2483
rect 2061 2424 2067 2477
rect 2077 2304 2083 2436
rect 2029 1964 2035 2256
rect 2077 2184 2083 2236
rect 2093 2223 2099 2616
rect 2109 2524 2115 2576
rect 2125 2524 2131 2677
rect 2157 2663 2163 2676
rect 2148 2657 2163 2663
rect 2173 2584 2179 2837
rect 2205 2744 2211 2856
rect 2285 2843 2291 2976
rect 2317 2924 2323 3036
rect 2349 2944 2355 3116
rect 2365 3104 2371 3116
rect 2381 3104 2387 3137
rect 2381 2944 2387 3076
rect 2333 2924 2339 2936
rect 2349 2904 2355 2936
rect 2413 2883 2419 3216
rect 2429 3104 2435 3296
rect 2589 3284 2595 3377
rect 2621 3284 2627 3356
rect 2445 3084 2451 3236
rect 2477 3084 2483 3096
rect 2525 3084 2531 3196
rect 2605 3104 2611 3116
rect 2612 3097 2627 3103
rect 2429 3024 2435 3036
rect 2445 2944 2451 3016
rect 2461 2944 2467 3076
rect 2477 3004 2483 3036
rect 2461 2903 2467 2916
rect 2445 2897 2467 2903
rect 2493 2903 2499 3036
rect 2509 2924 2515 2976
rect 2525 2944 2531 3016
rect 2570 3014 2582 3016
rect 2555 3006 2557 3014
rect 2565 3006 2567 3014
rect 2575 3006 2577 3014
rect 2585 3006 2587 3014
rect 2595 3006 2597 3014
rect 2570 3004 2582 3006
rect 2605 2904 2611 2936
rect 2493 2897 2515 2903
rect 2445 2883 2451 2897
rect 2413 2877 2451 2883
rect 2285 2837 2307 2843
rect 2253 2763 2259 2796
rect 2253 2757 2275 2763
rect 2189 2624 2195 2676
rect 2205 2584 2211 2696
rect 2221 2684 2227 2756
rect 2237 2704 2243 2716
rect 2157 2563 2163 2576
rect 2157 2557 2188 2563
rect 2141 2524 2147 2536
rect 2157 2524 2163 2557
rect 2125 2503 2131 2516
rect 2205 2504 2211 2516
rect 2125 2497 2147 2503
rect 2141 2383 2147 2497
rect 2237 2444 2243 2536
rect 2269 2504 2275 2757
rect 2285 2524 2291 2736
rect 2301 2704 2307 2837
rect 2317 2584 2323 2796
rect 2461 2784 2467 2796
rect 2333 2704 2339 2716
rect 2397 2704 2403 2776
rect 2356 2697 2371 2703
rect 2333 2544 2339 2696
rect 2365 2664 2371 2697
rect 2413 2683 2419 2696
rect 2381 2677 2419 2683
rect 2141 2377 2163 2383
rect 2141 2284 2147 2316
rect 2157 2304 2163 2377
rect 2173 2304 2179 2356
rect 2221 2304 2227 2436
rect 2237 2304 2243 2436
rect 2093 2217 2115 2223
rect 2093 2184 2099 2196
rect 2109 2124 2115 2217
rect 2125 2144 2131 2196
rect 2045 2004 2051 2116
rect 1997 1937 2019 1943
rect 1885 1844 1891 1896
rect 1949 1844 1955 1896
rect 1965 1884 1971 1896
rect 1981 1863 1987 1896
rect 1965 1857 1987 1863
rect 1885 1724 1891 1776
rect 1901 1604 1907 1716
rect 1917 1564 1923 1696
rect 1949 1664 1955 1816
rect 1949 1584 1955 1636
rect 1949 1504 1955 1516
rect 1885 1424 1891 1496
rect 1917 1464 1923 1496
rect 1869 1397 1891 1403
rect 1789 1364 1795 1376
rect 1693 1124 1699 1316
rect 1661 1104 1667 1116
rect 1693 1104 1699 1116
rect 1741 1104 1747 1316
rect 1757 1124 1763 1316
rect 1789 1244 1795 1316
rect 1837 1304 1843 1316
rect 1613 997 1651 1003
rect 1533 904 1539 916
rect 1581 883 1587 916
rect 1597 904 1603 916
rect 1613 903 1619 997
rect 1661 984 1667 1056
rect 1629 924 1635 976
rect 1613 897 1651 903
rect 1581 877 1628 883
rect 1469 704 1475 716
rect 1533 684 1539 856
rect 1581 724 1587 736
rect 1348 537 1363 543
rect 365 -23 387 -17
rect 477 -23 499 -17
rect 669 -23 691 -17
rect 781 -17 787 36
rect 1117 24 1123 36
rect 1066 14 1078 16
rect 1051 6 1053 14
rect 1061 6 1063 14
rect 1071 6 1073 14
rect 1081 6 1083 14
rect 1091 6 1093 14
rect 1066 4 1078 6
rect 781 -23 803 -17
rect 1133 -23 1139 36
rect 1165 -23 1171 16
rect 1229 -23 1235 516
rect 1245 304 1251 396
rect 1261 284 1267 516
rect 1293 444 1299 496
rect 1341 403 1347 516
rect 1325 397 1347 403
rect 1325 324 1331 397
rect 1341 304 1347 316
rect 1357 304 1363 537
rect 1357 284 1363 296
rect 1245 144 1251 236
rect 1293 124 1299 156
rect 1309 144 1315 236
rect 1373 184 1379 316
rect 1453 304 1459 536
rect 1485 526 1491 636
rect 1549 544 1555 696
rect 1581 624 1587 716
rect 1597 704 1603 716
rect 1645 684 1651 897
rect 1677 883 1683 956
rect 1693 884 1699 1076
rect 1773 1064 1779 1196
rect 1725 984 1731 1036
rect 1741 924 1747 976
rect 1757 964 1763 1036
rect 1773 924 1779 936
rect 1789 924 1795 1056
rect 1716 917 1731 923
rect 1725 903 1731 917
rect 1725 897 1788 903
rect 1668 877 1683 883
rect 1677 804 1683 836
rect 1693 704 1699 796
rect 1709 664 1715 676
rect 1597 544 1603 576
rect 1661 544 1667 636
rect 1709 543 1715 656
rect 1725 584 1731 676
rect 1741 604 1747 696
rect 1757 684 1763 756
rect 1773 624 1779 716
rect 1805 703 1811 1236
rect 1853 1144 1859 1236
rect 1821 963 1827 1136
rect 1837 1084 1843 1116
rect 1869 1104 1875 1356
rect 1885 1344 1891 1397
rect 1933 1384 1939 1476
rect 1965 1423 1971 1857
rect 1997 1824 2003 1937
rect 2045 1904 2051 1916
rect 2013 1804 2019 1856
rect 1981 1724 1987 1776
rect 2029 1724 2035 1876
rect 2061 1763 2067 1956
rect 2077 1784 2083 1876
rect 2045 1757 2067 1763
rect 2045 1724 2051 1757
rect 2093 1744 2099 2116
rect 2141 1984 2147 2276
rect 2157 2104 2163 2216
rect 2173 2204 2179 2296
rect 2205 2284 2211 2296
rect 2189 2277 2204 2283
rect 2189 2183 2195 2277
rect 2173 2177 2195 2183
rect 2173 2004 2179 2177
rect 2205 2124 2211 2216
rect 2221 2204 2227 2236
rect 2253 2144 2259 2296
rect 2269 2284 2275 2476
rect 2285 2304 2291 2316
rect 2301 2284 2307 2516
rect 2317 2444 2323 2476
rect 2109 1904 2115 1956
rect 2173 1924 2179 1976
rect 2205 1924 2211 2056
rect 2141 1884 2147 1896
rect 2125 1764 2131 1876
rect 2141 1744 2147 1776
rect 2013 1717 2028 1723
rect 1997 1703 2003 1716
rect 1981 1697 2003 1703
rect 1981 1664 1987 1697
rect 2013 1663 2019 1717
rect 1997 1657 2019 1663
rect 1997 1604 2003 1657
rect 2013 1604 2019 1636
rect 1997 1484 2003 1536
rect 2013 1524 2019 1536
rect 1956 1417 1971 1423
rect 1949 1384 1955 1416
rect 1885 1324 1891 1336
rect 1885 1124 1891 1136
rect 1869 963 1875 1076
rect 1885 1064 1891 1116
rect 1901 1084 1907 1236
rect 1917 1123 1923 1336
rect 1933 1324 1939 1336
rect 1917 1117 1939 1123
rect 1821 957 1843 963
rect 1837 944 1843 957
rect 1853 957 1875 963
rect 1853 944 1859 957
rect 1821 924 1827 936
rect 1853 924 1859 936
rect 1869 924 1875 936
rect 1901 924 1907 1036
rect 1933 963 1939 1117
rect 1949 1104 1955 1236
rect 1965 1104 1971 1316
rect 1981 1264 1987 1416
rect 1997 1344 2003 1376
rect 2013 1324 2019 1456
rect 1997 1264 2003 1316
rect 2029 1244 2035 1696
rect 2061 1664 2067 1736
rect 2045 1344 2051 1556
rect 2061 1344 2067 1376
rect 2077 1324 2083 1456
rect 2093 1324 2099 1736
rect 2157 1724 2163 1896
rect 2173 1884 2179 1916
rect 2221 1904 2227 2076
rect 2301 2064 2307 2256
rect 2317 2244 2323 2416
rect 2333 2304 2339 2536
rect 2349 2524 2355 2536
rect 2349 2283 2355 2356
rect 2365 2304 2371 2636
rect 2381 2564 2387 2677
rect 2381 2544 2387 2556
rect 2381 2484 2387 2536
rect 2397 2524 2403 2596
rect 2413 2424 2419 2616
rect 2429 2543 2435 2756
rect 2445 2664 2451 2696
rect 2477 2563 2483 2836
rect 2493 2784 2499 2796
rect 2493 2704 2499 2776
rect 2509 2744 2515 2897
rect 2573 2784 2579 2856
rect 2509 2604 2515 2716
rect 2525 2684 2531 2696
rect 2621 2644 2627 3097
rect 2637 3064 2643 3376
rect 2685 3304 2691 3416
rect 2797 3344 2803 3356
rect 2781 3324 2787 3336
rect 2845 3324 2851 3356
rect 2893 3324 2899 3336
rect 2685 3184 2691 3196
rect 2637 2964 2643 3036
rect 2653 2944 2659 3116
rect 2669 2964 2675 3136
rect 2685 3104 2691 3136
rect 2685 3044 2691 3096
rect 2637 2864 2643 2916
rect 2669 2904 2675 2936
rect 2653 2897 2668 2903
rect 2653 2783 2659 2897
rect 2685 2864 2691 3036
rect 2701 3004 2707 3076
rect 2717 3024 2723 3096
rect 2701 2924 2707 2956
rect 2717 2944 2723 2956
rect 2717 2903 2723 2916
rect 2701 2897 2723 2903
rect 2701 2884 2707 2897
rect 2644 2777 2659 2783
rect 2570 2614 2582 2616
rect 2555 2606 2557 2614
rect 2565 2606 2567 2614
rect 2575 2606 2577 2614
rect 2585 2606 2587 2614
rect 2595 2606 2597 2614
rect 2570 2604 2582 2606
rect 2461 2557 2483 2563
rect 2429 2537 2444 2543
rect 2461 2524 2467 2557
rect 2477 2537 2508 2543
rect 2477 2503 2483 2537
rect 2532 2517 2547 2523
rect 2429 2497 2483 2503
rect 2429 2484 2435 2497
rect 2509 2503 2515 2516
rect 2509 2497 2531 2503
rect 2445 2384 2451 2476
rect 2381 2304 2387 2356
rect 2340 2277 2355 2283
rect 2333 2204 2339 2276
rect 2381 2164 2387 2256
rect 2397 2224 2403 2236
rect 2429 2224 2435 2296
rect 2461 2244 2467 2476
rect 2493 2444 2499 2496
rect 2525 2484 2531 2497
rect 2477 2323 2483 2436
rect 2477 2317 2499 2323
rect 2477 2264 2483 2296
rect 2493 2284 2499 2317
rect 2493 2204 2499 2256
rect 2413 2184 2419 2196
rect 2445 2124 2451 2196
rect 2477 2103 2483 2196
rect 2509 2163 2515 2316
rect 2525 2304 2531 2436
rect 2541 2344 2547 2517
rect 2573 2484 2579 2516
rect 2589 2484 2595 2556
rect 2605 2524 2611 2556
rect 2621 2524 2627 2636
rect 2637 2564 2643 2616
rect 2653 2584 2659 2756
rect 2669 2564 2675 2616
rect 2685 2577 2723 2583
rect 2685 2543 2691 2577
rect 2717 2564 2723 2577
rect 2669 2537 2691 2543
rect 2669 2524 2675 2537
rect 2653 2444 2659 2476
rect 2541 2264 2547 2316
rect 2621 2224 2627 2296
rect 2525 2183 2531 2216
rect 2570 2214 2582 2216
rect 2555 2206 2557 2214
rect 2565 2206 2567 2214
rect 2575 2206 2577 2214
rect 2585 2206 2587 2214
rect 2595 2206 2597 2214
rect 2570 2204 2582 2206
rect 2525 2177 2547 2183
rect 2509 2157 2531 2163
rect 2493 2124 2499 2156
rect 2525 2144 2531 2157
rect 2477 2097 2524 2103
rect 2413 2077 2428 2083
rect 2173 1804 2179 1856
rect 2205 1824 2211 1896
rect 2237 1824 2243 1856
rect 2285 1844 2291 1916
rect 2301 1904 2307 1996
rect 2317 1964 2323 2056
rect 2317 1924 2323 1956
rect 2301 1824 2307 1896
rect 2317 1884 2323 1916
rect 2333 1904 2339 2076
rect 2413 1984 2419 2077
rect 2349 1844 2355 1896
rect 2365 1824 2371 1896
rect 2381 1864 2387 1956
rect 2429 1904 2435 1976
rect 2413 1883 2419 1896
rect 2461 1884 2467 2036
rect 2477 2004 2483 2076
rect 2493 1924 2499 2076
rect 2509 1884 2515 1976
rect 2541 1943 2547 2177
rect 2573 2137 2611 2143
rect 2573 2104 2579 2137
rect 2605 2124 2611 2137
rect 2637 2124 2643 2276
rect 2653 2264 2659 2296
rect 2653 2124 2659 2156
rect 2669 2144 2675 2496
rect 2685 2424 2691 2516
rect 2701 2504 2707 2556
rect 2717 2483 2723 2516
rect 2733 2484 2739 2516
rect 2701 2477 2723 2483
rect 2701 2303 2707 2477
rect 2717 2323 2723 2436
rect 2749 2324 2755 3276
rect 2765 3204 2771 3296
rect 2797 3144 2803 3316
rect 2797 3104 2803 3136
rect 2829 3104 2835 3136
rect 2909 3104 2915 3236
rect 2925 3143 2931 3376
rect 3469 3364 3475 3376
rect 3677 3364 3683 3463
rect 2941 3324 2947 3356
rect 3357 3344 3363 3356
rect 3677 3344 3683 3356
rect 3037 3324 3043 3336
rect 3133 3324 3139 3336
rect 3453 3324 3459 3336
rect 2973 3304 2979 3316
rect 2989 3284 2995 3316
rect 2925 3137 2947 3143
rect 2765 2924 2771 3096
rect 2781 3084 2787 3096
rect 2813 3083 2819 3096
rect 2829 3084 2835 3096
rect 2797 3077 2819 3083
rect 2797 2944 2803 3077
rect 2829 2944 2835 2956
rect 2781 2864 2787 2936
rect 2797 2924 2803 2936
rect 2820 2917 2835 2923
rect 2813 2904 2819 2916
rect 2765 2702 2771 2736
rect 2829 2684 2835 2917
rect 2845 2864 2851 2896
rect 2861 2864 2867 2936
rect 2877 2924 2883 3076
rect 2893 3024 2899 3096
rect 2925 3084 2931 3096
rect 2909 2964 2915 3076
rect 2941 2964 2947 3137
rect 3005 3124 3011 3236
rect 2957 3104 2963 3116
rect 2973 2944 2979 3076
rect 3021 3064 3027 3236
rect 2948 2937 2963 2943
rect 2957 2883 2963 2937
rect 3021 2924 3027 2996
rect 3053 2943 3059 3316
rect 3085 3284 3091 3316
rect 3069 2984 3075 3056
rect 3101 3023 3107 3236
rect 3085 3017 3107 3023
rect 3085 2964 3091 3017
rect 3044 2937 3059 2943
rect 3069 2937 3084 2943
rect 3037 2924 3043 2936
rect 2973 2904 2979 2916
rect 2957 2877 2979 2883
rect 2845 2724 2851 2756
rect 2909 2704 2915 2716
rect 2861 2564 2867 2696
rect 2909 2684 2915 2696
rect 2925 2684 2931 2716
rect 2941 2684 2947 2856
rect 2973 2844 2979 2877
rect 2989 2864 2995 2896
rect 3005 2844 3011 2916
rect 3053 2904 3059 2916
rect 3069 2904 3075 2937
rect 3117 2924 3123 3236
rect 3133 3124 3139 3316
rect 3293 3144 3299 3318
rect 3389 3304 3395 3316
rect 3229 3084 3235 3136
rect 3261 3104 3267 3116
rect 3133 2944 3139 3076
rect 3149 2924 3155 3056
rect 3165 2903 3171 3056
rect 3213 2924 3219 2956
rect 3229 2924 3235 2936
rect 3245 2904 3251 2936
rect 3277 2924 3283 3036
rect 3293 2944 3299 2956
rect 3149 2897 3171 2903
rect 2957 2784 2963 2836
rect 3021 2744 3027 2836
rect 3053 2744 3059 2896
rect 3069 2864 3075 2896
rect 2957 2704 2963 2716
rect 2989 2704 2995 2736
rect 3069 2724 3075 2856
rect 3101 2784 3107 2836
rect 3085 2763 3091 2776
rect 3085 2757 3107 2763
rect 3101 2744 3107 2757
rect 3021 2717 3036 2723
rect 3021 2704 3027 2717
rect 3044 2697 3059 2703
rect 2941 2537 2956 2543
rect 2925 2524 2931 2536
rect 2717 2317 2739 2323
rect 2685 2297 2707 2303
rect 2525 1937 2547 1943
rect 2413 1877 2435 1883
rect 2429 1823 2435 1877
rect 2445 1844 2451 1876
rect 2429 1817 2451 1823
rect 2173 1704 2179 1716
rect 2109 1303 2115 1636
rect 2173 1604 2179 1696
rect 2125 1504 2131 1576
rect 2173 1484 2179 1576
rect 2205 1504 2211 1736
rect 2237 1623 2243 1736
rect 2221 1617 2243 1623
rect 2221 1544 2227 1617
rect 2237 1584 2243 1596
rect 2237 1524 2243 1576
rect 2253 1524 2259 1656
rect 2285 1504 2291 1776
rect 2349 1743 2355 1816
rect 2445 1744 2451 1817
rect 2477 1784 2483 1876
rect 2493 1804 2499 1876
rect 2525 1783 2531 1937
rect 2557 1904 2563 1996
rect 2589 1844 2595 2116
rect 2669 2103 2675 2116
rect 2653 2097 2675 2103
rect 2637 2004 2643 2036
rect 2621 1917 2636 1923
rect 2570 1814 2582 1816
rect 2555 1806 2557 1814
rect 2565 1806 2567 1814
rect 2575 1806 2577 1814
rect 2585 1806 2587 1814
rect 2595 1806 2597 1814
rect 2570 1804 2582 1806
rect 2525 1777 2547 1783
rect 2509 1744 2515 1776
rect 2541 1744 2547 1777
rect 2557 1744 2563 1776
rect 2349 1737 2371 1743
rect 2317 1704 2323 1736
rect 2349 1644 2355 1716
rect 2093 1297 2115 1303
rect 2141 1337 2172 1343
rect 2045 1263 2051 1276
rect 2093 1264 2099 1297
rect 2045 1257 2067 1263
rect 2013 1124 2019 1236
rect 2045 1104 2051 1236
rect 2061 1144 2067 1257
rect 2029 1023 2035 1076
rect 2013 1017 2035 1023
rect 1917 957 1939 963
rect 1805 697 1820 703
rect 1917 684 1923 957
rect 1949 924 1955 956
rect 1965 924 1971 1016
rect 1981 944 1987 956
rect 1933 904 1939 916
rect 1837 664 1843 676
rect 1789 544 1795 636
rect 1709 537 1724 543
rect 1837 543 1843 656
rect 1853 564 1859 636
rect 1837 537 1852 543
rect 1613 524 1619 536
rect 1517 302 1523 516
rect 1549 464 1555 496
rect 1405 243 1411 256
rect 1396 237 1411 243
rect 1357 124 1363 176
rect 1405 124 1411 237
rect 1549 164 1555 276
rect 1581 264 1587 316
rect 1597 244 1603 516
rect 1613 384 1619 496
rect 1613 304 1619 316
rect 1629 304 1635 536
rect 1885 524 1891 656
rect 1965 644 1971 716
rect 2013 684 2019 1017
rect 2045 944 2051 1096
rect 2093 1044 2099 1256
rect 2109 1204 2115 1276
rect 2141 1144 2147 1337
rect 2189 1324 2195 1356
rect 2164 1317 2179 1323
rect 2061 924 2067 1016
rect 2093 944 2099 956
rect 2029 743 2035 836
rect 2029 737 2051 743
rect 2045 724 2051 737
rect 2093 684 2099 796
rect 2109 724 2115 976
rect 2141 964 2147 1036
rect 2157 1024 2163 1116
rect 2173 1104 2179 1317
rect 2189 1204 2195 1236
rect 2205 1144 2211 1496
rect 2253 1383 2259 1456
rect 2269 1404 2275 1436
rect 2285 1384 2291 1456
rect 2253 1377 2275 1383
rect 2221 1204 2227 1296
rect 2157 924 2163 936
rect 2173 804 2179 1076
rect 2189 1064 2195 1076
rect 2205 844 2211 1036
rect 2221 964 2227 1096
rect 2237 1064 2243 1076
rect 2269 1064 2275 1377
rect 2285 1264 2291 1316
rect 2301 1284 2307 1496
rect 2317 1364 2323 1576
rect 2333 1524 2339 1536
rect 2365 1383 2371 1737
rect 2397 1604 2403 1636
rect 2413 1584 2419 1736
rect 2445 1683 2451 1736
rect 2493 1724 2499 1736
rect 2532 1717 2547 1723
rect 2429 1677 2467 1683
rect 2429 1644 2435 1677
rect 2429 1504 2435 1596
rect 2445 1463 2451 1636
rect 2461 1604 2467 1677
rect 2461 1504 2467 1576
rect 2493 1504 2499 1596
rect 2541 1584 2547 1717
rect 2557 1524 2563 1716
rect 2573 1644 2579 1736
rect 2589 1664 2595 1736
rect 2621 1684 2627 1917
rect 2653 1904 2659 2097
rect 2685 2083 2691 2297
rect 2733 2284 2739 2317
rect 2749 2284 2755 2296
rect 2701 2084 2707 2236
rect 2717 2124 2723 2136
rect 2765 2124 2771 2416
rect 2797 2304 2803 2516
rect 2861 2484 2867 2518
rect 2941 2484 2947 2537
rect 2957 2504 2963 2516
rect 2845 2424 2851 2476
rect 2813 2304 2819 2316
rect 2797 2284 2803 2296
rect 2781 2144 2787 2156
rect 2813 2144 2819 2276
rect 2829 2224 2835 2336
rect 2845 2284 2851 2316
rect 2861 2244 2867 2276
rect 2877 2244 2883 2296
rect 2925 2284 2931 2316
rect 2973 2304 2979 2636
rect 3005 2524 3011 2676
rect 3021 2604 3027 2676
rect 3053 2664 3059 2697
rect 3069 2683 3075 2716
rect 3085 2704 3091 2736
rect 3092 2697 3107 2703
rect 3069 2677 3091 2683
rect 3037 2604 3043 2656
rect 3069 2584 3075 2656
rect 3085 2584 3091 2677
rect 3021 2503 3027 2536
rect 3021 2497 3043 2503
rect 2877 2144 2883 2216
rect 2893 2204 2899 2276
rect 2989 2263 2995 2316
rect 3005 2284 3011 2476
rect 3021 2304 3027 2416
rect 3037 2384 3043 2497
rect 3053 2424 3059 2496
rect 3101 2444 3107 2697
rect 3117 2664 3123 2776
rect 3133 2724 3139 2836
rect 3149 2704 3155 2897
rect 3133 2644 3139 2696
rect 3165 2664 3171 2776
rect 3181 2684 3187 2716
rect 3229 2704 3235 2896
rect 3133 2544 3139 2576
rect 3197 2524 3203 2696
rect 3245 2684 3251 2896
rect 3261 2684 3267 2716
rect 3293 2704 3299 2916
rect 3309 2744 3315 3096
rect 3325 3084 3331 3176
rect 3341 3084 3347 3276
rect 3389 3264 3395 3296
rect 3373 3104 3379 3116
rect 3325 2924 3331 3036
rect 3341 2844 3347 3016
rect 3373 2924 3379 3016
rect 3389 2864 3395 3256
rect 3405 3104 3411 3136
rect 3437 3084 3443 3136
rect 3453 3084 3459 3316
rect 3533 3104 3539 3316
rect 3581 3284 3587 3316
rect 3581 3084 3587 3094
rect 3421 2924 3427 3036
rect 3469 2924 3475 3016
rect 3501 2984 3507 2996
rect 3613 2944 3619 3076
rect 3645 3044 3651 3076
rect 3661 2964 3667 3316
rect 3789 3144 3795 3336
rect 3821 3304 3827 3318
rect 3885 3284 3891 3356
rect 3677 3104 3683 3116
rect 3725 3063 3731 3096
rect 3741 3084 3747 3136
rect 3949 3124 3955 3463
rect 3981 3324 3987 3396
rect 4301 3364 4307 3376
rect 3981 3304 3987 3316
rect 3949 3084 3955 3116
rect 3965 3104 3971 3256
rect 3981 3144 3987 3276
rect 3997 3264 4003 3316
rect 4109 3304 4115 3336
rect 4237 3324 4243 3336
rect 4125 3264 4131 3316
rect 3997 3224 4003 3236
rect 4074 3214 4086 3216
rect 4059 3206 4061 3214
rect 4069 3206 4071 3214
rect 4079 3206 4081 3214
rect 4089 3206 4091 3214
rect 4099 3206 4101 3214
rect 4074 3204 4086 3206
rect 3997 3184 4003 3196
rect 3725 3057 3747 3063
rect 3341 2783 3347 2836
rect 3332 2777 3347 2783
rect 3117 2444 3123 2516
rect 3213 2384 3219 2676
rect 3245 2664 3251 2676
rect 3309 2644 3315 2676
rect 3373 2524 3379 2536
rect 3085 2304 3091 2336
rect 3181 2304 3187 2336
rect 3037 2284 3043 2296
rect 2973 2257 2995 2263
rect 2893 2164 2899 2176
rect 2669 2077 2691 2083
rect 2669 1963 2675 2077
rect 2685 2003 2691 2036
rect 2733 2004 2739 2036
rect 2685 1997 2707 2003
rect 2669 1957 2691 1963
rect 2637 1824 2643 1836
rect 2653 1804 2659 1896
rect 2669 1884 2675 1936
rect 2685 1903 2691 1957
rect 2701 1924 2707 1997
rect 2685 1897 2707 1903
rect 2637 1764 2643 1776
rect 2653 1743 2659 1796
rect 2701 1763 2707 1897
rect 2717 1764 2723 1996
rect 2749 1924 2755 2016
rect 2749 1824 2755 1896
rect 2637 1737 2659 1743
rect 2685 1757 2707 1763
rect 2637 1724 2643 1737
rect 2669 1684 2675 1716
rect 2685 1663 2691 1757
rect 2669 1657 2691 1663
rect 2589 1524 2595 1536
rect 2605 1464 2611 1656
rect 2669 1623 2675 1657
rect 2660 1617 2675 1623
rect 2445 1457 2467 1463
rect 2365 1377 2387 1383
rect 2381 1324 2387 1377
rect 2420 1377 2428 1383
rect 2301 1103 2307 1256
rect 2317 1104 2323 1276
rect 2333 1104 2339 1116
rect 2292 1097 2307 1103
rect 2285 1064 2291 1076
rect 2237 963 2243 1056
rect 2253 984 2259 1036
rect 2237 957 2252 963
rect 2285 924 2291 1016
rect 2301 944 2307 956
rect 2301 924 2307 936
rect 2237 844 2243 916
rect 2253 717 2291 723
rect 2157 704 2163 716
rect 2253 703 2259 717
rect 2285 704 2291 717
rect 2244 697 2259 703
rect 2109 684 2115 696
rect 2173 684 2179 696
rect 2269 684 2275 696
rect 2301 684 2307 836
rect 2317 784 2323 1056
rect 2333 943 2339 1056
rect 2333 937 2355 943
rect 2333 904 2339 916
rect 2349 883 2355 937
rect 2381 924 2387 1216
rect 2445 1183 2451 1436
rect 2461 1324 2467 1457
rect 2493 1384 2499 1416
rect 2509 1404 2515 1436
rect 2477 1344 2483 1376
rect 2509 1323 2515 1396
rect 2500 1317 2515 1323
rect 2525 1304 2531 1436
rect 2570 1414 2582 1416
rect 2555 1406 2557 1414
rect 2565 1406 2567 1414
rect 2575 1406 2577 1414
rect 2585 1406 2587 1414
rect 2595 1406 2597 1414
rect 2570 1404 2582 1406
rect 2461 1204 2467 1296
rect 2525 1264 2531 1296
rect 2589 1284 2595 1336
rect 2605 1284 2611 1336
rect 2429 1177 2451 1183
rect 2397 984 2403 1116
rect 2429 1104 2435 1177
rect 2461 1163 2467 1176
rect 2445 1157 2467 1163
rect 2413 1084 2419 1096
rect 2445 1083 2451 1157
rect 2477 1143 2483 1196
rect 2461 1137 2483 1143
rect 2461 1124 2467 1137
rect 2621 1084 2627 1576
rect 2653 1504 2659 1616
rect 2685 1603 2691 1636
rect 2701 1624 2707 1696
rect 2685 1597 2707 1603
rect 2701 1544 2707 1597
rect 2749 1504 2755 1776
rect 2765 1764 2771 2116
rect 2813 2004 2819 2096
rect 2829 2024 2835 2136
rect 2781 1844 2787 1996
rect 2845 1964 2851 2096
rect 2877 2024 2883 2116
rect 2909 2003 2915 2216
rect 2877 1997 2915 2003
rect 2877 1984 2883 1997
rect 2765 1504 2771 1516
rect 2637 1324 2643 1456
rect 2653 1364 2659 1476
rect 2669 1444 2675 1496
rect 2669 1343 2675 1396
rect 2781 1384 2787 1836
rect 2797 1824 2803 1896
rect 2813 1744 2819 1856
rect 2845 1844 2851 1876
rect 2797 1584 2803 1716
rect 2813 1584 2819 1736
rect 2845 1704 2851 1796
rect 2877 1744 2883 1836
rect 2893 1724 2899 1976
rect 2925 1904 2931 1916
rect 2973 1904 2979 2257
rect 2989 2044 2995 2236
rect 3005 2104 3011 2116
rect 3021 2104 3027 2276
rect 3085 2124 3091 2156
rect 3101 2124 3107 2156
rect 3117 2104 3123 2296
rect 3133 2284 3139 2296
rect 3165 2124 3171 2236
rect 3197 2124 3203 2156
rect 3229 2123 3235 2236
rect 3245 2143 3251 2296
rect 3261 2244 3267 2256
rect 3245 2137 3267 2143
rect 3229 2117 3244 2123
rect 3181 2104 3187 2116
rect 2989 1984 2995 1996
rect 3021 1904 3027 2036
rect 3069 1904 3075 1936
rect 2909 1784 2915 1896
rect 2925 1824 2931 1836
rect 2925 1743 2931 1796
rect 2941 1784 2947 1796
rect 2957 1784 2963 1896
rect 2973 1884 2979 1896
rect 3085 1884 3091 1976
rect 2909 1737 2931 1743
rect 2893 1684 2899 1716
rect 2829 1504 2835 1616
rect 2845 1504 2851 1676
rect 2660 1337 2675 1343
rect 2685 1324 2691 1376
rect 2717 1344 2723 1376
rect 2653 1124 2659 1316
rect 2436 1077 2451 1083
rect 2413 964 2419 976
rect 2333 877 2355 883
rect 2333 784 2339 877
rect 2349 724 2355 856
rect 2397 804 2403 936
rect 1661 384 1667 496
rect 1677 464 1683 496
rect 1725 404 1731 516
rect 1741 444 1747 496
rect 1805 464 1811 496
rect 1629 284 1635 296
rect 1693 184 1699 316
rect 1773 304 1779 396
rect 1853 344 1859 516
rect 1869 324 1875 516
rect 1901 323 1907 556
rect 1981 544 1987 556
rect 1917 524 1923 536
rect 1965 524 1971 536
rect 1917 384 1923 476
rect 1901 317 1916 323
rect 1917 304 1923 316
rect 1949 304 1955 516
rect 1997 504 2003 616
rect 2013 463 2019 676
rect 2029 524 2035 636
rect 2093 624 2099 676
rect 2045 544 2051 576
rect 2013 457 2035 463
rect 2013 304 2019 316
rect 1549 126 1555 136
rect 1725 124 1731 276
rect 1949 264 1955 276
rect 1965 264 1971 296
rect 1821 124 1827 136
rect 1853 124 1859 256
rect 1901 184 1907 256
rect 1549 117 1555 118
rect 1245 44 1251 116
rect 1965 84 1971 116
rect 2013 104 2019 276
rect 2029 164 2035 457
rect 2045 404 2051 516
rect 2061 504 2067 516
rect 2077 504 2083 616
rect 2109 544 2115 616
rect 2173 544 2179 576
rect 2093 304 2099 536
rect 2189 524 2195 536
rect 2157 404 2163 516
rect 2205 504 2211 596
rect 2301 584 2307 656
rect 2221 524 2227 556
rect 2237 544 2243 576
rect 2317 564 2323 696
rect 2349 684 2355 716
rect 2381 703 2387 776
rect 2397 704 2403 716
rect 2372 697 2387 703
rect 2429 684 2435 1076
rect 2445 944 2451 996
rect 2477 823 2483 1056
rect 2570 1014 2582 1016
rect 2555 1006 2557 1014
rect 2565 1006 2567 1014
rect 2575 1006 2577 1014
rect 2585 1006 2587 1014
rect 2595 1006 2597 1014
rect 2570 1004 2582 1006
rect 2621 944 2627 996
rect 2637 984 2643 1116
rect 2653 1044 2659 1076
rect 2669 944 2675 1316
rect 2701 1124 2707 1336
rect 2797 1324 2803 1476
rect 2813 1404 2819 1476
rect 2797 1304 2803 1316
rect 2740 1277 2755 1283
rect 2701 944 2707 1056
rect 2717 984 2723 1116
rect 2749 1104 2755 1277
rect 2781 1184 2787 1276
rect 2733 1044 2739 1056
rect 2525 904 2531 916
rect 2468 817 2483 823
rect 2493 724 2499 856
rect 2541 723 2547 936
rect 2525 717 2547 723
rect 2477 704 2483 716
rect 2253 464 2259 536
rect 2365 524 2371 636
rect 2381 544 2387 676
rect 2484 637 2499 643
rect 2397 564 2403 576
rect 2493 563 2499 637
rect 2509 584 2515 696
rect 2477 557 2499 563
rect 2141 304 2147 316
rect 2100 297 2115 303
rect 2061 264 2067 296
rect 2077 184 2083 296
rect 2093 144 2099 256
rect 2029 126 2035 136
rect 2029 117 2035 118
rect 1325 -17 1331 36
rect 1373 -17 1379 36
rect 1613 -17 1619 36
rect 1885 -17 1891 36
rect 1325 -23 1347 -17
rect 1373 -23 1395 -17
rect 1613 -23 1635 -17
rect 1869 -23 1891 -17
rect 2109 -23 2115 297
rect 2157 284 2163 296
rect 2173 124 2179 436
rect 2221 324 2227 456
rect 2317 384 2323 516
rect 2333 464 2339 496
rect 2333 344 2339 456
rect 2365 304 2371 516
rect 2381 384 2387 536
rect 2445 524 2451 536
rect 2429 304 2435 516
rect 2461 384 2467 476
rect 2189 244 2195 296
rect 2301 284 2307 296
rect 2189 144 2195 196
rect 2205 144 2211 256
rect 2269 124 2275 276
rect 2125 104 2131 116
rect 2221 104 2227 116
rect 2253 104 2259 116
rect 2285 104 2291 256
rect 2349 164 2355 296
rect 2429 263 2435 296
rect 2445 284 2451 296
rect 2429 257 2451 263
rect 2365 184 2371 196
rect 2381 184 2387 256
rect 2365 143 2371 176
rect 2381 164 2387 176
rect 2356 137 2371 143
rect 2333 124 2339 136
rect 2349 84 2355 96
rect 2413 84 2419 136
rect 2445 104 2451 257
rect 2477 124 2483 557
rect 2525 544 2531 717
rect 2557 684 2563 836
rect 2573 704 2579 716
rect 2589 684 2595 696
rect 2605 683 2611 936
rect 2749 924 2755 1096
rect 2797 924 2803 1296
rect 2813 1283 2819 1396
rect 2829 1344 2835 1376
rect 2829 1304 2835 1336
rect 2845 1324 2851 1496
rect 2861 1444 2867 1676
rect 2909 1524 2915 1737
rect 2973 1724 2979 1856
rect 3053 1726 3059 1796
rect 2925 1644 2931 1676
rect 2925 1503 2931 1636
rect 3021 1564 3027 1636
rect 2957 1543 2963 1556
rect 2941 1537 2963 1543
rect 2941 1504 2947 1537
rect 2909 1497 2931 1503
rect 2877 1404 2883 1436
rect 2893 1424 2899 1496
rect 2909 1464 2915 1497
rect 2925 1424 2931 1476
rect 2877 1364 2883 1396
rect 2893 1324 2899 1416
rect 2925 1364 2931 1396
rect 2941 1344 2947 1476
rect 2957 1424 2963 1516
rect 3005 1484 3011 1516
rect 2957 1324 2963 1396
rect 2973 1344 2979 1416
rect 2989 1324 2995 1476
rect 3021 1324 3027 1556
rect 3037 1364 3043 1556
rect 3085 1523 3091 1876
rect 3101 1704 3107 2096
rect 3261 1984 3267 2137
rect 3172 1917 3187 1923
rect 3117 1904 3123 1916
rect 3181 1904 3187 1917
rect 3117 1704 3123 1716
rect 3117 1584 3123 1696
rect 3149 1603 3155 1876
rect 3165 1784 3171 1896
rect 3277 1844 3283 2056
rect 3293 1844 3299 1876
rect 3165 1637 3180 1643
rect 3165 1624 3171 1637
rect 3149 1597 3171 1603
rect 3108 1537 3139 1543
rect 3085 1517 3123 1523
rect 3069 1484 3075 1516
rect 3085 1504 3091 1517
rect 3053 1384 3059 1476
rect 2845 1284 2851 1316
rect 3005 1303 3011 1316
rect 3069 1304 3075 1476
rect 3101 1324 3107 1496
rect 3117 1484 3123 1517
rect 3133 1484 3139 1537
rect 3149 1504 3155 1576
rect 3117 1344 3123 1396
rect 3133 1364 3139 1396
rect 3165 1383 3171 1597
rect 3197 1503 3203 1796
rect 3293 1744 3299 1836
rect 3309 1744 3315 1876
rect 3229 1644 3235 1716
rect 3325 1704 3331 1856
rect 3357 1843 3363 2436
rect 3389 2284 3395 2696
rect 3405 2524 3411 2736
rect 3421 2544 3427 2856
rect 3437 2724 3443 2836
rect 3517 2724 3523 2836
rect 3453 2702 3459 2716
rect 3565 2704 3571 2816
rect 3581 2784 3587 2816
rect 3405 2504 3411 2516
rect 3421 2404 3427 2536
rect 3501 2524 3507 2616
rect 3517 2544 3523 2656
rect 3549 2644 3555 2696
rect 3565 2664 3571 2676
rect 3533 2564 3539 2616
rect 3549 2584 3555 2636
rect 3533 2504 3539 2556
rect 3565 2504 3571 2656
rect 3581 2644 3587 2716
rect 3597 2704 3603 2716
rect 3613 2704 3619 2836
rect 3613 2544 3619 2696
rect 3629 2684 3635 2956
rect 3693 2944 3699 2996
rect 3645 2684 3651 2696
rect 3661 2544 3667 2936
rect 3741 2724 3747 3057
rect 3757 2984 3763 3036
rect 3789 2944 3795 2956
rect 3821 2944 3827 3076
rect 3917 2944 3923 3076
rect 3789 2904 3795 2916
rect 3789 2764 3795 2896
rect 3949 2864 3955 2936
rect 3837 2824 3843 2836
rect 3677 2684 3683 2716
rect 3725 2684 3731 2696
rect 3741 2684 3747 2696
rect 3693 2603 3699 2636
rect 3741 2604 3747 2656
rect 3789 2604 3795 2696
rect 3677 2597 3699 2603
rect 3677 2526 3683 2597
rect 3741 2584 3747 2596
rect 3709 2504 3715 2536
rect 3540 2497 3555 2503
rect 3469 2484 3475 2496
rect 3453 2284 3459 2376
rect 3469 2304 3475 2436
rect 3389 2144 3395 2276
rect 3469 2163 3475 2296
rect 3517 2264 3523 2316
rect 3549 2304 3555 2497
rect 3565 2284 3571 2396
rect 3613 2384 3619 2496
rect 3469 2157 3491 2163
rect 3485 2124 3491 2157
rect 3501 2144 3507 2216
rect 3565 2143 3571 2276
rect 3581 2163 3587 2296
rect 3597 2184 3603 2196
rect 3581 2157 3603 2163
rect 3565 2137 3580 2143
rect 3405 2104 3411 2118
rect 3492 2117 3507 2123
rect 3389 1984 3395 2076
rect 3389 1904 3395 1976
rect 3437 1904 3443 2036
rect 3357 1837 3379 1843
rect 3357 1784 3363 1816
rect 3341 1724 3347 1736
rect 3213 1584 3219 1636
rect 3245 1504 3251 1636
rect 3188 1497 3203 1503
rect 3181 1424 3187 1436
rect 3149 1377 3171 1383
rect 3005 1297 3027 1303
rect 2813 1277 2835 1283
rect 2813 1104 2819 1256
rect 2829 1184 2835 1277
rect 2813 1084 2819 1096
rect 2669 804 2675 896
rect 2685 783 2691 796
rect 2644 777 2691 783
rect 2621 704 2627 756
rect 2669 684 2675 716
rect 2605 677 2627 683
rect 2570 614 2582 616
rect 2555 606 2557 614
rect 2565 606 2567 614
rect 2575 606 2577 614
rect 2585 606 2587 614
rect 2595 606 2597 614
rect 2570 604 2582 606
rect 2621 584 2627 677
rect 2637 584 2643 676
rect 2685 664 2691 716
rect 2717 704 2723 836
rect 2701 684 2707 696
rect 2733 684 2739 816
rect 2765 804 2771 836
rect 2781 804 2787 916
rect 2813 904 2819 936
rect 2829 924 2835 1036
rect 2845 963 2851 1236
rect 2861 1124 2867 1256
rect 2877 1104 2883 1296
rect 2989 1204 2995 1296
rect 3021 1284 3027 1297
rect 3133 1204 3139 1276
rect 2893 1104 2899 1116
rect 3005 1104 3011 1136
rect 3037 1104 3043 1196
rect 3069 1104 3075 1116
rect 3117 1104 3123 1116
rect 3133 1104 3139 1196
rect 3149 1184 3155 1377
rect 3165 1324 3171 1356
rect 3181 1344 3187 1376
rect 3213 1364 3219 1496
rect 3261 1484 3267 1576
rect 3293 1544 3299 1636
rect 3325 1584 3331 1696
rect 3373 1564 3379 1837
rect 3389 1724 3395 1816
rect 3421 1784 3427 1836
rect 3437 1724 3443 1736
rect 3453 1723 3459 1996
rect 3469 1784 3475 1796
rect 3485 1764 3491 1896
rect 3501 1864 3507 2117
rect 3533 2064 3539 2076
rect 3565 2064 3571 2116
rect 3565 1944 3571 2016
rect 3581 1984 3587 2136
rect 3597 1964 3603 2157
rect 3565 1924 3571 1936
rect 3533 1884 3539 1896
rect 3533 1824 3539 1876
rect 3444 1717 3459 1723
rect 3501 1723 3507 1816
rect 3613 1804 3619 2216
rect 3645 2184 3651 2196
rect 3645 2164 3651 2176
rect 3661 2164 3667 2316
rect 3709 2304 3715 2496
rect 3805 2444 3811 2696
rect 3821 2677 3836 2683
rect 3821 2404 3827 2677
rect 3853 2624 3859 2656
rect 3885 2624 3891 2696
rect 3837 2504 3843 2536
rect 3869 2526 3875 2556
rect 3901 2483 3907 2756
rect 3917 2744 3923 2816
rect 3965 2784 3971 2918
rect 3933 2584 3939 2736
rect 3997 2704 4003 3136
rect 4077 3124 4083 3136
rect 4029 2984 4035 3096
rect 4157 2944 4163 3136
rect 4173 3004 4179 3276
rect 4253 3143 4259 3276
rect 4349 3224 4355 3316
rect 4253 3137 4275 3143
rect 4269 3124 4275 3137
rect 4205 3102 4211 3103
rect 4029 2783 4035 2896
rect 4061 2844 4067 2916
rect 4077 2884 4083 2936
rect 4077 2844 4083 2876
rect 4189 2864 4195 3076
rect 4205 2984 4211 3094
rect 4237 2924 4243 2936
rect 4269 2904 4275 2916
rect 4205 2884 4211 2896
rect 4228 2837 4243 2843
rect 4074 2814 4086 2816
rect 4059 2806 4061 2814
rect 4069 2806 4071 2814
rect 4079 2806 4081 2814
rect 4089 2806 4091 2814
rect 4099 2806 4101 2814
rect 4074 2804 4086 2806
rect 4029 2777 4051 2783
rect 3997 2664 4003 2676
rect 3901 2477 3923 2483
rect 3901 2324 3907 2436
rect 3917 2384 3923 2477
rect 4029 2324 4035 2716
rect 4045 2704 4051 2777
rect 4141 2704 4147 2716
rect 4157 2684 4163 2836
rect 4173 2684 4179 2736
rect 4205 2724 4211 2756
rect 4045 2564 4051 2636
rect 4189 2563 4195 2636
rect 4173 2557 4195 2563
rect 4093 2544 4099 2556
rect 4061 2504 4067 2518
rect 4173 2504 4179 2557
rect 4189 2504 4195 2536
rect 4205 2523 4211 2716
rect 4237 2544 4243 2837
rect 4269 2764 4275 2896
rect 4285 2724 4291 3116
rect 4301 3104 4307 3116
rect 4317 3104 4323 3216
rect 4349 3144 4355 3156
rect 4477 3144 4483 3416
rect 4557 3404 4563 3463
rect 4653 3457 4675 3463
rect 4349 3064 4355 3136
rect 4365 2963 4371 2976
rect 4356 2957 4371 2963
rect 4349 2944 4355 2956
rect 4324 2937 4339 2943
rect 4333 2923 4339 2937
rect 4333 2917 4348 2923
rect 4301 2704 4307 2876
rect 4253 2624 4259 2696
rect 4269 2644 4275 2676
rect 4317 2624 4323 2696
rect 4349 2684 4355 2856
rect 4333 2644 4339 2676
rect 4285 2564 4291 2576
rect 4205 2517 4220 2523
rect 4253 2424 4259 2436
rect 4269 2424 4275 2536
rect 4285 2464 4291 2556
rect 4074 2414 4086 2416
rect 4059 2406 4061 2414
rect 4069 2406 4071 2414
rect 4079 2406 4081 2414
rect 4089 2406 4091 2414
rect 4099 2406 4101 2414
rect 4074 2404 4086 2406
rect 4125 2384 4131 2416
rect 3981 2317 3996 2323
rect 3757 2302 3763 2316
rect 3709 2124 3715 2296
rect 3821 2244 3827 2256
rect 3837 2144 3843 2196
rect 3869 2124 3875 2296
rect 3949 2223 3955 2296
rect 3965 2264 3971 2276
rect 3965 2223 3971 2236
rect 3949 2217 3971 2223
rect 3933 2144 3939 2156
rect 3629 2044 3635 2116
rect 3773 2104 3779 2118
rect 3885 2104 3891 2136
rect 3869 2024 3875 2096
rect 3629 1904 3635 2016
rect 3645 1904 3651 1936
rect 3629 1844 3635 1876
rect 3533 1724 3539 1796
rect 3581 1724 3587 1736
rect 3613 1724 3619 1796
rect 3677 1744 3683 1976
rect 3757 1884 3763 1896
rect 3837 1864 3843 1876
rect 3773 1784 3779 1856
rect 3677 1724 3683 1736
rect 3709 1724 3715 1756
rect 3492 1717 3507 1723
rect 3309 1523 3315 1536
rect 3300 1517 3315 1523
rect 3245 1444 3251 1456
rect 3245 1324 3251 1336
rect 3172 1317 3187 1323
rect 3181 1204 3187 1317
rect 3197 1284 3203 1316
rect 3229 1264 3235 1316
rect 3245 1303 3251 1316
rect 3245 1297 3260 1303
rect 3277 1284 3283 1376
rect 3293 1324 3299 1516
rect 3309 1424 3315 1496
rect 3341 1484 3347 1556
rect 3373 1504 3379 1516
rect 3405 1483 3411 1716
rect 3517 1704 3523 1716
rect 3693 1704 3699 1716
rect 3533 1697 3548 1703
rect 3421 1503 3427 1636
rect 3437 1523 3443 1536
rect 3437 1517 3459 1523
rect 3453 1504 3459 1517
rect 3421 1497 3436 1503
rect 3396 1477 3411 1483
rect 3325 1463 3331 1476
rect 3325 1457 3347 1463
rect 3341 1303 3347 1457
rect 3373 1344 3379 1476
rect 3389 1344 3395 1476
rect 3405 1444 3411 1456
rect 3357 1324 3363 1336
rect 3332 1297 3347 1303
rect 2861 1064 2867 1096
rect 2957 1084 2963 1096
rect 2973 1084 2979 1096
rect 2957 1004 2963 1056
rect 2845 957 2867 963
rect 2861 924 2867 957
rect 2916 937 2947 943
rect 2797 843 2803 896
rect 2813 864 2819 896
rect 2893 864 2899 916
rect 2941 903 2947 937
rect 2957 924 2963 996
rect 2941 897 2956 903
rect 2909 877 2947 883
rect 2909 843 2915 877
rect 2941 844 2947 877
rect 2797 837 2915 843
rect 2973 824 2979 1076
rect 3053 1044 3059 1076
rect 3069 1064 3075 1076
rect 3005 903 3011 936
rect 3021 924 3027 996
rect 3085 924 3091 1056
rect 3101 1044 3107 1076
rect 3165 1064 3171 1176
rect 3245 1124 3251 1136
rect 3197 1104 3203 1116
rect 3229 1104 3235 1116
rect 3293 1104 3299 1236
rect 3325 1184 3331 1296
rect 3341 1184 3347 1276
rect 3389 1203 3395 1316
rect 3405 1284 3411 1436
rect 3437 1383 3443 1496
rect 3453 1444 3459 1476
rect 3437 1377 3459 1383
rect 3437 1344 3443 1356
rect 3453 1324 3459 1377
rect 3437 1303 3443 1316
rect 3437 1297 3459 1303
rect 3453 1284 3459 1297
rect 3373 1197 3395 1203
rect 3101 904 3107 956
rect 3117 924 3123 1036
rect 3165 963 3171 1056
rect 3181 1044 3187 1076
rect 3165 957 3180 963
rect 3213 943 3219 1076
rect 3261 944 3267 1096
rect 3204 937 3219 943
rect 2996 897 3011 903
rect 3133 864 3139 936
rect 3149 924 3155 936
rect 3245 924 3251 936
rect 3277 924 3283 1096
rect 2749 783 2755 796
rect 2749 777 2803 783
rect 2797 764 2803 777
rect 2916 757 2947 763
rect 2765 703 2771 716
rect 2756 697 2771 703
rect 2781 684 2787 756
rect 2941 724 2947 757
rect 2909 702 2915 703
rect 2653 604 2659 656
rect 2669 564 2675 636
rect 2605 544 2611 556
rect 2493 464 2499 496
rect 2509 304 2515 516
rect 2541 424 2547 536
rect 2573 344 2579 476
rect 2637 464 2643 496
rect 2653 484 2659 536
rect 2493 164 2499 296
rect 2509 204 2515 296
rect 2573 284 2579 336
rect 2605 304 2611 336
rect 2621 224 2627 416
rect 2637 344 2643 416
rect 2669 364 2675 516
rect 2701 504 2707 516
rect 2733 484 2739 496
rect 2653 284 2659 336
rect 2701 304 2707 336
rect 2717 324 2723 476
rect 2749 443 2755 656
rect 2765 524 2771 616
rect 2781 544 2787 656
rect 2797 584 2803 676
rect 2845 664 2851 696
rect 2813 644 2819 656
rect 2813 604 2819 636
rect 2829 524 2835 576
rect 2781 517 2819 523
rect 2781 504 2787 517
rect 2813 503 2819 517
rect 2845 523 2851 656
rect 2877 643 2883 676
rect 2861 637 2883 643
rect 2861 544 2867 637
rect 2909 564 2915 694
rect 2845 517 2860 523
rect 2861 503 2867 516
rect 2813 497 2851 503
rect 2861 497 2883 503
rect 2845 483 2851 497
rect 2845 477 2860 483
rect 2749 437 2771 443
rect 2765 304 2771 437
rect 2570 214 2582 216
rect 2555 206 2557 214
rect 2565 206 2567 214
rect 2575 206 2577 214
rect 2585 206 2587 214
rect 2595 206 2597 214
rect 2570 204 2582 206
rect 2621 184 2627 216
rect 2637 184 2643 256
rect 2669 104 2675 296
rect 2701 204 2707 256
rect 2701 164 2707 176
rect 2685 64 2691 116
rect 2637 -23 2643 56
rect 2765 24 2771 276
rect 2781 244 2787 276
rect 2781 124 2787 156
rect 2781 84 2787 116
rect 2797 104 2803 336
rect 2813 324 2819 456
rect 2877 344 2883 497
rect 2893 344 2899 556
rect 2941 544 2947 676
rect 2909 504 2915 536
rect 2957 524 2963 596
rect 2932 517 2947 523
rect 2861 164 2867 296
rect 2909 284 2915 456
rect 2925 404 2931 436
rect 2941 404 2947 517
rect 2973 504 2979 816
rect 3037 804 3043 836
rect 3053 684 3059 716
rect 3069 704 3075 716
rect 3133 704 3139 856
rect 3149 724 3155 796
rect 3149 704 3155 716
rect 3117 684 3123 696
rect 3165 684 3171 716
rect 3213 704 3219 716
rect 3261 704 3267 916
rect 3261 684 3267 696
rect 3037 644 3043 676
rect 2980 497 2988 503
rect 3005 364 3011 616
rect 3069 584 3075 596
rect 3021 544 3027 576
rect 3085 564 3091 596
rect 3021 524 3027 536
rect 3037 524 3043 556
rect 3053 544 3059 556
rect 3101 524 3107 536
rect 3117 524 3123 656
rect 3277 583 3283 776
rect 3293 764 3299 1096
rect 3373 1064 3379 1197
rect 3405 1084 3411 1236
rect 3469 1224 3475 1516
rect 3485 1424 3491 1656
rect 3501 1504 3507 1556
rect 3517 1504 3523 1696
rect 3533 1664 3539 1697
rect 3485 1244 3491 1356
rect 3517 1303 3523 1476
rect 3549 1364 3555 1676
rect 3565 1424 3571 1496
rect 3581 1484 3587 1496
rect 3597 1484 3603 1656
rect 3613 1504 3619 1676
rect 3629 1504 3635 1676
rect 3645 1564 3651 1636
rect 3661 1544 3667 1556
rect 3508 1297 3523 1303
rect 3549 1264 3555 1336
rect 3565 1324 3571 1416
rect 3597 1383 3603 1476
rect 3645 1404 3651 1516
rect 3725 1504 3731 1716
rect 3757 1704 3763 1776
rect 3757 1524 3763 1696
rect 3805 1664 3811 1836
rect 3773 1584 3779 1636
rect 3757 1504 3763 1516
rect 3773 1504 3779 1536
rect 3661 1484 3667 1496
rect 3597 1377 3619 1383
rect 3613 1364 3619 1377
rect 3597 1324 3603 1356
rect 3613 1344 3619 1356
rect 3629 1324 3635 1336
rect 3469 1102 3475 1116
rect 3533 1004 3539 1076
rect 3453 984 3459 996
rect 3565 963 3571 1236
rect 3581 1124 3587 1316
rect 3597 1104 3603 1116
rect 3613 1104 3619 1156
rect 3629 1124 3635 1316
rect 3661 1224 3667 1236
rect 3661 1104 3667 1136
rect 3629 963 3635 1036
rect 3556 957 3571 963
rect 3613 957 3635 963
rect 3357 944 3363 956
rect 3309 923 3315 936
rect 3437 924 3443 936
rect 3517 924 3523 956
rect 3565 924 3571 936
rect 3613 924 3619 957
rect 3645 924 3651 936
rect 3677 924 3683 1256
rect 3693 1104 3699 1416
rect 3709 1324 3715 1376
rect 3725 1324 3731 1416
rect 3741 1324 3747 1456
rect 3757 1424 3763 1476
rect 3757 1303 3763 1416
rect 3773 1384 3779 1396
rect 3789 1324 3795 1376
rect 3741 1297 3763 1303
rect 3709 1104 3715 1156
rect 3741 1004 3747 1297
rect 3757 1104 3763 1136
rect 3757 944 3763 1076
rect 3309 917 3324 923
rect 3309 684 3315 716
rect 3325 704 3331 916
rect 3341 744 3347 916
rect 3357 724 3363 736
rect 3332 697 3347 703
rect 3325 663 3331 676
rect 3300 657 3331 663
rect 3277 577 3299 583
rect 3181 524 3187 556
rect 3213 524 3219 576
rect 3229 557 3244 563
rect 3117 484 3123 516
rect 3005 304 3011 316
rect 2973 143 2979 276
rect 3021 164 3027 476
rect 3037 284 3043 316
rect 3069 304 3075 316
rect 3085 303 3091 396
rect 3117 304 3123 356
rect 3085 297 3107 303
rect 3101 284 3107 297
rect 3085 244 3091 276
rect 3133 164 3139 456
rect 3149 264 3155 496
rect 3229 344 3235 557
rect 3165 337 3219 343
rect 3165 324 3171 337
rect 3213 323 3219 337
rect 3245 324 3251 536
rect 3277 524 3283 556
rect 3293 504 3299 577
rect 3325 564 3331 596
rect 3341 544 3347 697
rect 3389 624 3395 916
rect 3485 744 3491 916
rect 3501 864 3507 916
rect 3437 684 3443 696
rect 3373 584 3379 616
rect 3341 524 3347 536
rect 3357 524 3363 576
rect 3293 343 3299 436
rect 3261 337 3299 343
rect 3213 317 3235 323
rect 3181 304 3187 316
rect 2973 137 2988 143
rect 2829 84 2835 118
rect 2861 84 2867 116
rect 2925 104 2931 116
rect 3005 84 3011 116
rect 3133 84 3139 118
rect 3165 84 3171 296
rect 3213 224 3219 296
rect 3229 224 3235 317
rect 3245 264 3251 316
rect 3261 304 3267 337
rect 3341 324 3347 516
rect 3389 444 3395 616
rect 3453 504 3459 516
rect 3469 464 3475 676
rect 3501 524 3507 576
rect 3517 564 3523 916
rect 3693 864 3699 936
rect 3597 724 3603 736
rect 3597 664 3603 676
rect 3373 384 3379 416
rect 3469 344 3475 456
rect 3533 364 3539 496
rect 3581 484 3587 636
rect 3613 524 3619 816
rect 3645 644 3651 656
rect 3709 624 3715 836
rect 3757 544 3763 936
rect 3773 924 3779 1296
rect 3805 1204 3811 1656
rect 3837 1624 3843 1856
rect 3869 1844 3875 1876
rect 3901 1784 3907 2056
rect 3917 2024 3923 2116
rect 3949 2044 3955 2116
rect 3965 2104 3971 2217
rect 3981 2184 3987 2317
rect 4045 2304 4051 2316
rect 4125 2284 4131 2376
rect 4301 2284 4307 2496
rect 4333 2384 4339 2436
rect 4141 2244 4147 2256
rect 4349 2183 4355 2676
rect 4397 2524 4403 2636
rect 4413 2504 4419 2536
rect 4445 2484 4451 2716
rect 4477 2684 4483 3136
rect 4493 2724 4499 3396
rect 4509 3324 4515 3336
rect 4525 3084 4531 3336
rect 4621 3324 4627 3336
rect 4653 3324 4659 3457
rect 4573 3084 4579 3096
rect 4525 2944 4531 3076
rect 4621 3064 4627 3316
rect 4653 3104 4659 3316
rect 4669 3264 4675 3316
rect 4557 2944 4563 3036
rect 4573 2924 4579 3056
rect 4589 2884 4595 2996
rect 4621 2964 4627 2976
rect 4669 2924 4675 3216
rect 4573 2744 4579 2756
rect 4589 2744 4595 2876
rect 4541 2724 4547 2736
rect 4573 2704 4579 2716
rect 4493 2584 4499 2676
rect 4653 2604 4659 2696
rect 4509 2524 4515 2576
rect 4365 2284 4371 2296
rect 4381 2184 4387 2316
rect 4429 2304 4435 2436
rect 4445 2324 4451 2476
rect 4525 2324 4531 2596
rect 4669 2524 4675 2916
rect 4685 2863 4691 3276
rect 4701 3124 4707 3236
rect 4749 3224 4755 3316
rect 4797 3284 4803 3356
rect 4797 3244 4803 3276
rect 4925 3184 4931 3336
rect 4701 2884 4707 2896
rect 4749 2884 4755 3076
rect 4861 3044 4867 3056
rect 4829 2924 4835 2936
rect 4685 2857 4700 2863
rect 4701 2784 4707 2856
rect 4717 2744 4723 2776
rect 4701 2564 4707 2576
rect 4765 2564 4771 2596
rect 4493 2304 4499 2316
rect 4509 2304 4515 2316
rect 4413 2284 4419 2296
rect 4397 2184 4403 2236
rect 4333 2177 4355 2183
rect 3997 2144 4003 2176
rect 4333 2144 4339 2177
rect 4381 2144 4387 2176
rect 3949 1964 3955 2036
rect 3997 1984 4003 2136
rect 4029 2064 4035 2096
rect 4029 2024 4035 2056
rect 4125 2043 4131 2136
rect 4157 2064 4163 2116
rect 4285 2104 4291 2116
rect 4381 2104 4387 2136
rect 4125 2037 4147 2043
rect 4074 2014 4086 2016
rect 4059 2006 4061 2014
rect 4069 2006 4071 2014
rect 4079 2006 4081 2014
rect 4089 2006 4091 2014
rect 4099 2006 4101 2014
rect 4074 2004 4086 2006
rect 4141 1984 4147 2037
rect 4173 1924 4179 2016
rect 4189 1904 4195 2076
rect 4301 1984 4307 2076
rect 4397 1984 4403 2096
rect 4237 1904 4243 1956
rect 4317 1944 4323 1976
rect 3997 1824 4003 1894
rect 4109 1884 4115 1896
rect 3901 1744 3907 1776
rect 4029 1744 4035 1876
rect 4173 1824 4179 1836
rect 3837 1504 3843 1576
rect 3885 1504 3891 1716
rect 3933 1684 3939 1736
rect 3933 1544 3939 1676
rect 3965 1524 3971 1676
rect 4013 1484 4019 1676
rect 4109 1663 4115 1736
rect 4141 1724 4147 1736
rect 4221 1723 4227 1836
rect 4269 1784 4275 1936
rect 4301 1923 4307 1936
rect 4301 1917 4323 1923
rect 4285 1864 4291 1896
rect 4301 1784 4307 1896
rect 4221 1717 4236 1723
rect 4109 1657 4131 1663
rect 4074 1614 4086 1616
rect 4059 1606 4061 1614
rect 4069 1606 4071 1614
rect 4079 1606 4081 1614
rect 4089 1606 4091 1614
rect 4099 1606 4101 1614
rect 4074 1604 4086 1606
rect 4125 1544 4131 1657
rect 3805 1064 3811 1196
rect 3821 1084 3827 1236
rect 3837 1183 3843 1476
rect 3853 1324 3859 1436
rect 3869 1184 3875 1276
rect 3901 1263 3907 1456
rect 3917 1344 3923 1356
rect 4013 1344 4019 1476
rect 4029 1324 4035 1496
rect 4221 1404 4227 1717
rect 4253 1684 4259 1736
rect 4317 1524 4323 1917
rect 4333 1917 4348 1923
rect 4333 1784 4339 1917
rect 4381 1904 4387 1956
rect 4397 1944 4403 1976
rect 4381 1864 4387 1876
rect 4333 1764 4339 1776
rect 4349 1764 4355 1836
rect 4365 1784 4371 1836
rect 4397 1764 4403 1936
rect 4413 1924 4419 2156
rect 4429 2144 4435 2296
rect 4461 2084 4467 2236
rect 4525 2184 4531 2316
rect 4541 2304 4547 2516
rect 4573 2504 4579 2516
rect 4637 2504 4643 2518
rect 4589 2344 4595 2356
rect 4477 2124 4483 2136
rect 4461 2064 4467 2076
rect 4461 2024 4467 2036
rect 4509 1924 4515 1936
rect 4429 1884 4435 1916
rect 4541 1904 4547 2296
rect 4589 2264 4595 2336
rect 4717 2264 4723 2296
rect 4765 2284 4771 2556
rect 4781 2504 4787 2776
rect 4797 2704 4803 2916
rect 4845 2764 4851 2976
rect 4877 2964 4883 3056
rect 4893 2984 4899 3036
rect 4909 2763 4915 2956
rect 4925 2944 4931 3036
rect 4941 2864 4947 2876
rect 4925 2784 4931 2836
rect 4909 2757 4931 2763
rect 4797 2604 4803 2696
rect 4845 2664 4851 2694
rect 4797 2564 4803 2576
rect 4861 2524 4867 2596
rect 4829 2324 4835 2356
rect 4845 2324 4851 2416
rect 4589 2164 4595 2176
rect 4877 2144 4883 2756
rect 4909 2664 4915 2736
rect 4909 2524 4915 2576
rect 4893 2304 4899 2356
rect 4893 2124 4899 2296
rect 4909 2244 4915 2436
rect 4925 2204 4931 2757
rect 4957 2704 4963 3096
rect 4989 2924 4995 3256
rect 5005 2964 5011 3356
rect 4989 2883 4995 2916
rect 4989 2877 5011 2883
rect 4973 2864 4979 2876
rect 4973 2704 4979 2856
rect 4989 2724 4995 2836
rect 5005 2784 5011 2877
rect 4941 2344 4947 2376
rect 4957 2364 4963 2696
rect 4973 2664 4979 2676
rect 5005 2484 5011 2696
rect 5021 2604 5027 3236
rect 5037 3084 5043 3136
rect 5053 3084 5059 3096
rect 5069 3084 5075 3316
rect 5085 3284 5091 3336
rect 5053 2904 5059 2916
rect 5037 2744 5043 2896
rect 5037 2684 5043 2696
rect 5021 2524 5027 2536
rect 5069 2504 5075 2876
rect 5085 2864 5091 3036
rect 5037 2484 5043 2496
rect 5037 2424 5043 2476
rect 5053 2464 5059 2496
rect 5085 2384 5091 2836
rect 5101 2784 5107 3316
rect 5133 3104 5139 3236
rect 5101 2724 5107 2776
rect 4941 2264 4947 2336
rect 4925 2143 4931 2196
rect 4941 2184 4947 2236
rect 4925 2137 4947 2143
rect 4717 2104 4723 2118
rect 4797 2104 4803 2116
rect 4781 2084 4787 2096
rect 4429 1824 4435 1856
rect 4429 1764 4435 1816
rect 4445 1804 4451 1836
rect 4461 1804 4467 1876
rect 4365 1684 4371 1756
rect 4477 1744 4483 1896
rect 4493 1784 4499 1856
rect 4541 1844 4547 1876
rect 4525 1784 4531 1816
rect 4493 1764 4499 1776
rect 4525 1764 4531 1776
rect 4557 1743 4563 2036
rect 4573 1944 4579 2056
rect 4653 1984 4659 2076
rect 4717 1984 4723 2056
rect 4749 1944 4755 1996
rect 4589 1904 4595 1916
rect 4605 1883 4611 1916
rect 4653 1904 4659 1916
rect 4669 1884 4675 1916
rect 4717 1904 4723 1916
rect 4589 1877 4611 1883
rect 4589 1844 4595 1877
rect 4733 1844 4739 1916
rect 4749 1864 4755 1936
rect 4813 1903 4819 2116
rect 4925 2064 4931 2096
rect 4829 1924 4835 1956
rect 4804 1897 4819 1903
rect 4813 1844 4819 1897
rect 4589 1824 4595 1836
rect 4541 1737 4563 1743
rect 4397 1724 4403 1736
rect 4541 1724 4547 1737
rect 4557 1724 4563 1737
rect 4589 1724 4595 1816
rect 4733 1804 4739 1836
rect 4653 1724 4659 1756
rect 4797 1724 4803 1836
rect 4813 1724 4819 1736
rect 4381 1704 4387 1716
rect 4477 1704 4483 1716
rect 4605 1704 4611 1716
rect 4781 1704 4787 1716
rect 4685 1684 4691 1696
rect 4861 1684 4867 1716
rect 4877 1684 4883 1936
rect 4125 1364 4131 1376
rect 4253 1364 4259 1476
rect 3917 1304 3923 1316
rect 3901 1257 3923 1263
rect 3837 1177 3859 1183
rect 3853 924 3859 1177
rect 3901 1124 3907 1236
rect 3901 1084 3907 1096
rect 3917 1084 3923 1257
rect 3981 1244 3987 1276
rect 3981 1184 3987 1236
rect 4013 1124 4019 1316
rect 4029 1103 4035 1316
rect 4317 1304 4323 1516
rect 4557 1504 4563 1516
rect 4509 1484 4515 1496
rect 4573 1484 4579 1676
rect 4477 1444 4483 1476
rect 4074 1214 4086 1216
rect 4059 1206 4061 1214
rect 4069 1206 4071 1214
rect 4079 1206 4081 1214
rect 4089 1206 4091 1214
rect 4099 1206 4101 1214
rect 4074 1204 4086 1206
rect 4125 1164 4131 1236
rect 4333 1124 4339 1396
rect 4349 1344 4355 1356
rect 4397 1304 4403 1316
rect 4429 1184 4435 1336
rect 4445 1324 4451 1396
rect 4493 1324 4499 1336
rect 4445 1304 4451 1316
rect 4221 1104 4227 1116
rect 4020 1097 4035 1103
rect 3869 944 3875 1056
rect 3773 824 3779 916
rect 3805 804 3811 896
rect 3853 864 3859 916
rect 3949 903 3955 996
rect 3949 897 3971 903
rect 3885 804 3891 836
rect 3773 702 3779 716
rect 3837 684 3843 716
rect 3853 704 3859 716
rect 3892 697 3907 703
rect 3901 684 3907 697
rect 3773 544 3779 656
rect 3885 543 3891 676
rect 3901 604 3907 676
rect 3885 537 3900 543
rect 3565 364 3571 436
rect 3629 324 3635 356
rect 3277 224 3283 316
rect 3341 304 3347 316
rect 3293 297 3308 303
rect 3293 224 3299 297
rect 3565 302 3571 316
rect 3645 304 3651 316
rect 3693 304 3699 516
rect 3309 144 3315 276
rect 3325 264 3331 276
rect 3357 264 3363 296
rect 3325 144 3331 256
rect 3421 244 3427 296
rect 3357 184 3363 216
rect 3421 157 3452 163
rect 3197 124 3203 136
rect 3309 124 3315 136
rect 3421 124 3427 157
rect 3469 143 3475 216
rect 3485 204 3491 216
rect 3485 164 3491 196
rect 3460 137 3475 143
rect 3437 124 3443 136
rect 3501 124 3507 256
rect 3533 184 3539 256
rect 3597 204 3603 276
rect 3677 244 3683 276
rect 3741 264 3747 316
rect 3757 284 3763 536
rect 3821 464 3827 536
rect 3853 524 3859 536
rect 3853 484 3859 496
rect 3853 344 3859 456
rect 3661 164 3667 236
rect 3693 164 3699 176
rect 3661 124 3667 156
rect 3773 124 3779 276
rect 3805 144 3811 276
rect 3853 204 3859 336
rect 3885 304 3891 516
rect 3917 384 3923 536
rect 3949 524 3955 596
rect 3965 544 3971 897
rect 4077 864 4083 1076
rect 4141 984 4147 996
rect 4237 944 4243 1056
rect 4301 1004 4307 1076
rect 4333 904 4339 1036
rect 4397 964 4403 976
rect 4365 937 4380 943
rect 4074 814 4086 816
rect 4059 806 4061 814
rect 4069 806 4071 814
rect 4079 806 4081 814
rect 4089 806 4091 814
rect 4099 806 4101 814
rect 4074 804 4086 806
rect 4077 702 4083 716
rect 4141 684 4147 736
rect 4237 704 4243 716
rect 4253 684 4259 716
rect 4301 684 4307 856
rect 4365 784 4371 937
rect 4109 604 4115 676
rect 4301 624 4307 676
rect 4333 604 4339 636
rect 4093 564 4099 576
rect 4093 524 4099 556
rect 4221 526 4227 556
rect 4253 544 4259 596
rect 4365 564 4371 776
rect 4381 544 4387 576
rect 4221 517 4227 518
rect 3949 504 3955 516
rect 3949 324 3955 496
rect 3981 304 3987 436
rect 4074 414 4086 416
rect 4059 406 4061 414
rect 4069 406 4071 414
rect 4079 406 4081 414
rect 4089 406 4091 414
rect 4099 406 4101 414
rect 4074 404 4086 406
rect 4013 384 4019 396
rect 4013 284 4019 376
rect 4157 324 4163 356
rect 4157 304 4163 316
rect 4253 304 4259 536
rect 4285 524 4291 536
rect 4397 524 4403 836
rect 4429 563 4435 1176
rect 4477 944 4483 1056
rect 4509 984 4515 1436
rect 4525 1284 4531 1336
rect 4525 1264 4531 1276
rect 4573 1124 4579 1296
rect 4573 1084 4579 1096
rect 4541 1044 4547 1076
rect 4605 1064 4611 1636
rect 4621 1144 4627 1676
rect 4781 1524 4787 1636
rect 4701 1344 4707 1476
rect 4701 1324 4707 1336
rect 4621 1104 4627 1116
rect 4525 926 4531 936
rect 4557 804 4563 936
rect 4605 884 4611 1036
rect 4621 924 4627 1096
rect 4669 1084 4675 1216
rect 4701 1084 4707 1196
rect 4717 1144 4723 1156
rect 4845 1144 4851 1636
rect 4861 1584 4867 1676
rect 4877 1484 4883 1676
rect 4893 1504 4899 1696
rect 4941 1584 4947 2137
rect 5005 2124 5011 2136
rect 5005 1884 5011 2116
rect 4861 1444 4867 1456
rect 4877 1404 4883 1476
rect 4925 1364 4931 1376
rect 4861 1326 4867 1336
rect 4893 1324 4899 1336
rect 4957 1324 4963 1836
rect 4973 1744 4979 1856
rect 5037 1783 5043 2376
rect 5101 2043 5107 2516
rect 5117 2323 5123 3076
rect 5117 2317 5139 2323
rect 5085 2037 5107 2043
rect 5085 1943 5091 2037
rect 5085 1937 5107 1943
rect 5069 1884 5075 1896
rect 5085 1864 5091 1896
rect 5021 1777 5043 1783
rect 4973 1544 4979 1736
rect 4989 1726 4995 1736
rect 4957 1143 4963 1316
rect 4941 1137 4963 1143
rect 4717 1124 4723 1136
rect 4637 1004 4643 1076
rect 4909 1064 4915 1116
rect 4941 1104 4947 1137
rect 4957 1104 4963 1116
rect 4685 944 4691 976
rect 4685 904 4691 936
rect 4813 926 4819 956
rect 4845 944 4851 1056
rect 4941 983 4947 1096
rect 4973 1003 4979 1496
rect 5021 1364 5027 1777
rect 5053 1724 5059 1756
rect 5069 1724 5075 1836
rect 5101 1724 5107 1937
rect 5133 1904 5139 2317
rect 5149 2124 5155 2176
rect 5133 1804 5139 1836
rect 5117 1764 5123 1796
rect 5149 1724 5155 1856
rect 5101 1504 5107 1716
rect 5133 1704 5139 1716
rect 5037 1324 5043 1496
rect 5053 1324 5059 1476
rect 5069 1384 5075 1494
rect 5012 1297 5027 1303
rect 5021 1184 5027 1297
rect 4989 1124 4995 1176
rect 5005 1124 5011 1156
rect 5021 1104 5027 1136
rect 4925 977 4947 983
rect 4957 997 4979 1003
rect 4925 924 4931 977
rect 4941 944 4947 956
rect 4669 884 4675 896
rect 4749 864 4755 916
rect 4621 804 4627 856
rect 4445 684 4451 776
rect 4621 704 4627 796
rect 4685 702 4691 716
rect 4509 684 4515 696
rect 4461 644 4467 656
rect 4461 583 4467 636
rect 4452 577 4467 583
rect 4429 557 4451 563
rect 4429 524 4435 536
rect 4317 504 4323 516
rect 4253 284 4259 296
rect 3853 144 3859 196
rect 3981 144 3987 276
rect 4173 244 4179 276
rect 4013 126 4019 156
rect 4237 144 4243 196
rect 4349 144 4355 276
rect 4381 244 4387 256
rect 4445 244 4451 557
rect 4541 524 4547 636
rect 4621 623 4627 696
rect 4749 664 4755 736
rect 4781 704 4787 916
rect 4861 744 4867 796
rect 4877 784 4883 896
rect 4829 724 4835 736
rect 4605 617 4627 623
rect 4605 544 4611 617
rect 4637 584 4643 616
rect 4717 544 4723 656
rect 4717 524 4723 536
rect 4765 524 4771 696
rect 4381 224 4387 236
rect 4445 144 4451 236
rect 4013 117 4019 118
rect 3229 104 3235 116
rect 3325 24 3331 116
rect 3389 64 3395 116
rect 3565 84 3571 116
rect 3613 104 3619 116
rect 4141 104 4147 136
rect 4173 104 4179 116
rect 3885 84 3891 96
rect 4253 84 4259 136
rect 4461 124 4467 516
rect 4493 304 4499 316
rect 4509 284 4515 516
rect 4861 484 4867 736
rect 4877 704 4883 716
rect 4893 704 4899 716
rect 4957 704 4963 997
rect 4989 924 4995 1096
rect 5053 944 5059 1316
rect 5069 1284 5075 1296
rect 5069 1124 5075 1216
rect 5085 1204 5091 1296
rect 5117 1284 5123 1396
rect 5101 1264 5107 1276
rect 5117 1143 5123 1276
rect 5108 1137 5123 1143
rect 5149 1124 5155 1196
rect 4957 684 4963 696
rect 4909 604 4915 656
rect 4909 583 4915 596
rect 4909 577 4924 583
rect 4909 524 4915 536
rect 4868 477 4876 483
rect 4573 324 4579 356
rect 4557 144 4563 196
rect 4573 124 4579 316
rect 4605 243 4611 276
rect 4605 237 4627 243
rect 4381 104 4387 118
rect 4477 104 4483 116
rect 4509 104 4515 116
rect 4589 103 4595 236
rect 4621 184 4627 237
rect 4637 204 4643 436
rect 4701 324 4707 436
rect 4765 304 4771 376
rect 4781 323 4787 436
rect 4781 317 4796 323
rect 4685 144 4691 276
rect 4813 264 4819 336
rect 4861 304 4867 376
rect 4893 324 4899 436
rect 4957 384 4963 676
rect 4973 664 4979 896
rect 4989 864 4995 876
rect 5005 804 5011 876
rect 5021 784 5027 936
rect 5069 924 5075 1096
rect 4989 724 4995 756
rect 5037 744 5043 836
rect 5053 804 5059 876
rect 5069 724 5075 916
rect 5149 904 5155 1116
rect 5133 684 5139 776
rect 4989 523 4995 636
rect 4989 517 5004 523
rect 5021 284 5027 536
rect 4717 184 4723 256
rect 4797 204 4803 236
rect 4701 124 4707 136
rect 4925 124 4931 196
rect 4973 144 4979 276
rect 5021 184 5027 276
rect 5133 144 5139 676
rect 4589 97 4604 103
rect 4074 14 4086 16
rect 4059 6 4061 14
rect 4069 6 4071 14
rect 4079 6 4081 14
rect 4089 6 4091 14
rect 4099 6 4101 14
rect 4074 4 4086 6
<< m3contact >>
rect 140 3356 148 3364
rect 364 3356 372 3364
rect 12 3316 20 3324
rect 348 3336 356 3344
rect 476 3336 484 3344
rect 668 3336 676 3344
rect 236 3316 244 3324
rect 300 3316 308 3324
rect 348 3316 356 3324
rect 332 3296 340 3304
rect 60 3136 68 3144
rect 92 3136 100 3144
rect 252 3136 260 3144
rect 12 3096 20 3104
rect 236 3076 244 3084
rect 12 2996 20 3004
rect 44 2996 52 3004
rect 364 3296 372 3304
rect 396 3276 404 3284
rect 364 3256 372 3264
rect 348 3096 356 3104
rect 460 3296 468 3304
rect 492 3316 500 3324
rect 524 3316 532 3324
rect 412 3236 420 3244
rect 380 3156 388 3164
rect 444 3136 452 3144
rect 476 3116 484 3124
rect 476 3096 484 3104
rect 268 2976 276 2984
rect 396 2976 404 2984
rect 124 2916 132 2924
rect 268 2916 276 2924
rect 204 2776 212 2784
rect 140 2736 148 2744
rect 44 2716 52 2724
rect 172 2716 180 2724
rect 12 2696 20 2704
rect 172 2696 180 2704
rect 44 2676 52 2684
rect 60 2636 68 2644
rect 60 2536 68 2544
rect 12 2496 20 2504
rect 12 2336 20 2344
rect 44 2316 52 2324
rect 60 2296 68 2304
rect 108 2656 116 2664
rect 124 2456 132 2464
rect 108 2436 116 2444
rect 108 2356 116 2364
rect 460 2916 468 2924
rect 332 2816 340 2824
rect 524 3296 532 3304
rect 924 3396 932 3404
rect 1308 3376 1316 3384
rect 1500 3376 1508 3384
rect 1948 3376 1956 3384
rect 1932 3356 1940 3364
rect 2547 3406 2555 3414
rect 2557 3406 2565 3414
rect 2567 3406 2575 3414
rect 2577 3406 2585 3414
rect 2587 3406 2595 3414
rect 2597 3406 2605 3414
rect 2284 3396 2292 3404
rect 2524 3396 2532 3404
rect 2252 3356 2260 3364
rect 2428 3356 2436 3364
rect 732 3336 740 3344
rect 1068 3336 1076 3344
rect 1228 3336 1236 3344
rect 1292 3336 1300 3344
rect 1596 3336 1604 3344
rect 1836 3336 1844 3344
rect 2172 3336 2180 3344
rect 2220 3336 2228 3344
rect 732 3316 740 3324
rect 652 3276 660 3284
rect 700 3276 708 3284
rect 732 3276 740 3284
rect 604 3256 612 3264
rect 588 3236 596 3244
rect 716 3236 724 3244
rect 540 3156 548 3164
rect 668 3156 676 3164
rect 556 3136 564 3144
rect 508 3116 516 3124
rect 540 3096 548 3104
rect 636 3116 644 3124
rect 508 3076 516 3084
rect 476 2756 484 2764
rect 380 2696 388 2704
rect 204 2676 212 2684
rect 316 2676 324 2684
rect 380 2676 388 2684
rect 428 2676 436 2684
rect 412 2616 420 2624
rect 492 2656 500 2664
rect 444 2596 452 2604
rect 476 2596 484 2604
rect 332 2556 340 2564
rect 268 2536 276 2544
rect 316 2536 324 2544
rect 236 2518 244 2524
rect 236 2516 244 2518
rect 300 2516 308 2524
rect 300 2456 308 2464
rect 156 2436 164 2444
rect 188 2336 196 2344
rect 220 2316 228 2324
rect 364 2536 372 2544
rect 348 2516 356 2524
rect 364 2316 372 2324
rect 124 2296 132 2304
rect 140 2296 148 2304
rect 188 2296 196 2304
rect 316 2296 324 2304
rect 604 3016 612 3024
rect 588 2956 596 2964
rect 620 2936 628 2944
rect 652 3096 660 3104
rect 700 3036 708 3044
rect 860 3256 868 3264
rect 780 3236 788 3244
rect 812 3176 820 3184
rect 828 3176 836 3184
rect 812 3136 820 3144
rect 780 3116 788 3124
rect 732 3096 740 3104
rect 700 2956 708 2964
rect 716 2956 724 2964
rect 684 2936 692 2944
rect 908 3116 916 3124
rect 1004 3296 1012 3304
rect 1004 3256 1012 3264
rect 1228 3316 1236 3324
rect 1276 3316 1284 3324
rect 1436 3318 1444 3324
rect 1436 3316 1444 3318
rect 1532 3316 1540 3324
rect 1372 3296 1380 3304
rect 1564 3296 1572 3304
rect 1196 3276 1204 3284
rect 1292 3276 1300 3284
rect 1180 3256 1188 3264
rect 940 3236 948 3244
rect 1164 3236 1172 3244
rect 1043 3206 1051 3214
rect 1053 3206 1061 3214
rect 1063 3206 1071 3214
rect 1073 3206 1081 3214
rect 1083 3206 1091 3214
rect 1093 3206 1101 3214
rect 1148 3116 1156 3124
rect 1132 3096 1140 3104
rect 924 3076 932 3084
rect 748 3056 756 3064
rect 1004 3056 1012 3064
rect 796 3036 804 3044
rect 844 2996 852 3004
rect 732 2936 740 2944
rect 748 2936 756 2944
rect 860 2936 868 2944
rect 780 2916 788 2924
rect 828 2916 836 2924
rect 636 2876 644 2884
rect 764 2876 772 2884
rect 732 2836 740 2844
rect 652 2816 660 2824
rect 556 2776 564 2784
rect 588 2736 596 2744
rect 540 2716 548 2724
rect 524 2696 532 2704
rect 636 2716 644 2724
rect 700 2756 708 2764
rect 732 2756 740 2764
rect 668 2736 676 2744
rect 796 2736 804 2744
rect 764 2716 772 2724
rect 716 2696 724 2704
rect 748 2696 756 2704
rect 604 2676 612 2684
rect 572 2636 580 2644
rect 572 2616 580 2624
rect 604 2616 612 2624
rect 588 2596 596 2604
rect 508 2536 516 2544
rect 556 2536 564 2544
rect 508 2496 516 2504
rect 556 2496 564 2504
rect 540 2476 548 2484
rect 492 2376 500 2384
rect 476 2356 484 2364
rect 492 2336 500 2344
rect 460 2316 468 2324
rect 108 2276 116 2284
rect 172 2276 180 2284
rect 428 2276 436 2284
rect 44 2116 52 2124
rect 156 2116 164 2124
rect 12 2096 20 2104
rect 60 2096 68 2104
rect 108 2096 116 2104
rect 44 1916 52 1924
rect 140 2096 148 2104
rect 396 2156 404 2164
rect 300 2118 308 2124
rect 300 2116 308 2118
rect 140 2036 148 2044
rect 172 2036 180 2044
rect 284 1936 292 1944
rect 204 1916 212 1924
rect 12 1896 20 1904
rect 92 1896 100 1904
rect 124 1896 132 1904
rect 172 1896 180 1904
rect 60 1856 68 1864
rect 92 1696 100 1704
rect 44 1516 52 1524
rect 204 1876 212 1884
rect 220 1816 228 1824
rect 412 2136 420 2144
rect 364 2116 372 2124
rect 412 2116 420 2124
rect 364 2096 372 2104
rect 476 2276 484 2284
rect 476 2156 484 2164
rect 524 2156 532 2164
rect 508 2076 516 2084
rect 540 1976 548 1984
rect 684 2636 692 2644
rect 636 2596 644 2604
rect 620 2576 628 2584
rect 860 2896 868 2904
rect 940 2956 948 2964
rect 956 2936 964 2944
rect 972 2936 980 2944
rect 1036 3036 1044 3044
rect 1036 2936 1044 2944
rect 1180 3096 1188 3104
rect 1228 3176 1236 3184
rect 1308 3156 1316 3164
rect 1260 3096 1268 3104
rect 1212 3076 1220 3084
rect 1180 2996 1188 3004
rect 1196 2976 1204 2984
rect 908 2916 916 2924
rect 988 2916 996 2924
rect 1020 2916 1028 2924
rect 1164 2916 1172 2924
rect 972 2896 980 2904
rect 1004 2896 1012 2904
rect 892 2816 900 2824
rect 860 2776 868 2784
rect 844 2756 852 2764
rect 828 2716 836 2724
rect 780 2696 788 2704
rect 812 2696 820 2704
rect 924 2796 932 2804
rect 876 2736 884 2744
rect 908 2736 916 2744
rect 892 2716 900 2724
rect 908 2716 916 2724
rect 796 2676 804 2684
rect 812 2676 820 2684
rect 876 2676 884 2684
rect 924 2676 932 2684
rect 732 2556 740 2564
rect 764 2556 772 2564
rect 876 2556 884 2564
rect 636 2536 644 2544
rect 764 2536 772 2544
rect 908 2536 916 2544
rect 620 2516 628 2524
rect 620 2356 628 2364
rect 604 2336 612 2344
rect 908 2516 916 2524
rect 668 2496 676 2504
rect 684 2296 692 2304
rect 748 2302 756 2304
rect 748 2296 756 2302
rect 684 2256 692 2264
rect 860 2436 868 2444
rect 828 2296 836 2304
rect 908 2316 916 2324
rect 812 2276 820 2284
rect 1132 2856 1140 2864
rect 1148 2856 1156 2864
rect 1020 2816 1028 2824
rect 1004 2702 1012 2704
rect 1004 2696 1012 2702
rect 1043 2806 1051 2814
rect 1053 2806 1061 2814
rect 1063 2806 1071 2814
rect 1073 2806 1081 2814
rect 1083 2806 1091 2814
rect 1093 2806 1101 2814
rect 1116 2796 1124 2804
rect 1036 2696 1044 2704
rect 1148 2776 1156 2784
rect 1148 2736 1156 2744
rect 1116 2676 1124 2684
rect 1036 2656 1044 2664
rect 956 2516 964 2524
rect 1004 2556 1012 2564
rect 1292 3076 1300 3084
rect 1228 2976 1236 2984
rect 1532 3216 1540 3224
rect 1580 3216 1588 3224
rect 1468 3096 1476 3104
rect 1324 3056 1332 3064
rect 1244 2956 1252 2964
rect 1260 2936 1268 2944
rect 1228 2916 1236 2924
rect 1260 2916 1268 2924
rect 1212 2736 1220 2744
rect 1420 3056 1428 3064
rect 1372 3036 1380 3044
rect 1356 2956 1364 2964
rect 1340 2936 1348 2944
rect 1388 2976 1396 2984
rect 1404 2976 1412 2984
rect 1484 3076 1492 3084
rect 1500 2996 1508 3004
rect 1468 2976 1476 2984
rect 1516 2976 1524 2984
rect 1436 2916 1444 2924
rect 1388 2836 1396 2844
rect 1292 2796 1300 2804
rect 1324 2796 1332 2804
rect 1260 2776 1268 2784
rect 1276 2776 1284 2784
rect 1532 2956 1540 2964
rect 1548 2916 1556 2924
rect 1500 2896 1508 2904
rect 1452 2776 1460 2784
rect 1452 2736 1460 2744
rect 1420 2716 1428 2724
rect 1436 2716 1444 2724
rect 1212 2676 1220 2684
rect 1228 2676 1236 2684
rect 1244 2676 1252 2684
rect 1196 2656 1204 2664
rect 1500 2796 1508 2804
rect 1500 2756 1508 2764
rect 1468 2716 1476 2724
rect 1484 2716 1492 2724
rect 1468 2696 1476 2704
rect 1612 3276 1620 3284
rect 1740 3318 1748 3324
rect 1740 3316 1748 3318
rect 1836 3296 1844 3304
rect 1804 3276 1812 3284
rect 1868 3316 1876 3324
rect 1900 3316 1908 3324
rect 1868 3296 1876 3304
rect 2076 3296 2084 3304
rect 2028 3276 2036 3284
rect 2140 3276 2148 3284
rect 2252 3316 2260 3324
rect 1852 3236 1860 3244
rect 2156 3236 2164 3244
rect 1948 3216 1956 3224
rect 2012 3216 2020 3224
rect 2108 3216 2116 3224
rect 1804 3196 1812 3204
rect 1724 3136 1732 3144
rect 1708 3096 1716 3104
rect 1596 3076 1604 3084
rect 1580 2976 1588 2984
rect 1692 3056 1700 3064
rect 1756 3096 1764 3104
rect 1708 2996 1716 3004
rect 1724 2996 1732 3004
rect 1628 2976 1636 2984
rect 1692 2976 1700 2984
rect 1628 2936 1636 2944
rect 1644 2936 1652 2944
rect 1692 2936 1700 2944
rect 1644 2916 1652 2924
rect 1612 2896 1620 2904
rect 1628 2896 1636 2904
rect 1660 2896 1668 2904
rect 1580 2776 1588 2784
rect 1612 2696 1620 2704
rect 1292 2656 1300 2664
rect 1308 2656 1316 2664
rect 1340 2656 1348 2664
rect 1356 2656 1364 2664
rect 1404 2656 1412 2664
rect 1372 2636 1380 2644
rect 1260 2616 1268 2624
rect 1356 2616 1364 2624
rect 1324 2596 1332 2604
rect 1244 2576 1252 2584
rect 1260 2576 1268 2584
rect 1132 2536 1140 2544
rect 1164 2536 1172 2544
rect 1228 2536 1236 2544
rect 1132 2516 1140 2524
rect 1116 2496 1124 2504
rect 1196 2496 1204 2504
rect 1043 2406 1051 2414
rect 1053 2406 1061 2414
rect 1063 2406 1071 2414
rect 1073 2406 1081 2414
rect 1083 2406 1091 2414
rect 1093 2406 1101 2414
rect 1404 2596 1412 2604
rect 1388 2536 1396 2544
rect 1292 2516 1300 2524
rect 1340 2496 1348 2504
rect 1164 2476 1172 2484
rect 1212 2476 1220 2484
rect 1372 2476 1380 2484
rect 1132 2456 1140 2464
rect 1116 2396 1124 2404
rect 988 2376 996 2384
rect 924 2276 932 2284
rect 876 2256 884 2264
rect 924 2256 932 2264
rect 908 2176 916 2184
rect 620 2156 628 2164
rect 668 2156 676 2164
rect 572 2136 580 2144
rect 620 2136 628 2144
rect 956 2296 964 2304
rect 1116 2302 1124 2304
rect 1116 2296 1124 2302
rect 812 2136 820 2144
rect 716 2116 724 2124
rect 620 2056 628 2064
rect 588 1996 596 2004
rect 460 1956 468 1964
rect 524 1956 532 1964
rect 556 1956 564 1964
rect 588 1956 596 1964
rect 412 1916 420 1924
rect 348 1902 356 1904
rect 348 1896 356 1902
rect 348 1776 356 1784
rect 476 1896 484 1904
rect 508 1896 516 1904
rect 636 1896 644 1904
rect 460 1876 468 1884
rect 572 1876 580 1884
rect 636 1876 644 1884
rect 412 1856 420 1864
rect 460 1856 468 1864
rect 556 1856 564 1864
rect 236 1736 244 1744
rect 124 1716 132 1724
rect 204 1716 212 1724
rect 332 1716 340 1724
rect 156 1696 164 1704
rect 172 1696 180 1704
rect 300 1696 308 1704
rect 188 1676 196 1684
rect 284 1676 292 1684
rect 204 1516 212 1524
rect 12 1496 20 1504
rect 92 1496 100 1504
rect 172 1496 180 1504
rect 332 1496 340 1504
rect 108 1396 116 1404
rect 44 1376 52 1384
rect 108 1376 116 1384
rect 12 1336 20 1344
rect 236 1356 244 1364
rect 140 1336 148 1344
rect 60 1296 68 1304
rect 92 1296 100 1304
rect 44 1116 52 1124
rect 12 1096 20 1104
rect 300 1376 308 1384
rect 428 1516 436 1524
rect 348 1336 356 1344
rect 220 1156 228 1164
rect 268 1136 276 1144
rect 300 1116 308 1124
rect 332 1276 340 1284
rect 332 1256 340 1264
rect 268 1096 276 1104
rect 316 1096 324 1104
rect 252 1076 260 1084
rect 60 936 68 944
rect 156 936 164 944
rect 236 936 244 944
rect 44 916 52 924
rect 108 916 116 924
rect 140 916 148 924
rect 252 916 260 924
rect 412 1316 420 1324
rect 412 1296 420 1304
rect 364 1116 372 1124
rect 348 1076 356 1084
rect 284 916 292 924
rect 12 896 20 904
rect 92 896 100 904
rect 140 876 148 884
rect 172 876 180 884
rect 284 896 292 904
rect 428 936 436 944
rect 332 836 340 844
rect 220 756 228 764
rect 12 736 20 744
rect 44 736 52 744
rect 156 736 164 744
rect 348 716 356 724
rect 60 696 68 704
rect 108 696 116 704
rect 284 702 292 704
rect 284 696 292 702
rect 60 676 68 684
rect 92 636 100 644
rect 140 616 148 624
rect 332 556 340 564
rect 396 736 404 744
rect 428 736 436 744
rect 556 1836 564 1844
rect 588 1716 596 1724
rect 684 1956 692 1964
rect 924 2116 932 2124
rect 812 1996 820 2004
rect 780 1896 788 1904
rect 684 1876 692 1884
rect 668 1756 676 1764
rect 668 1716 676 1724
rect 652 1636 660 1644
rect 540 1616 548 1624
rect 588 1576 596 1584
rect 476 1556 484 1564
rect 524 1476 532 1484
rect 620 1476 628 1484
rect 652 1476 660 1484
rect 668 1436 676 1444
rect 652 1396 660 1404
rect 620 1356 628 1364
rect 492 1102 500 1104
rect 492 1096 500 1102
rect 748 1836 756 1844
rect 764 1756 772 1764
rect 716 1736 724 1744
rect 700 1536 708 1544
rect 700 1476 708 1484
rect 684 1416 692 1424
rect 684 1336 692 1344
rect 620 1296 628 1304
rect 556 1276 564 1284
rect 556 1136 564 1144
rect 588 1136 596 1144
rect 556 1096 564 1104
rect 604 1076 612 1084
rect 636 1076 644 1084
rect 556 1016 564 1024
rect 604 1016 612 1024
rect 588 956 596 964
rect 492 936 500 944
rect 524 936 532 944
rect 732 1296 740 1304
rect 716 1136 724 1144
rect 716 1116 724 1124
rect 700 1016 708 1024
rect 684 976 692 984
rect 732 936 740 944
rect 492 916 500 924
rect 636 916 644 924
rect 732 916 740 924
rect 556 876 564 884
rect 508 736 516 744
rect 460 716 468 724
rect 524 696 532 704
rect 652 836 660 844
rect 572 676 580 684
rect 380 656 388 664
rect 428 656 436 664
rect 284 516 292 524
rect 540 656 548 664
rect 444 636 452 644
rect 12 496 20 504
rect 44 476 52 484
rect 204 476 212 484
rect 140 356 148 364
rect 12 336 20 344
rect 428 496 436 504
rect 396 476 404 484
rect 428 476 436 484
rect 348 276 356 284
rect 60 136 68 144
rect 332 196 340 204
rect 220 136 228 144
rect 428 296 436 304
rect 460 516 468 524
rect 460 476 468 484
rect 476 456 484 464
rect 460 336 468 344
rect 524 556 532 564
rect 508 536 516 544
rect 508 516 516 524
rect 524 496 532 504
rect 492 376 500 384
rect 588 636 596 644
rect 556 576 564 584
rect 636 736 644 744
rect 748 896 756 904
rect 684 796 692 804
rect 716 736 724 744
rect 572 536 580 544
rect 620 536 628 544
rect 652 536 660 544
rect 748 836 756 844
rect 796 1716 804 1724
rect 972 2216 980 2224
rect 972 2176 980 2184
rect 1052 2156 1060 2164
rect 1004 2136 1012 2144
rect 1116 2136 1124 2144
rect 1004 2096 1012 2104
rect 1052 2096 1060 2104
rect 940 2036 948 2044
rect 1068 2036 1076 2044
rect 876 1916 884 1924
rect 844 1756 852 1764
rect 876 1736 884 1744
rect 812 1696 820 1704
rect 780 1676 788 1684
rect 796 1416 804 1424
rect 828 1676 836 1684
rect 860 1676 868 1684
rect 828 1476 836 1484
rect 780 1376 788 1384
rect 828 1396 836 1404
rect 844 1376 852 1384
rect 796 1356 804 1364
rect 812 1356 820 1364
rect 780 1336 788 1344
rect 844 1296 852 1304
rect 828 1256 836 1264
rect 812 1156 820 1164
rect 1043 2006 1051 2014
rect 1053 2006 1061 2014
rect 1063 2006 1071 2014
rect 1073 2006 1081 2014
rect 1083 2006 1091 2014
rect 1093 2006 1101 2014
rect 1004 1916 1012 1924
rect 1052 1916 1060 1924
rect 972 1896 980 1904
rect 940 1756 948 1764
rect 940 1716 948 1724
rect 876 1496 884 1504
rect 908 1536 916 1544
rect 940 1536 948 1544
rect 924 1496 932 1504
rect 892 1476 900 1484
rect 892 1336 900 1344
rect 908 1316 916 1324
rect 1004 1876 1012 1884
rect 1036 1876 1044 1884
rect 1052 1876 1060 1884
rect 988 1516 996 1524
rect 972 1476 980 1484
rect 1036 1776 1044 1784
rect 1228 2316 1236 2324
rect 1244 2316 1252 2324
rect 1148 2276 1156 2284
rect 1308 2416 1316 2424
rect 1372 2416 1380 2424
rect 1356 2356 1364 2364
rect 1260 2296 1268 2304
rect 1340 2296 1348 2304
rect 1244 2256 1252 2264
rect 1196 2196 1204 2204
rect 1308 2136 1316 2144
rect 1212 2116 1220 2124
rect 1260 2116 1268 2124
rect 1148 2096 1156 2104
rect 1180 2076 1188 2084
rect 1228 2096 1236 2104
rect 1228 1896 1236 1904
rect 1372 2316 1380 2324
rect 1420 2516 1428 2524
rect 1404 2496 1412 2504
rect 1500 2676 1508 2684
rect 1532 2676 1540 2684
rect 1484 2616 1492 2624
rect 1452 2416 1460 2424
rect 1420 2296 1428 2304
rect 1580 2556 1588 2564
rect 1548 2518 1556 2524
rect 1548 2516 1556 2518
rect 1500 2496 1508 2504
rect 1500 2476 1508 2484
rect 1532 2436 1540 2444
rect 1516 2336 1524 2344
rect 1372 2096 1380 2104
rect 1292 1916 1300 1924
rect 1308 1916 1316 1924
rect 1340 1916 1348 1924
rect 1468 2196 1476 2204
rect 1516 2256 1524 2264
rect 1516 2196 1524 2204
rect 1548 2156 1556 2164
rect 1580 2416 1588 2424
rect 1660 2856 1668 2864
rect 1644 2576 1652 2584
rect 1676 2536 1684 2544
rect 1660 2516 1668 2524
rect 1628 2496 1636 2504
rect 1644 2496 1652 2504
rect 1916 3176 1924 3184
rect 1820 3136 1828 3144
rect 1980 3116 1988 3124
rect 1996 3116 2004 3124
rect 1948 3096 1956 3104
rect 1996 3096 2004 3104
rect 2044 3176 2052 3184
rect 2076 3116 2084 3124
rect 2044 3096 2052 3104
rect 1884 3056 1892 3064
rect 1900 3056 1908 3064
rect 2044 3076 2052 3084
rect 2092 3076 2100 3084
rect 1980 2976 1988 2984
rect 1772 2956 1780 2964
rect 1948 2956 1956 2964
rect 2012 2956 2020 2964
rect 1756 2936 1764 2944
rect 2060 2976 2068 2984
rect 2076 2976 2084 2984
rect 2140 3116 2148 3124
rect 2204 3276 2212 3284
rect 2188 3236 2196 3244
rect 2108 2956 2116 2964
rect 1980 2936 1988 2944
rect 2044 2936 2052 2944
rect 2092 2936 2100 2944
rect 2108 2936 2116 2944
rect 1804 2896 1812 2904
rect 1708 2856 1716 2864
rect 1740 2856 1748 2864
rect 1980 2816 1988 2824
rect 1996 2816 2004 2824
rect 1820 2756 1828 2764
rect 1804 2716 1812 2724
rect 1852 2736 1860 2744
rect 1868 2736 1876 2744
rect 1740 2676 1748 2684
rect 1724 2576 1732 2584
rect 1708 2556 1716 2564
rect 1964 2736 1972 2744
rect 1980 2736 1988 2744
rect 1932 2716 1940 2724
rect 1948 2716 1956 2724
rect 2172 2976 2180 2984
rect 2156 2936 2164 2944
rect 2028 2876 2036 2884
rect 2076 2876 2084 2884
rect 2092 2876 2100 2884
rect 2060 2836 2068 2844
rect 2076 2836 2084 2844
rect 2060 2816 2068 2824
rect 1868 2696 1876 2704
rect 1964 2696 1972 2704
rect 1980 2696 1988 2704
rect 1820 2656 1828 2664
rect 1756 2616 1764 2624
rect 1852 2656 1860 2664
rect 1884 2656 1892 2664
rect 1772 2576 1780 2584
rect 1836 2556 1844 2564
rect 2140 2856 2148 2864
rect 2140 2816 2148 2824
rect 2108 2776 2116 2784
rect 2092 2756 2100 2764
rect 1916 2656 1924 2664
rect 1980 2656 1988 2664
rect 1948 2616 1956 2624
rect 1932 2576 1940 2584
rect 1820 2536 1828 2544
rect 1900 2536 1908 2544
rect 1788 2516 1796 2524
rect 1692 2456 1700 2464
rect 1724 2456 1732 2464
rect 1644 2436 1652 2444
rect 1772 2436 1780 2444
rect 1820 2436 1828 2444
rect 1612 2376 1620 2384
rect 1596 2296 1604 2304
rect 1676 2296 1684 2304
rect 1564 2136 1572 2144
rect 1772 2296 1780 2304
rect 1788 2296 1796 2304
rect 1660 2276 1668 2284
rect 1756 2276 1764 2284
rect 1772 2276 1780 2284
rect 1660 2256 1668 2264
rect 1676 2236 1684 2244
rect 1596 2176 1604 2184
rect 1628 2176 1636 2184
rect 1692 2136 1700 2144
rect 1548 2116 1556 2124
rect 1580 2116 1588 2124
rect 1660 2116 1668 2124
rect 1484 2096 1492 2104
rect 1548 2096 1556 2104
rect 1468 2076 1476 2084
rect 1532 2036 1540 2044
rect 1484 2016 1492 2024
rect 1388 1896 1396 1904
rect 1132 1876 1140 1884
rect 1196 1876 1204 1884
rect 1244 1876 1252 1884
rect 1276 1876 1284 1884
rect 1452 1916 1460 1924
rect 1468 1916 1476 1924
rect 1500 1956 1508 1964
rect 1420 1876 1428 1884
rect 1196 1836 1204 1844
rect 1292 1856 1300 1864
rect 1228 1796 1236 1804
rect 1276 1796 1284 1804
rect 1212 1776 1220 1784
rect 1116 1736 1124 1744
rect 1148 1716 1156 1724
rect 1020 1616 1028 1624
rect 1043 1606 1051 1614
rect 1053 1606 1061 1614
rect 1063 1606 1071 1614
rect 1073 1606 1081 1614
rect 1083 1606 1091 1614
rect 1093 1606 1101 1614
rect 1132 1676 1140 1684
rect 1180 1676 1188 1684
rect 1116 1536 1124 1544
rect 1084 1516 1092 1524
rect 1004 1456 1012 1464
rect 1036 1476 1044 1484
rect 1020 1436 1028 1444
rect 956 1416 964 1424
rect 972 1336 980 1344
rect 940 1316 948 1324
rect 940 1276 948 1284
rect 924 1176 932 1184
rect 796 1136 804 1144
rect 876 1156 884 1164
rect 860 1116 868 1124
rect 844 1096 852 1104
rect 892 1096 900 1104
rect 956 1096 964 1104
rect 780 1076 788 1084
rect 796 1056 804 1064
rect 876 976 884 984
rect 892 936 900 944
rect 828 916 836 924
rect 780 816 788 824
rect 764 696 772 704
rect 748 656 756 664
rect 764 616 772 624
rect 732 556 740 564
rect 684 516 692 524
rect 620 476 628 484
rect 588 456 596 464
rect 572 356 580 364
rect 620 336 628 344
rect 540 296 548 304
rect 444 276 452 284
rect 508 276 516 284
rect 428 196 436 204
rect 444 176 452 184
rect 460 156 468 164
rect 636 296 644 304
rect 828 876 836 884
rect 812 716 820 724
rect 1004 1316 1012 1324
rect 1020 1296 1028 1304
rect 988 1276 996 1284
rect 1052 1456 1060 1464
rect 1116 1496 1124 1504
rect 1084 1416 1092 1424
rect 1100 1416 1108 1424
rect 1100 1356 1108 1364
rect 1340 1836 1348 1844
rect 1324 1796 1332 1804
rect 1516 1836 1524 1844
rect 1580 2076 1588 2084
rect 1564 2016 1572 2024
rect 1564 1936 1572 1944
rect 1548 1916 1556 1924
rect 1548 1856 1556 1864
rect 1468 1796 1476 1804
rect 1324 1736 1332 1744
rect 1356 1718 1364 1724
rect 1356 1716 1364 1718
rect 1468 1716 1476 1724
rect 1292 1696 1300 1704
rect 1244 1636 1252 1644
rect 1212 1496 1220 1504
rect 1228 1496 1236 1504
rect 1276 1596 1284 1604
rect 1404 1676 1412 1684
rect 1356 1556 1364 1564
rect 1356 1536 1364 1544
rect 1308 1516 1316 1524
rect 1340 1516 1348 1524
rect 1436 1556 1444 1564
rect 1404 1516 1412 1524
rect 1420 1516 1428 1524
rect 1164 1436 1172 1444
rect 1180 1436 1188 1444
rect 1132 1356 1140 1364
rect 1100 1316 1108 1324
rect 988 1136 996 1144
rect 972 1056 980 1064
rect 940 1016 948 1024
rect 988 1016 996 1024
rect 1004 1016 1012 1024
rect 988 916 996 924
rect 1068 1236 1076 1244
rect 1043 1206 1051 1214
rect 1053 1206 1061 1214
rect 1063 1206 1071 1214
rect 1073 1206 1081 1214
rect 1083 1206 1091 1214
rect 1093 1206 1101 1214
rect 1116 1196 1124 1204
rect 1148 1336 1156 1344
rect 1180 1296 1188 1304
rect 1132 1176 1140 1184
rect 1116 1156 1124 1164
rect 1100 1096 1108 1104
rect 1084 1076 1092 1084
rect 1100 1056 1108 1064
rect 1116 1056 1124 1064
rect 1036 936 1044 944
rect 1116 916 1124 924
rect 908 856 916 864
rect 1004 856 1012 864
rect 1043 806 1051 814
rect 1053 806 1061 814
rect 1063 806 1071 814
rect 1073 806 1081 814
rect 1083 806 1091 814
rect 1093 806 1101 814
rect 1020 796 1028 804
rect 1004 776 1012 784
rect 924 736 932 744
rect 1052 736 1060 744
rect 1068 736 1076 744
rect 940 716 948 724
rect 1036 716 1044 724
rect 812 656 820 664
rect 844 656 852 664
rect 892 576 900 584
rect 844 556 852 564
rect 892 556 900 564
rect 908 556 916 564
rect 876 536 884 544
rect 1212 1336 1220 1344
rect 1212 1276 1220 1284
rect 1196 1156 1204 1164
rect 1244 1136 1252 1144
rect 1212 1116 1220 1124
rect 1164 1076 1172 1084
rect 1180 1076 1188 1084
rect 1228 1096 1236 1104
rect 1196 1016 1204 1024
rect 1196 976 1204 984
rect 1180 936 1188 944
rect 1228 1016 1236 1024
rect 1164 916 1172 924
rect 1180 916 1188 924
rect 1212 916 1220 924
rect 1148 796 1156 804
rect 1132 716 1140 724
rect 1020 676 1028 684
rect 1004 576 1012 584
rect 1052 536 1060 544
rect 908 496 916 504
rect 924 496 932 504
rect 828 456 836 464
rect 956 496 964 504
rect 988 496 996 504
rect 1068 496 1076 504
rect 972 456 980 464
rect 1020 456 1028 464
rect 1132 456 1140 464
rect 940 376 948 384
rect 956 376 964 384
rect 1116 436 1124 444
rect 1043 406 1051 414
rect 1053 406 1061 414
rect 1063 406 1071 414
rect 1073 406 1081 414
rect 1083 406 1091 414
rect 1093 406 1101 414
rect 956 356 964 364
rect 1020 356 1028 364
rect 988 336 996 344
rect 940 316 948 324
rect 716 276 724 284
rect 764 276 772 284
rect 588 136 596 144
rect 700 236 708 244
rect 236 118 244 124
rect 236 116 244 118
rect 412 116 420 124
rect 540 116 548 124
rect 12 96 20 104
rect 108 96 116 104
rect 300 96 308 104
rect 332 96 340 104
rect 412 96 420 104
rect 796 236 804 244
rect 732 116 740 124
rect 764 116 772 124
rect 940 276 948 284
rect 892 236 900 244
rect 1004 236 1012 244
rect 988 216 996 224
rect 812 136 820 144
rect 844 136 852 144
rect 924 136 932 144
rect 1132 196 1140 204
rect 1196 836 1204 844
rect 1212 836 1220 844
rect 1180 776 1188 784
rect 1196 696 1204 704
rect 1164 596 1172 604
rect 1196 236 1204 244
rect 1196 196 1204 204
rect 1148 156 1156 164
rect 764 96 772 104
rect 1004 96 1012 104
rect 1132 136 1140 144
rect 1180 136 1188 144
rect 1132 116 1140 124
rect 1452 1496 1460 1504
rect 1324 1416 1332 1424
rect 1340 1416 1348 1424
rect 1420 1416 1428 1424
rect 1324 1376 1332 1384
rect 1340 1336 1348 1344
rect 1452 1356 1460 1364
rect 1308 1316 1316 1324
rect 1276 1296 1284 1304
rect 1292 1296 1300 1304
rect 1276 1276 1284 1284
rect 1292 1056 1300 1064
rect 1356 1276 1364 1284
rect 1340 1216 1348 1224
rect 1420 1336 1428 1344
rect 1388 1316 1396 1324
rect 1404 1216 1412 1224
rect 1340 1116 1348 1124
rect 1324 1096 1332 1104
rect 1340 1056 1348 1064
rect 1308 1016 1316 1024
rect 1292 976 1300 984
rect 1324 956 1332 964
rect 1260 896 1268 904
rect 1292 896 1300 904
rect 1308 736 1316 744
rect 1436 1276 1444 1284
rect 1628 2096 1636 2104
rect 1628 2016 1636 2024
rect 1612 1896 1620 1904
rect 1580 1776 1588 1784
rect 1708 1956 1716 1964
rect 1740 2136 1748 2144
rect 1644 1916 1652 1924
rect 1724 1916 1732 1924
rect 1756 2036 1764 2044
rect 1500 1716 1508 1724
rect 1596 1716 1604 1724
rect 1596 1636 1604 1644
rect 1532 1596 1540 1604
rect 1564 1576 1572 1584
rect 1500 1496 1508 1504
rect 1580 1496 1588 1504
rect 1628 1836 1636 1844
rect 1644 1776 1652 1784
rect 1644 1736 1652 1744
rect 1644 1656 1652 1664
rect 1676 1756 1684 1764
rect 1692 1756 1700 1764
rect 1900 2496 1908 2504
rect 1868 2276 1876 2284
rect 1788 2256 1796 2264
rect 1788 2196 1796 2204
rect 1772 1936 1780 1944
rect 1772 1916 1780 1924
rect 1772 1896 1780 1904
rect 1740 1796 1748 1804
rect 1820 2096 1828 2104
rect 1804 1956 1812 1964
rect 1900 2256 1908 2264
rect 1852 2196 1860 2204
rect 1868 2196 1876 2204
rect 1884 2196 1892 2204
rect 1852 2156 1860 2164
rect 1868 2116 1876 2124
rect 1836 2076 1844 2084
rect 1900 2156 1908 2164
rect 1996 2576 2004 2584
rect 1964 2556 1972 2564
rect 1980 2556 1988 2564
rect 1980 2516 1988 2524
rect 1964 2496 1972 2504
rect 1932 2356 1940 2364
rect 1948 2356 1956 2364
rect 1948 2316 1956 2324
rect 1916 2116 1924 2124
rect 1900 2076 1908 2084
rect 1884 2016 1892 2024
rect 2172 2856 2180 2864
rect 2348 3316 2356 3324
rect 2412 3316 2420 3324
rect 2492 3316 2500 3324
rect 2684 3416 2692 3424
rect 2556 3336 2564 3344
rect 2348 3296 2356 3304
rect 2428 3296 2436 3304
rect 2524 3296 2532 3304
rect 2332 3276 2340 3284
rect 2284 3236 2292 3244
rect 2204 3176 2212 3184
rect 2268 3176 2276 3184
rect 2236 3136 2244 3144
rect 2332 3136 2340 3144
rect 2236 3096 2244 3104
rect 2252 3076 2260 3084
rect 2220 3056 2228 3064
rect 2252 3036 2260 3044
rect 2252 2976 2260 2984
rect 2236 2936 2244 2944
rect 2252 2936 2260 2944
rect 2220 2916 2228 2924
rect 2412 3216 2420 3224
rect 2348 3116 2356 3124
rect 2364 3116 2372 3124
rect 2284 2976 2292 2984
rect 2268 2916 2276 2924
rect 2204 2856 2212 2864
rect 2124 2696 2132 2704
rect 2156 2696 2164 2704
rect 2028 2656 2036 2664
rect 2108 2656 2116 2664
rect 2044 2636 2052 2644
rect 2092 2616 2100 2624
rect 2044 2596 2052 2604
rect 2012 2436 2020 2444
rect 2028 2296 2036 2304
rect 1964 2256 1972 2264
rect 1980 2256 1988 2264
rect 2012 2276 2020 2284
rect 1932 2036 1940 2044
rect 1916 1996 1924 2004
rect 1948 1996 1956 2004
rect 1868 1956 1876 1964
rect 1900 1956 1908 1964
rect 1916 1956 1924 1964
rect 1836 1916 1844 1924
rect 1852 1916 1860 1924
rect 1804 1856 1812 1864
rect 1820 1836 1828 1844
rect 1804 1696 1812 1704
rect 1660 1636 1668 1644
rect 1676 1616 1684 1624
rect 1644 1596 1652 1604
rect 1644 1496 1652 1504
rect 1692 1556 1700 1564
rect 1708 1556 1716 1564
rect 1756 1556 1764 1564
rect 1708 1516 1716 1524
rect 1740 1516 1748 1524
rect 1708 1496 1716 1504
rect 1724 1496 1732 1504
rect 1516 1376 1524 1384
rect 1500 1356 1508 1364
rect 1612 1316 1620 1324
rect 1484 1276 1492 1284
rect 1516 1276 1524 1284
rect 1468 1216 1476 1224
rect 1372 1136 1380 1144
rect 1420 1136 1428 1144
rect 1372 1076 1380 1084
rect 1356 976 1364 984
rect 1420 1036 1428 1044
rect 1388 976 1396 984
rect 1388 936 1396 944
rect 1340 916 1348 924
rect 1372 916 1380 924
rect 1388 896 1396 904
rect 1404 896 1412 904
rect 1356 816 1364 824
rect 1404 736 1412 744
rect 1340 716 1348 724
rect 1276 696 1284 704
rect 1324 696 1332 704
rect 1340 696 1348 704
rect 1260 676 1268 684
rect 1244 656 1252 664
rect 1228 576 1236 584
rect 1356 676 1364 684
rect 1420 676 1428 684
rect 1324 656 1332 664
rect 1340 616 1348 624
rect 1452 916 1460 924
rect 1484 1176 1492 1184
rect 1484 1156 1492 1164
rect 1596 1276 1604 1284
rect 1580 1196 1588 1204
rect 1564 1156 1572 1164
rect 1580 1156 1588 1164
rect 1548 1136 1556 1144
rect 1596 1136 1604 1144
rect 1516 1102 1524 1104
rect 1516 1096 1524 1102
rect 1516 1056 1524 1064
rect 1484 1016 1492 1024
rect 1500 976 1508 984
rect 1580 976 1588 984
rect 1612 1116 1620 1124
rect 1612 1096 1620 1104
rect 1676 1416 1684 1424
rect 1724 1416 1732 1424
rect 1724 1376 1732 1384
rect 1740 1376 1748 1384
rect 1740 1336 1748 1344
rect 1804 1596 1812 1604
rect 1852 1816 1860 1824
rect 1836 1736 1844 1744
rect 1852 1576 1860 1584
rect 1852 1556 1860 1564
rect 1820 1516 1828 1524
rect 1836 1516 1844 1524
rect 1836 1496 1844 1504
rect 1804 1416 1812 1424
rect 1996 2136 2004 2144
rect 1996 1996 2004 2004
rect 1980 1956 1988 1964
rect 1996 1956 2004 1964
rect 2076 2576 2084 2584
rect 2060 2496 2068 2504
rect 2060 2416 2068 2424
rect 2060 2276 2068 2284
rect 2028 2256 2036 2264
rect 2108 2576 2116 2584
rect 2140 2656 2148 2664
rect 2332 2936 2340 2944
rect 2380 2936 2388 2944
rect 2316 2916 2324 2924
rect 2348 2896 2356 2904
rect 2636 3376 2644 3384
rect 2620 3356 2628 3364
rect 2588 3276 2596 3284
rect 2620 3276 2628 3284
rect 2444 3236 2452 3244
rect 2524 3196 2532 3204
rect 2604 3116 2612 3124
rect 2444 3076 2452 3084
rect 2476 3076 2484 3084
rect 2428 3016 2436 3024
rect 2444 3016 2452 3024
rect 2492 3036 2500 3044
rect 2476 2996 2484 3004
rect 2444 2936 2452 2944
rect 2460 2936 2468 2944
rect 2444 2916 2452 2924
rect 2524 3016 2532 3024
rect 2508 2976 2516 2984
rect 2547 3006 2555 3014
rect 2557 3006 2565 3014
rect 2567 3006 2575 3014
rect 2577 3006 2585 3014
rect 2587 3006 2595 3014
rect 2597 3006 2605 3014
rect 2604 2936 2612 2944
rect 2252 2796 2260 2804
rect 2220 2756 2228 2764
rect 2268 2776 2276 2784
rect 2204 2736 2212 2744
rect 2188 2616 2196 2624
rect 2236 2716 2244 2724
rect 2252 2696 2260 2704
rect 2156 2576 2164 2584
rect 2172 2576 2180 2584
rect 2204 2576 2212 2584
rect 2140 2536 2148 2544
rect 2188 2556 2196 2564
rect 2204 2496 2212 2504
rect 2252 2516 2260 2524
rect 2284 2736 2292 2744
rect 2316 2796 2324 2804
rect 2460 2796 2468 2804
rect 2396 2776 2404 2784
rect 2332 2716 2340 2724
rect 2380 2716 2388 2724
rect 2428 2756 2436 2764
rect 2316 2576 2324 2584
rect 2364 2656 2372 2664
rect 2364 2636 2372 2644
rect 2332 2536 2340 2544
rect 2348 2536 2356 2544
rect 2300 2516 2308 2524
rect 2268 2496 2276 2504
rect 2252 2476 2260 2484
rect 2268 2476 2276 2484
rect 2188 2436 2196 2444
rect 2220 2436 2228 2444
rect 2236 2436 2244 2444
rect 2108 2296 2116 2304
rect 2172 2356 2180 2364
rect 2156 2296 2164 2304
rect 2188 2296 2196 2304
rect 2204 2296 2212 2304
rect 2236 2296 2244 2304
rect 2140 2276 2148 2284
rect 2092 2196 2100 2204
rect 2076 2176 2084 2184
rect 2076 2156 2084 2164
rect 2060 2136 2068 2144
rect 2124 2196 2132 2204
rect 2092 2116 2100 2124
rect 2044 1996 2052 2004
rect 2028 1956 2036 1964
rect 2060 1956 2068 1964
rect 1964 1916 1972 1924
rect 1884 1896 1892 1904
rect 1964 1896 1972 1904
rect 1884 1836 1892 1844
rect 1948 1836 1956 1844
rect 1948 1816 1956 1824
rect 1884 1776 1892 1784
rect 1900 1716 1908 1724
rect 1932 1716 1940 1724
rect 1916 1696 1924 1704
rect 1900 1596 1908 1604
rect 1948 1656 1956 1664
rect 1948 1576 1956 1584
rect 1916 1556 1924 1564
rect 1884 1516 1892 1524
rect 1900 1496 1908 1504
rect 1948 1496 1956 1504
rect 1916 1456 1924 1464
rect 1884 1416 1892 1424
rect 1788 1376 1796 1384
rect 1804 1356 1812 1364
rect 1868 1356 1876 1364
rect 1708 1316 1716 1324
rect 1740 1316 1748 1324
rect 1772 1316 1780 1324
rect 1788 1316 1796 1324
rect 1676 1296 1684 1304
rect 1660 1116 1668 1124
rect 1692 1116 1700 1124
rect 1836 1296 1844 1304
rect 1788 1236 1796 1244
rect 1804 1236 1812 1244
rect 1772 1196 1780 1204
rect 1756 1116 1764 1124
rect 1740 1096 1748 1104
rect 1660 1056 1668 1064
rect 1516 916 1524 924
rect 1596 916 1604 924
rect 1532 896 1540 904
rect 1596 896 1604 904
rect 1628 976 1636 984
rect 1660 976 1668 984
rect 1660 956 1668 964
rect 1676 956 1684 964
rect 1644 936 1652 944
rect 1628 876 1636 884
rect 1532 856 1540 864
rect 1468 696 1476 704
rect 1516 696 1524 704
rect 1580 716 1588 724
rect 1260 516 1268 524
rect 1212 136 1220 144
rect 1196 96 1204 104
rect 1036 36 1044 44
rect 1132 36 1140 44
rect 1116 16 1124 24
rect 1043 6 1051 14
rect 1053 6 1061 14
rect 1063 6 1071 14
rect 1073 6 1081 14
rect 1083 6 1091 14
rect 1093 6 1101 14
rect 1164 16 1172 24
rect 1244 396 1252 404
rect 1292 436 1300 444
rect 1324 436 1332 444
rect 1340 376 1348 384
rect 1324 316 1332 324
rect 1340 316 1348 324
rect 1420 516 1428 524
rect 1356 296 1364 304
rect 1324 276 1332 284
rect 1356 276 1364 284
rect 1244 236 1252 244
rect 1308 236 1316 244
rect 1260 176 1268 184
rect 1292 156 1300 164
rect 1596 696 1604 704
rect 1628 696 1636 704
rect 1660 876 1668 884
rect 1788 1096 1796 1104
rect 1724 1056 1732 1064
rect 1772 1056 1780 1064
rect 1708 1036 1716 1044
rect 1724 1036 1732 1044
rect 1724 976 1732 984
rect 1740 976 1748 984
rect 1756 956 1764 964
rect 1756 936 1764 944
rect 1708 896 1716 904
rect 1772 916 1780 924
rect 1692 876 1700 884
rect 1740 836 1748 844
rect 1676 796 1684 804
rect 1692 796 1700 804
rect 1660 716 1668 724
rect 1740 756 1748 764
rect 1756 756 1764 764
rect 1660 676 1668 684
rect 1708 656 1716 664
rect 1596 636 1604 644
rect 1660 636 1668 644
rect 1580 616 1588 624
rect 1596 576 1604 584
rect 1548 536 1556 544
rect 1628 536 1636 544
rect 1756 676 1764 684
rect 1788 696 1796 704
rect 1820 1136 1828 1144
rect 1852 1136 1860 1144
rect 1836 1116 1844 1124
rect 1948 1416 1956 1424
rect 2044 1916 2052 1924
rect 1996 1816 2004 1824
rect 2012 1796 2020 1804
rect 1980 1776 1988 1784
rect 2076 1916 2084 1924
rect 2076 1876 2084 1884
rect 2156 2216 2164 2224
rect 2172 2196 2180 2204
rect 2204 2216 2212 2224
rect 2220 2196 2228 2204
rect 2284 2296 2292 2304
rect 2316 2436 2324 2444
rect 2316 2416 2324 2424
rect 2268 2276 2276 2284
rect 2300 2276 2308 2284
rect 2300 2256 2308 2264
rect 2284 2156 2292 2164
rect 2220 2136 2228 2144
rect 2252 2136 2260 2144
rect 2188 2116 2196 2124
rect 2284 2118 2292 2124
rect 2284 2116 2292 2118
rect 2220 2076 2228 2084
rect 2204 2056 2212 2064
rect 2172 1996 2180 2004
rect 2140 1976 2148 1984
rect 2172 1976 2180 1984
rect 2108 1956 2116 1964
rect 2188 1956 2196 1964
rect 2172 1916 2180 1924
rect 2204 1916 2212 1924
rect 2156 1896 2164 1904
rect 2140 1876 2148 1884
rect 2140 1776 2148 1784
rect 2124 1756 2132 1764
rect 2092 1736 2100 1744
rect 1980 1656 1988 1664
rect 2028 1716 2036 1724
rect 2028 1696 2036 1704
rect 1996 1596 2004 1604
rect 2012 1596 2020 1604
rect 1980 1576 1988 1584
rect 1996 1536 2004 1544
rect 1980 1496 1988 1504
rect 2012 1516 2020 1524
rect 2012 1456 2020 1464
rect 1980 1416 1988 1424
rect 1932 1376 1940 1384
rect 1884 1336 1892 1344
rect 1916 1336 1924 1344
rect 1932 1336 1940 1344
rect 1884 1136 1892 1144
rect 1884 1116 1892 1124
rect 1868 1076 1876 1084
rect 1836 1056 1844 1064
rect 1852 1036 1860 1044
rect 1964 1316 1972 1324
rect 1932 1136 1940 1144
rect 1916 1096 1924 1104
rect 1900 1076 1908 1084
rect 1820 936 1828 944
rect 1868 936 1876 944
rect 1996 1376 2004 1384
rect 1980 1256 1988 1264
rect 1996 1256 2004 1264
rect 2060 1656 2068 1664
rect 2044 1556 2052 1564
rect 2076 1456 2084 1464
rect 2060 1376 2068 1384
rect 2044 1336 2052 1344
rect 2348 2356 2356 2364
rect 2412 2616 2420 2624
rect 2396 2596 2404 2604
rect 2380 2556 2388 2564
rect 2380 2476 2388 2484
rect 2396 2476 2404 2484
rect 2444 2656 2452 2664
rect 2492 2796 2500 2804
rect 2492 2776 2500 2784
rect 2572 2856 2580 2864
rect 2508 2736 2516 2744
rect 2508 2716 2516 2724
rect 2524 2676 2532 2684
rect 2924 3376 2932 3384
rect 2796 3356 2804 3364
rect 2844 3356 2852 3364
rect 2748 3336 2756 3344
rect 2780 3336 2788 3344
rect 2892 3336 2900 3344
rect 2732 3316 2740 3324
rect 2796 3316 2804 3324
rect 2860 3316 2868 3324
rect 2684 3296 2692 3304
rect 2748 3276 2756 3284
rect 2684 3196 2692 3204
rect 2668 3136 2676 3144
rect 2684 3136 2692 3144
rect 2636 3036 2644 3044
rect 2636 2956 2644 2964
rect 2684 3036 2692 3044
rect 2652 2936 2660 2944
rect 2636 2856 2644 2864
rect 2668 2896 2676 2904
rect 2732 3076 2740 3084
rect 2716 3016 2724 3024
rect 2700 2996 2708 3004
rect 2700 2956 2708 2964
rect 2716 2956 2724 2964
rect 2684 2856 2692 2864
rect 2732 2836 2740 2844
rect 2652 2756 2660 2764
rect 2620 2636 2628 2644
rect 2547 2606 2555 2614
rect 2557 2606 2565 2614
rect 2567 2606 2575 2614
rect 2577 2606 2585 2614
rect 2587 2606 2595 2614
rect 2597 2606 2605 2614
rect 2508 2596 2516 2604
rect 2588 2556 2596 2564
rect 2604 2556 2612 2564
rect 2492 2496 2500 2504
rect 2428 2476 2436 2484
rect 2444 2476 2452 2484
rect 2460 2476 2468 2484
rect 2412 2416 2420 2424
rect 2380 2356 2388 2364
rect 2364 2296 2372 2304
rect 2316 2236 2324 2244
rect 2348 2256 2356 2264
rect 2332 2196 2340 2204
rect 2492 2436 2500 2444
rect 2524 2436 2532 2444
rect 2492 2356 2500 2364
rect 2508 2316 2516 2324
rect 2492 2276 2500 2284
rect 2476 2256 2484 2264
rect 2492 2256 2500 2264
rect 2460 2236 2468 2244
rect 2396 2216 2404 2224
rect 2428 2216 2436 2224
rect 2412 2196 2420 2204
rect 2444 2196 2452 2204
rect 2476 2196 2484 2204
rect 2492 2196 2500 2204
rect 2380 2156 2388 2164
rect 2492 2156 2500 2164
rect 2556 2516 2564 2524
rect 2572 2516 2580 2524
rect 2636 2616 2644 2624
rect 2700 2696 2708 2704
rect 2668 2616 2676 2624
rect 2700 2556 2708 2564
rect 2716 2556 2724 2564
rect 2668 2516 2676 2524
rect 2668 2496 2676 2504
rect 2572 2476 2580 2484
rect 2588 2476 2596 2484
rect 2652 2476 2660 2484
rect 2652 2436 2660 2444
rect 2540 2336 2548 2344
rect 2540 2316 2548 2324
rect 2604 2276 2612 2284
rect 2540 2256 2548 2264
rect 2524 2216 2532 2224
rect 2620 2216 2628 2224
rect 2547 2206 2555 2214
rect 2557 2206 2565 2214
rect 2567 2206 2575 2214
rect 2577 2206 2585 2214
rect 2587 2206 2595 2214
rect 2597 2206 2605 2214
rect 2524 2136 2532 2144
rect 2332 2076 2340 2084
rect 2300 2056 2308 2064
rect 2316 2056 2324 2064
rect 2300 1996 2308 2004
rect 2252 1956 2260 1964
rect 2284 1916 2292 1924
rect 2236 1856 2244 1864
rect 2316 1956 2324 1964
rect 2316 1916 2324 1924
rect 2268 1836 2276 1844
rect 2284 1836 2292 1844
rect 2428 2076 2436 2084
rect 2476 2076 2484 2084
rect 2492 2076 2500 2084
rect 2412 1976 2420 1984
rect 2428 1976 2436 1984
rect 2380 1956 2388 1964
rect 2348 1896 2356 1904
rect 2332 1836 2340 1844
rect 2348 1836 2356 1844
rect 2396 1916 2404 1924
rect 2412 1896 2420 1904
rect 2444 1896 2452 1904
rect 2476 1996 2484 2004
rect 2508 1976 2516 1984
rect 2492 1916 2500 1924
rect 2492 1896 2500 1904
rect 2524 1956 2532 1964
rect 2652 2256 2660 2264
rect 2652 2156 2660 2164
rect 2716 2516 2724 2524
rect 2732 2516 2740 2524
rect 2700 2496 2708 2504
rect 2684 2416 2692 2424
rect 2684 2316 2692 2324
rect 2716 2436 2724 2444
rect 2764 3196 2772 3204
rect 2796 3136 2804 3144
rect 2828 3136 2836 3144
rect 2940 3356 2948 3364
rect 3356 3356 3364 3364
rect 3468 3356 3476 3364
rect 3676 3356 3684 3364
rect 3036 3336 3044 3344
rect 3132 3336 3140 3344
rect 3324 3336 3332 3344
rect 3628 3336 3636 3344
rect 3788 3336 3796 3344
rect 2956 3316 2964 3324
rect 3052 3316 3060 3324
rect 2972 3296 2980 3304
rect 2988 3276 2996 3284
rect 3020 3236 3028 3244
rect 2924 3116 2932 3124
rect 2764 3096 2772 3104
rect 2908 3096 2916 3104
rect 2780 3076 2788 3084
rect 2828 3076 2836 3084
rect 2828 2956 2836 2964
rect 2796 2916 2804 2924
rect 2812 2896 2820 2904
rect 2780 2856 2788 2864
rect 2764 2736 2772 2744
rect 2924 3076 2932 3084
rect 2892 3016 2900 3024
rect 2956 3116 2964 3124
rect 3004 3116 3012 3124
rect 2988 3096 2996 3104
rect 2988 3076 2996 3084
rect 2908 2956 2916 2964
rect 3036 3136 3044 3144
rect 3020 2996 3028 3004
rect 2876 2876 2884 2884
rect 2972 2936 2980 2944
rect 3084 3276 3092 3284
rect 3100 3236 3108 3244
rect 3068 3056 3076 3064
rect 3036 2916 3044 2924
rect 2972 2896 2980 2904
rect 2844 2856 2852 2864
rect 2860 2856 2868 2864
rect 2940 2856 2948 2864
rect 2844 2756 2852 2764
rect 2908 2736 2916 2744
rect 2844 2716 2852 2724
rect 2860 2716 2868 2724
rect 2908 2716 2916 2724
rect 2924 2716 2932 2724
rect 2860 2696 2868 2704
rect 2988 2856 2996 2864
rect 3164 3276 3172 3284
rect 3388 3316 3396 3324
rect 3436 3316 3444 3324
rect 3452 3316 3460 3324
rect 3660 3316 3668 3324
rect 3340 3276 3348 3284
rect 3324 3176 3332 3184
rect 3228 3136 3236 3144
rect 3292 3136 3300 3144
rect 3132 3116 3140 3124
rect 3164 3102 3172 3104
rect 3164 3096 3172 3102
rect 3260 3096 3268 3104
rect 3308 3096 3316 3104
rect 3132 3076 3140 3084
rect 3276 3076 3284 3084
rect 3148 3056 3156 3064
rect 3052 2896 3060 2904
rect 3068 2896 3076 2904
rect 3276 3036 3284 3044
rect 3212 2956 3220 2964
rect 3244 2936 3252 2944
rect 3228 2916 3236 2924
rect 3292 2956 3300 2964
rect 3292 2936 3300 2944
rect 2956 2836 2964 2844
rect 2972 2836 2980 2844
rect 3004 2836 3012 2844
rect 3020 2836 3028 2844
rect 3068 2856 3076 2864
rect 2988 2736 2996 2744
rect 3020 2736 3028 2744
rect 3052 2736 3060 2744
rect 2956 2716 2964 2724
rect 3100 2836 3108 2844
rect 3132 2836 3140 2844
rect 3084 2776 3092 2784
rect 3116 2776 3124 2784
rect 3084 2736 3092 2744
rect 3100 2736 3108 2744
rect 2908 2676 2916 2684
rect 3004 2676 3012 2684
rect 2972 2636 2980 2644
rect 2796 2516 2804 2524
rect 2764 2416 2772 2424
rect 2668 2136 2676 2144
rect 2636 2116 2644 2124
rect 2556 1996 2564 2004
rect 2380 1856 2388 1864
rect 2204 1816 2212 1824
rect 2236 1816 2244 1824
rect 2300 1816 2308 1824
rect 2348 1816 2356 1824
rect 2364 1816 2372 1824
rect 2460 1876 2468 1884
rect 2492 1876 2500 1884
rect 2444 1836 2452 1844
rect 2172 1796 2180 1804
rect 2252 1776 2260 1784
rect 2284 1776 2292 1784
rect 2204 1736 2212 1744
rect 2156 1716 2164 1724
rect 2172 1716 2180 1724
rect 2092 1316 2100 1324
rect 2172 1596 2180 1604
rect 2124 1576 2132 1584
rect 2172 1576 2180 1584
rect 2220 1716 2228 1724
rect 2220 1636 2228 1644
rect 2252 1656 2260 1664
rect 2236 1596 2244 1604
rect 2220 1536 2228 1544
rect 2236 1516 2244 1524
rect 2252 1516 2260 1524
rect 2316 1736 2324 1744
rect 2492 1796 2500 1804
rect 2460 1776 2468 1784
rect 2476 1776 2484 1784
rect 2508 1776 2516 1784
rect 2636 1996 2644 2004
rect 2588 1836 2596 1844
rect 2547 1806 2555 1814
rect 2557 1806 2565 1814
rect 2567 1806 2575 1814
rect 2577 1806 2585 1814
rect 2587 1806 2595 1814
rect 2597 1806 2605 1814
rect 2556 1776 2564 1784
rect 2316 1696 2324 1704
rect 2348 1636 2356 1644
rect 2316 1576 2324 1584
rect 2300 1496 2308 1504
rect 2188 1356 2196 1364
rect 2028 1236 2036 1244
rect 2044 1236 2052 1244
rect 2012 1116 2020 1124
rect 2092 1256 2100 1264
rect 2060 1136 2068 1144
rect 1948 1096 1956 1104
rect 1964 1096 1972 1104
rect 2044 1096 2052 1104
rect 2060 1102 2068 1104
rect 2060 1096 2068 1102
rect 1964 1016 1972 1024
rect 1852 916 1860 924
rect 1868 896 1876 904
rect 1948 956 1956 964
rect 1980 956 1988 964
rect 1932 916 1940 924
rect 1948 916 1956 924
rect 1996 896 2004 904
rect 1964 716 1972 724
rect 1916 676 1924 684
rect 1836 656 1844 664
rect 1884 656 1892 664
rect 1788 636 1796 644
rect 1772 616 1780 624
rect 1740 596 1748 604
rect 1724 576 1732 584
rect 1852 556 1860 564
rect 1868 536 1876 544
rect 1516 516 1524 524
rect 1612 516 1620 524
rect 1580 476 1588 484
rect 1548 456 1556 464
rect 1548 276 1556 284
rect 1404 256 1412 264
rect 1356 176 1364 184
rect 1372 176 1380 184
rect 1420 176 1428 184
rect 1580 256 1588 264
rect 1612 316 1620 324
rect 1980 702 1988 704
rect 1980 696 1988 702
rect 2108 1196 2116 1204
rect 2156 1316 2164 1324
rect 2156 1256 2164 1264
rect 2140 1136 2148 1144
rect 2124 1116 2132 1124
rect 2156 1116 2164 1124
rect 2124 1096 2132 1104
rect 2092 1036 2100 1044
rect 2140 1036 2148 1044
rect 2060 1016 2068 1024
rect 2108 976 2116 984
rect 2092 936 2100 944
rect 2028 916 2036 924
rect 2076 916 2084 924
rect 2092 796 2100 804
rect 2060 696 2068 704
rect 2076 696 2084 704
rect 2188 1316 2196 1324
rect 2188 1196 2196 1204
rect 2284 1456 2292 1464
rect 2268 1396 2276 1404
rect 2220 1296 2228 1304
rect 2220 1196 2228 1204
rect 2204 1136 2212 1144
rect 2188 1076 2196 1084
rect 2156 1016 2164 1024
rect 2140 956 2148 964
rect 2156 936 2164 944
rect 2188 896 2196 904
rect 2236 1076 2244 1084
rect 2284 1376 2292 1384
rect 2332 1516 2340 1524
rect 2492 1736 2500 1744
rect 2524 1736 2532 1744
rect 2540 1736 2548 1744
rect 2572 1736 2580 1744
rect 2588 1736 2596 1744
rect 2396 1636 2404 1644
rect 2396 1596 2404 1604
rect 2460 1716 2468 1724
rect 2428 1636 2436 1644
rect 2444 1636 2452 1644
rect 2428 1596 2436 1604
rect 2412 1576 2420 1584
rect 2460 1596 2468 1604
rect 2492 1596 2500 1604
rect 2460 1576 2468 1584
rect 2636 1916 2644 1924
rect 2716 2296 2724 2304
rect 2748 2316 2756 2324
rect 2748 2276 2756 2284
rect 2748 2256 2756 2264
rect 2700 2236 2708 2244
rect 2716 2136 2724 2144
rect 2924 2516 2932 2524
rect 2956 2516 2964 2524
rect 2844 2476 2852 2484
rect 2860 2476 2868 2484
rect 2940 2476 2948 2484
rect 2844 2416 2852 2424
rect 2828 2336 2836 2344
rect 2812 2316 2820 2324
rect 2796 2296 2804 2304
rect 2812 2276 2820 2284
rect 2780 2256 2788 2264
rect 2780 2156 2788 2164
rect 2844 2316 2852 2324
rect 2924 2316 2932 2324
rect 3036 2656 3044 2664
rect 3052 2656 3060 2664
rect 3068 2656 3076 2664
rect 3020 2596 3028 2604
rect 3036 2596 3044 2604
rect 3004 2516 3012 2524
rect 3036 2516 3044 2524
rect 3004 2476 3012 2484
rect 2988 2316 2996 2324
rect 2860 2236 2868 2244
rect 2876 2236 2884 2244
rect 2828 2216 2836 2224
rect 2876 2216 2884 2224
rect 2940 2256 2948 2264
rect 3020 2416 3028 2424
rect 3052 2496 3060 2504
rect 3132 2716 3140 2724
rect 3180 2896 3188 2904
rect 3228 2896 3236 2904
rect 3164 2776 3172 2784
rect 3148 2696 3156 2704
rect 3196 2736 3204 2744
rect 3180 2716 3188 2724
rect 3196 2696 3204 2704
rect 3132 2636 3140 2644
rect 3132 2536 3140 2544
rect 3276 2856 3284 2864
rect 3260 2716 3268 2724
rect 3436 3276 3444 3284
rect 3388 3256 3396 3264
rect 3372 3096 3380 3104
rect 3324 3076 3332 3084
rect 3324 3036 3332 3044
rect 3340 3016 3348 3024
rect 3372 3016 3380 3024
rect 3356 2896 3364 2904
rect 3404 3136 3412 3144
rect 3436 3136 3444 3144
rect 3420 3096 3428 3104
rect 3580 3276 3588 3284
rect 3452 3076 3460 3084
rect 3580 3076 3588 3084
rect 3420 3036 3428 3044
rect 3452 3036 3460 3044
rect 3468 3016 3476 3024
rect 3500 2996 3508 3004
rect 3644 3036 3652 3044
rect 3692 3276 3700 3284
rect 3820 3296 3828 3304
rect 3932 3316 3940 3324
rect 3932 3296 3940 3304
rect 3884 3276 3892 3284
rect 3740 3136 3748 3144
rect 3676 3096 3684 3104
rect 3724 3096 3732 3104
rect 3676 3076 3684 3084
rect 4476 3416 4484 3424
rect 3980 3396 3988 3404
rect 4300 3376 4308 3384
rect 4396 3376 4404 3384
rect 4108 3336 4116 3344
rect 4236 3336 4244 3344
rect 4380 3336 4388 3344
rect 3980 3316 3988 3324
rect 3964 3296 3972 3304
rect 3980 3276 3988 3284
rect 3964 3256 3972 3264
rect 3884 3102 3892 3104
rect 3884 3096 3892 3102
rect 4172 3316 4180 3324
rect 4188 3316 4196 3324
rect 4252 3316 4260 3324
rect 4012 3276 4020 3284
rect 4156 3296 4164 3304
rect 4300 3296 4308 3304
rect 4140 3276 4148 3284
rect 4172 3276 4180 3284
rect 4268 3276 4276 3284
rect 3996 3256 4004 3264
rect 4124 3256 4132 3264
rect 3996 3216 4004 3224
rect 4051 3206 4059 3214
rect 4061 3206 4069 3214
rect 4071 3206 4079 3214
rect 4081 3206 4089 3214
rect 4091 3206 4099 3214
rect 4101 3206 4109 3214
rect 3996 3196 4004 3204
rect 3996 3136 4004 3144
rect 4156 3136 4164 3144
rect 3820 3076 3828 3084
rect 3948 3076 3956 3084
rect 3692 2996 3700 3004
rect 3628 2956 3636 2964
rect 3660 2956 3668 2964
rect 3404 2916 3412 2924
rect 3612 2916 3620 2924
rect 3388 2856 3396 2864
rect 3420 2856 3428 2864
rect 3340 2836 3348 2844
rect 3308 2736 3316 2744
rect 3404 2736 3412 2744
rect 3388 2696 3396 2704
rect 3212 2676 3220 2684
rect 3100 2436 3108 2444
rect 3116 2436 3124 2444
rect 3052 2416 3060 2424
rect 3244 2656 3252 2664
rect 3308 2636 3316 2644
rect 3324 2536 3332 2544
rect 3260 2518 3268 2524
rect 3260 2516 3268 2518
rect 3372 2516 3380 2524
rect 3356 2496 3364 2504
rect 3356 2436 3364 2444
rect 3036 2376 3044 2384
rect 3052 2336 3060 2344
rect 3084 2336 3092 2344
rect 3180 2336 3188 2344
rect 3244 2296 3252 2304
rect 3020 2276 3028 2284
rect 3036 2276 3044 2284
rect 2908 2216 2916 2224
rect 2892 2196 2900 2204
rect 2892 2156 2900 2164
rect 2812 2136 2820 2144
rect 2828 2136 2836 2144
rect 2700 2076 2708 2084
rect 2748 2016 2756 2024
rect 2684 1976 2692 1984
rect 2652 1896 2660 1904
rect 2636 1816 2644 1824
rect 2716 1996 2724 2004
rect 2732 1996 2740 2004
rect 2700 1916 2708 1924
rect 2652 1796 2660 1804
rect 2636 1776 2644 1784
rect 2684 1776 2692 1784
rect 2748 1916 2756 1924
rect 2748 1896 2756 1904
rect 2748 1816 2756 1824
rect 2748 1776 2756 1784
rect 2620 1676 2628 1684
rect 2668 1676 2676 1684
rect 2588 1656 2596 1664
rect 2604 1656 2612 1664
rect 2716 1756 2724 1764
rect 2700 1696 2708 1704
rect 2572 1636 2580 1644
rect 2556 1516 2564 1524
rect 2588 1516 2596 1524
rect 2492 1496 2500 1504
rect 2652 1616 2660 1624
rect 2620 1576 2628 1584
rect 2444 1436 2452 1444
rect 2428 1376 2436 1384
rect 2300 1276 2308 1284
rect 2316 1276 2324 1284
rect 2284 1256 2292 1264
rect 2300 1256 2308 1264
rect 2412 1236 2420 1244
rect 2428 1236 2436 1244
rect 2380 1216 2388 1224
rect 2332 1116 2340 1124
rect 2364 1096 2372 1104
rect 2284 1076 2292 1084
rect 2268 1056 2276 1064
rect 2364 1056 2372 1064
rect 2220 956 2228 964
rect 2284 1016 2292 1024
rect 2252 976 2260 984
rect 2300 956 2308 964
rect 2220 916 2228 924
rect 2300 916 2308 924
rect 2268 856 2276 864
rect 2204 836 2212 844
rect 2236 836 2244 844
rect 2300 836 2308 844
rect 2172 796 2180 804
rect 2108 716 2116 724
rect 2156 716 2164 724
rect 2236 716 2244 724
rect 2332 916 2340 924
rect 2604 1456 2612 1464
rect 2508 1436 2516 1444
rect 2492 1416 2500 1424
rect 2508 1396 2516 1404
rect 2476 1376 2484 1384
rect 2492 1376 2500 1384
rect 2547 1406 2555 1414
rect 2557 1406 2565 1414
rect 2567 1406 2575 1414
rect 2577 1406 2585 1414
rect 2587 1406 2595 1414
rect 2597 1406 2605 1414
rect 2604 1336 2612 1344
rect 2460 1296 2468 1304
rect 2588 1276 2596 1284
rect 2604 1276 2612 1284
rect 2524 1256 2532 1264
rect 2460 1196 2468 1204
rect 2476 1196 2484 1204
rect 2396 1116 2404 1124
rect 2460 1176 2468 1184
rect 2412 1076 2420 1084
rect 2460 1116 2468 1124
rect 2476 1116 2484 1124
rect 2460 1096 2468 1104
rect 2604 1102 2612 1104
rect 2604 1096 2612 1102
rect 2700 1616 2708 1624
rect 2844 2096 2852 2104
rect 2860 2096 2868 2104
rect 2828 2016 2836 2024
rect 2780 1996 2788 2004
rect 2812 1996 2820 2004
rect 2876 2016 2884 2024
rect 2876 1976 2884 1984
rect 2892 1976 2900 1984
rect 2844 1956 2852 1964
rect 2780 1836 2788 1844
rect 2764 1756 2772 1764
rect 2700 1496 2708 1504
rect 2764 1496 2772 1504
rect 2652 1476 2660 1484
rect 2636 1456 2644 1464
rect 2716 1476 2724 1484
rect 2668 1436 2676 1444
rect 2668 1396 2676 1404
rect 2652 1356 2660 1364
rect 2844 1876 2852 1884
rect 2796 1816 2804 1824
rect 2844 1836 2852 1844
rect 2844 1796 2852 1804
rect 2876 1736 2884 1744
rect 3084 2156 3092 2164
rect 3100 2156 3108 2164
rect 3052 2136 3060 2144
rect 3132 2276 3140 2284
rect 3148 2236 3156 2244
rect 3164 2236 3172 2244
rect 3228 2236 3236 2244
rect 3196 2156 3204 2164
rect 3260 2256 3268 2264
rect 3004 2096 3012 2104
rect 3020 2096 3028 2104
rect 3100 2096 3108 2104
rect 3116 2096 3124 2104
rect 3180 2096 3188 2104
rect 2988 2036 2996 2044
rect 3020 2036 3028 2044
rect 2988 1996 2996 2004
rect 3036 1976 3044 1984
rect 3084 1976 3092 1984
rect 3068 1936 3076 1944
rect 2924 1896 2932 1904
rect 2972 1896 2980 1904
rect 2924 1816 2932 1824
rect 2924 1796 2932 1804
rect 2940 1796 2948 1804
rect 2908 1776 2916 1784
rect 2972 1856 2980 1864
rect 2956 1776 2964 1784
rect 2844 1696 2852 1704
rect 2844 1676 2852 1684
rect 2860 1676 2868 1684
rect 2892 1676 2900 1684
rect 2828 1616 2836 1624
rect 2812 1576 2820 1584
rect 2796 1496 2804 1504
rect 2844 1496 2852 1504
rect 2796 1476 2804 1484
rect 2684 1376 2692 1384
rect 2716 1376 2724 1384
rect 2780 1376 2788 1384
rect 2700 1356 2708 1364
rect 2700 1336 2708 1344
rect 2652 1316 2660 1324
rect 2668 1316 2676 1324
rect 2684 1316 2692 1324
rect 2636 1116 2644 1124
rect 2652 1116 2660 1124
rect 2396 976 2404 984
rect 2412 956 2420 964
rect 2380 916 2388 924
rect 2380 896 2388 904
rect 2348 856 2356 864
rect 2316 776 2324 784
rect 2332 776 2340 784
rect 2396 796 2404 804
rect 2380 776 2388 784
rect 2364 756 2372 764
rect 2348 716 2356 724
rect 2316 696 2324 704
rect 2332 696 2340 704
rect 2108 676 2116 684
rect 2172 676 2180 684
rect 2268 676 2276 684
rect 1964 636 1972 644
rect 1996 616 2004 624
rect 1900 556 1908 564
rect 1980 556 1988 564
rect 1708 516 1716 524
rect 1884 516 1892 524
rect 1660 496 1668 504
rect 1676 456 1684 464
rect 1804 456 1812 464
rect 1740 436 1748 444
rect 1724 396 1732 404
rect 1772 396 1780 404
rect 1628 296 1636 304
rect 1596 236 1604 244
rect 1852 336 1860 344
rect 1884 376 1892 384
rect 1868 316 1876 324
rect 1964 536 1972 544
rect 1916 516 1924 524
rect 1932 496 1940 504
rect 1916 376 1924 384
rect 1916 316 1924 324
rect 2028 636 2036 644
rect 2172 656 2180 664
rect 2076 616 2084 624
rect 2092 616 2100 624
rect 2108 616 2116 624
rect 2044 576 2052 584
rect 2060 516 2068 524
rect 2028 476 2036 484
rect 2012 316 2020 324
rect 1948 296 1956 304
rect 1980 296 1988 304
rect 1724 276 1732 284
rect 1948 276 1956 284
rect 1660 176 1668 184
rect 1692 176 1700 184
rect 1548 136 1556 144
rect 1900 256 1908 264
rect 1964 256 1972 264
rect 1788 118 1796 124
rect 1788 116 1796 118
rect 1820 116 1828 124
rect 1964 116 1972 124
rect 1260 96 1268 104
rect 2204 596 2212 604
rect 2172 576 2180 584
rect 2124 556 2132 564
rect 2092 536 2100 544
rect 2076 496 2084 504
rect 2044 396 2052 404
rect 2108 516 2116 524
rect 2188 516 2196 524
rect 2124 496 2132 504
rect 2236 576 2244 584
rect 2300 576 2308 584
rect 2220 556 2228 564
rect 2396 716 2404 724
rect 2476 1056 2484 1064
rect 2444 996 2452 1004
rect 2444 936 2452 944
rect 2460 816 2468 824
rect 2547 1006 2555 1014
rect 2557 1006 2565 1014
rect 2567 1006 2575 1014
rect 2577 1006 2585 1014
rect 2587 1006 2595 1014
rect 2597 1006 2605 1014
rect 2620 996 2628 1004
rect 2652 1076 2660 1084
rect 2652 1036 2660 1044
rect 2812 1396 2820 1404
rect 2796 1296 2804 1304
rect 2732 1276 2740 1284
rect 2700 1116 2708 1124
rect 2716 1116 2724 1124
rect 2780 1276 2788 1284
rect 2732 1056 2740 1064
rect 2620 936 2628 944
rect 2524 896 2532 904
rect 2492 856 2500 864
rect 2556 836 2564 844
rect 2444 696 2452 704
rect 2476 696 2484 704
rect 2508 696 2516 704
rect 2380 676 2388 684
rect 2412 676 2420 684
rect 2492 676 2500 684
rect 2364 636 2372 644
rect 2268 556 2276 564
rect 2316 556 2324 564
rect 2188 496 2196 504
rect 2204 496 2212 504
rect 2396 576 2404 584
rect 2476 576 2484 584
rect 2444 536 2452 544
rect 2268 516 2276 524
rect 2316 516 2324 524
rect 2332 516 2340 524
rect 2220 456 2228 464
rect 2252 456 2260 464
rect 2172 436 2180 444
rect 2156 396 2164 404
rect 2140 316 2148 324
rect 2060 256 2068 264
rect 2092 256 2100 264
rect 2076 176 2084 184
rect 2028 136 2036 144
rect 2012 96 2020 104
rect 1964 76 1972 84
rect 1244 36 1252 44
rect 2156 276 2164 284
rect 2156 236 2164 244
rect 2140 136 2148 144
rect 2332 456 2340 464
rect 2332 336 2340 344
rect 2220 316 2228 324
rect 2396 516 2404 524
rect 2380 376 2388 384
rect 2460 476 2468 484
rect 2252 296 2260 304
rect 2364 296 2372 304
rect 2300 276 2308 284
rect 2204 256 2212 264
rect 2188 236 2196 244
rect 2188 196 2196 204
rect 2220 156 2228 164
rect 2284 256 2292 264
rect 2124 116 2132 124
rect 2172 116 2180 124
rect 2268 116 2276 124
rect 2444 276 2452 284
rect 2364 196 2372 204
rect 2396 236 2404 244
rect 2364 176 2372 184
rect 2380 176 2388 184
rect 2348 156 2356 164
rect 2332 136 2340 144
rect 2316 116 2324 124
rect 2220 96 2228 104
rect 2252 96 2260 104
rect 2348 96 2356 104
rect 2572 716 2580 724
rect 2588 696 2596 704
rect 2828 1376 2836 1384
rect 3052 1796 3060 1804
rect 2988 1736 2996 1744
rect 2924 1636 2932 1644
rect 3020 1636 3028 1644
rect 2908 1516 2916 1524
rect 2876 1496 2884 1504
rect 2892 1496 2900 1504
rect 2940 1556 2948 1564
rect 2956 1556 2964 1564
rect 3020 1556 3028 1564
rect 3036 1556 3044 1564
rect 2956 1516 2964 1524
rect 3004 1516 3012 1524
rect 2876 1476 2884 1484
rect 2860 1436 2868 1444
rect 2876 1436 2884 1444
rect 2940 1496 2948 1504
rect 2940 1476 2948 1484
rect 2892 1416 2900 1424
rect 2924 1416 2932 1424
rect 2876 1396 2884 1404
rect 2924 1396 2932 1404
rect 2972 1496 2980 1504
rect 2956 1416 2964 1424
rect 2972 1416 2980 1424
rect 2956 1396 2964 1404
rect 2972 1336 2980 1344
rect 3004 1336 3012 1344
rect 3212 2076 3220 2084
rect 3116 2056 3124 2064
rect 3276 2056 3284 2064
rect 3196 1976 3204 1984
rect 3260 1976 3268 1984
rect 3116 1896 3124 1904
rect 3164 1896 3172 1904
rect 3180 1896 3188 1904
rect 3148 1876 3156 1884
rect 3100 1696 3108 1704
rect 3116 1696 3124 1704
rect 3180 1876 3188 1884
rect 3308 1896 3316 1904
rect 3292 1876 3300 1884
rect 3308 1876 3316 1884
rect 3276 1836 3284 1844
rect 3292 1836 3300 1844
rect 3196 1796 3204 1804
rect 3164 1776 3172 1784
rect 3164 1616 3172 1624
rect 3116 1576 3124 1584
rect 3148 1576 3156 1584
rect 3052 1496 3060 1504
rect 3084 1496 3092 1504
rect 3100 1496 3108 1504
rect 3068 1476 3076 1484
rect 3052 1376 3060 1384
rect 3036 1356 3044 1364
rect 3052 1356 3060 1364
rect 3052 1336 3060 1344
rect 2972 1316 2980 1324
rect 2988 1316 2996 1324
rect 2828 1296 2836 1304
rect 2876 1296 2884 1304
rect 2908 1296 2916 1304
rect 2988 1296 2996 1304
rect 3116 1396 3124 1404
rect 3132 1396 3140 1404
rect 3292 1736 3300 1744
rect 3276 1716 3284 1724
rect 3372 2296 3380 2304
rect 3516 2836 3524 2844
rect 3612 2836 3620 2844
rect 3564 2816 3572 2824
rect 3580 2816 3588 2824
rect 3436 2716 3444 2724
rect 3452 2716 3460 2724
rect 3580 2776 3588 2784
rect 3596 2716 3604 2724
rect 3532 2696 3540 2704
rect 3548 2696 3556 2704
rect 3516 2656 3524 2664
rect 3500 2616 3508 2624
rect 3484 2536 3492 2544
rect 3404 2496 3412 2504
rect 3564 2656 3572 2664
rect 3548 2636 3556 2644
rect 3532 2616 3540 2624
rect 3436 2516 3444 2524
rect 3500 2516 3508 2524
rect 3580 2636 3588 2644
rect 3644 2696 3652 2704
rect 3724 2896 3732 2904
rect 3756 2976 3764 2984
rect 3788 2956 3796 2964
rect 3756 2916 3764 2924
rect 3788 2896 3796 2904
rect 3804 2856 3812 2864
rect 3948 2856 3956 2864
rect 3836 2816 3844 2824
rect 3916 2816 3924 2824
rect 3788 2756 3796 2764
rect 3900 2756 3908 2764
rect 3756 2736 3764 2744
rect 3740 2716 3748 2724
rect 3740 2696 3748 2704
rect 3804 2696 3812 2704
rect 3676 2676 3684 2684
rect 3724 2676 3732 2684
rect 3740 2656 3748 2664
rect 3612 2536 3620 2544
rect 3740 2596 3748 2604
rect 3788 2596 3796 2604
rect 3468 2496 3476 2504
rect 3532 2496 3540 2504
rect 3468 2436 3476 2444
rect 3420 2396 3428 2404
rect 3452 2376 3460 2384
rect 3484 2296 3492 2304
rect 3564 2496 3572 2504
rect 3612 2496 3620 2504
rect 3708 2496 3716 2504
rect 3564 2396 3572 2404
rect 3660 2316 3668 2324
rect 3516 2256 3524 2264
rect 3500 2216 3508 2224
rect 3388 2136 3396 2144
rect 3468 2136 3476 2144
rect 3500 2136 3508 2144
rect 3628 2236 3636 2244
rect 3612 2216 3620 2224
rect 3596 2196 3604 2204
rect 3404 2096 3412 2104
rect 3484 2096 3492 2104
rect 3388 2076 3396 2084
rect 3436 2036 3444 2044
rect 3388 1976 3396 1984
rect 3452 1996 3460 2004
rect 3356 1816 3364 1824
rect 3340 1736 3348 1744
rect 3324 1696 3332 1704
rect 3228 1636 3236 1644
rect 3212 1576 3220 1584
rect 3260 1576 3268 1584
rect 3244 1496 3252 1504
rect 3196 1476 3204 1484
rect 3180 1416 3188 1424
rect 3132 1356 3140 1364
rect 2812 1256 2820 1264
rect 2844 1276 2852 1284
rect 2860 1256 2868 1264
rect 2828 1176 2836 1184
rect 2812 1076 2820 1084
rect 2780 916 2788 924
rect 2796 916 2804 924
rect 2668 796 2676 804
rect 2684 796 2692 804
rect 2636 776 2644 784
rect 2620 756 2628 764
rect 2684 716 2692 724
rect 2620 696 2628 704
rect 2547 606 2555 614
rect 2557 606 2565 614
rect 2567 606 2575 614
rect 2577 606 2585 614
rect 2587 606 2595 614
rect 2597 606 2605 614
rect 2636 676 2644 684
rect 2668 676 2676 684
rect 2732 816 2740 824
rect 2716 696 2724 704
rect 2860 1116 2868 1124
rect 3132 1276 3140 1284
rect 2988 1196 2996 1204
rect 3036 1196 3044 1204
rect 3132 1196 3140 1204
rect 3004 1156 3012 1164
rect 2940 1136 2948 1144
rect 3004 1136 3012 1144
rect 2892 1116 2900 1124
rect 3068 1116 3076 1124
rect 3180 1376 3188 1384
rect 3164 1356 3172 1364
rect 3276 1556 3284 1564
rect 3324 1576 3332 1584
rect 3388 1816 3396 1824
rect 3420 1776 3428 1784
rect 3436 1736 3444 1744
rect 3404 1716 3412 1724
rect 3468 1936 3476 1944
rect 3468 1796 3476 1804
rect 3532 2056 3540 2064
rect 3564 2056 3572 2064
rect 3564 2016 3572 2024
rect 3516 1976 3524 1984
rect 3580 1976 3588 1984
rect 3596 1956 3604 1964
rect 3564 1936 3572 1944
rect 3532 1896 3540 1904
rect 3596 1876 3604 1884
rect 3500 1856 3508 1864
rect 3500 1816 3508 1824
rect 3532 1816 3540 1824
rect 3484 1756 3492 1764
rect 3644 2196 3652 2204
rect 3804 2436 3812 2444
rect 3852 2616 3860 2624
rect 3884 2616 3892 2624
rect 3868 2556 3876 2564
rect 3836 2496 3844 2504
rect 3932 2736 3940 2744
rect 4076 3116 4084 3124
rect 4028 3096 4036 3104
rect 4380 3296 4388 3304
rect 4316 3216 4324 3224
rect 4348 3216 4356 3224
rect 4284 3116 4292 3124
rect 4172 2996 4180 3004
rect 4156 2936 4164 2944
rect 4076 2876 4084 2884
rect 4252 2936 4260 2944
rect 4236 2916 4244 2924
rect 4268 2896 4276 2904
rect 4204 2876 4212 2884
rect 4188 2856 4196 2864
rect 4060 2836 4068 2844
rect 4076 2836 4084 2844
rect 4156 2836 4164 2844
rect 4220 2836 4228 2844
rect 4051 2806 4059 2814
rect 4061 2806 4069 2814
rect 4071 2806 4079 2814
rect 4081 2806 4089 2814
rect 4091 2806 4099 2814
rect 4101 2806 4109 2814
rect 4028 2716 4036 2724
rect 3964 2696 3972 2704
rect 3996 2656 4004 2664
rect 3900 2436 3908 2444
rect 3820 2396 3828 2404
rect 4140 2716 4148 2724
rect 4044 2696 4052 2704
rect 4204 2756 4212 2764
rect 4172 2736 4180 2744
rect 4220 2716 4228 2724
rect 4044 2556 4052 2564
rect 4092 2556 4100 2564
rect 4220 2696 4228 2704
rect 4268 2756 4276 2764
rect 4348 3156 4356 3164
rect 4492 3396 4500 3404
rect 4556 3396 4564 3404
rect 4476 3136 4484 3144
rect 4300 3096 4308 3104
rect 4460 3096 4468 3104
rect 4348 2956 4356 2964
rect 4348 2916 4356 2924
rect 4444 2916 4452 2924
rect 4316 2896 4324 2904
rect 4300 2876 4308 2884
rect 4348 2856 4356 2864
rect 4268 2636 4276 2644
rect 4444 2716 4452 2724
rect 4332 2636 4340 2644
rect 4252 2616 4260 2624
rect 4316 2616 4324 2624
rect 4284 2556 4292 2564
rect 4060 2496 4068 2504
rect 4188 2496 4196 2504
rect 4300 2496 4308 2504
rect 4284 2456 4292 2464
rect 4124 2416 4132 2424
rect 4252 2416 4260 2424
rect 4268 2416 4276 2424
rect 4051 2406 4059 2414
rect 4061 2406 4069 2414
rect 4071 2406 4079 2414
rect 4081 2406 4089 2414
rect 4091 2406 4099 2414
rect 4101 2406 4109 2414
rect 4124 2376 4132 2384
rect 3756 2316 3764 2324
rect 3868 2316 3876 2324
rect 3644 2156 3652 2164
rect 3660 2156 3668 2164
rect 3868 2296 3876 2304
rect 3820 2236 3828 2244
rect 3836 2196 3844 2204
rect 3964 2276 3972 2284
rect 3964 2256 3972 2264
rect 3964 2236 3972 2244
rect 3932 2156 3940 2164
rect 3868 2116 3876 2124
rect 3772 2096 3780 2104
rect 3884 2096 3892 2104
rect 3628 2036 3636 2044
rect 3900 2056 3908 2064
rect 3628 2016 3636 2024
rect 3868 2016 3876 2024
rect 3676 1976 3684 1984
rect 3644 1896 3652 1904
rect 3628 1836 3636 1844
rect 3532 1796 3540 1804
rect 3612 1796 3620 1804
rect 3580 1736 3588 1744
rect 3852 1896 3860 1904
rect 3756 1876 3764 1884
rect 3836 1876 3844 1884
rect 3868 1876 3876 1884
rect 3804 1836 3812 1844
rect 3756 1776 3764 1784
rect 3708 1756 3716 1764
rect 3676 1736 3684 1744
rect 3596 1716 3604 1724
rect 3724 1716 3732 1724
rect 3340 1556 3348 1564
rect 3372 1556 3380 1564
rect 3292 1536 3300 1544
rect 3308 1536 3316 1544
rect 3292 1516 3300 1524
rect 3244 1436 3252 1444
rect 3260 1376 3268 1384
rect 3276 1376 3284 1384
rect 3212 1356 3220 1364
rect 3164 1276 3172 1284
rect 3244 1316 3252 1324
rect 3196 1276 3204 1284
rect 3260 1296 3268 1304
rect 3372 1516 3380 1524
rect 3372 1476 3380 1484
rect 3516 1696 3524 1704
rect 3484 1656 3492 1664
rect 3420 1636 3428 1644
rect 3308 1416 3316 1424
rect 3308 1336 3316 1344
rect 3324 1316 3332 1324
rect 3324 1296 3332 1304
rect 3404 1436 3412 1444
rect 3388 1336 3396 1344
rect 3356 1316 3364 1324
rect 3276 1276 3284 1284
rect 3228 1256 3236 1264
rect 3196 1236 3204 1244
rect 3292 1236 3300 1244
rect 3180 1196 3188 1204
rect 3148 1176 3156 1184
rect 3164 1176 3172 1184
rect 2860 1096 2868 1104
rect 2908 1096 2916 1104
rect 2972 1096 2980 1104
rect 3116 1096 3124 1104
rect 2956 1076 2964 1084
rect 2860 1056 2868 1064
rect 2956 1056 2964 1064
rect 2956 996 2964 1004
rect 2844 936 2852 944
rect 2876 936 2884 944
rect 2908 936 2916 944
rect 2876 916 2884 924
rect 2892 916 2900 924
rect 2796 896 2804 904
rect 2812 896 2820 904
rect 2812 856 2820 864
rect 2892 856 2900 864
rect 2924 856 2932 864
rect 2940 836 2948 844
rect 3068 1056 3076 1064
rect 3084 1056 3092 1064
rect 3052 1036 3060 1044
rect 3020 996 3028 1004
rect 2988 896 2996 904
rect 3196 1116 3204 1124
rect 3244 1116 3252 1124
rect 3340 1276 3348 1284
rect 3452 1436 3460 1444
rect 3436 1356 3444 1364
rect 3404 1276 3412 1284
rect 3228 1096 3236 1104
rect 3260 1096 3268 1104
rect 3276 1096 3284 1104
rect 3132 1056 3140 1064
rect 3100 1036 3108 1044
rect 3116 1036 3124 1044
rect 3100 956 3108 964
rect 3180 1036 3188 1044
rect 3148 936 3156 944
rect 3244 936 3252 944
rect 3084 896 3092 904
rect 3100 896 3108 904
rect 3228 916 3236 924
rect 3260 916 3268 924
rect 3132 856 3140 864
rect 3020 836 3028 844
rect 3036 836 3044 844
rect 2972 816 2980 824
rect 2748 796 2756 804
rect 2764 796 2772 804
rect 2780 796 2788 804
rect 2780 756 2788 764
rect 2796 756 2804 764
rect 2908 756 2916 764
rect 2748 716 2756 724
rect 2764 716 2772 724
rect 2940 716 2948 724
rect 2700 676 2708 684
rect 2716 676 2724 684
rect 2780 676 2788 684
rect 2684 656 2692 664
rect 2748 656 2756 664
rect 2780 656 2788 664
rect 2652 596 2660 604
rect 2620 576 2628 584
rect 2604 556 2612 564
rect 2668 556 2676 564
rect 2524 536 2532 544
rect 2508 516 2516 524
rect 2492 456 2500 464
rect 2572 476 2580 484
rect 2540 416 2548 424
rect 2652 476 2660 484
rect 2636 456 2644 464
rect 2620 416 2628 424
rect 2636 416 2644 424
rect 2604 356 2612 364
rect 2572 336 2580 344
rect 2604 336 2612 344
rect 2684 496 2692 504
rect 2700 496 2708 504
rect 2716 476 2724 484
rect 2732 476 2740 484
rect 2668 356 2676 364
rect 2636 336 2644 344
rect 2652 336 2660 344
rect 2700 336 2708 344
rect 2636 296 2644 304
rect 2764 616 2772 624
rect 2876 676 2884 684
rect 2844 656 2852 664
rect 2812 636 2820 644
rect 2812 596 2820 604
rect 2828 576 2836 584
rect 2780 496 2788 504
rect 2796 496 2804 504
rect 2908 556 2916 564
rect 2812 456 2820 464
rect 2796 336 2804 344
rect 2684 296 2692 304
rect 2748 296 2756 304
rect 2764 296 2772 304
rect 2636 256 2644 264
rect 2620 216 2628 224
rect 2547 206 2555 214
rect 2557 206 2565 214
rect 2567 206 2575 214
rect 2577 206 2585 214
rect 2587 206 2595 214
rect 2597 206 2605 214
rect 2508 196 2516 204
rect 2492 156 2500 164
rect 2780 276 2788 284
rect 2700 196 2708 204
rect 2700 156 2708 164
rect 2444 96 2452 104
rect 2668 96 2676 104
rect 2412 76 2420 84
rect 2636 56 2644 64
rect 2684 56 2692 64
rect 2780 156 2788 164
rect 2956 596 2964 604
rect 2940 536 2948 544
rect 2908 496 2916 504
rect 2908 456 2916 464
rect 2876 336 2884 344
rect 2892 336 2900 344
rect 2812 316 2820 324
rect 2860 296 2868 304
rect 2892 296 2900 304
rect 3036 796 3044 804
rect 3052 716 3060 724
rect 3068 716 3076 724
rect 3148 796 3156 804
rect 3180 756 3188 764
rect 3148 716 3156 724
rect 3164 716 3172 724
rect 3212 716 3220 724
rect 3276 776 3284 784
rect 3228 696 3236 704
rect 3036 676 3044 684
rect 3116 676 3124 684
rect 3164 676 3172 684
rect 3244 676 3252 684
rect 3260 676 3268 684
rect 3116 656 3124 664
rect 3004 616 3012 624
rect 2972 496 2980 504
rect 2924 396 2932 404
rect 2940 396 2948 404
rect 3068 596 3076 604
rect 3084 596 3092 604
rect 3020 576 3028 584
rect 3036 556 3044 564
rect 3052 556 3060 564
rect 3020 536 3028 544
rect 3212 576 3220 584
rect 3500 1556 3508 1564
rect 3692 1696 3700 1704
rect 3548 1676 3556 1684
rect 3612 1676 3620 1684
rect 3628 1676 3636 1684
rect 3532 1656 3540 1664
rect 3516 1496 3524 1504
rect 3516 1476 3524 1484
rect 3484 1416 3492 1424
rect 3500 1356 3508 1364
rect 3532 1436 3540 1444
rect 3596 1656 3604 1664
rect 3564 1496 3572 1504
rect 3580 1496 3588 1504
rect 3644 1556 3652 1564
rect 3660 1556 3668 1564
rect 3692 1516 3700 1524
rect 3564 1416 3572 1424
rect 3548 1356 3556 1364
rect 3756 1696 3764 1704
rect 3740 1656 3748 1664
rect 3804 1656 3812 1664
rect 3772 1576 3780 1584
rect 3756 1516 3764 1524
rect 3660 1496 3668 1504
rect 3772 1496 3780 1504
rect 3740 1456 3748 1464
rect 3692 1416 3700 1424
rect 3724 1416 3732 1424
rect 3644 1396 3652 1404
rect 3596 1356 3604 1364
rect 3612 1356 3620 1364
rect 3628 1336 3636 1344
rect 3644 1316 3652 1324
rect 3564 1276 3572 1284
rect 3548 1256 3556 1264
rect 3484 1236 3492 1244
rect 3564 1236 3572 1244
rect 3468 1216 3476 1224
rect 3468 1116 3476 1124
rect 3548 1116 3556 1124
rect 3548 1096 3556 1104
rect 3404 1076 3412 1084
rect 3468 1076 3476 1084
rect 3372 1056 3380 1064
rect 3452 996 3460 1004
rect 3532 996 3540 1004
rect 3516 956 3524 964
rect 3612 1156 3620 1164
rect 3596 1116 3604 1124
rect 3676 1256 3684 1264
rect 3660 1216 3668 1224
rect 3660 1136 3668 1144
rect 3628 1116 3636 1124
rect 3356 936 3364 944
rect 3436 936 3444 944
rect 3628 936 3636 944
rect 3708 1376 3716 1384
rect 3756 1416 3764 1424
rect 3740 1316 3748 1324
rect 3772 1396 3780 1404
rect 3788 1376 3796 1384
rect 3708 1156 3716 1164
rect 3724 1056 3732 1064
rect 3772 1296 3780 1304
rect 3756 1136 3764 1144
rect 3756 1076 3764 1084
rect 3740 996 3748 1004
rect 3388 916 3396 924
rect 3564 916 3572 924
rect 3644 916 3652 924
rect 3292 756 3300 764
rect 3340 736 3348 744
rect 3356 716 3364 724
rect 3324 696 3332 704
rect 3308 676 3316 684
rect 3324 676 3332 684
rect 3324 596 3332 604
rect 3180 556 3188 564
rect 3100 516 3108 524
rect 3180 496 3188 504
rect 3020 476 3028 484
rect 3116 476 3124 484
rect 3004 356 3012 364
rect 3004 316 3012 324
rect 2988 296 2996 304
rect 2860 156 2868 164
rect 2892 136 2900 144
rect 2940 136 2948 144
rect 3132 456 3140 464
rect 3084 396 3092 404
rect 3068 316 3076 324
rect 3116 356 3124 364
rect 3036 276 3044 284
rect 3084 236 3092 244
rect 3260 556 3268 564
rect 3276 556 3284 564
rect 3164 316 3172 324
rect 3180 316 3188 324
rect 3228 336 3236 344
rect 3500 856 3508 864
rect 3484 736 3492 744
rect 3436 676 3444 684
rect 3372 616 3380 624
rect 3388 616 3396 624
rect 3356 576 3364 584
rect 3340 536 3348 544
rect 3292 496 3300 504
rect 3148 256 3156 264
rect 3020 156 3028 164
rect 2988 136 2996 144
rect 2796 96 2804 104
rect 2860 116 2868 124
rect 2924 116 2932 124
rect 2972 116 2980 124
rect 3004 116 3012 124
rect 3196 276 3204 284
rect 3420 536 3428 544
rect 3452 496 3460 504
rect 3500 576 3508 584
rect 3740 916 3748 924
rect 3692 856 3700 864
rect 3580 836 3588 844
rect 3612 816 3620 824
rect 3596 716 3604 724
rect 3548 696 3556 704
rect 3596 656 3604 664
rect 3516 556 3524 564
rect 3516 516 3524 524
rect 3468 456 3476 464
rect 3388 436 3396 444
rect 3372 416 3380 424
rect 3436 356 3444 364
rect 3596 536 3604 544
rect 3628 716 3636 724
rect 3628 676 3636 684
rect 3644 656 3652 664
rect 3708 616 3716 624
rect 3996 2316 4004 2324
rect 4028 2316 4036 2324
rect 4044 2316 4052 2324
rect 4028 2296 4036 2304
rect 4252 2296 4260 2304
rect 4332 2436 4340 2444
rect 4140 2256 4148 2264
rect 3996 2176 4004 2184
rect 4172 2176 4180 2184
rect 4396 2636 4404 2644
rect 4412 2496 4420 2504
rect 4508 3336 4516 3344
rect 4620 3336 4628 3344
rect 4620 3316 4628 3324
rect 4732 3316 4740 3324
rect 4588 3296 4596 3304
rect 4572 3096 4580 3104
rect 4524 3076 4532 3084
rect 4716 3296 4724 3304
rect 4684 3276 4692 3284
rect 4668 3256 4676 3264
rect 4668 3216 4676 3224
rect 4652 3096 4660 3104
rect 4652 3076 4660 3084
rect 4572 3056 4580 3064
rect 4620 3056 4628 3064
rect 4556 2936 4564 2944
rect 4588 3036 4596 3044
rect 4588 2996 4596 3004
rect 4556 2916 4564 2924
rect 4572 2916 4580 2924
rect 4620 2976 4628 2984
rect 4620 2876 4628 2884
rect 4540 2736 4548 2744
rect 4572 2736 4580 2744
rect 4588 2736 4596 2744
rect 4620 2736 4628 2744
rect 4492 2716 4500 2724
rect 4556 2716 4564 2724
rect 4572 2716 4580 2724
rect 4508 2696 4516 2704
rect 4540 2636 4548 2644
rect 4524 2596 4532 2604
rect 4652 2596 4660 2604
rect 4508 2576 4516 2584
rect 4476 2556 4484 2564
rect 4508 2516 4516 2524
rect 4444 2476 4452 2484
rect 4428 2436 4436 2444
rect 4364 2336 4372 2344
rect 4412 2336 4420 2344
rect 4364 2276 4372 2284
rect 4636 2556 4644 2564
rect 4540 2516 4548 2524
rect 4908 3316 4916 3324
rect 4796 3236 4804 3244
rect 4748 3216 4756 3224
rect 4988 3256 4996 3264
rect 4700 3116 4708 3124
rect 4780 3116 4788 3124
rect 4716 3102 4724 3104
rect 4716 3096 4724 3102
rect 4780 3096 4788 3104
rect 4828 3096 4836 3104
rect 4956 3096 4964 3104
rect 4716 2976 4724 2984
rect 4700 2936 4708 2944
rect 4860 3036 4868 3044
rect 4844 2976 4852 2984
rect 4828 2936 4836 2944
rect 4700 2876 4708 2884
rect 4700 2856 4708 2864
rect 4716 2776 4724 2784
rect 4780 2776 4788 2784
rect 4716 2736 4724 2744
rect 4764 2596 4772 2604
rect 4700 2576 4708 2584
rect 4764 2556 4772 2564
rect 4492 2316 4500 2324
rect 4524 2316 4532 2324
rect 4412 2296 4420 2304
rect 4508 2296 4516 2304
rect 4396 2236 4404 2244
rect 4380 2176 4388 2184
rect 4364 2156 4372 2164
rect 4412 2156 4420 2164
rect 4124 2136 4132 2144
rect 4156 2136 4164 2144
rect 3964 2096 3972 2104
rect 3948 2036 3956 2044
rect 3916 2016 3924 2024
rect 4028 2056 4036 2064
rect 4140 2096 4148 2104
rect 4284 2096 4292 2104
rect 4380 2096 4388 2104
rect 4188 2076 4196 2084
rect 4300 2076 4308 2084
rect 4156 2056 4164 2064
rect 4028 2016 4036 2024
rect 4051 2006 4059 2014
rect 4061 2006 4069 2014
rect 4071 2006 4079 2014
rect 4081 2006 4089 2014
rect 4091 2006 4099 2014
rect 4101 2006 4109 2014
rect 4172 2016 4180 2024
rect 3996 1976 4004 1984
rect 4140 1976 4148 1984
rect 3948 1956 3956 1964
rect 4316 1976 4324 1984
rect 4396 1976 4404 1984
rect 4236 1956 4244 1964
rect 4380 1956 4388 1964
rect 4268 1936 4276 1944
rect 4108 1896 4116 1904
rect 4140 1896 4148 1904
rect 3996 1816 4004 1824
rect 3900 1776 3908 1784
rect 4172 1816 4180 1824
rect 3884 1716 3892 1724
rect 3836 1616 3844 1624
rect 3836 1576 3844 1584
rect 3900 1696 3908 1704
rect 3916 1696 3924 1704
rect 4076 1718 4084 1724
rect 4076 1716 4084 1718
rect 3964 1676 3972 1684
rect 4012 1676 4020 1684
rect 3932 1536 3940 1544
rect 3980 1496 3988 1504
rect 4140 1716 4148 1724
rect 4284 1856 4292 1864
rect 4300 1776 4308 1784
rect 4300 1736 4308 1744
rect 4204 1696 4212 1704
rect 4051 1606 4059 1614
rect 4061 1606 4069 1614
rect 4071 1606 4079 1614
rect 4081 1606 4089 1614
rect 4091 1606 4099 1614
rect 4101 1606 4109 1614
rect 4092 1556 4100 1564
rect 4204 1496 4212 1504
rect 3836 1476 3844 1484
rect 3804 1196 3812 1204
rect 3788 1176 3796 1184
rect 3852 1436 3860 1444
rect 3916 1356 3924 1364
rect 4012 1336 4020 1344
rect 4268 1696 4276 1704
rect 4300 1696 4308 1704
rect 4252 1676 4260 1684
rect 4380 1856 4388 1864
rect 4364 1836 4372 1844
rect 4332 1776 4340 1784
rect 4508 2256 4516 2264
rect 4428 2136 4436 2144
rect 4428 2096 4436 2104
rect 4668 2516 4676 2524
rect 4748 2516 4756 2524
rect 4572 2496 4580 2504
rect 4636 2496 4644 2504
rect 4748 2496 4756 2504
rect 4588 2356 4596 2364
rect 4476 2136 4484 2144
rect 4508 2136 4516 2144
rect 4460 2056 4468 2064
rect 4460 2016 4468 2024
rect 4412 1916 4420 1924
rect 4428 1916 4436 1924
rect 4508 1916 4516 1924
rect 4892 2976 4900 2984
rect 4876 2956 4884 2964
rect 4908 2956 4916 2964
rect 4876 2936 4884 2944
rect 4844 2756 4852 2764
rect 4876 2756 4884 2764
rect 4924 2936 4932 2944
rect 4924 2916 4932 2924
rect 4924 2896 4932 2904
rect 4940 2856 4948 2864
rect 4924 2776 4932 2784
rect 4844 2656 4852 2664
rect 4796 2596 4804 2604
rect 4860 2596 4868 2604
rect 4796 2556 4804 2564
rect 4844 2416 4852 2424
rect 4812 2336 4820 2344
rect 4828 2316 4836 2324
rect 4860 2316 4868 2324
rect 4828 2296 4836 2304
rect 4860 2296 4868 2304
rect 4764 2276 4772 2284
rect 4716 2256 4724 2264
rect 4588 2156 4596 2164
rect 4844 2156 4852 2164
rect 4908 2736 4916 2744
rect 4908 2576 4916 2584
rect 4908 2436 4916 2444
rect 4892 2356 4900 2364
rect 4748 2136 4756 2144
rect 4908 2236 4916 2244
rect 5036 3336 5044 3344
rect 5004 2956 5012 2964
rect 4972 2896 4980 2904
rect 4972 2856 4980 2864
rect 4956 2696 4964 2704
rect 4972 2696 4980 2704
rect 5004 2696 5012 2704
rect 4940 2376 4948 2384
rect 4972 2656 4980 2664
rect 5036 3136 5044 3144
rect 5084 3276 5092 3284
rect 5052 3076 5060 3084
rect 5068 3076 5076 3084
rect 5052 2896 5060 2904
rect 5036 2736 5044 2744
rect 5036 2676 5044 2684
rect 5020 2596 5028 2604
rect 5052 2576 5060 2584
rect 5020 2536 5028 2544
rect 5084 2856 5092 2864
rect 5068 2496 5076 2504
rect 5036 2476 5044 2484
rect 5020 2456 5028 2464
rect 5052 2456 5060 2464
rect 5036 2416 5044 2424
rect 5132 3096 5140 3104
rect 5116 3076 5124 3084
rect 5100 2716 5108 2724
rect 5100 2516 5108 2524
rect 5036 2376 5044 2384
rect 5084 2376 5092 2384
rect 4956 2356 4964 2364
rect 4940 2336 4948 2344
rect 5004 2302 5012 2304
rect 5004 2296 5012 2302
rect 4972 2276 4980 2284
rect 4940 2236 4948 2244
rect 4924 2196 4932 2204
rect 4812 2116 4820 2124
rect 4892 2116 4900 2124
rect 4924 2116 4932 2124
rect 4716 2096 4724 2104
rect 4796 2096 4804 2104
rect 4652 2076 4660 2084
rect 4780 2076 4788 2084
rect 4572 2056 4580 2064
rect 4540 1896 4548 1904
rect 4428 1856 4436 1864
rect 4428 1816 4436 1824
rect 4444 1796 4452 1804
rect 4460 1796 4468 1804
rect 4348 1756 4356 1764
rect 4364 1756 4372 1764
rect 4396 1756 4404 1764
rect 4492 1856 4500 1864
rect 4524 1836 4532 1844
rect 4540 1836 4548 1844
rect 4524 1816 4532 1824
rect 4492 1776 4500 1784
rect 4524 1776 4532 1784
rect 4508 1756 4516 1764
rect 4396 1736 4404 1744
rect 4476 1736 4484 1744
rect 4716 2056 4724 2064
rect 4748 1996 4756 2004
rect 4588 1956 4596 1964
rect 4572 1936 4580 1944
rect 4636 1936 4644 1944
rect 4700 1936 4708 1944
rect 4748 1936 4756 1944
rect 4588 1916 4596 1924
rect 4652 1916 4660 1924
rect 4716 1916 4724 1924
rect 4668 1876 4676 1884
rect 4924 2056 4932 2064
rect 4828 1956 4836 1964
rect 4844 1936 4852 1944
rect 4876 1936 4884 1944
rect 4828 1896 4836 1904
rect 4588 1836 4596 1844
rect 4732 1836 4740 1844
rect 4796 1836 4804 1844
rect 4812 1836 4820 1844
rect 4588 1816 4596 1824
rect 4732 1796 4740 1804
rect 4652 1756 4660 1764
rect 4812 1736 4820 1744
rect 4556 1716 4564 1724
rect 4700 1716 4708 1724
rect 4860 1716 4868 1724
rect 4380 1696 4388 1704
rect 4476 1696 4484 1704
rect 4604 1696 4612 1704
rect 4684 1696 4692 1704
rect 4780 1696 4788 1704
rect 4924 1896 4932 1904
rect 4892 1696 4900 1704
rect 4572 1676 4580 1684
rect 4732 1676 4740 1684
rect 4764 1676 4772 1684
rect 4876 1676 4884 1684
rect 4316 1516 4324 1524
rect 4508 1516 4516 1524
rect 4556 1516 4564 1524
rect 4252 1476 4260 1484
rect 4220 1396 4228 1404
rect 4284 1436 4292 1444
rect 4124 1356 4132 1364
rect 4044 1336 4052 1344
rect 4252 1318 4260 1324
rect 4252 1316 4260 1318
rect 3916 1296 3924 1304
rect 3820 1076 3828 1084
rect 3804 1056 3812 1064
rect 3868 1176 3876 1184
rect 3900 1116 3908 1124
rect 3980 1236 3988 1244
rect 3980 1176 3988 1184
rect 3980 1116 3988 1124
rect 4012 1116 4020 1124
rect 4012 1096 4020 1104
rect 4412 1502 4420 1504
rect 4412 1496 4420 1502
rect 4508 1496 4516 1504
rect 4444 1476 4452 1484
rect 4476 1436 4484 1444
rect 4508 1436 4516 1444
rect 4588 1436 4596 1444
rect 4332 1396 4340 1404
rect 4444 1396 4452 1404
rect 4316 1296 4324 1304
rect 4051 1206 4059 1214
rect 4061 1206 4069 1214
rect 4071 1206 4079 1214
rect 4081 1206 4089 1214
rect 4091 1206 4099 1214
rect 4101 1206 4109 1214
rect 4044 1176 4052 1184
rect 4124 1156 4132 1164
rect 4348 1356 4356 1364
rect 4428 1336 4436 1344
rect 4348 1316 4356 1324
rect 4396 1296 4404 1304
rect 4492 1316 4500 1324
rect 4444 1296 4452 1304
rect 4492 1296 4500 1304
rect 4428 1176 4436 1184
rect 4220 1116 4228 1124
rect 3900 1076 3908 1084
rect 3980 1076 3988 1084
rect 3868 1056 3876 1064
rect 3948 996 3956 1004
rect 3836 916 3844 924
rect 3772 816 3780 824
rect 4044 936 4052 944
rect 3964 916 3972 924
rect 3852 856 3860 864
rect 3804 796 3812 804
rect 3884 796 3892 804
rect 3948 736 3956 744
rect 3772 716 3780 724
rect 3852 716 3860 724
rect 3932 696 3940 704
rect 3836 676 3844 684
rect 3884 676 3892 684
rect 3756 536 3764 544
rect 3900 596 3908 604
rect 3948 596 3956 604
rect 3900 536 3908 544
rect 3612 516 3620 524
rect 3692 516 3700 524
rect 3644 496 3652 504
rect 3580 476 3588 484
rect 3612 476 3620 484
rect 3532 356 3540 364
rect 3564 356 3572 364
rect 3628 356 3636 364
rect 3340 316 3348 324
rect 3564 316 3572 324
rect 3644 316 3652 324
rect 3244 256 3252 264
rect 3308 276 3316 284
rect 3212 216 3220 224
rect 3228 216 3236 224
rect 3276 216 3284 224
rect 3292 216 3300 224
rect 3324 256 3332 264
rect 3356 256 3364 264
rect 3660 296 3668 304
rect 3692 276 3700 284
rect 3532 256 3540 264
rect 3420 236 3428 244
rect 3356 216 3364 224
rect 3468 216 3476 224
rect 3484 216 3492 224
rect 3244 136 3252 144
rect 3292 136 3300 144
rect 3324 136 3332 144
rect 3372 136 3380 144
rect 3436 136 3444 144
rect 3484 196 3492 204
rect 3788 518 3796 524
rect 3788 516 3796 518
rect 3852 516 3860 524
rect 3884 516 3892 524
rect 3852 476 3860 484
rect 3820 456 3828 464
rect 3852 456 3860 464
rect 3820 376 3828 384
rect 3788 296 3796 304
rect 3756 276 3764 284
rect 3740 256 3748 264
rect 3660 236 3668 244
rect 3676 236 3684 244
rect 3596 196 3604 204
rect 3660 156 3668 164
rect 3692 156 3700 164
rect 4140 996 4148 1004
rect 4348 1036 4356 1044
rect 4300 996 4308 1004
rect 4300 936 4308 944
rect 4268 918 4276 924
rect 4268 916 4276 918
rect 4396 956 4404 964
rect 4348 916 4356 924
rect 4076 856 4084 864
rect 4300 856 4308 864
rect 4051 806 4059 814
rect 4061 806 4069 814
rect 4071 806 4079 814
rect 4081 806 4089 814
rect 4091 806 4099 814
rect 4101 806 4109 814
rect 4140 736 4148 744
rect 4076 716 4084 724
rect 4252 716 4260 724
rect 4236 696 4244 704
rect 4284 696 4292 704
rect 4380 916 4388 924
rect 4396 836 4404 844
rect 4364 776 4372 784
rect 4300 616 4308 624
rect 4108 596 4116 604
rect 4252 596 4260 604
rect 4332 596 4340 604
rect 4092 556 4100 564
rect 4220 556 4228 564
rect 4380 576 4388 584
rect 4332 556 4340 564
rect 4364 556 4372 564
rect 4380 536 4388 544
rect 4092 516 4100 524
rect 3932 496 3940 504
rect 4012 496 4020 504
rect 3916 376 3924 384
rect 3948 316 3956 324
rect 4051 406 4059 414
rect 4061 406 4069 414
rect 4071 406 4079 414
rect 4081 406 4089 414
rect 4091 406 4099 414
rect 4101 406 4109 414
rect 4012 396 4020 404
rect 4012 376 4020 384
rect 4188 376 4196 384
rect 3884 296 3892 304
rect 3948 302 3956 304
rect 3948 296 3956 302
rect 3980 296 3988 304
rect 4156 356 4164 364
rect 4044 316 4052 324
rect 4156 316 4164 324
rect 4476 1102 4484 1104
rect 4476 1096 4484 1102
rect 4572 1296 4580 1304
rect 4524 1256 4532 1264
rect 4572 1116 4580 1124
rect 4572 1096 4580 1104
rect 4716 1502 4724 1504
rect 4716 1496 4724 1502
rect 4780 1496 4788 1504
rect 4812 1496 4820 1504
rect 4700 1476 4708 1484
rect 4732 1376 4740 1384
rect 4636 1316 4644 1324
rect 4700 1316 4708 1324
rect 4668 1216 4676 1224
rect 4652 1176 4660 1184
rect 4620 1136 4628 1144
rect 4620 1116 4628 1124
rect 4604 1056 4612 1064
rect 4540 1036 4548 1044
rect 4604 1036 4612 1044
rect 4508 976 4516 984
rect 4588 956 4596 964
rect 4476 936 4484 944
rect 4524 936 4532 944
rect 4700 1196 4708 1204
rect 4716 1156 4724 1164
rect 4860 1576 4868 1584
rect 5004 2136 5012 2144
rect 4956 1836 4964 1844
rect 4924 1496 4932 1504
rect 4860 1436 4868 1444
rect 4876 1396 4884 1404
rect 4924 1376 4932 1384
rect 4860 1336 4868 1344
rect 5052 2116 5060 2124
rect 5132 2556 5140 2564
rect 5132 2336 5140 2344
rect 5052 1936 5060 1944
rect 5100 1956 5108 1964
rect 5068 1876 5076 1884
rect 5084 1856 5092 1864
rect 4988 1736 4996 1744
rect 4972 1496 4980 1504
rect 4892 1316 4900 1324
rect 4844 1136 4852 1144
rect 4716 1116 4724 1124
rect 4908 1116 4916 1124
rect 4844 1102 4852 1104
rect 4844 1096 4852 1102
rect 4956 1096 4964 1104
rect 4684 1036 4692 1044
rect 4636 996 4644 1004
rect 4812 956 4820 964
rect 4652 936 4660 944
rect 4684 936 4692 944
rect 4620 916 4628 924
rect 4636 916 4644 924
rect 5148 2176 5156 2184
rect 5148 2116 5156 2124
rect 5132 1896 5140 1904
rect 5148 1856 5156 1864
rect 5132 1836 5140 1844
rect 5116 1796 5124 1804
rect 5132 1796 5140 1804
rect 5116 1756 5124 1764
rect 5116 1736 5124 1744
rect 5052 1716 5060 1724
rect 5068 1716 5076 1724
rect 5132 1716 5140 1724
rect 5148 1716 5156 1724
rect 5036 1496 5044 1504
rect 5020 1356 5028 1364
rect 4988 1336 4996 1344
rect 5020 1336 5028 1344
rect 5100 1496 5108 1504
rect 5116 1396 5124 1404
rect 5052 1316 5060 1324
rect 5100 1316 5108 1324
rect 4988 1176 4996 1184
rect 5004 1156 5012 1164
rect 5020 1136 5028 1144
rect 5036 1136 5044 1144
rect 5004 1116 5012 1124
rect 4988 1096 4996 1104
rect 5020 1096 5028 1104
rect 4876 956 4884 964
rect 4780 916 4788 924
rect 4940 936 4948 944
rect 4924 916 4932 924
rect 4684 896 4692 904
rect 4604 876 4612 884
rect 4668 876 4676 884
rect 4620 856 4628 864
rect 4748 856 4756 864
rect 4556 796 4564 804
rect 4620 796 4628 804
rect 4444 776 4452 784
rect 4556 736 4564 744
rect 4540 716 4548 724
rect 4748 736 4756 744
rect 4684 716 4692 724
rect 4444 676 4452 684
rect 4508 676 4516 684
rect 4460 636 4468 644
rect 4284 516 4292 524
rect 4316 516 4324 524
rect 4364 516 4372 524
rect 4428 516 4436 524
rect 4140 296 4148 304
rect 4268 296 4276 304
rect 3980 276 3988 284
rect 4252 276 4260 284
rect 3852 196 3860 204
rect 4172 236 4180 244
rect 4236 196 4244 204
rect 4012 156 4020 164
rect 4188 156 4196 164
rect 3804 136 3812 144
rect 4380 256 4388 264
rect 4860 796 4868 804
rect 4828 736 4836 744
rect 4796 716 4804 724
rect 4764 696 4772 704
rect 4716 656 4724 664
rect 4636 616 4644 624
rect 4732 556 4740 564
rect 4652 536 4660 544
rect 4716 536 4724 544
rect 4828 576 4836 584
rect 4844 536 4852 544
rect 4460 516 4468 524
rect 4700 516 4708 524
rect 4780 516 4788 524
rect 4444 236 4452 244
rect 4380 216 4388 224
rect 4236 136 4244 144
rect 4252 136 4260 144
rect 3196 116 3204 124
rect 3228 116 3236 124
rect 3276 116 3284 124
rect 3308 116 3316 124
rect 3580 116 3588 124
rect 3228 96 3236 104
rect 2780 76 2788 84
rect 2828 76 2836 84
rect 2860 76 2868 84
rect 3004 76 3012 84
rect 3132 76 3140 84
rect 3164 76 3172 84
rect 4172 116 4180 124
rect 4220 116 4228 124
rect 3612 96 3620 104
rect 3884 96 3892 104
rect 4140 96 4148 104
rect 4492 316 4500 324
rect 4876 716 4884 724
rect 5068 1276 5076 1284
rect 5068 1216 5076 1224
rect 5100 1276 5108 1284
rect 5084 1196 5092 1204
rect 5084 1176 5092 1184
rect 5100 1136 5108 1144
rect 5148 1196 5156 1204
rect 5148 1116 5156 1124
rect 5068 1096 5076 1104
rect 5084 1096 5092 1104
rect 5020 936 5028 944
rect 5052 936 5060 944
rect 4972 896 4980 904
rect 4892 696 4900 704
rect 4956 676 4964 684
rect 4908 596 4916 604
rect 4908 536 4916 544
rect 4892 516 4900 524
rect 4684 476 4692 484
rect 4796 476 4804 484
rect 4860 476 4868 484
rect 4572 356 4580 364
rect 4540 276 4548 284
rect 4556 196 4564 204
rect 4540 136 4548 144
rect 4620 256 4628 264
rect 4460 116 4468 124
rect 4508 116 4516 124
rect 4380 96 4388 104
rect 4476 96 4484 104
rect 4764 376 4772 384
rect 4668 316 4676 324
rect 4860 376 4868 384
rect 4812 336 4820 344
rect 4668 296 4676 304
rect 4764 296 4772 304
rect 4684 276 4692 284
rect 4636 196 4644 204
rect 4988 876 4996 884
rect 5004 796 5012 804
rect 4988 756 4996 764
rect 5052 796 5060 804
rect 5036 736 5044 744
rect 5132 776 5140 784
rect 5068 716 5076 724
rect 4972 656 4980 664
rect 4956 376 4964 384
rect 4908 336 4916 344
rect 4892 296 4900 304
rect 5004 296 5012 304
rect 4796 196 4804 204
rect 4924 196 4932 204
rect 4716 176 4724 184
rect 4812 176 4820 184
rect 4604 136 4612 144
rect 4700 136 4708 144
rect 4780 136 4788 144
rect 4876 136 4884 144
rect 5132 136 5140 144
rect 3564 76 3572 84
rect 4252 76 4260 84
rect 3388 56 3396 64
rect 3628 56 3636 64
rect 3388 36 3396 44
rect 4620 36 4628 44
rect 2764 16 2772 24
rect 3324 16 3332 24
rect 4051 6 4059 14
rect 4061 6 4069 14
rect 4071 6 4079 14
rect 4081 6 4089 14
rect 4091 6 4099 14
rect 4101 6 4109 14
<< metal3 >>
rect 2692 3417 3852 3423
rect 3860 3417 4476 3423
rect 2546 3414 2606 3416
rect 2546 3406 2547 3414
rect 2556 3406 2557 3414
rect 2595 3406 2596 3414
rect 2605 3406 2606 3414
rect 2546 3404 2606 3406
rect 932 3397 2284 3403
rect 2292 3397 2524 3403
rect 2621 3397 3980 3403
rect 1316 3377 1500 3383
rect 1508 3377 1516 3383
rect 2621 3383 2627 3397
rect 4500 3397 4556 3403
rect 1956 3377 2627 3383
rect 2644 3377 2924 3383
rect 2932 3377 4300 3383
rect 4308 3377 4396 3383
rect 148 3357 364 3363
rect 1597 3357 1644 3363
rect 1597 3344 1603 3357
rect 1652 3357 1932 3363
rect 2436 3357 2620 3363
rect 2644 3357 2796 3363
rect 2852 3357 2940 3363
rect 2948 3357 3356 3363
rect 3364 3357 3468 3363
rect 3684 3357 4115 3363
rect 4109 3344 4115 3357
rect 356 3337 476 3343
rect 676 3337 732 3343
rect 1076 3337 1228 3343
rect 1300 3337 1596 3343
rect 1844 3337 2172 3343
rect 2196 3337 2220 3343
rect 2564 3337 2748 3343
rect 2788 3337 2892 3343
rect 2900 3337 2988 3343
rect 3044 3337 3132 3343
rect 3332 3337 3628 3343
rect 3636 3337 3788 3343
rect 4116 3337 4236 3343
rect 4388 3337 4508 3343
rect 4628 3337 5036 3343
rect 20 3317 236 3323
rect 244 3317 300 3323
rect 356 3317 492 3323
rect 532 3317 732 3323
rect 1236 3317 1276 3323
rect 1284 3317 1292 3323
rect 1444 3317 1532 3323
rect 1748 3317 1868 3323
rect 1908 3317 2252 3323
rect 2356 3317 2412 3323
rect 2420 3317 2492 3323
rect 2509 3317 2636 3323
rect 340 3297 364 3303
rect 468 3297 524 3303
rect 1012 3297 1372 3303
rect 1380 3297 1564 3303
rect 1844 3297 1868 3303
rect 2084 3297 2348 3303
rect 2509 3303 2515 3317
rect 2804 3317 2860 3323
rect 2964 3317 3052 3323
rect 3396 3317 3436 3323
rect 3460 3317 3660 3323
rect 3924 3317 3932 3323
rect 3988 3317 4172 3323
rect 4196 3317 4252 3323
rect 4260 3317 4620 3323
rect 4740 3317 4908 3323
rect 2436 3297 2515 3303
rect 2532 3297 2684 3303
rect 2861 3303 2867 3316
rect 2861 3297 2972 3303
rect 2996 3297 3699 3303
rect 3693 3284 3699 3297
rect 3828 3297 3932 3303
rect 3972 3297 4156 3303
rect 4308 3297 4380 3303
rect 4596 3297 4716 3303
rect 404 3277 652 3283
rect 708 3277 732 3283
rect 1204 3277 1292 3283
rect 1620 3277 1804 3283
rect 2036 3277 2124 3283
rect 2148 3277 2204 3283
rect 2212 3277 2332 3283
rect 2484 3277 2588 3283
rect 2628 3277 2748 3283
rect 2996 3277 3084 3283
rect 3092 3277 3164 3283
rect 3172 3277 3340 3283
rect 3444 3277 3580 3283
rect 3700 3277 3884 3283
rect 3988 3277 4012 3283
rect 4020 3277 4140 3283
rect 4148 3277 4172 3283
rect 4180 3277 4268 3283
rect 4692 3277 5084 3283
rect 372 3257 604 3263
rect 612 3257 860 3263
rect 868 3257 1004 3263
rect 1188 3257 3388 3263
rect 3972 3257 3996 3263
rect 4004 3257 4124 3263
rect 4132 3257 4668 3263
rect 4676 3257 4988 3263
rect 420 3237 588 3243
rect 724 3237 780 3243
rect 948 3237 1164 3243
rect 1860 3237 2156 3243
rect 2164 3237 2188 3243
rect 2292 3237 2435 3243
rect 1540 3217 1580 3223
rect 1588 3217 1948 3223
rect 2020 3217 2108 3223
rect 2116 3217 2284 3223
rect 2381 3217 2412 3223
rect 1042 3214 1102 3216
rect 1042 3206 1043 3214
rect 1052 3206 1053 3214
rect 1091 3206 1092 3214
rect 1101 3206 1102 3214
rect 1042 3204 1102 3206
rect 1812 3197 2156 3203
rect 2381 3203 2387 3217
rect 2429 3223 2435 3237
rect 2452 3237 2892 3243
rect 3028 3237 3100 3243
rect 3108 3237 4796 3243
rect 2429 3217 3996 3223
rect 4324 3217 4348 3223
rect 4356 3217 4668 3223
rect 4676 3217 4748 3223
rect 4050 3214 4110 3216
rect 4050 3206 4051 3214
rect 4060 3206 4061 3214
rect 4099 3206 4100 3214
rect 4109 3206 4110 3214
rect 4050 3204 4110 3206
rect 2164 3197 2387 3203
rect 2532 3197 2684 3203
rect 2772 3197 3996 3203
rect 724 3177 812 3183
rect 836 3177 1228 3183
rect 1924 3177 2044 3183
rect 2052 3177 2204 3183
rect 2276 3177 2924 3183
rect 2932 3177 3324 3183
rect 388 3157 540 3163
rect 676 3157 835 3163
rect -35 3137 60 3143
rect 100 3137 252 3143
rect 260 3137 444 3143
rect 564 3137 812 3143
rect 829 3143 835 3157
rect 1316 3157 4348 3163
rect 829 3137 1724 3143
rect 1828 3137 2236 3143
rect 2340 3137 2668 3143
rect 2692 3137 2796 3143
rect 2836 3137 3036 3143
rect 3044 3137 3228 3143
rect 3300 3137 3404 3143
rect 3444 3137 3724 3143
rect 3732 3137 3740 3143
rect 3748 3137 3996 3143
rect 4004 3137 4156 3143
rect 4484 3137 5036 3143
rect 484 3117 508 3123
rect 644 3117 780 3123
rect 916 3117 1148 3123
rect 1172 3117 1388 3123
rect 1492 3117 1980 3123
rect 2004 3117 2076 3123
rect 2148 3117 2348 3123
rect 2372 3117 2604 3123
rect 2644 3117 2924 3123
rect 2964 3117 3004 3123
rect 3140 3117 4076 3123
rect 4084 3117 4284 3123
rect 4708 3117 4780 3123
rect -35 3097 12 3103
rect 356 3097 476 3103
rect 548 3097 652 3103
rect 740 3097 812 3103
rect 1140 3097 1180 3103
rect 1188 3097 1196 3103
rect 1268 3097 1468 3103
rect 1620 3097 1708 3103
rect 1716 3097 1756 3103
rect 1956 3097 1996 3103
rect 2052 3097 2060 3103
rect 2244 3097 2732 3103
rect 2772 3097 2908 3103
rect 3172 3097 3251 3103
rect 244 3077 508 3083
rect 516 3077 924 3083
rect 941 3077 1164 3083
rect 941 3063 947 3077
rect 1220 3077 1292 3083
rect 1492 3077 1596 3083
rect 2036 3077 2044 3083
rect 2100 3077 2252 3083
rect 2292 3077 2444 3083
rect 2484 3077 2732 3083
rect 2788 3077 2828 3083
rect 2932 3077 2988 3083
rect 3005 3077 3132 3083
rect 756 3057 947 3063
rect 1012 3057 1324 3063
rect 1428 3057 1692 3063
rect 1700 3057 1884 3063
rect 1908 3057 2220 3063
rect 2237 3057 2636 3063
rect 708 3037 796 3043
rect 1044 3037 1372 3043
rect 2237 3043 2243 3057
rect 3005 3063 3011 3077
rect 3245 3083 3251 3097
rect 3268 3097 3308 3103
rect 3316 3097 3372 3103
rect 3380 3097 3420 3103
rect 3684 3097 3724 3103
rect 3892 3097 4028 3103
rect 4308 3097 4460 3103
rect 4580 3097 4652 3103
rect 4724 3097 4780 3103
rect 4836 3097 4956 3103
rect 4964 3097 5132 3103
rect 3245 3077 3276 3083
rect 3332 3077 3452 3083
rect 3588 3077 3676 3083
rect 3828 3077 3948 3083
rect 3956 3077 4460 3083
rect 4532 3077 4652 3083
rect 5060 3077 5068 3083
rect 5076 3077 5116 3083
rect 2653 3057 3011 3063
rect 1396 3037 2243 3043
rect 2260 3037 2492 3043
rect 2653 3043 2659 3057
rect 3076 3057 3148 3063
rect 4580 3057 4620 3063
rect 2644 3037 2659 3043
rect 2692 3037 3276 3043
rect 3332 3037 3420 3043
rect 3428 3037 3452 3043
rect 3460 3037 3644 3043
rect 4596 3037 4860 3043
rect 612 3017 2428 3023
rect 2452 3017 2524 3023
rect 2724 3017 2892 3023
rect 2900 3017 3340 3023
rect 3380 3017 3468 3023
rect 4589 3023 4595 3036
rect 3476 3017 4595 3023
rect 2546 3014 2606 3016
rect 2546 3006 2547 3014
rect 2556 3006 2557 3014
rect 2595 3006 2596 3014
rect 2605 3006 2606 3014
rect 2546 3004 2606 3006
rect 20 2997 44 3003
rect 852 2997 1171 3003
rect 276 2977 396 2983
rect 1165 2983 1171 2997
rect 1188 2997 1500 3003
rect 1508 2997 1708 3003
rect 1732 2997 2476 3003
rect 2708 2997 3020 3003
rect 3028 2997 3500 3003
rect 3508 2997 3692 3003
rect 4180 2997 4588 3003
rect 1165 2977 1196 2983
rect 1236 2977 1388 2983
rect 1412 2977 1468 2983
rect 1524 2977 1580 2983
rect 1636 2977 1692 2983
rect 1716 2977 1980 2983
rect 1997 2977 2060 2983
rect 596 2957 620 2963
rect 628 2957 700 2963
rect 724 2957 899 2963
rect 628 2937 684 2943
rect 692 2937 732 2943
rect 756 2937 860 2943
rect 868 2937 876 2943
rect 893 2943 899 2957
rect 948 2957 1059 2963
rect 893 2937 956 2943
rect 980 2937 1036 2943
rect 1053 2943 1059 2957
rect 1252 2957 1356 2963
rect 1364 2957 1532 2963
rect 1540 2957 1772 2963
rect 1997 2963 2003 2977
rect 2084 2977 2131 2983
rect 1956 2957 2003 2963
rect 2020 2957 2108 2963
rect 2125 2963 2131 2977
rect 2180 2977 2252 2983
rect 2292 2977 2508 2983
rect 2516 2977 3756 2983
rect 3764 2977 4172 2983
rect 4308 2977 4620 2983
rect 4628 2977 4716 2983
rect 4852 2977 4892 2983
rect 2125 2957 2636 2963
rect 2676 2957 2700 2963
rect 2724 2957 2828 2963
rect 2916 2957 3084 2963
rect 3220 2957 3292 2963
rect 3636 2957 3660 2963
rect 3668 2957 3788 2963
rect 4141 2957 4348 2963
rect 1053 2937 1260 2943
rect 1348 2937 1628 2943
rect 1700 2937 1756 2943
rect 1764 2937 1868 2943
rect 1988 2937 2028 2943
rect 2052 2937 2092 2943
rect 2116 2937 2156 2943
rect 2228 2937 2236 2943
rect 2260 2937 2332 2943
rect 2388 2937 2444 2943
rect 2468 2937 2604 2943
rect 2612 2937 2652 2943
rect 2660 2937 2972 2943
rect 2980 2937 3244 2943
rect 4141 2943 4147 2957
rect 4916 2957 5004 2963
rect 3300 2937 4147 2943
rect 4164 2937 4252 2943
rect 4260 2937 4556 2943
rect 4708 2937 4828 2943
rect 4884 2937 4924 2943
rect 132 2917 268 2923
rect 276 2917 460 2923
rect 788 2917 828 2923
rect 836 2917 844 2923
rect 916 2917 988 2923
rect 1028 2917 1164 2923
rect 1172 2917 1228 2923
rect 1268 2917 1324 2923
rect 1332 2917 1436 2923
rect 1524 2917 1548 2923
rect 1652 2917 2220 2923
rect 2260 2917 2268 2923
rect 2324 2917 2444 2923
rect 2452 2917 2796 2923
rect 2804 2917 3036 2923
rect 3044 2917 3228 2923
rect 3236 2917 3404 2923
rect 3620 2917 3756 2923
rect 4244 2917 4339 2923
rect 868 2897 972 2903
rect 980 2897 1004 2903
rect 1508 2897 1612 2903
rect 1636 2897 1644 2903
rect 1668 2897 1708 2903
rect 2253 2903 2259 2916
rect 1812 2897 2259 2903
rect 2356 2897 2444 2903
rect 2676 2897 2812 2903
rect 2980 2897 3052 2903
rect 3076 2897 3180 2903
rect 3236 2897 3356 2903
rect 3732 2897 3788 2903
rect 4276 2897 4316 2903
rect 4333 2903 4339 2917
rect 4356 2917 4444 2923
rect 4468 2917 4556 2923
rect 4580 2917 4924 2923
rect 4973 2917 5187 2923
rect 4973 2904 4979 2917
rect 4333 2897 4924 2903
rect 4932 2897 4972 2903
rect 5060 2897 5100 2903
rect 5181 2897 5187 2917
rect 644 2877 764 2883
rect 980 2877 1292 2883
rect 1300 2877 2028 2883
rect 2036 2877 2076 2883
rect 2100 2877 2764 2883
rect 2804 2877 2876 2883
rect 2893 2883 2899 2896
rect 2893 2877 4076 2883
rect 4212 2877 4300 2883
rect 4628 2877 4700 2883
rect 884 2857 1132 2863
rect 1156 2857 1660 2863
rect 1716 2857 1740 2863
rect 1748 2857 2140 2863
rect 2180 2857 2188 2863
rect 2212 2857 2508 2863
rect 2580 2857 2636 2863
rect 2644 2857 2684 2863
rect 2788 2857 2844 2863
rect 2852 2857 2860 2863
rect 2868 2857 2940 2863
rect 2948 2857 2988 2863
rect 2996 2857 3068 2863
rect 3092 2857 3276 2863
rect 3348 2857 3388 2863
rect 3428 2857 3804 2863
rect 3956 2857 4188 2863
rect 4196 2857 4348 2863
rect 4708 2857 4940 2863
rect 4948 2857 4972 2863
rect 5076 2857 5084 2863
rect 740 2837 1123 2843
rect 340 2817 652 2823
rect 900 2817 1020 2823
rect 1117 2823 1123 2837
rect 1396 2837 2060 2843
rect 2084 2837 2732 2843
rect 2772 2837 2956 2843
rect 2980 2837 3004 2843
rect 3028 2837 3100 2843
rect 3140 2837 3276 2843
rect 3348 2837 3516 2843
rect 3620 2837 4060 2843
rect 4084 2837 4156 2843
rect 4164 2837 4220 2843
rect 1117 2817 1980 2823
rect 2004 2817 2060 2823
rect 2148 2817 3564 2823
rect 3588 2817 3836 2823
rect 3844 2817 3916 2823
rect 1042 2814 1102 2816
rect 1042 2806 1043 2814
rect 1052 2806 1053 2814
rect 1091 2806 1092 2814
rect 1101 2806 1102 2814
rect 1042 2804 1102 2806
rect 4050 2814 4110 2816
rect 4050 2806 4051 2814
rect 4060 2806 4061 2814
rect 4099 2806 4100 2814
rect 4109 2806 4110 2814
rect 4050 2804 4110 2806
rect 932 2797 1004 2803
rect 1124 2797 1292 2803
rect 1332 2797 1500 2803
rect 1716 2797 1900 2803
rect 1940 2797 1996 2803
rect 2004 2797 2252 2803
rect 2324 2797 2460 2803
rect 2500 2797 3603 2803
rect 212 2777 556 2783
rect 868 2777 1148 2783
rect 1268 2777 1276 2783
rect 1284 2777 1452 2783
rect 1460 2777 1580 2783
rect 1588 2777 1843 2783
rect 1837 2764 1843 2777
rect 1876 2777 2108 2783
rect 2132 2777 2268 2783
rect 2404 2777 2492 2783
rect 2516 2777 3084 2783
rect 3124 2777 3164 2783
rect 3172 2777 3580 2783
rect 3597 2783 3603 2797
rect 3597 2777 4716 2783
rect 4788 2777 4924 2783
rect 484 2757 700 2763
rect 740 2757 819 2763
rect 148 2737 588 2743
rect 676 2737 796 2743
rect 813 2743 819 2757
rect 852 2757 1484 2763
rect 1508 2757 1820 2763
rect 1844 2757 2092 2763
rect 2100 2757 2220 2763
rect 2228 2757 2428 2763
rect 2445 2757 2652 2763
rect 813 2737 876 2743
rect 916 2737 1148 2743
rect 1156 2737 1212 2743
rect 1220 2737 1452 2743
rect 1460 2737 1852 2743
rect 1876 2737 1964 2743
rect 1988 2737 2204 2743
rect 2445 2743 2451 2757
rect 2669 2757 2796 2763
rect 2292 2737 2451 2743
rect 2669 2743 2675 2757
rect 2852 2757 3779 2763
rect 2516 2737 2675 2743
rect 2772 2737 2908 2743
rect 2996 2737 3020 2743
rect 3060 2737 3084 2743
rect 3108 2737 3196 2743
rect 3316 2737 3404 2743
rect 3412 2737 3756 2743
rect 3773 2743 3779 2757
rect 3796 2757 3900 2763
rect 3908 2757 4204 2763
rect 4212 2757 4268 2763
rect 4852 2757 4876 2763
rect 3773 2737 3932 2743
rect 3940 2737 4172 2743
rect 4548 2737 4572 2743
rect 4596 2737 4620 2743
rect 4724 2737 4908 2743
rect 4980 2737 5036 2743
rect 52 2717 172 2723
rect 548 2717 636 2723
rect 772 2717 828 2723
rect 836 2717 892 2723
rect 916 2717 1420 2723
rect 1444 2717 1468 2723
rect 1492 2717 1804 2723
rect 1876 2717 1932 2723
rect 1956 2717 2156 2723
rect 2244 2717 2332 2723
rect 2356 2717 2380 2723
rect 2516 2717 2844 2723
rect 2868 2717 2908 2723
rect 2964 2717 3132 2723
rect 3188 2717 3260 2723
rect 3284 2717 3436 2723
rect 3460 2717 3596 2723
rect 3748 2717 4028 2723
rect 4036 2717 4140 2723
rect 4180 2717 4220 2723
rect 4452 2717 4492 2723
rect 4500 2717 4556 2723
rect 4580 2717 4748 2723
rect 4756 2717 5100 2723
rect -35 2697 12 2703
rect 180 2697 380 2703
rect 532 2697 716 2703
rect 756 2697 780 2703
rect 820 2697 1004 2703
rect 1044 2697 1468 2703
rect 1620 2697 1868 2703
rect 1908 2697 1964 2703
rect 1988 2697 2060 2703
rect 2068 2697 2124 2703
rect 2164 2697 2252 2703
rect 2292 2697 2444 2703
rect 2452 2697 2700 2703
rect 2708 2697 2860 2703
rect 2868 2697 3148 2703
rect 3156 2697 3196 2703
rect 3204 2697 3388 2703
rect 3556 2697 3644 2703
rect 3732 2697 3740 2703
rect 3812 2697 3964 2703
rect 4052 2697 4220 2703
rect 4516 2697 4956 2703
rect 4980 2697 5004 2703
rect 52 2677 204 2683
rect 324 2677 380 2683
rect 436 2677 515 2683
rect 116 2657 492 2663
rect 509 2663 515 2677
rect 612 2677 796 2683
rect 820 2677 876 2683
rect 884 2677 924 2683
rect 1012 2677 1116 2683
rect 1220 2677 1228 2683
rect 1236 2677 1244 2683
rect 1300 2677 1500 2683
rect 1540 2677 1740 2683
rect 1748 2677 2476 2683
rect 2484 2677 2524 2683
rect 2916 2677 3004 2683
rect 3012 2677 3212 2683
rect 3220 2677 3676 2683
rect 3684 2677 3724 2683
rect 4788 2677 5036 2683
rect 509 2657 1036 2663
rect 1204 2657 1292 2663
rect 1316 2657 1340 2663
rect 1364 2657 1404 2663
rect 1412 2657 1420 2663
rect 1828 2657 1836 2663
rect 1860 2657 1884 2663
rect 1924 2657 1980 2663
rect 2116 2657 2140 2663
rect 2164 2657 2348 2663
rect 2372 2657 2444 2663
rect 2452 2657 3036 2663
rect 3076 2657 3244 2663
rect 3524 2657 3564 2663
rect 3572 2657 3731 2663
rect 68 2637 572 2643
rect 692 2637 1372 2643
rect 1421 2643 1427 2656
rect 1421 2637 2044 2643
rect 2052 2637 2060 2643
rect 2100 2637 2364 2643
rect 2516 2637 2620 2643
rect 2628 2637 2972 2643
rect 2980 2637 2988 2643
rect 2996 2637 3132 2643
rect 3156 2637 3308 2643
rect 3316 2637 3548 2643
rect 3572 2637 3580 2643
rect 3725 2643 3731 2657
rect 3748 2657 3996 2663
rect 4852 2657 4972 2663
rect 3725 2637 4268 2643
rect 4276 2637 4332 2643
rect 4404 2637 4540 2643
rect 420 2617 572 2623
rect 612 2617 1260 2623
rect 1332 2617 1356 2623
rect 1364 2617 1484 2623
rect 1492 2617 1756 2623
rect 1764 2617 1772 2623
rect 1780 2617 1948 2623
rect 2100 2617 2188 2623
rect 2260 2617 2412 2623
rect 2644 2617 2668 2623
rect 2676 2617 3500 2623
rect 3540 2617 3852 2623
rect 3860 2617 3884 2623
rect 3892 2617 4252 2623
rect 4260 2617 4316 2623
rect 4324 2617 4492 2623
rect 2546 2614 2606 2616
rect 2546 2606 2547 2614
rect 2556 2606 2557 2614
rect 2595 2606 2596 2614
rect 2605 2606 2606 2614
rect 2546 2604 2606 2606
rect 452 2597 476 2603
rect 596 2597 620 2603
rect 628 2597 636 2603
rect 653 2597 1292 2603
rect 653 2583 659 2597
rect 1332 2597 1404 2603
rect 1412 2597 2019 2603
rect 628 2577 659 2583
rect 1005 2577 1244 2583
rect 1005 2564 1011 2577
rect 1268 2577 1644 2583
rect 1732 2577 1772 2583
rect 1780 2577 1932 2583
rect 1940 2577 1996 2583
rect 2013 2583 2019 2597
rect 2052 2597 2355 2603
rect 2349 2584 2355 2597
rect 2404 2597 2508 2603
rect 2676 2597 2764 2603
rect 3044 2597 3740 2603
rect 3796 2597 3820 2603
rect 4532 2597 4652 2603
rect 4772 2597 4796 2603
rect 4804 2597 4860 2603
rect 5028 2597 5036 2603
rect 2013 2577 2076 2583
rect 2116 2577 2156 2583
rect 2212 2577 2316 2583
rect 2356 2577 4300 2583
rect 4516 2577 4700 2583
rect 4916 2577 5052 2583
rect 340 2557 387 2563
rect -35 2537 60 2543
rect 276 2537 316 2543
rect 324 2537 364 2543
rect 381 2543 387 2557
rect 724 2557 732 2563
rect 756 2557 764 2563
rect 884 2557 1004 2563
rect 1588 2557 1612 2563
rect 1716 2557 1836 2563
rect 1844 2557 1964 2563
rect 2173 2563 2179 2576
rect 1988 2557 2179 2563
rect 2196 2557 2371 2563
rect 381 2537 508 2543
rect 564 2537 636 2543
rect 772 2537 908 2543
rect 1140 2537 1164 2543
rect 1236 2537 1388 2543
rect 1421 2537 1676 2543
rect 1421 2524 1427 2537
rect 1828 2537 1900 2543
rect 1908 2537 2140 2543
rect 2148 2537 2332 2543
rect 2340 2537 2348 2543
rect 2365 2543 2371 2557
rect 2388 2557 2588 2563
rect 2612 2557 2700 2563
rect 2724 2557 3651 2563
rect 2365 2537 3132 2543
rect 3140 2537 3324 2543
rect 3492 2537 3612 2543
rect 3620 2537 3628 2543
rect 3645 2543 3651 2557
rect 3876 2557 4044 2563
rect 4100 2557 4204 2563
rect 4292 2557 4476 2563
rect 4644 2557 4764 2563
rect 4804 2557 5132 2563
rect 4797 2543 4803 2556
rect 3645 2537 4803 2543
rect 4820 2537 5020 2543
rect 5028 2537 5068 2543
rect 244 2517 300 2523
rect 356 2517 620 2523
rect 916 2517 956 2523
rect 964 2517 972 2523
rect 1140 2517 1292 2523
rect 1300 2517 1420 2523
rect 1556 2517 1660 2523
rect 1796 2517 1804 2523
rect 1876 2517 1955 2523
rect -35 2497 12 2503
rect 516 2497 556 2503
rect 676 2497 1116 2503
rect 1204 2497 1340 2503
rect 1357 2497 1404 2503
rect 548 2477 1164 2483
rect 1357 2483 1363 2497
rect 1492 2497 1500 2503
rect 1620 2497 1628 2503
rect 1652 2497 1891 2503
rect 1220 2477 1363 2483
rect 1380 2477 1500 2483
rect 1508 2477 1644 2483
rect 1652 2477 1868 2483
rect 1885 2483 1891 2497
rect 1908 2497 1932 2503
rect 1949 2503 1955 2517
rect 1972 2517 1980 2523
rect 2132 2517 2252 2523
rect 2308 2517 2556 2523
rect 2580 2517 2668 2523
rect 2692 2517 2716 2523
rect 2740 2517 2796 2523
rect 2804 2517 2924 2523
rect 2964 2517 3004 2523
rect 3044 2517 3052 2523
rect 3268 2517 3372 2523
rect 3508 2517 4508 2523
rect 4548 2517 4668 2523
rect 4676 2517 4748 2523
rect 4756 2517 5100 2523
rect 1949 2497 1964 2503
rect 2068 2497 2188 2503
rect 2196 2497 2204 2503
rect 2276 2497 2451 2503
rect 2445 2484 2451 2497
rect 2500 2497 2668 2503
rect 2708 2497 3052 2503
rect 3364 2497 3404 2503
rect 3476 2497 3532 2503
rect 3572 2497 3612 2503
rect 3716 2497 3836 2503
rect 4068 2497 4188 2503
rect 4212 2497 4300 2503
rect 4308 2497 4412 2503
rect 4420 2497 4572 2503
rect 4644 2497 4748 2503
rect 1885 2477 2252 2483
rect 2276 2477 2380 2483
rect 2404 2477 2428 2483
rect 2468 2477 2572 2483
rect 2596 2477 2652 2483
rect 2660 2477 2844 2483
rect 2868 2477 2940 2483
rect 3012 2477 4444 2483
rect 4916 2477 4972 2483
rect 5181 2483 5187 2503
rect 5044 2477 5187 2483
rect 132 2457 300 2463
rect 1140 2457 1692 2463
rect 1700 2457 1724 2463
rect 1732 2457 1900 2463
rect 1972 2457 1996 2463
rect 2036 2457 4284 2463
rect 5028 2457 5052 2463
rect 116 2437 156 2443
rect 868 2437 1532 2443
rect 1652 2437 1772 2443
rect 1780 2437 1820 2443
rect 1876 2437 2012 2443
rect 2196 2437 2220 2443
rect 2244 2437 2316 2443
rect 2452 2437 2492 2443
rect 2532 2437 2636 2443
rect 2660 2437 2716 2443
rect 2772 2437 3100 2443
rect 3124 2437 3356 2443
rect 3476 2437 3804 2443
rect 3908 2437 4332 2443
rect 4436 2437 4812 2443
rect 4884 2437 4908 2443
rect 1316 2417 1372 2423
rect 1588 2417 2028 2423
rect 2068 2417 2316 2423
rect 2420 2417 2684 2423
rect 2692 2417 2764 2423
rect 2852 2417 3020 2423
rect 3060 2417 3820 2423
rect 4132 2417 4252 2423
rect 4276 2417 4844 2423
rect 4852 2417 5036 2423
rect 1042 2414 1102 2416
rect 1042 2406 1043 2414
rect 1052 2406 1053 2414
rect 1091 2406 1092 2414
rect 1101 2406 1102 2414
rect 1042 2404 1102 2406
rect 4050 2414 4110 2416
rect 4050 2406 4051 2414
rect 4060 2406 4061 2414
rect 4099 2406 4100 2414
rect 4109 2406 4110 2414
rect 4050 2404 4110 2406
rect 1124 2397 2092 2403
rect 2228 2397 2892 2403
rect 2900 2397 3420 2403
rect 3428 2397 3468 2403
rect 3572 2397 3820 2403
rect 996 2377 1612 2383
rect 1620 2377 3036 2383
rect 3044 2377 3452 2383
rect 3460 2377 4124 2383
rect 4148 2377 4940 2383
rect 5044 2377 5084 2383
rect 116 2357 476 2363
rect 484 2357 620 2363
rect 1364 2357 1932 2363
rect 1956 2357 2156 2363
rect 2180 2357 2348 2363
rect 2388 2357 2492 2363
rect 2500 2357 2508 2363
rect 2525 2357 4588 2363
rect -35 2337 12 2343
rect 196 2337 492 2343
rect 612 2337 1395 2343
rect 52 2317 220 2323
rect 372 2317 460 2323
rect 916 2317 1228 2323
rect 1252 2317 1372 2323
rect 1389 2323 1395 2337
rect 2525 2343 2531 2357
rect 4900 2357 4956 2363
rect 1524 2337 2531 2343
rect 2548 2337 2764 2343
rect 2836 2337 3052 2343
rect 3092 2337 3180 2343
rect 3188 2337 4140 2343
rect 4372 2337 4412 2343
rect 4420 2337 4812 2343
rect 4948 2337 5132 2343
rect 1389 2317 1948 2323
rect 2125 2317 2508 2323
rect 2125 2304 2131 2317
rect 2548 2317 2659 2323
rect -35 2297 60 2303
rect 132 2297 140 2303
rect 148 2297 188 2303
rect 324 2297 684 2303
rect 756 2297 828 2303
rect 964 2297 1116 2303
rect 1268 2297 1340 2303
rect 1364 2297 1420 2303
rect 1428 2297 1484 2303
rect 1604 2297 1676 2303
rect 1796 2297 1964 2303
rect 2036 2297 2108 2303
rect 2164 2297 2188 2303
rect 2212 2297 2236 2303
rect 2244 2297 2284 2303
rect 2372 2297 2636 2303
rect 2653 2303 2659 2317
rect 2676 2317 2684 2323
rect 2701 2317 2748 2323
rect 2701 2303 2707 2317
rect 2820 2317 2828 2323
rect 2852 2317 2924 2323
rect 2996 2317 3660 2323
rect 3764 2317 3868 2323
rect 4004 2317 4028 2323
rect 4036 2317 4044 2323
rect 4500 2317 4524 2323
rect 4836 2317 4860 2323
rect 2653 2297 2707 2303
rect 2724 2297 2796 2303
rect 2813 2297 3244 2303
rect 116 2277 172 2283
rect 180 2277 428 2283
rect 484 2277 812 2283
rect 932 2277 940 2283
rect 1156 2277 1660 2283
rect 1716 2277 1756 2283
rect 1780 2277 1868 2283
rect 1908 2277 2012 2283
rect 2068 2277 2140 2283
rect 2189 2283 2195 2296
rect 2813 2284 2819 2297
rect 3380 2297 3484 2303
rect 3876 2297 3916 2303
rect 4036 2297 4252 2303
rect 4420 2297 4508 2303
rect 4756 2297 4828 2303
rect 4868 2297 5004 2303
rect 2189 2277 2268 2283
rect 2285 2277 2300 2283
rect 692 2257 748 2263
rect 756 2257 876 2263
rect 932 2257 1244 2263
rect 1428 2257 1516 2263
rect 1668 2257 1788 2263
rect 1908 2257 1964 2263
rect 1988 2257 2028 2263
rect 2285 2263 2291 2277
rect 2317 2277 2492 2283
rect 2036 2257 2291 2263
rect 2317 2263 2323 2277
rect 2612 2277 2668 2283
rect 2756 2277 2764 2283
rect 2836 2277 3020 2283
rect 3044 2277 3132 2283
rect 3140 2277 3964 2283
rect 4749 2283 4755 2296
rect 4372 2277 4755 2283
rect 4772 2277 4972 2283
rect 2308 2257 2323 2263
rect 2452 2257 2476 2263
rect 2500 2257 2540 2263
rect 2660 2257 2748 2263
rect 2788 2257 2940 2263
rect 2948 2257 3260 2263
rect 3268 2257 3516 2263
rect 3972 2257 4140 2263
rect 4516 2257 4716 2263
rect 628 2237 1676 2243
rect 1780 2237 2252 2243
rect 2324 2237 2460 2243
rect 2516 2237 2700 2243
rect 2884 2237 3148 2243
rect 3172 2237 3228 2243
rect 3236 2237 3628 2243
rect 3636 2237 3820 2243
rect 3972 2237 4396 2243
rect 4916 2237 4940 2243
rect 852 2217 972 2223
rect 980 2217 1548 2223
rect 1556 2217 2156 2223
rect 2164 2217 2204 2223
rect 2212 2217 2396 2223
rect 2436 2217 2524 2223
rect 2628 2217 2828 2223
rect 2884 2217 2892 2223
rect 2916 2217 3500 2223
rect 4909 2223 4915 2236
rect 3620 2217 4915 2223
rect 2546 2214 2606 2216
rect 2546 2206 2547 2214
rect 2556 2206 2557 2214
rect 2595 2206 2596 2214
rect 2605 2206 2606 2214
rect 2546 2204 2606 2206
rect 1204 2197 1468 2203
rect 1796 2197 1852 2203
rect 1892 2197 2092 2203
rect 2132 2197 2172 2203
rect 2196 2197 2220 2203
rect 2237 2197 2316 2203
rect 916 2177 972 2183
rect 980 2177 1596 2183
rect 1604 2177 1628 2183
rect 1652 2177 2076 2183
rect 2237 2183 2243 2197
rect 2340 2197 2412 2203
rect 2452 2197 2476 2203
rect 2484 2197 2492 2203
rect 2644 2197 2892 2203
rect 2964 2197 3052 2203
rect 3092 2197 3340 2203
rect 3348 2197 3596 2203
rect 3652 2197 3836 2203
rect 3853 2197 4924 2203
rect 2100 2177 2243 2183
rect 3853 2183 3859 2197
rect 2260 2177 3859 2183
rect 4004 2177 4172 2183
rect 4388 2177 5148 2183
rect 404 2157 476 2163
rect 532 2157 620 2163
rect 676 2157 812 2163
rect 1060 2157 1196 2163
rect 1556 2157 1836 2163
rect 1860 2157 1900 2163
rect 1940 2157 2028 2163
rect 2068 2157 2076 2163
rect 2301 2157 2380 2163
rect 420 2137 572 2143
rect 820 2137 1004 2143
rect 1124 2137 1308 2143
rect 1316 2137 1564 2143
rect 1572 2137 1692 2143
rect 1748 2137 1996 2143
rect 2068 2137 2220 2143
rect 2301 2143 2307 2157
rect 2500 2157 2652 2163
rect 2660 2157 2780 2163
rect 2788 2157 2892 2163
rect 2957 2157 3084 2163
rect 2260 2137 2307 2143
rect 2356 2137 2508 2143
rect 2532 2137 2659 2143
rect 52 2117 156 2123
rect 308 2117 364 2123
rect 420 2117 716 2123
rect 932 2117 940 2123
rect 1220 2117 1260 2123
rect 1268 2117 1356 2123
rect 1556 2117 1580 2123
rect 1668 2117 1804 2123
rect 1812 2117 1868 2123
rect 1924 2117 2092 2123
rect 2196 2117 2284 2123
rect 2324 2117 2636 2123
rect 2653 2123 2659 2137
rect 2676 2137 2716 2143
rect 2724 2137 2812 2143
rect 2957 2143 2963 2157
rect 3108 2157 3196 2163
rect 3204 2157 3644 2163
rect 3668 2157 3932 2163
rect 3940 2157 4364 2163
rect 4420 2157 4588 2163
rect 4596 2157 4844 2163
rect 2836 2137 2963 2143
rect 3060 2137 3388 2143
rect 3508 2137 4124 2143
rect 4148 2137 4156 2143
rect 4436 2137 4476 2143
rect 4500 2137 4508 2143
rect 4756 2137 5004 2143
rect 2653 2117 2700 2123
rect 2740 2117 3868 2123
rect 3876 2117 4812 2123
rect 4820 2117 4892 2123
rect 4932 2117 5052 2123
rect 5156 2117 5187 2123
rect -35 2097 12 2103
rect 68 2097 108 2103
rect 148 2097 364 2103
rect 1012 2097 1052 2103
rect 1156 2097 1228 2103
rect 1380 2097 1484 2103
rect 1556 2097 1628 2103
rect 1828 2097 1996 2103
rect 2004 2097 2380 2103
rect 2452 2097 2844 2103
rect 2868 2097 3004 2103
rect 3028 2097 3100 2103
rect 3108 2097 3116 2103
rect 3124 2097 3180 2103
rect 3412 2097 3484 2103
rect 3780 2097 3884 2103
rect 3956 2097 3964 2103
rect 4148 2097 4284 2103
rect 4388 2097 4428 2103
rect 4724 2097 4796 2103
rect 516 2077 1180 2083
rect 1476 2077 1580 2083
rect 1588 2077 1836 2083
rect 1860 2077 1884 2083
rect 1908 2077 2220 2083
rect 2340 2077 2412 2083
rect 2436 2077 2476 2083
rect 2500 2077 2691 2083
rect 628 2057 1644 2063
rect 1748 2057 2204 2063
rect 2292 2057 2300 2063
rect 2324 2057 2668 2063
rect 2685 2063 2691 2077
rect 2708 2077 3212 2083
rect 3396 2077 4188 2083
rect 4196 2077 4300 2083
rect 4660 2077 4780 2083
rect 2685 2057 3116 2063
rect 3284 2057 3532 2063
rect 3860 2057 3900 2063
rect 4036 2057 4156 2063
rect 4468 2057 4572 2063
rect 4724 2057 4924 2063
rect 148 2037 172 2043
rect 948 2037 1068 2043
rect 1076 2037 1532 2043
rect 1540 2037 1756 2043
rect 1764 2037 1932 2043
rect 1940 2037 2988 2043
rect 3028 2037 3436 2043
rect 3444 2037 3628 2043
rect 3636 2037 3948 2043
rect 1492 2017 1564 2023
rect 1636 2017 1884 2023
rect 1940 2017 2748 2023
rect 2781 2017 2828 2023
rect 1042 2014 1102 2016
rect 1042 2006 1043 2014
rect 1052 2006 1053 2014
rect 1091 2006 1092 2014
rect 1101 2006 1102 2014
rect 1042 2004 1102 2006
rect 2781 2004 2787 2017
rect 2884 2017 3084 2023
rect 3572 2017 3628 2023
rect 3636 2017 3868 2023
rect 3876 2017 3916 2023
rect 3924 2017 4028 2023
rect 4180 2017 4460 2023
rect 4050 2014 4110 2016
rect 4050 2006 4051 2014
rect 4060 2006 4061 2014
rect 4099 2006 4100 2014
rect 4109 2006 4110 2014
rect 4050 2004 4110 2006
rect 596 1997 812 2003
rect 1117 1997 1916 2003
rect 1117 1983 1123 1997
rect 1956 1997 1964 2003
rect 2004 1997 2044 2003
rect 2052 1997 2060 2003
rect 2180 1997 2220 2003
rect 2308 1997 2444 2003
rect 2484 1997 2556 2003
rect 2644 1997 2716 2003
rect 2740 1997 2780 2003
rect 2820 1997 2828 2003
rect 2836 1997 2988 2003
rect 3460 1997 4019 2003
rect 548 1977 1123 1983
rect 1140 1977 2124 1983
rect 2148 1977 2172 1983
rect 2180 1977 2211 1983
rect 468 1957 524 1963
rect 532 1957 556 1963
rect 564 1957 588 1963
rect 692 1957 1500 1963
rect 1716 1957 1804 1963
rect 1876 1957 1900 1963
rect 1924 1957 1980 1963
rect 2036 1957 2060 1963
rect 2116 1957 2188 1963
rect 2205 1963 2211 1977
rect 2260 1977 2412 1983
rect 2436 1977 2508 1983
rect 2516 1977 2684 1983
rect 2708 1977 2876 1983
rect 2900 1977 3036 1983
rect 3092 1977 3196 1983
rect 3268 1977 3388 1983
rect 3524 1977 3580 1983
rect 3684 1977 3996 1983
rect 4013 1983 4019 1997
rect 4125 1997 4748 2003
rect 4125 1983 4131 1997
rect 4013 1977 4131 1983
rect 4148 1977 4316 1983
rect 4324 1977 4396 1983
rect 2205 1957 2252 1963
rect 2260 1957 2316 1963
rect 2388 1957 2524 1963
rect 2532 1957 2764 1963
rect 2852 1957 3596 1963
rect 3956 1957 4236 1963
rect 4244 1957 4380 1963
rect 4596 1957 4828 1963
rect 292 1937 1564 1943
rect 1572 1937 1772 1943
rect 1780 1937 3068 1943
rect 3076 1937 3308 1943
rect 3316 1937 3436 1943
rect 3476 1937 3564 1943
rect 3597 1943 3603 1956
rect 3597 1937 3852 1943
rect 3860 1937 4268 1943
rect 4580 1937 4636 1943
rect 4644 1937 4700 1943
rect 4756 1937 4844 1943
rect 4884 1937 5052 1943
rect 5060 1937 5068 1943
rect 52 1917 204 1923
rect 372 1917 412 1923
rect 884 1917 1004 1923
rect 1012 1917 1052 1923
rect 1060 1917 1292 1923
rect 1316 1917 1340 1923
rect 1460 1917 1468 1923
rect 1476 1917 1548 1923
rect 1652 1917 1724 1923
rect 1732 1917 1772 1923
rect 1844 1917 1852 1923
rect 1860 1917 1964 1923
rect 1972 1917 2044 1923
rect 2084 1917 2172 1923
rect 2212 1917 2284 1923
rect 2324 1917 2396 1923
rect 2420 1917 2492 1923
rect 2644 1917 2700 1923
rect 2756 1917 4412 1923
rect 4436 1917 4508 1923
rect 4516 1917 4588 1923
rect 4596 1917 4652 1923
rect 4660 1917 4716 1923
rect -35 1897 12 1903
rect 100 1897 124 1903
rect 132 1897 172 1903
rect 356 1897 476 1903
rect 516 1897 636 1903
rect 788 1897 972 1903
rect 1236 1897 1388 1903
rect 1620 1897 1772 1903
rect 1892 1897 1964 1903
rect 1972 1897 2092 1903
rect 2164 1897 2348 1903
rect 2420 1897 2444 1903
rect 2500 1897 2652 1903
rect 2756 1897 2924 1903
rect 2980 1897 3107 1903
rect 212 1877 460 1883
rect 580 1877 636 1883
rect 644 1877 684 1883
rect 1012 1877 1036 1883
rect 1060 1877 1132 1883
rect 1204 1877 1244 1883
rect 1284 1877 1420 1883
rect 1453 1877 1836 1883
rect 1453 1864 1459 1877
rect 2004 1877 2076 1883
rect 2148 1877 2460 1883
rect 2500 1877 2844 1883
rect 2964 1877 2988 1883
rect 3101 1883 3107 1897
rect 3124 1897 3164 1903
rect 3188 1897 3308 1903
rect 3540 1897 3644 1903
rect 3860 1897 4108 1903
rect 4148 1897 4540 1903
rect 4836 1897 4924 1903
rect 4948 1897 5132 1903
rect 3101 1877 3148 1883
rect 3188 1877 3292 1883
rect 3316 1877 3523 1883
rect 68 1857 412 1863
rect 420 1857 460 1863
rect 564 1857 1219 1863
rect 564 1837 748 1843
rect 756 1837 1196 1843
rect 1213 1843 1219 1857
rect 1300 1857 1452 1863
rect 1556 1857 1804 1863
rect 1972 1857 2220 1863
rect 2244 1857 2380 1863
rect 2420 1857 2796 1863
rect 2804 1857 2972 1863
rect 2980 1857 3436 1863
rect 3444 1857 3500 1863
rect 3517 1863 3523 1877
rect 3604 1877 3756 1883
rect 3844 1877 3868 1883
rect 4029 1877 4668 1883
rect 4029 1863 4035 1877
rect 4676 1877 5027 1883
rect 3517 1857 4035 1863
rect 4292 1857 4380 1863
rect 4388 1857 4428 1863
rect 5021 1863 5027 1877
rect 5181 1883 5187 1903
rect 5140 1877 5187 1883
rect 4500 1857 5011 1863
rect 5021 1857 5084 1863
rect 1805 1844 1811 1856
rect 1213 1837 1340 1843
rect 1524 1837 1628 1843
rect 1828 1837 1884 1843
rect 1956 1837 2156 1843
rect 2173 1837 2268 1843
rect 228 1817 1132 1823
rect 1716 1817 1852 1823
rect 1860 1817 1948 1823
rect 2173 1823 2179 1837
rect 2292 1837 2332 1843
rect 2356 1837 2444 1843
rect 2452 1837 2588 1843
rect 2596 1837 2780 1843
rect 2852 1837 3276 1843
rect 3300 1837 3628 1843
rect 3636 1837 3804 1843
rect 3828 1837 4364 1843
rect 4548 1837 4588 1843
rect 4740 1837 4796 1843
rect 4820 1837 4956 1843
rect 5005 1843 5011 1857
rect 5092 1857 5148 1863
rect 5005 1837 5132 1843
rect 2004 1817 2179 1823
rect 2212 1817 2236 1823
rect 2308 1817 2348 1823
rect 2372 1817 2515 1823
rect 1236 1797 1276 1803
rect 1332 1797 1468 1803
rect 1748 1797 1996 1803
rect 2020 1797 2172 1803
rect 2180 1797 2492 1803
rect 2509 1803 2515 1817
rect 2644 1817 2748 1823
rect 2804 1817 2924 1823
rect 2964 1817 3356 1823
rect 3396 1817 3500 1823
rect 3508 1817 3532 1823
rect 4004 1817 4172 1823
rect 4436 1817 4524 1823
rect 4596 1817 5132 1823
rect 5181 1823 5187 1843
rect 5181 1817 5203 1823
rect 2546 1814 2606 1816
rect 2546 1806 2547 1814
rect 2556 1806 2557 1814
rect 2595 1806 2596 1814
rect 2605 1806 2606 1814
rect 2546 1804 2606 1806
rect 2509 1797 2531 1803
rect 356 1777 963 1783
rect 676 1757 764 1763
rect 852 1757 940 1763
rect 957 1763 963 1777
rect 1044 1777 1212 1783
rect 1588 1777 1644 1783
rect 1892 1777 1980 1783
rect 1988 1777 2140 1783
rect 2148 1777 2252 1783
rect 2292 1777 2460 1783
rect 2484 1777 2508 1783
rect 2525 1783 2531 1797
rect 2660 1797 2844 1803
rect 2868 1797 2924 1803
rect 2948 1797 3052 1803
rect 3204 1797 3468 1803
rect 3540 1797 3612 1803
rect 4148 1797 4444 1803
rect 4468 1797 4732 1803
rect 4740 1797 5116 1803
rect 5140 1797 5187 1803
rect 2525 1777 2556 1783
rect 2644 1777 2684 1783
rect 2756 1777 2908 1783
rect 2964 1777 3164 1783
rect 3172 1777 3420 1783
rect 3428 1777 3756 1783
rect 3908 1777 4236 1783
rect 4308 1777 4332 1783
rect 4340 1777 4492 1783
rect 5197 1783 5203 1817
rect 4532 1777 5203 1783
rect 957 1757 1676 1763
rect 1700 1757 2124 1763
rect 2164 1757 2716 1763
rect 2909 1763 2915 1776
rect 2909 1757 3484 1763
rect 3492 1757 3708 1763
rect 3716 1757 4348 1763
rect 4372 1757 4396 1763
rect 4516 1757 4652 1763
rect 4660 1757 4940 1763
rect 5124 1757 5187 1763
rect -35 1737 236 1743
rect 724 1737 876 1743
rect 884 1737 1116 1743
rect 1124 1737 1324 1743
rect 1332 1737 1644 1743
rect 1844 1737 1939 1743
rect 1933 1724 1939 1737
rect 2100 1737 2204 1743
rect 2212 1737 2316 1743
rect 2500 1737 2524 1743
rect 2548 1737 2572 1743
rect 2596 1737 2876 1743
rect 2996 1737 3292 1743
rect 3348 1737 3436 1743
rect 3588 1737 3676 1743
rect 4308 1737 4396 1743
rect 4484 1737 4780 1743
rect 4788 1737 4812 1743
rect 4996 1737 5116 1743
rect 132 1717 204 1723
rect 340 1717 588 1723
rect 676 1717 796 1723
rect 948 1717 1148 1723
rect 1364 1717 1468 1723
rect 1508 1717 1548 1723
rect 1604 1717 1900 1723
rect 2036 1717 2156 1723
rect 2180 1717 2220 1723
rect 2356 1717 2460 1723
rect 2484 1717 3276 1723
rect 3412 1717 3596 1723
rect 3732 1717 3884 1723
rect 4084 1717 4140 1723
rect 4564 1717 4700 1723
rect 4868 1717 5052 1723
rect 5076 1717 5132 1723
rect 5156 1717 5187 1723
rect -35 1697 92 1703
rect 100 1697 156 1703
rect 180 1697 300 1703
rect 500 1697 556 1703
rect 820 1697 1292 1703
rect 1812 1697 1916 1703
rect 2036 1697 2284 1703
rect 2324 1697 2700 1703
rect 2852 1697 3100 1703
rect 3124 1697 3324 1703
rect 3524 1697 3692 1703
rect 3764 1697 3900 1703
rect 3924 1697 4204 1703
rect 4276 1697 4300 1703
rect 4308 1697 4380 1703
rect 4388 1697 4476 1703
rect 4612 1697 4684 1703
rect 4692 1697 4780 1703
rect 4788 1697 4892 1703
rect 4900 1697 5068 1703
rect 196 1677 284 1683
rect 788 1677 828 1683
rect 836 1677 860 1683
rect 868 1677 1132 1683
rect 1140 1677 1180 1683
rect 1412 1677 1580 1683
rect 1588 1677 2060 1683
rect 2068 1677 2620 1683
rect 2676 1677 2844 1683
rect 2868 1677 2892 1683
rect 2900 1677 3548 1683
rect 3556 1677 3564 1683
rect 3572 1677 3612 1683
rect 3636 1677 3964 1683
rect 4020 1677 4252 1683
rect 4260 1677 4572 1683
rect 4740 1677 4764 1683
rect 4772 1677 4876 1683
rect 820 1657 1644 1663
rect 1956 1657 1980 1663
rect 1988 1657 2060 1663
rect 2068 1657 2252 1663
rect 2388 1657 2588 1663
rect 2612 1657 2860 1663
rect 2877 1657 3443 1663
rect 660 1637 1244 1643
rect 1252 1637 1324 1643
rect 1332 1637 1516 1643
rect 1524 1637 1596 1643
rect 1604 1637 1660 1643
rect 1668 1637 2188 1643
rect 2228 1637 2348 1643
rect 2404 1637 2428 1643
rect 2452 1637 2572 1643
rect 2877 1643 2883 1657
rect 2580 1637 2883 1643
rect 2932 1637 3011 1643
rect 548 1617 1020 1623
rect 1684 1617 2515 1623
rect 1042 1614 1102 1616
rect 1042 1606 1043 1614
rect 1052 1606 1053 1614
rect 1091 1606 1092 1614
rect 1101 1606 1102 1614
rect 1042 1604 1102 1606
rect 1284 1597 1532 1603
rect 1652 1597 1740 1603
rect 1812 1597 1875 1603
rect 596 1577 1443 1583
rect 1437 1564 1443 1577
rect 1572 1577 1852 1583
rect 1869 1583 1875 1597
rect 1908 1597 1996 1603
rect 2020 1597 2028 1603
rect 2180 1597 2220 1603
rect 2244 1597 2396 1603
rect 2436 1597 2444 1603
rect 2468 1597 2492 1603
rect 2509 1603 2515 1617
rect 2644 1617 2652 1623
rect 2708 1617 2828 1623
rect 2836 1617 2988 1623
rect 3005 1623 3011 1637
rect 3028 1637 3228 1643
rect 3236 1637 3420 1643
rect 3437 1643 3443 1657
rect 3492 1657 3532 1663
rect 3604 1657 3740 1663
rect 3812 1657 4524 1663
rect 3437 1637 3948 1643
rect 3005 1617 3164 1623
rect 3188 1617 3836 1623
rect 4050 1614 4110 1616
rect 4050 1606 4051 1614
rect 4060 1606 4061 1614
rect 4099 1606 4100 1614
rect 4109 1606 4110 1614
rect 4050 1604 4110 1606
rect 2509 1597 3859 1603
rect 1869 1577 1948 1583
rect 1988 1577 2124 1583
rect 2180 1577 2316 1583
rect 2324 1577 2412 1583
rect 2420 1577 2460 1583
rect 2468 1577 2620 1583
rect 2628 1577 2812 1583
rect 2820 1577 3116 1583
rect 3156 1577 3212 1583
rect 3268 1577 3299 1583
rect 484 1557 1356 1563
rect 1444 1557 1692 1563
rect 1716 1557 1740 1563
rect 1764 1557 1852 1563
rect 1924 1557 2044 1563
rect 2068 1557 2284 1563
rect 2388 1557 2940 1563
rect 2964 1557 3020 1563
rect 3044 1557 3276 1563
rect 3293 1563 3299 1577
rect 3332 1577 3468 1583
rect 3476 1577 3772 1583
rect 3780 1577 3836 1583
rect 3853 1583 3859 1597
rect 3853 1577 4860 1583
rect 3293 1557 3340 1563
rect 3508 1557 3644 1563
rect 3668 1557 4092 1563
rect 708 1537 908 1543
rect 948 1537 1116 1543
rect 1124 1537 1356 1543
rect 1364 1537 1996 1543
rect 2004 1537 2220 1543
rect 2228 1537 3292 1543
rect 3316 1537 3932 1543
rect 52 1517 204 1523
rect 436 1517 988 1523
rect 1092 1517 1308 1523
rect 1348 1517 1404 1523
rect 1428 1517 1708 1523
rect 1748 1517 1820 1523
rect 1844 1517 1884 1523
rect 1892 1517 2012 1523
rect 2100 1517 2236 1523
rect 2260 1517 2332 1523
rect 2340 1517 2556 1523
rect 2596 1517 2668 1523
rect 2685 1517 2908 1523
rect -35 1497 12 1503
rect 100 1497 172 1503
rect 180 1497 332 1503
rect 884 1497 924 1503
rect 1124 1497 1212 1503
rect 1236 1497 1452 1503
rect 1508 1497 1580 1503
rect 1732 1497 1836 1503
rect 1908 1497 1948 1503
rect 1988 1497 1996 1503
rect 2004 1497 2156 1503
rect 2308 1497 2476 1503
rect 2685 1503 2691 1517
rect 2964 1517 3004 1523
rect 3124 1517 3292 1523
rect 3380 1517 3587 1523
rect 3581 1504 3587 1517
rect 3700 1517 3756 1523
rect 4324 1517 4508 1523
rect 4516 1517 4556 1523
rect 2500 1497 2691 1503
rect 2708 1497 2764 1503
rect 2852 1497 2876 1503
rect 2900 1497 2940 1503
rect 2964 1497 2972 1503
rect 3060 1497 3084 1503
rect 3108 1497 3244 1503
rect 3252 1497 3516 1503
rect 3524 1497 3564 1503
rect 3588 1497 3660 1503
rect 3668 1497 3772 1503
rect 3988 1497 4204 1503
rect 4420 1497 4508 1503
rect 4724 1497 4780 1503
rect 4820 1497 4924 1503
rect 4932 1497 4972 1503
rect 4980 1497 5036 1503
rect 5044 1497 5100 1503
rect 532 1477 620 1483
rect 660 1477 700 1483
rect 836 1477 892 1483
rect 900 1477 940 1483
rect 980 1477 1036 1483
rect 1044 1477 1612 1483
rect 1620 1477 2092 1483
rect 2100 1477 2643 1483
rect 2637 1464 2643 1477
rect 2660 1477 2716 1483
rect 2772 1477 2796 1483
rect 2884 1477 2940 1483
rect 2948 1477 3068 1483
rect 3076 1477 3196 1483
rect 3204 1477 3372 1483
rect 3380 1477 3516 1483
rect 3636 1477 3836 1483
rect 4260 1477 4444 1483
rect 4452 1477 4700 1483
rect 1012 1457 1052 1463
rect 1060 1457 1164 1463
rect 1172 1457 1804 1463
rect 1812 1457 1916 1463
rect 1924 1457 2012 1463
rect 2020 1457 2076 1463
rect 2164 1457 2284 1463
rect 2356 1457 2604 1463
rect 3629 1463 3635 1476
rect 2644 1457 3635 1463
rect 3748 1457 4291 1463
rect 4285 1444 4291 1457
rect 676 1437 876 1443
rect 1028 1437 1164 1443
rect 1188 1437 2028 1443
rect 2036 1437 2444 1443
rect 2516 1437 2668 1443
rect 2676 1437 2860 1443
rect 2884 1437 3180 1443
rect 3252 1437 3404 1443
rect 3460 1437 3532 1443
rect 4292 1437 4476 1443
rect 4516 1437 4588 1443
rect 4596 1437 4860 1443
rect 692 1417 796 1423
rect 964 1417 1084 1423
rect 1108 1417 1324 1423
rect 1348 1417 1420 1423
rect 1684 1417 1724 1423
rect 1748 1417 1804 1423
rect 1892 1417 1948 1423
rect 1988 1417 2492 1423
rect 2676 1417 2892 1423
rect 2932 1417 2956 1423
rect 2980 1417 3180 1423
rect 3316 1417 3484 1423
rect 3572 1417 3692 1423
rect 3700 1417 3724 1423
rect 3764 1417 4140 1423
rect 2546 1414 2606 1416
rect 2546 1406 2547 1414
rect 2556 1406 2557 1414
rect 2595 1406 2596 1414
rect 2605 1406 2606 1414
rect 2546 1404 2606 1406
rect 20 1397 108 1403
rect 660 1397 828 1403
rect 884 1397 2268 1403
rect 2292 1397 2508 1403
rect 2676 1397 2812 1403
rect 2884 1397 2924 1403
rect 2964 1397 3020 1403
rect 3140 1397 3644 1403
rect 3661 1397 3772 1403
rect 52 1377 108 1383
rect 116 1377 300 1383
rect 788 1377 844 1383
rect 852 1377 1324 1383
rect 1332 1377 1516 1383
rect 1556 1377 1724 1383
rect 1748 1377 1772 1383
rect 1780 1377 1788 1383
rect 1940 1377 1996 1383
rect 2004 1377 2060 1383
rect 2068 1377 2275 1383
rect 244 1357 620 1363
rect 756 1357 796 1363
rect 820 1357 1100 1363
rect 1140 1357 1443 1363
rect -35 1337 12 1343
rect 148 1337 348 1343
rect 692 1337 780 1343
rect 900 1337 972 1343
rect 1156 1337 1212 1343
rect 1348 1337 1420 1343
rect 1437 1343 1443 1357
rect 1460 1357 1500 1363
rect 1508 1357 1804 1363
rect 1876 1357 2188 1363
rect 2269 1363 2275 1377
rect 2292 1377 2412 1383
rect 2436 1377 2476 1383
rect 2500 1377 2684 1383
rect 2724 1377 2780 1383
rect 2836 1377 3052 1383
rect 3060 1377 3084 1383
rect 3188 1377 3260 1383
rect 3661 1383 3667 1397
rect 4228 1397 4332 1403
rect 4340 1397 4444 1403
rect 4884 1397 5116 1403
rect 3284 1377 3667 1383
rect 3716 1377 3788 1383
rect 3796 1377 4732 1383
rect 4740 1377 4924 1383
rect 2269 1357 2652 1363
rect 2708 1357 2924 1363
rect 2964 1357 3036 1363
rect 3060 1357 3132 1363
rect 3172 1357 3212 1363
rect 3444 1357 3500 1363
rect 3556 1357 3596 1363
rect 3620 1357 3916 1363
rect 4132 1357 4348 1363
rect 5028 1357 5068 1363
rect 1437 1337 1740 1343
rect 1892 1337 1916 1343
rect 1940 1337 1987 1343
rect 420 1317 908 1323
rect 948 1317 1004 1323
rect 1108 1317 1308 1323
rect 1396 1317 1548 1323
rect 1620 1317 1644 1323
rect 1652 1317 1708 1323
rect 1716 1317 1740 1323
rect 1748 1317 1772 1323
rect 1796 1317 1964 1323
rect 1981 1323 1987 1337
rect 2052 1337 2252 1343
rect 2260 1337 2604 1343
rect 2644 1337 2675 1343
rect 2669 1324 2675 1337
rect 2708 1337 2972 1343
rect 3012 1337 3052 1343
rect 3092 1337 3308 1343
rect 3316 1337 3388 1343
rect 3396 1337 3628 1343
rect 3988 1337 4012 1343
rect 4052 1337 4428 1343
rect 4868 1337 4988 1343
rect 5028 1337 5036 1343
rect 1981 1317 2092 1323
rect 2196 1317 2652 1323
rect 2692 1317 2972 1323
rect 2996 1317 3244 1323
rect 3316 1317 3324 1323
rect 3364 1317 3635 1323
rect -35 1297 60 1303
rect 100 1297 412 1303
rect 541 1297 620 1303
rect 541 1283 547 1297
rect 740 1297 844 1303
rect 852 1297 1020 1303
rect 1188 1297 1276 1303
rect 1300 1297 1676 1303
rect 1844 1297 2220 1303
rect 2468 1297 2796 1303
rect 2836 1297 2876 1303
rect 2916 1297 2988 1303
rect 3028 1297 3219 1303
rect 340 1277 547 1283
rect 564 1277 940 1283
rect 996 1277 1212 1283
rect 1284 1277 1356 1283
rect 1428 1277 1436 1283
rect 1492 1277 1516 1283
rect 1604 1277 2300 1283
rect 2324 1277 2380 1283
rect 2445 1283 2451 1296
rect 2445 1277 2588 1283
rect 2612 1277 2732 1283
rect 2788 1277 2844 1283
rect 2852 1277 3132 1283
rect 3172 1277 3196 1283
rect 3213 1283 3219 1297
rect 3268 1297 3324 1303
rect 3332 1297 3596 1303
rect 3629 1303 3635 1317
rect 3652 1317 3740 1323
rect 4260 1317 4348 1323
rect 4500 1317 4636 1323
rect 4708 1317 4892 1323
rect 4900 1317 5052 1323
rect 3629 1297 3772 1303
rect 3780 1297 3916 1303
rect 4308 1297 4316 1303
rect 4324 1297 4396 1303
rect 4452 1297 4492 1303
rect 4500 1297 4572 1303
rect 3213 1277 3276 1283
rect 3348 1277 3404 1283
rect 3412 1277 3564 1283
rect 5076 1277 5100 1283
rect 340 1257 364 1263
rect 836 1257 1980 1263
rect 2004 1257 2092 1263
rect 2164 1257 2284 1263
rect 2308 1257 2467 1263
rect 1076 1237 1196 1243
rect 1204 1237 1788 1243
rect 1812 1237 2028 1243
rect 2052 1237 2412 1243
rect 2436 1237 2444 1243
rect 2461 1243 2467 1257
rect 2532 1257 2812 1263
rect 2868 1257 3180 1263
rect 3236 1257 3500 1263
rect 3556 1257 3676 1263
rect 3684 1257 4524 1263
rect 2461 1237 3196 1243
rect 3300 1237 3372 1243
rect 3492 1237 3564 1243
rect 3572 1237 3980 1243
rect 4884 1237 5100 1243
rect 1348 1217 1404 1223
rect 1476 1217 2220 1223
rect 2228 1217 2380 1223
rect 2388 1217 2828 1223
rect 2868 1217 3468 1223
rect 3508 1217 3660 1223
rect 4676 1217 4908 1223
rect 4916 1217 5068 1223
rect 5076 1217 5187 1223
rect 1042 1214 1102 1216
rect 1042 1206 1043 1214
rect 1052 1206 1053 1214
rect 1091 1206 1092 1214
rect 1101 1206 1102 1214
rect 1042 1204 1102 1206
rect 4050 1214 4110 1216
rect 4050 1206 4051 1214
rect 4060 1206 4061 1214
rect 4099 1206 4100 1214
rect 4109 1206 4110 1214
rect 4050 1204 4110 1206
rect 1124 1197 1580 1203
rect 1780 1197 2108 1203
rect 2116 1197 2188 1203
rect 2228 1197 2460 1203
rect 2484 1197 2956 1203
rect 2996 1197 3036 1203
rect 3140 1197 3180 1203
rect 3220 1197 3804 1203
rect 4708 1197 5084 1203
rect 5092 1197 5148 1203
rect 5181 1197 5187 1217
rect 932 1177 1132 1183
rect 1140 1177 1484 1183
rect 1492 1177 2444 1183
rect 2468 1177 2828 1183
rect 2836 1177 3148 1183
rect 3172 1177 3788 1183
rect 3796 1177 3868 1183
rect 3988 1177 4044 1183
rect 4436 1177 4652 1183
rect 4996 1177 5084 1183
rect 228 1157 812 1163
rect 884 1157 1116 1163
rect 1204 1157 1420 1163
rect 1492 1157 1564 1163
rect 1588 1157 3004 1163
rect 3620 1157 3708 1163
rect 3716 1157 4124 1163
rect 4141 1157 4716 1163
rect 276 1137 556 1143
rect 596 1137 716 1143
rect 804 1137 988 1143
rect 996 1137 1244 1143
rect 1380 1137 1420 1143
rect 1428 1137 1548 1143
rect 1556 1137 1596 1143
rect 1604 1137 1820 1143
rect 1828 1137 1852 1143
rect 1892 1137 1932 1143
rect 1940 1137 2060 1143
rect 2148 1137 2156 1143
rect 2212 1137 2252 1143
rect 2269 1137 2764 1143
rect 52 1117 300 1123
rect 308 1117 364 1123
rect 724 1117 860 1123
rect 1220 1117 1340 1123
rect 1364 1117 1548 1123
rect 1588 1117 1612 1123
rect 1620 1117 1660 1123
rect 1700 1117 1756 1123
rect 1764 1117 1811 1123
rect -35 1097 12 1103
rect 276 1097 316 1103
rect 500 1097 556 1103
rect 852 1097 892 1103
rect 964 1097 1100 1103
rect 1236 1097 1324 1103
rect 1332 1097 1452 1103
rect 1524 1097 1612 1103
rect 1748 1097 1788 1103
rect 1805 1103 1811 1117
rect 1844 1117 1884 1123
rect 2020 1117 2124 1123
rect 2269 1123 2275 1137
rect 2948 1137 3004 1143
rect 3668 1137 3756 1143
rect 4141 1143 4147 1157
rect 5012 1157 5187 1163
rect 3764 1137 4147 1143
rect 4628 1137 4652 1143
rect 4852 1137 5020 1143
rect 5044 1137 5100 1143
rect 2164 1117 2275 1123
rect 2340 1117 2348 1123
rect 2404 1117 2460 1123
rect 2484 1117 2636 1123
rect 2660 1117 2700 1123
rect 2724 1117 2860 1123
rect 2900 1117 3068 1123
rect 3076 1117 3196 1123
rect 3204 1117 3244 1123
rect 3476 1117 3548 1123
rect 3604 1117 3628 1123
rect 3908 1117 3980 1123
rect 4020 1117 4220 1123
rect 4580 1117 4620 1123
rect 4724 1117 4908 1123
rect 4948 1117 5004 1123
rect 5156 1117 5187 1123
rect 1805 1097 1916 1103
rect 1924 1097 1948 1103
rect 1972 1097 2044 1103
rect 2068 1097 2124 1103
rect 2141 1097 2364 1103
rect 260 1077 348 1083
rect 612 1077 636 1083
rect 788 1077 995 1083
rect 804 1057 972 1063
rect 989 1063 995 1077
rect 1092 1077 1164 1083
rect 1172 1077 1180 1083
rect 1188 1077 1372 1083
rect 1380 1077 1868 1083
rect 1876 1077 1900 1083
rect 2141 1083 2147 1097
rect 2468 1097 2604 1103
rect 2868 1097 2908 1103
rect 2980 1097 3116 1103
rect 3124 1097 3228 1103
rect 3236 1097 3260 1103
rect 3444 1097 3548 1103
rect 3556 1097 4012 1103
rect 4484 1097 4572 1103
rect 4852 1097 4956 1103
rect 4996 1097 5020 1103
rect 5028 1097 5068 1103
rect 5076 1097 5084 1103
rect 1972 1077 2147 1083
rect 2196 1077 2236 1083
rect 2244 1077 2284 1083
rect 2420 1077 2652 1083
rect 2820 1077 2956 1083
rect 2996 1077 3404 1083
rect 3764 1077 3820 1083
rect 3908 1077 3980 1083
rect 989 1057 1100 1063
rect 1124 1057 1292 1063
rect 1348 1057 1516 1063
rect 1556 1057 1660 1063
rect 1732 1057 1772 1063
rect 1844 1057 2268 1063
rect 2276 1057 2364 1063
rect 2484 1057 2636 1063
rect 2740 1057 2860 1063
rect 2964 1057 3068 1063
rect 3092 1057 3132 1063
rect 3380 1057 3724 1063
rect 3812 1057 3868 1063
rect 4564 1057 4604 1063
rect 532 1037 1356 1043
rect 1428 1037 1708 1043
rect 1732 1037 1852 1043
rect 2068 1037 2083 1043
rect 564 1017 604 1023
rect 612 1017 700 1023
rect 708 1017 748 1023
rect 948 1017 988 1023
rect 1012 1017 1196 1023
rect 1204 1017 1228 1023
rect 1236 1017 1308 1023
rect 1316 1017 1484 1023
rect 1492 1017 1964 1023
rect 1972 1017 2060 1023
rect 2077 1023 2083 1037
rect 2100 1037 2124 1043
rect 2148 1037 2627 1043
rect 2077 1017 2156 1023
rect 2292 1017 2476 1023
rect 2621 1023 2627 1037
rect 2660 1037 2988 1043
rect 3060 1037 3100 1043
rect 3124 1037 3180 1043
rect 3188 1037 4348 1043
rect 4356 1037 4540 1043
rect 4612 1037 4684 1043
rect 2621 1017 4147 1023
rect 2546 1014 2606 1016
rect 2546 1006 2547 1014
rect 2556 1006 2557 1014
rect 2595 1006 2596 1014
rect 2605 1006 2606 1014
rect 2546 1004 2606 1006
rect 4141 1004 4147 1017
rect 692 997 2444 1003
rect 2628 997 2828 1003
rect 2868 997 2956 1003
rect 3028 997 3452 1003
rect 3540 997 3740 1003
rect 3748 997 3948 1003
rect 4148 997 4300 1003
rect 4628 997 4636 1003
rect 692 977 876 983
rect 980 977 1196 983
rect 1300 977 1356 983
rect 1396 977 1500 983
rect 1508 977 1580 983
rect 1588 977 1628 983
rect 1668 977 1724 983
rect 1748 977 1987 983
rect 1981 964 1987 977
rect 2116 977 2252 983
rect 2269 977 2396 983
rect 596 957 1219 963
rect -35 937 60 943
rect 164 937 236 943
rect 436 937 492 943
rect 532 937 732 943
rect 900 937 1036 943
rect 1188 937 1196 943
rect 1213 943 1219 957
rect 1332 957 1660 963
rect 1684 957 1756 963
rect 1821 957 1948 963
rect 1821 944 1827 957
rect 1988 957 2140 963
rect 2269 963 2275 977
rect 2420 977 4508 983
rect 2228 957 2275 963
rect 2308 957 2412 963
rect 2429 957 3100 963
rect 1213 937 1388 943
rect 1460 937 1644 943
rect 1652 937 1756 943
rect 1876 937 2092 943
rect 2429 943 2435 957
rect 3188 957 3516 963
rect 3533 957 4396 963
rect 2164 937 2435 943
rect 2452 937 2620 943
rect 2772 937 2844 943
rect 2884 937 2908 943
rect 2932 937 2956 943
rect 2964 937 3148 943
rect 3252 937 3356 943
rect 3533 943 3539 957
rect 4404 957 4588 963
rect 4820 957 4876 963
rect 3444 937 3539 943
rect 3604 937 3628 943
rect 4052 937 4300 943
rect 4308 937 4476 943
rect 4532 937 4652 943
rect 4692 937 4940 943
rect 5028 937 5052 943
rect 52 917 108 923
rect 148 917 252 923
rect 292 917 492 923
rect 644 917 684 923
rect 740 917 828 923
rect 996 917 1116 923
rect 1188 917 1212 923
rect 1236 917 1340 923
rect 1380 917 1452 923
rect 1524 917 1596 923
rect 1620 917 1731 923
rect -35 897 12 903
rect 100 897 284 903
rect 756 897 1260 903
rect 1300 897 1388 903
rect 1412 897 1532 903
rect 1604 897 1708 903
rect 1725 903 1731 917
rect 1748 917 1772 923
rect 1860 917 1932 923
rect 1956 917 2019 923
rect 1725 897 1868 903
rect 1940 897 1996 903
rect 2013 903 2019 917
rect 2084 917 2220 923
rect 2228 917 2300 923
rect 2340 917 2380 923
rect 2484 917 2547 923
rect 2013 897 2188 903
rect 2388 897 2524 903
rect 2541 903 2547 917
rect 2644 917 2780 923
rect 2804 917 2876 923
rect 2900 917 3228 923
rect 3268 917 3388 923
rect 3572 917 3644 923
rect 3748 917 3820 923
rect 3844 917 3964 923
rect 4276 917 4348 923
rect 4388 917 4620 923
rect 4644 917 4780 923
rect 4788 917 4924 923
rect 2541 897 2796 903
rect 2820 897 2988 903
rect 2996 897 3084 903
rect 3108 897 4684 903
rect 4980 897 5187 903
rect 148 877 172 883
rect 564 877 812 883
rect 836 877 1612 883
rect 1636 877 1660 883
rect 1677 877 1692 883
rect 916 857 1004 863
rect 1012 857 1532 863
rect 1677 863 1683 877
rect 1700 877 2156 883
rect 2164 877 4604 883
rect 4676 877 4988 883
rect 1540 857 1683 863
rect 1693 857 2268 863
rect 340 837 652 843
rect 756 837 1196 843
rect 1693 843 1699 857
rect 2356 857 2492 863
rect 2500 857 2812 863
rect 2836 857 2892 863
rect 2932 857 3132 863
rect 3140 857 3500 863
rect 3508 857 3692 863
rect 3860 857 3884 863
rect 4084 857 4300 863
rect 4628 857 4748 863
rect 1220 837 1699 843
rect 1780 837 2204 843
rect 2244 837 2300 843
rect 2308 837 2556 843
rect 2925 843 2931 856
rect 2564 837 2931 843
rect 2948 837 3020 843
rect 3044 837 3580 843
rect 3828 837 4396 843
rect 788 817 972 823
rect 1364 817 2460 823
rect 2484 817 2732 823
rect 2740 817 2972 823
rect 3092 817 3612 823
rect 3620 817 3772 823
rect 1042 814 1102 816
rect 1042 806 1043 814
rect 1052 806 1053 814
rect 1091 806 1092 814
rect 1101 806 1102 814
rect 1042 804 1102 806
rect 4050 814 4110 816
rect 4050 806 4051 814
rect 4060 806 4061 814
rect 4099 806 4100 814
rect 4109 806 4110 814
rect 4050 804 4110 806
rect 692 797 1020 803
rect 1156 797 1676 803
rect 1700 797 2060 803
rect 2100 797 2172 803
rect 2180 797 2396 803
rect 2404 797 2659 803
rect 1012 777 1180 783
rect 1204 777 2316 783
rect 2340 777 2348 783
rect 2388 777 2636 783
rect 2653 783 2659 797
rect 2692 797 2748 803
rect 2788 797 3036 803
rect 3156 797 3804 803
rect 3812 797 3884 803
rect 4564 797 4620 803
rect 4660 797 4860 803
rect 4868 797 5004 803
rect 5012 797 5052 803
rect 2653 777 3276 783
rect 3284 777 4364 783
rect 4452 777 5132 783
rect 228 757 1740 763
rect 1764 757 2364 763
rect 2388 757 2620 763
rect 2644 757 2780 763
rect 2804 757 2908 763
rect 2932 757 3180 763
rect 3252 757 3292 763
rect 3309 757 4563 763
rect -35 737 12 743
rect 52 737 156 743
rect 164 737 396 743
rect 436 737 508 743
rect 644 737 716 743
rect 932 737 1052 743
rect 1076 737 1228 743
rect 1316 737 1404 743
rect 3309 743 3315 757
rect 4557 744 4563 757
rect 4996 757 5068 763
rect 1412 737 3315 743
rect 3348 737 3484 743
rect 3492 737 3948 743
rect 3956 737 4140 743
rect 4564 737 4748 743
rect 4836 737 5036 743
rect 356 717 460 723
rect 820 717 940 723
rect 1044 717 1132 723
rect 1300 717 1340 723
rect 1588 717 1660 723
rect 1972 717 2108 723
rect 2164 717 2236 723
rect 2244 717 2348 723
rect 2404 717 2531 723
rect -35 697 12 703
rect 20 697 60 703
rect 68 697 108 703
rect 292 697 524 703
rect 772 697 1196 703
rect 1284 697 1324 703
rect 1348 697 1452 703
rect 1476 697 1516 703
rect 1533 697 1596 703
rect 68 677 556 683
rect 564 677 572 683
rect 1012 677 1020 683
rect 1268 677 1356 683
rect 1364 677 1420 683
rect 1533 683 1539 697
rect 1636 697 1788 703
rect 1988 697 2060 703
rect 2084 697 2092 703
rect 2132 697 2316 703
rect 2340 697 2380 703
rect 2484 697 2508 703
rect 2525 703 2531 717
rect 2580 717 2636 723
rect 2692 717 2748 723
rect 2772 717 2924 723
rect 2948 717 3052 723
rect 3076 717 3148 723
rect 3172 717 3212 723
rect 3220 717 3356 723
rect 3604 717 3628 723
rect 3780 717 3852 723
rect 4084 717 4252 723
rect 4548 717 4556 723
rect 4692 717 4796 723
rect 4884 717 5068 723
rect 2525 697 2588 703
rect 2628 697 2716 703
rect 2733 697 3219 703
rect 1492 677 1539 683
rect 1556 677 1660 683
rect 1684 677 1756 683
rect 1924 677 2108 683
rect 2116 677 2156 683
rect 2180 677 2188 683
rect 2276 677 2380 683
rect 2420 677 2492 683
rect 2644 677 2668 683
rect 2733 683 2739 697
rect 3213 684 3219 697
rect 3236 697 3324 703
rect 3556 697 3932 703
rect 3940 697 3948 703
rect 4244 697 4284 703
rect 4292 697 4300 703
rect 4772 697 4892 703
rect 4900 697 5187 703
rect 2724 677 2739 683
rect 2788 677 2876 683
rect 2884 677 3036 683
rect 3124 677 3164 683
rect 3220 677 3244 683
rect 3268 677 3308 683
rect 3332 677 3436 683
rect 3636 677 3836 683
rect 3892 677 3980 683
rect 4244 677 4444 683
rect 4516 677 4956 683
rect 388 657 428 663
rect 436 657 540 663
rect 548 657 748 663
rect 820 657 844 663
rect 948 657 1244 663
rect 1332 657 1708 663
rect 1716 657 1836 663
rect 1892 657 2172 663
rect 2189 657 2684 663
rect 100 637 444 643
rect 596 637 1548 643
rect 1588 637 1596 643
rect 1668 637 1772 643
rect 1796 637 1964 643
rect 2189 643 2195 657
rect 2756 657 2780 663
rect 2852 657 2956 663
rect 3124 657 3596 663
rect 3604 657 3644 663
rect 4724 657 4972 663
rect 2036 637 2195 643
rect 2372 637 2771 643
rect 2765 624 2771 637
rect 2820 637 4460 643
rect 148 617 764 623
rect 772 617 1340 623
rect 1588 617 1772 623
rect 1780 617 1996 623
rect 2004 617 2076 623
rect 2116 617 2348 623
rect 2772 617 2892 623
rect 3012 617 3372 623
rect 3396 617 3708 623
rect 4308 617 4620 623
rect 4628 617 4636 623
rect 2546 614 2606 616
rect 2546 606 2547 614
rect 2556 606 2557 614
rect 2595 606 2596 614
rect 2605 606 2606 614
rect 2546 604 2606 606
rect 1172 597 1676 603
rect 1748 597 2204 603
rect 2660 597 2812 603
rect 2964 597 3068 603
rect 3092 597 3324 603
rect 3332 597 3891 603
rect 564 577 892 583
rect 1012 577 1196 583
rect 1236 577 1596 583
rect 1604 577 1724 583
rect 1732 577 2044 583
rect 2052 577 2172 583
rect 2180 577 2236 583
rect 2308 577 2396 583
rect 2404 577 2412 583
rect 2589 577 2620 583
rect 340 557 524 563
rect 740 557 844 563
rect 852 557 892 563
rect 916 557 1740 563
rect 1860 557 1900 563
rect 1908 557 1932 563
rect 1972 557 1980 563
rect 1997 557 2124 563
rect 516 537 524 543
rect 580 537 620 543
rect 660 537 876 543
rect 884 537 1052 543
rect 1060 537 1548 543
rect 1636 537 1868 543
rect 1997 543 2003 557
rect 2228 557 2268 563
rect 2589 563 2595 577
rect 2740 577 2828 583
rect 2836 577 3020 583
rect 3220 577 3340 583
rect 3364 577 3500 583
rect 3885 583 3891 597
rect 3908 597 3948 603
rect 4116 597 4252 603
rect 4260 597 4332 603
rect 4349 597 4908 603
rect 4349 583 4355 597
rect 3508 577 3811 583
rect 3885 577 4355 583
rect 2324 557 2595 563
rect 2612 557 2636 563
rect 2676 557 2908 563
rect 2964 557 3036 563
rect 3060 557 3148 563
rect 3188 557 3260 563
rect 3284 557 3436 563
rect 3444 557 3516 563
rect 3805 563 3811 577
rect 4388 577 4828 583
rect 3805 557 4092 563
rect 4228 557 4332 563
rect 4372 557 4732 563
rect 1972 537 2003 543
rect 2100 537 2252 543
rect 2260 537 2444 543
rect 2532 537 2828 543
rect 2836 537 2940 543
rect 3028 537 3340 543
rect 3380 537 3420 543
rect 3604 537 3756 543
rect 3908 537 4380 543
rect 4660 537 4716 543
rect 4852 537 4908 543
rect 4916 537 4940 543
rect 292 517 460 523
rect 516 517 547 523
rect -35 497 12 503
rect 436 497 524 503
rect 541 503 547 517
rect 692 517 1260 523
rect 1268 517 1420 523
rect 1524 517 1612 523
rect 1716 517 1884 523
rect 1924 517 2060 523
rect 2116 517 2188 523
rect 2276 517 2316 523
rect 2340 517 2396 523
rect 2516 517 2764 523
rect 2772 517 3100 523
rect 3108 517 3180 523
rect 3188 517 3516 523
rect 3620 517 3692 523
rect 3796 517 3852 523
rect 4100 517 4284 523
rect 4324 517 4364 523
rect 4372 517 4428 523
rect 4436 517 4460 523
rect 4708 517 4780 523
rect 4788 517 4876 523
rect 4884 517 4892 523
rect 541 497 908 503
rect 932 497 956 503
rect 996 497 1068 503
rect 1668 497 1932 503
rect 2084 497 2124 503
rect 2132 497 2188 503
rect 2212 497 2684 503
rect 2708 497 2780 503
rect 2804 497 2908 503
rect 2916 497 2972 503
rect 2989 497 3180 503
rect 52 477 204 483
rect 212 477 396 483
rect 436 477 460 483
rect 628 477 1580 483
rect 1748 477 2028 483
rect 2196 477 2460 483
rect 2580 477 2652 483
rect 2660 477 2716 483
rect 2724 477 2732 483
rect 2989 483 2995 497
rect 3300 497 3308 503
rect 3460 497 3644 503
rect 3940 497 4012 503
rect 2772 477 2995 483
rect 3028 477 3116 483
rect 3252 477 3580 483
rect 3620 477 3852 483
rect 4692 477 4796 483
rect 4804 477 4860 483
rect 484 457 588 463
rect 836 457 972 463
rect 1028 457 1132 463
rect 1140 457 1548 463
rect 1556 457 1676 463
rect 1684 457 1804 463
rect 2228 457 2252 463
rect 2260 457 2332 463
rect 2500 457 2636 463
rect 2644 457 2700 463
rect 2708 457 2812 463
rect 2916 457 3132 463
rect 3140 457 3468 463
rect 3828 457 3852 463
rect 1124 437 1292 443
rect 1332 437 1740 443
rect 2180 437 2668 443
rect 2676 437 2988 443
rect 2996 437 3388 443
rect 2548 417 2620 423
rect 2644 417 3372 423
rect 1042 414 1102 416
rect 1042 406 1043 414
rect 1052 406 1053 414
rect 1091 406 1092 414
rect 1101 406 1102 414
rect 1042 404 1102 406
rect 4050 414 4110 416
rect 4050 406 4051 414
rect 4060 406 4061 414
rect 4099 406 4100 414
rect 4109 406 4110 414
rect 4050 404 4110 406
rect 1252 397 1724 403
rect 1780 397 2044 403
rect 2164 397 2924 403
rect 2948 397 3084 403
rect 3156 397 4012 403
rect 500 377 940 383
rect 964 377 1043 383
rect 148 357 572 363
rect 964 357 1020 363
rect 1037 363 1043 377
rect 1348 377 1484 383
rect 1892 377 1916 383
rect 2388 377 3820 383
rect 3828 377 3916 383
rect 4020 377 4188 383
rect 4772 377 4860 383
rect 4868 377 4956 383
rect 1037 357 2604 363
rect 2676 357 3004 363
rect 3124 357 3436 363
rect 3444 357 3532 363
rect 3572 357 3628 363
rect 4164 357 4572 363
rect 20 337 460 343
rect 628 337 988 343
rect 1860 337 2243 343
rect 948 317 1324 323
rect 1332 317 1340 323
rect 1348 317 1612 323
rect 1620 317 1868 323
rect 1924 317 2012 323
rect 2148 317 2220 323
rect 2237 323 2243 337
rect 2340 337 2572 343
rect 2612 337 2636 343
rect 2660 337 2700 343
rect 2804 337 2876 343
rect 2900 337 3228 343
rect 3236 337 4812 343
rect 4820 337 4908 343
rect 2237 317 2764 323
rect 2820 317 2892 323
rect 2973 317 3004 323
rect 436 297 540 303
rect 644 297 1292 303
rect 1364 297 1628 303
rect 1812 297 1948 303
rect 1988 297 2252 303
rect 2260 297 2364 303
rect 2644 297 2684 303
rect 2740 297 2748 303
rect 2772 297 2860 303
rect 2973 303 2979 317
rect 3076 317 3084 323
rect 3124 317 3164 323
rect 3188 317 3340 323
rect 3572 317 3644 323
rect 3956 317 4044 323
rect 4052 317 4156 323
rect 4500 317 4668 323
rect 2900 297 2979 303
rect 2996 297 3660 303
rect 3668 297 3788 303
rect 3796 297 3884 303
rect 3956 297 3980 303
rect 4148 297 4268 303
rect 4676 297 4764 303
rect 4900 297 5004 303
rect 356 277 444 283
rect 452 277 508 283
rect 516 277 716 283
rect 772 277 940 283
rect 1332 277 1356 283
rect 1556 277 1724 283
rect 1956 277 2156 283
rect 2308 277 2444 283
rect 2452 277 2780 283
rect 2788 277 3036 283
rect 3188 277 3196 283
rect 3204 277 3308 283
rect 3348 277 3395 283
rect 1412 257 1580 263
rect 1908 257 1964 263
rect 1972 257 2060 263
rect 2068 257 2092 263
rect 2212 257 2284 263
rect 2292 257 2636 263
rect 2644 257 3148 263
rect 3156 257 3244 263
rect 3252 257 3324 263
rect 3364 257 3372 263
rect 3389 263 3395 277
rect 3412 277 3692 283
rect 3700 277 3756 283
rect 3988 277 4252 283
rect 4548 277 4684 283
rect 3389 257 3532 263
rect 3661 257 3740 263
rect 3661 244 3667 257
rect 4388 257 4620 263
rect 708 237 796 243
rect 804 237 892 243
rect 1012 237 1196 243
rect 1204 237 1244 243
rect 1252 237 1308 243
rect 1604 237 2156 243
rect 2196 237 2396 243
rect 2413 237 2883 243
rect 2413 223 2419 237
rect 996 217 2419 223
rect 2628 217 2860 223
rect 2877 223 2883 237
rect 3092 237 3404 243
rect 3428 237 3660 243
rect 3684 237 4172 243
rect 4180 237 4444 243
rect 2877 217 3116 223
rect 3156 217 3212 223
rect 3236 217 3276 223
rect 3300 217 3340 223
rect 3364 217 3468 223
rect 3492 217 4380 223
rect 2546 214 2606 216
rect 2546 206 2547 214
rect 2556 206 2557 214
rect 2595 206 2596 214
rect 2605 206 2606 214
rect 2546 204 2606 206
rect 340 197 428 203
rect 1140 197 1196 203
rect 2100 197 2188 203
rect 2372 197 2508 203
rect 2708 197 3484 203
rect 3604 197 3852 203
rect 4244 197 4556 203
rect 4564 197 4636 203
rect 4804 197 4924 203
rect 452 177 1260 183
rect 1364 177 1372 183
rect 1380 177 1420 183
rect 1668 177 1692 183
rect 2084 177 2364 183
rect 2388 177 4716 183
rect 4724 177 4812 183
rect 468 157 1148 163
rect 1300 157 2220 163
rect 2356 157 2492 163
rect 2500 157 2700 163
rect 2788 157 2828 163
rect 2868 157 3020 163
rect 3053 157 3532 163
rect -35 137 60 143
rect 228 137 588 143
rect 596 137 812 143
rect 820 137 844 143
rect 932 137 1132 143
rect 1188 137 1212 143
rect 1556 137 1580 143
rect 2036 137 2140 143
rect 2340 137 2380 143
rect 2701 143 2707 156
rect 2701 137 2892 143
rect 2909 137 2940 143
rect 244 117 412 123
rect 548 117 732 123
rect 772 117 1132 123
rect 1796 117 1804 123
rect 1828 117 1964 123
rect 2132 117 2172 123
rect 2276 117 2316 123
rect 2324 117 2851 123
rect -35 97 12 103
rect 116 97 300 103
rect 340 97 412 103
rect 772 97 1004 103
rect 1204 97 1260 103
rect 2020 97 2220 103
rect 2260 97 2348 103
rect 2452 97 2668 103
rect 2676 97 2796 103
rect 2845 103 2851 117
rect 2909 123 2915 137
rect 3053 143 3059 157
rect 3668 157 3692 163
rect 4020 157 4188 163
rect 2996 137 3059 143
rect 3188 137 3244 143
rect 3300 137 3308 143
rect 3332 137 3372 143
rect 3812 137 4236 143
rect 4260 137 4540 143
rect 4612 137 4700 143
rect 4788 137 4876 143
rect 5140 137 5187 143
rect 2868 117 2915 123
rect 2932 117 2972 123
rect 2980 117 2988 123
rect 3012 117 3196 123
rect 3236 117 3244 123
rect 3252 117 3276 123
rect 3316 117 3580 123
rect 4180 117 4220 123
rect 4228 117 4460 123
rect 4468 117 4508 123
rect 2845 97 2883 103
rect 1972 77 2412 83
rect 2420 77 2780 83
rect 2836 77 2860 83
rect 2877 83 2883 97
rect 2900 97 3228 103
rect 3380 97 3612 103
rect 3620 97 3884 103
rect 3892 97 4140 103
rect 4388 97 4476 103
rect 2877 77 3004 83
rect 3140 77 3148 83
rect 3172 77 3564 83
rect 3572 77 4252 83
rect 2164 57 2636 63
rect 2644 57 2684 63
rect 2692 57 3212 63
rect 3396 57 3628 63
rect 1044 37 1132 43
rect 1252 37 3388 43
rect 3933 37 4620 43
rect 1124 17 1164 23
rect 2772 17 3324 23
rect 3933 23 3939 37
rect 3332 17 3939 23
rect 1042 14 1102 16
rect 1042 6 1043 14
rect 1052 6 1053 14
rect 1091 6 1092 14
rect 1101 6 1102 14
rect 1042 4 1102 6
rect 4050 14 4110 16
rect 4050 6 4051 14
rect 4060 6 4061 14
rect 4099 6 4100 14
rect 4109 6 4110 14
rect 4050 4 4110 6
<< m4contact >>
rect 3852 3416 3860 3424
rect 2548 3406 2555 3414
rect 2555 3406 2556 3414
rect 2560 3406 2565 3414
rect 2565 3406 2567 3414
rect 2567 3406 2568 3414
rect 2572 3406 2575 3414
rect 2575 3406 2577 3414
rect 2577 3406 2580 3414
rect 2584 3406 2585 3414
rect 2585 3406 2587 3414
rect 2587 3406 2592 3414
rect 2596 3406 2597 3414
rect 2597 3406 2604 3414
rect 1516 3376 1524 3384
rect 1644 3356 1652 3364
rect 2252 3356 2260 3364
rect 2636 3356 2644 3364
rect 2188 3336 2196 3344
rect 2988 3336 2996 3344
rect 1292 3316 1300 3324
rect 1900 3316 1908 3324
rect 2636 3316 2644 3324
rect 2732 3316 2740 3324
rect 3916 3316 3924 3324
rect 2988 3296 2996 3304
rect 2124 3276 2132 3284
rect 2476 3276 2484 3284
rect 2284 3216 2292 3224
rect 1044 3206 1051 3214
rect 1051 3206 1052 3214
rect 1056 3206 1061 3214
rect 1061 3206 1063 3214
rect 1063 3206 1064 3214
rect 1068 3206 1071 3214
rect 1071 3206 1073 3214
rect 1073 3206 1076 3214
rect 1080 3206 1081 3214
rect 1081 3206 1083 3214
rect 1083 3206 1088 3214
rect 1092 3206 1093 3214
rect 1093 3206 1100 3214
rect 2156 3196 2164 3204
rect 2892 3236 2900 3244
rect 4052 3206 4059 3214
rect 4059 3206 4060 3214
rect 4064 3206 4069 3214
rect 4069 3206 4071 3214
rect 4071 3206 4072 3214
rect 4076 3206 4079 3214
rect 4079 3206 4081 3214
rect 4081 3206 4084 3214
rect 4088 3206 4089 3214
rect 4089 3206 4091 3214
rect 4091 3206 4096 3214
rect 4100 3206 4101 3214
rect 4101 3206 4108 3214
rect 716 3176 724 3184
rect 2924 3176 2932 3184
rect 3724 3136 3732 3144
rect 1164 3116 1172 3124
rect 1388 3116 1396 3124
rect 1484 3116 1492 3124
rect 2636 3116 2644 3124
rect 812 3096 820 3104
rect 1196 3096 1204 3104
rect 1612 3096 1620 3104
rect 1996 3096 2004 3104
rect 2060 3096 2068 3104
rect 2732 3096 2740 3104
rect 2988 3096 2996 3104
rect 1164 3076 1172 3084
rect 2028 3076 2036 3084
rect 2284 3076 2292 3084
rect 1388 3036 1396 3044
rect 2636 3056 2644 3064
rect 4460 3076 4468 3084
rect 2548 3006 2555 3014
rect 2555 3006 2556 3014
rect 2560 3006 2565 3014
rect 2565 3006 2567 3014
rect 2567 3006 2568 3014
rect 2572 3006 2575 3014
rect 2575 3006 2577 3014
rect 2577 3006 2580 3014
rect 2584 3006 2585 3014
rect 2585 3006 2587 3014
rect 2587 3006 2592 3014
rect 2596 3006 2597 3014
rect 2597 3006 2604 3014
rect 1708 2976 1716 2984
rect 620 2956 628 2964
rect 876 2936 884 2944
rect 4172 2976 4180 2984
rect 4300 2976 4308 2984
rect 2668 2956 2676 2964
rect 3084 2956 3092 2964
rect 1644 2936 1652 2944
rect 1868 2936 1876 2944
rect 2028 2936 2036 2944
rect 2156 2936 2164 2944
rect 2220 2936 2228 2944
rect 4876 2956 4884 2964
rect 844 2916 852 2924
rect 1324 2916 1332 2924
rect 1516 2916 1524 2924
rect 2252 2916 2260 2924
rect 1644 2896 1652 2904
rect 1708 2896 1716 2904
rect 2444 2896 2452 2904
rect 2892 2896 2900 2904
rect 4460 2916 4468 2924
rect 5100 2896 5108 2904
rect 972 2876 980 2884
rect 1292 2876 1300 2884
rect 2028 2876 2036 2884
rect 2764 2876 2772 2884
rect 2796 2876 2804 2884
rect 876 2856 884 2864
rect 2188 2856 2196 2864
rect 2508 2856 2516 2864
rect 3084 2856 3092 2864
rect 3340 2856 3348 2864
rect 5068 2856 5076 2864
rect 2764 2836 2772 2844
rect 3276 2836 3284 2844
rect 1044 2806 1051 2814
rect 1051 2806 1052 2814
rect 1056 2806 1061 2814
rect 1061 2806 1063 2814
rect 1063 2806 1064 2814
rect 1068 2806 1071 2814
rect 1071 2806 1073 2814
rect 1073 2806 1076 2814
rect 1080 2806 1081 2814
rect 1081 2806 1083 2814
rect 1083 2806 1088 2814
rect 1092 2806 1093 2814
rect 1093 2806 1100 2814
rect 4052 2806 4059 2814
rect 4059 2806 4060 2814
rect 4064 2806 4069 2814
rect 4069 2806 4071 2814
rect 4071 2806 4072 2814
rect 4076 2806 4079 2814
rect 4079 2806 4081 2814
rect 4081 2806 4084 2814
rect 4088 2806 4089 2814
rect 4089 2806 4091 2814
rect 4091 2806 4096 2814
rect 4100 2806 4101 2814
rect 4101 2806 4108 2814
rect 1004 2796 1012 2804
rect 1708 2796 1716 2804
rect 1900 2796 1908 2804
rect 1932 2796 1940 2804
rect 1996 2796 2004 2804
rect 1868 2776 1876 2784
rect 2124 2776 2132 2784
rect 2508 2776 2516 2784
rect 1484 2756 1492 2764
rect 1836 2756 1844 2764
rect 2796 2756 2804 2764
rect 4972 2736 4980 2744
rect 1868 2716 1876 2724
rect 2156 2716 2164 2724
rect 2348 2716 2356 2724
rect 2924 2716 2932 2724
rect 3276 2716 3284 2724
rect 4172 2716 4180 2724
rect 4748 2716 4756 2724
rect 1900 2696 1908 2704
rect 2060 2696 2068 2704
rect 2284 2696 2292 2704
rect 2444 2696 2452 2704
rect 3532 2696 3540 2704
rect 3724 2696 3732 2704
rect 1004 2676 1012 2684
rect 1292 2676 1300 2684
rect 2476 2676 2484 2684
rect 4780 2676 4788 2684
rect 1420 2656 1428 2664
rect 1836 2656 1844 2664
rect 2028 2656 2036 2664
rect 2156 2656 2164 2664
rect 2348 2656 2356 2664
rect 3052 2656 3060 2664
rect 2060 2636 2068 2644
rect 2092 2636 2100 2644
rect 2508 2636 2516 2644
rect 2988 2636 2996 2644
rect 3148 2636 3156 2644
rect 3564 2636 3572 2644
rect 1324 2616 1332 2624
rect 1772 2616 1780 2624
rect 2252 2616 2260 2624
rect 4492 2616 4500 2624
rect 2548 2606 2555 2614
rect 2555 2606 2556 2614
rect 2560 2606 2565 2614
rect 2565 2606 2567 2614
rect 2567 2606 2568 2614
rect 2572 2606 2575 2614
rect 2575 2606 2577 2614
rect 2577 2606 2580 2614
rect 2584 2606 2585 2614
rect 2585 2606 2587 2614
rect 2587 2606 2592 2614
rect 2596 2606 2597 2614
rect 2597 2606 2604 2614
rect 620 2596 628 2604
rect 1292 2596 1300 2604
rect 2668 2596 2676 2604
rect 2764 2596 2772 2604
rect 3020 2596 3028 2604
rect 3820 2596 3828 2604
rect 5036 2596 5044 2604
rect 2348 2576 2356 2584
rect 4300 2576 4308 2584
rect 716 2556 724 2564
rect 748 2556 756 2564
rect 1612 2556 1620 2564
rect 3628 2536 3636 2544
rect 4204 2556 4212 2564
rect 4812 2536 4820 2544
rect 5068 2536 5076 2544
rect 972 2516 980 2524
rect 1804 2516 1812 2524
rect 1868 2516 1876 2524
rect 1484 2496 1492 2504
rect 1612 2496 1620 2504
rect 1644 2476 1652 2484
rect 1868 2476 1876 2484
rect 1932 2496 1940 2504
rect 1964 2516 1972 2524
rect 2124 2516 2132 2524
rect 2684 2516 2692 2524
rect 3052 2516 3060 2524
rect 3436 2516 3444 2524
rect 2188 2496 2196 2504
rect 4204 2496 4212 2504
rect 5068 2496 5076 2504
rect 4908 2476 4916 2484
rect 4972 2476 4980 2484
rect 1900 2456 1908 2464
rect 1964 2456 1972 2464
rect 1996 2456 2004 2464
rect 2028 2456 2036 2464
rect 1868 2436 1876 2444
rect 2444 2436 2452 2444
rect 2636 2436 2644 2444
rect 2764 2436 2772 2444
rect 4812 2436 4820 2444
rect 4876 2436 4884 2444
rect 1452 2416 1460 2424
rect 2028 2416 2036 2424
rect 3020 2416 3028 2424
rect 3820 2416 3828 2424
rect 1044 2406 1051 2414
rect 1051 2406 1052 2414
rect 1056 2406 1061 2414
rect 1061 2406 1063 2414
rect 1063 2406 1064 2414
rect 1068 2406 1071 2414
rect 1071 2406 1073 2414
rect 1073 2406 1076 2414
rect 1080 2406 1081 2414
rect 1081 2406 1083 2414
rect 1083 2406 1088 2414
rect 1092 2406 1093 2414
rect 1093 2406 1100 2414
rect 4052 2406 4059 2414
rect 4059 2406 4060 2414
rect 4064 2406 4069 2414
rect 4069 2406 4071 2414
rect 4071 2406 4072 2414
rect 4076 2406 4079 2414
rect 4079 2406 4081 2414
rect 4081 2406 4084 2414
rect 4088 2406 4089 2414
rect 4089 2406 4091 2414
rect 4091 2406 4096 2414
rect 4100 2406 4101 2414
rect 4101 2406 4108 2414
rect 2092 2396 2100 2404
rect 2220 2396 2228 2404
rect 2892 2396 2900 2404
rect 3468 2396 3476 2404
rect 492 2376 500 2384
rect 4140 2376 4148 2384
rect 2156 2356 2164 2364
rect 2508 2356 2516 2364
rect 2764 2336 2772 2344
rect 4140 2336 4148 2344
rect 1356 2296 1364 2304
rect 1484 2296 1492 2304
rect 1772 2296 1780 2304
rect 1964 2296 1972 2304
rect 2124 2296 2132 2304
rect 2636 2296 2644 2304
rect 2668 2316 2676 2324
rect 2828 2316 2836 2324
rect 940 2276 948 2284
rect 1708 2276 1716 2284
rect 1900 2276 1908 2284
rect 3916 2296 3924 2304
rect 4748 2296 4756 2304
rect 748 2256 756 2264
rect 1420 2256 1428 2264
rect 2668 2276 2676 2284
rect 2764 2276 2772 2284
rect 2828 2276 2836 2284
rect 2348 2256 2356 2264
rect 2444 2256 2452 2264
rect 620 2236 628 2244
rect 1772 2236 1780 2244
rect 2252 2236 2260 2244
rect 2508 2236 2516 2244
rect 2860 2236 2868 2244
rect 844 2216 852 2224
rect 1548 2216 1556 2224
rect 2892 2216 2900 2224
rect 2548 2206 2555 2214
rect 2555 2206 2556 2214
rect 2560 2206 2565 2214
rect 2565 2206 2567 2214
rect 2567 2206 2568 2214
rect 2572 2206 2575 2214
rect 2575 2206 2577 2214
rect 2577 2206 2580 2214
rect 2584 2206 2585 2214
rect 2585 2206 2587 2214
rect 2587 2206 2592 2214
rect 2596 2206 2597 2214
rect 2597 2206 2604 2214
rect 1516 2196 1524 2204
rect 1868 2196 1876 2204
rect 2188 2196 2196 2204
rect 1644 2176 1652 2184
rect 2092 2176 2100 2184
rect 2316 2196 2324 2204
rect 2636 2196 2644 2204
rect 2956 2196 2964 2204
rect 3052 2196 3060 2204
rect 3084 2196 3092 2204
rect 3340 2196 3348 2204
rect 2252 2176 2260 2184
rect 812 2156 820 2164
rect 1196 2156 1204 2164
rect 1836 2156 1844 2164
rect 1932 2156 1940 2164
rect 2028 2156 2036 2164
rect 2060 2156 2068 2164
rect 2284 2156 2292 2164
rect 620 2136 628 2144
rect 2220 2136 2228 2144
rect 2348 2136 2356 2144
rect 2508 2136 2516 2144
rect 940 2116 948 2124
rect 1356 2116 1364 2124
rect 1804 2116 1812 2124
rect 2316 2116 2324 2124
rect 3468 2136 3476 2144
rect 4140 2136 4148 2144
rect 4492 2136 4500 2144
rect 2700 2116 2708 2124
rect 2732 2116 2740 2124
rect 1996 2096 2004 2104
rect 2380 2096 2388 2104
rect 2444 2096 2452 2104
rect 3948 2096 3956 2104
rect 1852 2076 1860 2084
rect 1884 2076 1892 2084
rect 2412 2076 2420 2084
rect 1644 2056 1652 2064
rect 1740 2056 1748 2064
rect 2284 2056 2292 2064
rect 2668 2056 2676 2064
rect 3564 2056 3572 2064
rect 3852 2056 3860 2064
rect 1932 2016 1940 2024
rect 1044 2006 1051 2014
rect 1051 2006 1052 2014
rect 1056 2006 1061 2014
rect 1061 2006 1063 2014
rect 1063 2006 1064 2014
rect 1068 2006 1071 2014
rect 1071 2006 1073 2014
rect 1073 2006 1076 2014
rect 1080 2006 1081 2014
rect 1081 2006 1083 2014
rect 1083 2006 1088 2014
rect 1092 2006 1093 2014
rect 1093 2006 1100 2014
rect 3084 2016 3092 2024
rect 4052 2006 4059 2014
rect 4059 2006 4060 2014
rect 4064 2006 4069 2014
rect 4069 2006 4071 2014
rect 4071 2006 4072 2014
rect 4076 2006 4079 2014
rect 4079 2006 4081 2014
rect 4081 2006 4084 2014
rect 4088 2006 4089 2014
rect 4089 2006 4091 2014
rect 4091 2006 4096 2014
rect 4100 2006 4101 2014
rect 4101 2006 4108 2014
rect 1964 1996 1972 2004
rect 2060 1996 2068 2004
rect 2220 1996 2228 2004
rect 2444 1996 2452 2004
rect 2828 1996 2836 2004
rect 1132 1976 1140 1984
rect 2124 1976 2132 1984
rect 1996 1956 2004 1964
rect 2252 1976 2260 1984
rect 2700 1976 2708 1984
rect 2764 1956 2772 1964
rect 5100 1956 5108 1964
rect 3308 1936 3316 1944
rect 3436 1936 3444 1944
rect 3852 1936 3860 1944
rect 5068 1936 5076 1944
rect 364 1916 372 1924
rect 2412 1916 2420 1924
rect 2092 1896 2100 1904
rect 1836 1876 1844 1884
rect 1996 1876 2004 1884
rect 2956 1876 2964 1884
rect 2988 1876 2996 1884
rect 4940 1896 4948 1904
rect 1452 1856 1460 1864
rect 1964 1856 1972 1864
rect 2220 1856 2228 1864
rect 2412 1856 2420 1864
rect 2796 1856 2804 1864
rect 3436 1856 3444 1864
rect 5068 1876 5076 1884
rect 5132 1876 5140 1884
rect 1804 1836 1812 1844
rect 2156 1836 2164 1844
rect 1132 1816 1140 1824
rect 1708 1816 1716 1824
rect 3820 1836 3828 1844
rect 4524 1836 4532 1844
rect 1996 1796 2004 1804
rect 2956 1816 2964 1824
rect 5132 1816 5140 1824
rect 2548 1806 2555 1814
rect 2555 1806 2556 1814
rect 2560 1806 2565 1814
rect 2565 1806 2567 1814
rect 2567 1806 2568 1814
rect 2572 1806 2575 1814
rect 2575 1806 2577 1814
rect 2577 1806 2580 1814
rect 2584 1806 2585 1814
rect 2585 1806 2587 1814
rect 2587 1806 2592 1814
rect 2596 1806 2597 1814
rect 2597 1806 2604 1814
rect 2860 1796 2868 1804
rect 4140 1796 4148 1804
rect 4236 1776 4244 1784
rect 2156 1756 2164 1764
rect 2764 1756 2772 1764
rect 4940 1756 4948 1764
rect 4780 1736 4788 1744
rect 1548 1716 1556 1724
rect 1932 1716 1940 1724
rect 2348 1716 2356 1724
rect 2476 1716 2484 1724
rect 3276 1716 3284 1724
rect 492 1696 500 1704
rect 556 1696 564 1704
rect 2284 1696 2292 1704
rect 5068 1696 5076 1704
rect 1580 1676 1588 1684
rect 2060 1676 2068 1684
rect 3564 1676 3572 1684
rect 812 1656 820 1664
rect 2380 1656 2388 1664
rect 2860 1656 2868 1664
rect 1324 1636 1332 1644
rect 1516 1636 1524 1644
rect 2188 1636 2196 1644
rect 1044 1606 1051 1614
rect 1051 1606 1052 1614
rect 1056 1606 1061 1614
rect 1061 1606 1063 1614
rect 1063 1606 1064 1614
rect 1068 1606 1071 1614
rect 1071 1606 1073 1614
rect 1073 1606 1076 1614
rect 1080 1606 1081 1614
rect 1081 1606 1083 1614
rect 1083 1606 1088 1614
rect 1092 1606 1093 1614
rect 1093 1606 1100 1614
rect 1740 1596 1748 1604
rect 2028 1596 2036 1604
rect 2220 1596 2228 1604
rect 2444 1596 2452 1604
rect 2636 1616 2644 1624
rect 2988 1616 2996 1624
rect 4524 1656 4532 1664
rect 3948 1636 3956 1644
rect 3180 1616 3188 1624
rect 4052 1606 4059 1614
rect 4059 1606 4060 1614
rect 4064 1606 4069 1614
rect 4069 1606 4071 1614
rect 4071 1606 4072 1614
rect 4076 1606 4079 1614
rect 4079 1606 4081 1614
rect 4081 1606 4084 1614
rect 4088 1606 4089 1614
rect 4089 1606 4091 1614
rect 4091 1606 4096 1614
rect 4100 1606 4101 1614
rect 4101 1606 4108 1614
rect 1740 1556 1748 1564
rect 2060 1556 2068 1564
rect 2284 1556 2292 1564
rect 2380 1556 2388 1564
rect 3468 1576 3476 1584
rect 3372 1556 3380 1564
rect 2092 1516 2100 1524
rect 2668 1516 2676 1524
rect 1644 1496 1652 1504
rect 1708 1496 1716 1504
rect 1996 1496 2004 1504
rect 2156 1496 2164 1504
rect 2476 1496 2484 1504
rect 3116 1516 3124 1524
rect 2796 1496 2804 1504
rect 2956 1496 2964 1504
rect 940 1476 948 1484
rect 1612 1476 1620 1484
rect 2092 1476 2100 1484
rect 2764 1476 2772 1484
rect 3628 1476 3636 1484
rect 1164 1456 1172 1464
rect 1804 1456 1812 1464
rect 2156 1456 2164 1464
rect 2348 1456 2356 1464
rect 876 1436 884 1444
rect 2028 1436 2036 1444
rect 3180 1436 3188 1444
rect 3852 1436 3860 1444
rect 1740 1416 1748 1424
rect 2668 1416 2676 1424
rect 4140 1416 4148 1424
rect 2548 1406 2555 1414
rect 2555 1406 2556 1414
rect 2560 1406 2565 1414
rect 2565 1406 2567 1414
rect 2567 1406 2568 1414
rect 2572 1406 2575 1414
rect 2575 1406 2577 1414
rect 2577 1406 2580 1414
rect 2584 1406 2585 1414
rect 2585 1406 2587 1414
rect 2587 1406 2592 1414
rect 2596 1406 2597 1414
rect 2597 1406 2604 1414
rect 12 1396 20 1404
rect 876 1396 884 1404
rect 2284 1396 2292 1404
rect 3020 1396 3028 1404
rect 3116 1396 3124 1404
rect 1548 1376 1556 1384
rect 1772 1376 1780 1384
rect 748 1356 756 1364
rect 1452 1356 1460 1364
rect 2412 1376 2420 1384
rect 3084 1376 3092 1384
rect 2924 1356 2932 1364
rect 2956 1356 2964 1364
rect 5068 1356 5076 1364
rect 1548 1316 1556 1324
rect 1644 1316 1652 1324
rect 2252 1336 2260 1344
rect 2636 1336 2644 1344
rect 3084 1336 3092 1344
rect 3980 1336 3988 1344
rect 5036 1336 5044 1344
rect 2156 1316 2164 1324
rect 3308 1316 3316 1324
rect 2444 1296 2452 1304
rect 3020 1296 3028 1304
rect 1420 1276 1428 1284
rect 2380 1276 2388 1284
rect 3596 1296 3604 1304
rect 5100 1316 5108 1324
rect 4300 1296 4308 1304
rect 364 1256 372 1264
rect 1196 1236 1204 1244
rect 2444 1236 2452 1244
rect 3180 1256 3188 1264
rect 3500 1256 3508 1264
rect 3372 1236 3380 1244
rect 4876 1236 4884 1244
rect 5100 1236 5108 1244
rect 2220 1216 2228 1224
rect 2828 1216 2836 1224
rect 2860 1216 2868 1224
rect 3500 1216 3508 1224
rect 4908 1216 4916 1224
rect 1044 1206 1051 1214
rect 1051 1206 1052 1214
rect 1056 1206 1061 1214
rect 1061 1206 1063 1214
rect 1063 1206 1064 1214
rect 1068 1206 1071 1214
rect 1071 1206 1073 1214
rect 1073 1206 1076 1214
rect 1080 1206 1081 1214
rect 1081 1206 1083 1214
rect 1083 1206 1088 1214
rect 1092 1206 1093 1214
rect 1093 1206 1100 1214
rect 4052 1206 4059 1214
rect 4059 1206 4060 1214
rect 4064 1206 4069 1214
rect 4069 1206 4071 1214
rect 4071 1206 4072 1214
rect 4076 1206 4079 1214
rect 4079 1206 4081 1214
rect 4081 1206 4084 1214
rect 4088 1206 4089 1214
rect 4089 1206 4091 1214
rect 4091 1206 4096 1214
rect 4100 1206 4101 1214
rect 4101 1206 4108 1214
rect 2956 1196 2964 1204
rect 3212 1196 3220 1204
rect 2444 1176 2452 1184
rect 1420 1156 1428 1164
rect 2156 1136 2164 1144
rect 2252 1136 2260 1144
rect 1356 1116 1364 1124
rect 1548 1116 1556 1124
rect 1580 1116 1588 1124
rect 1452 1096 1460 1104
rect 2764 1136 2772 1144
rect 4652 1136 4660 1144
rect 2348 1116 2356 1124
rect 2892 1116 2900 1124
rect 4940 1116 4948 1124
rect 1964 1076 1972 1084
rect 3276 1096 3284 1104
rect 3436 1096 3444 1104
rect 2188 1076 2196 1084
rect 2988 1076 2996 1084
rect 3468 1076 3476 1084
rect 1548 1056 1556 1064
rect 1836 1056 1844 1064
rect 2636 1056 2644 1064
rect 4556 1056 4564 1064
rect 524 1036 532 1044
rect 1356 1036 1364 1044
rect 2060 1036 2068 1044
rect 748 1016 756 1024
rect 2124 1036 2132 1044
rect 2476 1016 2484 1024
rect 2988 1036 2996 1044
rect 2548 1006 2555 1014
rect 2555 1006 2556 1014
rect 2560 1006 2565 1014
rect 2565 1006 2567 1014
rect 2567 1006 2568 1014
rect 2572 1006 2575 1014
rect 2575 1006 2577 1014
rect 2577 1006 2580 1014
rect 2584 1006 2585 1014
rect 2585 1006 2587 1014
rect 2587 1006 2592 1014
rect 2596 1006 2597 1014
rect 2597 1006 2604 1014
rect 684 996 692 1004
rect 2828 996 2836 1004
rect 2860 996 2868 1004
rect 3532 996 3540 1004
rect 4620 996 4628 1004
rect 972 976 980 984
rect 1196 936 1204 944
rect 1324 956 1332 964
rect 2412 976 2420 984
rect 1452 936 1460 944
rect 3180 956 3188 964
rect 2764 936 2772 944
rect 2924 936 2932 944
rect 2956 936 2964 944
rect 3596 936 3604 944
rect 684 916 692 924
rect 1164 916 1172 924
rect 1228 916 1236 924
rect 1612 916 1620 924
rect 1740 916 1748 924
rect 1932 896 1940 904
rect 2028 916 2036 924
rect 2476 916 2484 924
rect 2636 916 2644 924
rect 3820 916 3828 924
rect 812 876 820 884
rect 1612 876 1620 884
rect 1004 856 1012 864
rect 2156 876 2164 884
rect 2828 856 2836 864
rect 3884 856 3892 864
rect 1740 836 1748 844
rect 1772 836 1780 844
rect 3820 836 3828 844
rect 972 816 980 824
rect 2476 816 2484 824
rect 3084 816 3092 824
rect 1044 806 1051 814
rect 1051 806 1052 814
rect 1056 806 1061 814
rect 1061 806 1063 814
rect 1063 806 1064 814
rect 1068 806 1071 814
rect 1071 806 1073 814
rect 1073 806 1076 814
rect 1080 806 1081 814
rect 1081 806 1083 814
rect 1083 806 1088 814
rect 1092 806 1093 814
rect 1093 806 1100 814
rect 4052 806 4059 814
rect 4059 806 4060 814
rect 4064 806 4069 814
rect 4069 806 4071 814
rect 4071 806 4072 814
rect 4076 806 4079 814
rect 4079 806 4081 814
rect 4081 806 4084 814
rect 4088 806 4089 814
rect 4089 806 4091 814
rect 4091 806 4096 814
rect 4100 806 4101 814
rect 4101 806 4108 814
rect 2060 796 2068 804
rect 1196 776 1204 784
rect 2348 776 2356 784
rect 2668 796 2676 804
rect 2764 796 2772 804
rect 4652 796 4660 804
rect 2380 756 2388 764
rect 2636 756 2644 764
rect 2924 756 2932 764
rect 3244 756 3252 764
rect 1228 736 1236 744
rect 5068 756 5076 764
rect 1292 716 1300 724
rect 12 696 20 704
rect 1452 696 1460 704
rect 556 676 564 684
rect 1004 676 1012 684
rect 1484 676 1492 684
rect 2092 696 2100 704
rect 2124 696 2132 704
rect 2380 696 2388 704
rect 2444 696 2452 704
rect 2636 716 2644 724
rect 2924 716 2932 724
rect 4556 716 4564 724
rect 1548 676 1556 684
rect 1676 676 1684 684
rect 2156 676 2164 684
rect 2188 676 2196 684
rect 2700 676 2708 684
rect 3948 696 3956 704
rect 4300 696 4308 704
rect 3212 676 3220 684
rect 3980 676 3988 684
rect 4236 676 4244 684
rect 940 656 948 664
rect 1548 636 1556 644
rect 1580 636 1588 644
rect 1772 636 1780 644
rect 2956 656 2964 664
rect 2092 616 2100 624
rect 2348 616 2356 624
rect 2892 616 2900 624
rect 4620 616 4628 624
rect 2548 606 2555 614
rect 2555 606 2556 614
rect 2560 606 2565 614
rect 2565 606 2567 614
rect 2567 606 2568 614
rect 2572 606 2575 614
rect 2575 606 2577 614
rect 2577 606 2580 614
rect 2584 606 2585 614
rect 2585 606 2587 614
rect 2587 606 2592 614
rect 2596 606 2597 614
rect 2597 606 2604 614
rect 1676 596 1684 604
rect 1196 576 1204 584
rect 2412 576 2420 584
rect 2476 576 2484 584
rect 1740 556 1748 564
rect 1932 556 1940 564
rect 1964 556 1972 564
rect 524 536 532 544
rect 2732 576 2740 584
rect 3340 576 3348 584
rect 2636 556 2644 564
rect 2956 556 2964 564
rect 3148 556 3156 564
rect 3436 556 3444 564
rect 2252 536 2260 544
rect 2828 536 2836 544
rect 3372 536 3380 544
rect 4940 536 4948 544
rect 2764 516 2772 524
rect 3180 516 3188 524
rect 3884 516 3892 524
rect 4876 516 4884 524
rect 1740 476 1748 484
rect 2188 476 2196 484
rect 2764 476 2772 484
rect 3308 496 3316 504
rect 3244 476 3252 484
rect 2700 456 2708 464
rect 2668 436 2676 444
rect 2988 436 2996 444
rect 1044 406 1051 414
rect 1051 406 1052 414
rect 1056 406 1061 414
rect 1061 406 1063 414
rect 1063 406 1064 414
rect 1068 406 1071 414
rect 1071 406 1073 414
rect 1073 406 1076 414
rect 1080 406 1081 414
rect 1081 406 1083 414
rect 1083 406 1088 414
rect 1092 406 1093 414
rect 1093 406 1100 414
rect 4052 406 4059 414
rect 4059 406 4060 414
rect 4064 406 4069 414
rect 4069 406 4071 414
rect 4071 406 4072 414
rect 4076 406 4079 414
rect 4079 406 4081 414
rect 4081 406 4084 414
rect 4088 406 4089 414
rect 4089 406 4091 414
rect 4091 406 4096 414
rect 4100 406 4101 414
rect 4101 406 4108 414
rect 3148 396 3156 404
rect 1484 376 1492 384
rect 2764 316 2772 324
rect 2892 316 2900 324
rect 1292 296 1300 304
rect 1804 296 1812 304
rect 2732 296 2740 304
rect 3084 316 3092 324
rect 3116 316 3124 324
rect 3180 276 3188 284
rect 3340 276 3348 284
rect 3372 256 3380 264
rect 3404 276 3412 284
rect 2860 216 2868 224
rect 3404 236 3412 244
rect 3116 216 3124 224
rect 3148 216 3156 224
rect 3340 216 3348 224
rect 2548 206 2555 214
rect 2555 206 2556 214
rect 2560 206 2565 214
rect 2565 206 2567 214
rect 2567 206 2568 214
rect 2572 206 2575 214
rect 2575 206 2577 214
rect 2577 206 2580 214
rect 2584 206 2585 214
rect 2585 206 2587 214
rect 2587 206 2592 214
rect 2596 206 2597 214
rect 2597 206 2604 214
rect 2092 196 2100 204
rect 2828 156 2836 164
rect 1580 136 1588 144
rect 2380 136 2388 144
rect 1804 116 1812 124
rect 3532 156 3540 164
rect 3180 136 3188 144
rect 3308 136 3316 144
rect 3436 136 3444 144
rect 2988 116 2996 124
rect 3244 116 3252 124
rect 2892 96 2900 104
rect 3372 96 3380 104
rect 3148 76 3156 84
rect 2156 56 2164 64
rect 3212 56 3220 64
rect 1044 6 1051 14
rect 1051 6 1052 14
rect 1056 6 1061 14
rect 1061 6 1063 14
rect 1063 6 1064 14
rect 1068 6 1071 14
rect 1071 6 1073 14
rect 1073 6 1076 14
rect 1080 6 1081 14
rect 1081 6 1083 14
rect 1083 6 1088 14
rect 1092 6 1093 14
rect 1093 6 1100 14
rect 4052 6 4059 14
rect 4059 6 4060 14
rect 4064 6 4069 14
rect 4069 6 4071 14
rect 4071 6 4072 14
rect 4076 6 4079 14
rect 4079 6 4081 14
rect 4081 6 4084 14
rect 4088 6 4089 14
rect 4089 6 4091 14
rect 4091 6 4096 14
rect 4100 6 4101 14
rect 4101 6 4108 14
<< metal4 >>
rect 3850 3424 3862 3426
rect 3850 3416 3852 3424
rect 3860 3416 3862 3424
rect 1040 3214 1104 3416
rect 2544 3414 2608 3416
rect 2544 3406 2548 3414
rect 2556 3406 2560 3414
rect 2568 3406 2572 3414
rect 2580 3406 2584 3414
rect 2592 3406 2596 3414
rect 2604 3406 2608 3414
rect 1514 3384 1526 3386
rect 1514 3376 1516 3384
rect 1524 3376 1526 3384
rect 1040 3206 1044 3214
rect 1052 3206 1056 3214
rect 1064 3206 1068 3214
rect 1076 3206 1080 3214
rect 1088 3206 1092 3214
rect 1100 3206 1104 3214
rect 714 3184 726 3186
rect 714 3176 716 3184
rect 724 3176 726 3184
rect 618 2964 630 2966
rect 618 2956 620 2964
rect 628 2956 630 2964
rect 618 2604 630 2956
rect 618 2596 620 2604
rect 628 2596 630 2604
rect 618 2594 630 2596
rect 714 2564 726 3176
rect 810 3104 822 3106
rect 810 3096 812 3104
rect 820 3096 822 3104
rect 714 2556 716 2564
rect 724 2556 726 2564
rect 714 2554 726 2556
rect 746 2564 758 2566
rect 746 2556 748 2564
rect 756 2556 758 2564
rect 490 2384 502 2386
rect 490 2376 492 2384
rect 500 2376 502 2384
rect 362 1924 374 1926
rect 362 1916 364 1924
rect 372 1916 374 1924
rect 10 1404 22 1406
rect 10 1396 12 1404
rect 20 1396 22 1404
rect 10 704 22 1396
rect 362 1264 374 1916
rect 490 1704 502 2376
rect 746 2264 758 2556
rect 746 2256 748 2264
rect 756 2256 758 2264
rect 746 2254 758 2256
rect 618 2244 630 2246
rect 618 2236 620 2244
rect 628 2236 630 2244
rect 618 2144 630 2236
rect 810 2164 822 3096
rect 874 2944 886 2946
rect 874 2936 876 2944
rect 884 2936 886 2944
rect 842 2924 854 2926
rect 842 2916 844 2924
rect 852 2916 854 2924
rect 842 2224 854 2916
rect 874 2864 886 2936
rect 874 2856 876 2864
rect 884 2856 886 2864
rect 874 2854 886 2856
rect 970 2884 982 2886
rect 970 2876 972 2884
rect 980 2876 982 2884
rect 970 2524 982 2876
rect 1040 2814 1104 3206
rect 1290 3324 1302 3326
rect 1290 3316 1292 3324
rect 1300 3316 1302 3324
rect 1162 3124 1174 3126
rect 1162 3116 1164 3124
rect 1172 3116 1174 3124
rect 1162 3084 1174 3116
rect 1162 3076 1164 3084
rect 1172 3076 1174 3084
rect 1162 3074 1174 3076
rect 1194 3104 1206 3106
rect 1194 3096 1196 3104
rect 1204 3096 1206 3104
rect 1040 2806 1044 2814
rect 1052 2806 1056 2814
rect 1064 2806 1068 2814
rect 1076 2806 1080 2814
rect 1088 2806 1092 2814
rect 1100 2806 1104 2814
rect 1002 2804 1014 2806
rect 1002 2796 1004 2804
rect 1012 2796 1014 2804
rect 1002 2684 1014 2796
rect 1002 2676 1004 2684
rect 1012 2676 1014 2684
rect 1002 2674 1014 2676
rect 970 2516 972 2524
rect 980 2516 982 2524
rect 970 2514 982 2516
rect 1040 2414 1104 2806
rect 1040 2406 1044 2414
rect 1052 2406 1056 2414
rect 1064 2406 1068 2414
rect 1076 2406 1080 2414
rect 1088 2406 1092 2414
rect 1100 2406 1104 2414
rect 842 2216 844 2224
rect 852 2216 854 2224
rect 842 2214 854 2216
rect 938 2284 950 2286
rect 938 2276 940 2284
rect 948 2276 950 2284
rect 810 2156 812 2164
rect 820 2156 822 2164
rect 810 2154 822 2156
rect 618 2136 620 2144
rect 628 2136 630 2144
rect 618 2134 630 2136
rect 938 2124 950 2276
rect 938 2116 940 2124
rect 948 2116 950 2124
rect 938 2114 950 2116
rect 1040 2014 1104 2406
rect 1194 2164 1206 3096
rect 1290 2884 1302 3316
rect 1386 3124 1398 3126
rect 1386 3116 1388 3124
rect 1396 3116 1398 3124
rect 1386 3044 1398 3116
rect 1386 3036 1388 3044
rect 1396 3036 1398 3044
rect 1386 3034 1398 3036
rect 1482 3124 1494 3126
rect 1482 3116 1484 3124
rect 1492 3116 1494 3124
rect 1290 2876 1292 2884
rect 1300 2876 1302 2884
rect 1290 2874 1302 2876
rect 1322 2924 1334 2926
rect 1322 2916 1324 2924
rect 1332 2916 1334 2924
rect 1290 2684 1302 2686
rect 1290 2676 1292 2684
rect 1300 2676 1302 2684
rect 1290 2604 1302 2676
rect 1322 2624 1334 2916
rect 1482 2764 1494 3116
rect 1514 2924 1526 3376
rect 1642 3364 1654 3366
rect 1642 3356 1644 3364
rect 1652 3356 1654 3364
rect 1514 2916 1516 2924
rect 1524 2916 1526 2924
rect 1514 2914 1526 2916
rect 1610 3104 1622 3106
rect 1610 3096 1612 3104
rect 1620 3096 1622 3104
rect 1482 2756 1484 2764
rect 1492 2756 1494 2764
rect 1482 2754 1494 2756
rect 1322 2616 1324 2624
rect 1332 2616 1334 2624
rect 1322 2614 1334 2616
rect 1418 2664 1430 2666
rect 1418 2656 1420 2664
rect 1428 2656 1430 2664
rect 1290 2596 1292 2604
rect 1300 2596 1302 2604
rect 1290 2594 1302 2596
rect 1194 2156 1196 2164
rect 1204 2156 1206 2164
rect 1194 2154 1206 2156
rect 1354 2304 1366 2306
rect 1354 2296 1356 2304
rect 1364 2296 1366 2304
rect 1354 2124 1366 2296
rect 1418 2264 1430 2656
rect 1610 2564 1622 3096
rect 1642 2944 1654 3356
rect 2250 3364 2262 3366
rect 2250 3356 2252 3364
rect 2260 3356 2262 3364
rect 2186 3344 2198 3346
rect 2186 3336 2188 3344
rect 2196 3336 2198 3344
rect 2186 3326 2198 3336
rect 1898 3324 1910 3326
rect 1898 3316 1900 3324
rect 1908 3316 1910 3324
rect 1642 2936 1644 2944
rect 1652 2936 1654 2944
rect 1642 2934 1654 2936
rect 1706 2984 1718 2986
rect 1706 2976 1708 2984
rect 1716 2976 1718 2984
rect 1610 2556 1612 2564
rect 1620 2556 1622 2564
rect 1610 2554 1622 2556
rect 1642 2904 1654 2906
rect 1642 2896 1644 2904
rect 1652 2896 1654 2904
rect 1482 2504 1494 2506
rect 1482 2496 1484 2504
rect 1492 2496 1494 2504
rect 1418 2256 1420 2264
rect 1428 2256 1430 2264
rect 1418 2254 1430 2256
rect 1450 2424 1462 2426
rect 1450 2416 1452 2424
rect 1460 2416 1462 2424
rect 1354 2116 1356 2124
rect 1364 2116 1366 2124
rect 1354 2114 1366 2116
rect 1040 2006 1044 2014
rect 1052 2006 1056 2014
rect 1064 2006 1068 2014
rect 1076 2006 1080 2014
rect 1088 2006 1092 2014
rect 1100 2006 1104 2014
rect 490 1696 492 1704
rect 500 1696 502 1704
rect 490 1694 502 1696
rect 554 1704 566 1706
rect 554 1696 556 1704
rect 564 1696 566 1704
rect 362 1256 364 1264
rect 372 1256 374 1264
rect 362 1254 374 1256
rect 10 696 12 704
rect 20 696 22 704
rect 10 694 22 696
rect 522 1044 534 1046
rect 522 1036 524 1044
rect 532 1036 534 1044
rect 522 544 534 1036
rect 554 684 566 1696
rect 810 1664 822 1666
rect 810 1656 812 1664
rect 820 1656 822 1664
rect 746 1364 758 1366
rect 746 1356 748 1364
rect 756 1356 758 1364
rect 746 1024 758 1356
rect 746 1016 748 1024
rect 756 1016 758 1024
rect 746 1014 758 1016
rect 682 1004 694 1006
rect 682 996 684 1004
rect 692 996 694 1004
rect 682 924 694 996
rect 682 916 684 924
rect 692 916 694 924
rect 682 914 694 916
rect 810 884 822 1656
rect 1040 1614 1104 2006
rect 1130 1984 1142 1986
rect 1130 1976 1132 1984
rect 1140 1976 1142 1984
rect 1130 1824 1142 1976
rect 1450 1864 1462 2416
rect 1482 2304 1494 2496
rect 1482 2296 1484 2304
rect 1492 2296 1494 2304
rect 1482 2294 1494 2296
rect 1610 2504 1622 2506
rect 1610 2496 1612 2504
rect 1620 2496 1622 2504
rect 1546 2224 1558 2226
rect 1546 2216 1548 2224
rect 1556 2216 1558 2224
rect 1450 1856 1452 1864
rect 1460 1856 1462 1864
rect 1450 1854 1462 1856
rect 1514 2204 1526 2206
rect 1514 2196 1516 2204
rect 1524 2196 1526 2204
rect 1130 1816 1132 1824
rect 1140 1816 1142 1824
rect 1130 1814 1142 1816
rect 1040 1606 1044 1614
rect 1052 1606 1056 1614
rect 1064 1606 1068 1614
rect 1076 1606 1080 1614
rect 1088 1606 1092 1614
rect 1100 1606 1104 1614
rect 938 1484 950 1486
rect 938 1476 940 1484
rect 948 1476 950 1484
rect 874 1444 886 1446
rect 874 1436 876 1444
rect 884 1436 886 1444
rect 874 1404 886 1436
rect 874 1396 876 1404
rect 884 1396 886 1404
rect 874 1394 886 1396
rect 810 876 812 884
rect 820 876 822 884
rect 810 874 822 876
rect 554 676 556 684
rect 564 676 566 684
rect 554 674 566 676
rect 938 664 950 1476
rect 1040 1214 1104 1606
rect 1322 1644 1334 1646
rect 1322 1636 1324 1644
rect 1332 1636 1334 1644
rect 1040 1206 1044 1214
rect 1052 1206 1056 1214
rect 1064 1206 1068 1214
rect 1076 1206 1080 1214
rect 1088 1206 1092 1214
rect 1100 1206 1104 1214
rect 970 984 982 986
rect 970 976 972 984
rect 980 976 982 984
rect 970 824 982 976
rect 970 816 972 824
rect 980 816 982 824
rect 970 814 982 816
rect 1002 864 1014 866
rect 1002 856 1004 864
rect 1012 856 1014 864
rect 1002 684 1014 856
rect 1002 676 1004 684
rect 1012 676 1014 684
rect 1002 674 1014 676
rect 1040 814 1104 1206
rect 1162 1464 1174 1466
rect 1162 1456 1164 1464
rect 1172 1456 1174 1464
rect 1162 924 1174 1456
rect 1194 1244 1206 1246
rect 1194 1236 1196 1244
rect 1204 1236 1206 1244
rect 1194 944 1206 1236
rect 1322 964 1334 1636
rect 1514 1644 1526 2196
rect 1546 1724 1558 2216
rect 1546 1716 1548 1724
rect 1556 1716 1558 1724
rect 1546 1714 1558 1716
rect 1514 1636 1516 1644
rect 1524 1636 1526 1644
rect 1514 1634 1526 1636
rect 1578 1684 1590 1686
rect 1578 1676 1580 1684
rect 1588 1676 1590 1684
rect 1546 1384 1558 1386
rect 1546 1376 1548 1384
rect 1556 1376 1558 1384
rect 1450 1364 1462 1366
rect 1450 1356 1452 1364
rect 1460 1356 1462 1364
rect 1418 1284 1430 1286
rect 1418 1276 1420 1284
rect 1428 1276 1430 1284
rect 1418 1164 1430 1276
rect 1418 1156 1420 1164
rect 1428 1156 1430 1164
rect 1418 1154 1430 1156
rect 1354 1124 1366 1126
rect 1354 1116 1356 1124
rect 1364 1116 1366 1124
rect 1354 1044 1366 1116
rect 1354 1036 1356 1044
rect 1364 1036 1366 1044
rect 1354 1034 1366 1036
rect 1450 1104 1462 1356
rect 1546 1324 1558 1376
rect 1546 1316 1548 1324
rect 1556 1316 1558 1324
rect 1546 1314 1558 1316
rect 1450 1096 1452 1104
rect 1460 1096 1462 1104
rect 1322 956 1324 964
rect 1332 956 1334 964
rect 1322 954 1334 956
rect 1194 936 1196 944
rect 1204 936 1206 944
rect 1194 934 1206 936
rect 1450 944 1462 1096
rect 1546 1124 1558 1126
rect 1546 1116 1548 1124
rect 1556 1116 1558 1124
rect 1546 1064 1558 1116
rect 1578 1124 1590 1676
rect 1610 1484 1622 2496
rect 1642 2484 1654 2896
rect 1706 2904 1718 2976
rect 1706 2896 1708 2904
rect 1716 2896 1718 2904
rect 1706 2894 1718 2896
rect 1866 2944 1878 2946
rect 1866 2936 1868 2944
rect 1876 2936 1878 2944
rect 1642 2476 1644 2484
rect 1652 2476 1654 2484
rect 1642 2474 1654 2476
rect 1706 2804 1718 2806
rect 1706 2796 1708 2804
rect 1716 2796 1718 2804
rect 1706 2284 1718 2796
rect 1866 2784 1878 2936
rect 1866 2776 1868 2784
rect 1876 2776 1878 2784
rect 1866 2774 1878 2776
rect 1898 2804 1910 3316
rect 2154 3314 2198 3326
rect 2154 3286 2166 3314
rect 2122 3284 2166 3286
rect 2122 3276 2124 3284
rect 2132 3276 2166 3284
rect 2122 3274 2166 3276
rect 2154 3204 2166 3206
rect 2154 3196 2156 3204
rect 2164 3196 2166 3204
rect 1994 3104 2006 3106
rect 1994 3096 1996 3104
rect 2004 3096 2006 3104
rect 1898 2796 1900 2804
rect 1908 2796 1910 2804
rect 1834 2764 1846 2766
rect 1834 2756 1836 2764
rect 1844 2756 1846 2764
rect 1834 2664 1846 2756
rect 1834 2656 1836 2664
rect 1844 2656 1846 2664
rect 1834 2654 1846 2656
rect 1866 2724 1878 2726
rect 1866 2716 1868 2724
rect 1876 2716 1878 2724
rect 1770 2624 1782 2626
rect 1770 2616 1772 2624
rect 1780 2616 1782 2624
rect 1770 2304 1782 2616
rect 1770 2296 1772 2304
rect 1780 2296 1782 2304
rect 1770 2294 1782 2296
rect 1802 2524 1814 2526
rect 1802 2516 1804 2524
rect 1812 2516 1814 2524
rect 1706 2276 1708 2284
rect 1716 2276 1718 2284
rect 1706 2274 1718 2276
rect 1770 2244 1782 2246
rect 1770 2236 1772 2244
rect 1780 2236 1782 2244
rect 1642 2184 1654 2186
rect 1642 2176 1644 2184
rect 1652 2176 1654 2184
rect 1642 2064 1654 2176
rect 1642 2056 1644 2064
rect 1652 2056 1654 2064
rect 1642 2054 1654 2056
rect 1738 2064 1750 2066
rect 1738 2056 1740 2064
rect 1748 2056 1750 2064
rect 1706 1824 1718 1826
rect 1706 1816 1708 1824
rect 1716 1816 1718 1824
rect 1610 1476 1612 1484
rect 1620 1476 1622 1484
rect 1610 1474 1622 1476
rect 1642 1504 1654 1506
rect 1642 1496 1644 1504
rect 1652 1496 1654 1504
rect 1642 1324 1654 1496
rect 1706 1504 1718 1816
rect 1738 1604 1750 2056
rect 1738 1596 1740 1604
rect 1748 1596 1750 1604
rect 1738 1594 1750 1596
rect 1706 1496 1708 1504
rect 1716 1496 1718 1504
rect 1706 1494 1718 1496
rect 1738 1564 1750 1566
rect 1738 1556 1740 1564
rect 1748 1556 1750 1564
rect 1738 1424 1750 1556
rect 1738 1416 1740 1424
rect 1748 1416 1750 1424
rect 1738 1414 1750 1416
rect 1770 1384 1782 2236
rect 1802 2124 1814 2516
rect 1866 2524 1878 2716
rect 1898 2704 1910 2796
rect 1898 2696 1900 2704
rect 1908 2696 1910 2704
rect 1898 2694 1910 2696
rect 1930 2804 1942 2806
rect 1930 2796 1932 2804
rect 1940 2796 1942 2804
rect 1866 2516 1868 2524
rect 1876 2516 1878 2524
rect 1866 2514 1878 2516
rect 1930 2504 1942 2796
rect 1994 2804 2006 3096
rect 2058 3104 2070 3106
rect 2058 3096 2060 3104
rect 2068 3096 2070 3104
rect 2026 3084 2038 3086
rect 2026 3076 2028 3084
rect 2036 3076 2038 3084
rect 2026 2944 2038 3076
rect 2026 2936 2028 2944
rect 2036 2936 2038 2944
rect 2026 2934 2038 2936
rect 1994 2796 1996 2804
rect 2004 2796 2006 2804
rect 1994 2794 2006 2796
rect 2026 2884 2038 2886
rect 2026 2876 2028 2884
rect 2036 2876 2038 2884
rect 2026 2664 2038 2876
rect 2058 2704 2070 3096
rect 2154 2944 2166 3196
rect 2154 2936 2156 2944
rect 2164 2936 2166 2944
rect 2154 2934 2166 2936
rect 2218 2944 2230 2946
rect 2218 2936 2220 2944
rect 2228 2936 2230 2944
rect 2186 2864 2198 2866
rect 2186 2856 2188 2864
rect 2196 2856 2198 2864
rect 2058 2696 2060 2704
rect 2068 2696 2070 2704
rect 2058 2694 2070 2696
rect 2122 2784 2134 2786
rect 2122 2776 2124 2784
rect 2132 2776 2134 2784
rect 2026 2656 2028 2664
rect 2036 2656 2038 2664
rect 2026 2654 2038 2656
rect 2058 2644 2070 2646
rect 2058 2636 2060 2644
rect 2068 2636 2070 2644
rect 1930 2496 1932 2504
rect 1940 2496 1942 2504
rect 1930 2494 1942 2496
rect 1962 2524 1974 2526
rect 1962 2516 1964 2524
rect 1972 2516 1974 2524
rect 1866 2484 1878 2486
rect 1866 2476 1868 2484
rect 1876 2476 1878 2484
rect 1866 2444 1878 2476
rect 1866 2436 1868 2444
rect 1876 2436 1878 2444
rect 1866 2204 1878 2436
rect 1898 2464 1910 2466
rect 1898 2456 1900 2464
rect 1908 2456 1910 2464
rect 1898 2284 1910 2456
rect 1962 2464 1974 2516
rect 1962 2456 1964 2464
rect 1972 2456 1974 2464
rect 1962 2454 1974 2456
rect 1994 2464 2006 2466
rect 1994 2456 1996 2464
rect 2004 2456 2006 2464
rect 1898 2276 1900 2284
rect 1908 2276 1910 2284
rect 1898 2274 1910 2276
rect 1962 2304 1974 2306
rect 1962 2296 1964 2304
rect 1972 2296 1974 2304
rect 1866 2196 1868 2204
rect 1876 2196 1878 2204
rect 1866 2194 1878 2196
rect 1802 2116 1804 2124
rect 1812 2116 1814 2124
rect 1802 2114 1814 2116
rect 1834 2164 1846 2166
rect 1834 2156 1836 2164
rect 1844 2156 1846 2164
rect 1834 2086 1846 2156
rect 1930 2164 1942 2166
rect 1930 2156 1932 2164
rect 1940 2156 1942 2164
rect 1930 2086 1942 2156
rect 1834 2084 1862 2086
rect 1834 2076 1852 2084
rect 1860 2076 1862 2084
rect 1834 2074 1862 2076
rect 1882 2084 1942 2086
rect 1882 2076 1884 2084
rect 1892 2076 1942 2084
rect 1882 2074 1942 2076
rect 1930 2024 1942 2026
rect 1930 2016 1932 2024
rect 1940 2016 1942 2024
rect 1834 1884 1846 1886
rect 1834 1876 1836 1884
rect 1844 1876 1846 1884
rect 1802 1844 1814 1846
rect 1802 1836 1804 1844
rect 1812 1836 1814 1844
rect 1802 1464 1814 1836
rect 1802 1456 1804 1464
rect 1812 1456 1814 1464
rect 1802 1454 1814 1456
rect 1770 1376 1772 1384
rect 1780 1376 1782 1384
rect 1770 1374 1782 1376
rect 1642 1316 1644 1324
rect 1652 1316 1654 1324
rect 1642 1314 1654 1316
rect 1578 1116 1580 1124
rect 1588 1116 1590 1124
rect 1578 1114 1590 1116
rect 1546 1056 1548 1064
rect 1556 1056 1558 1064
rect 1546 1054 1558 1056
rect 1834 1064 1846 1876
rect 1930 1724 1942 2016
rect 1962 2004 1974 2296
rect 1994 2104 2006 2456
rect 2026 2464 2038 2466
rect 2026 2456 2028 2464
rect 2036 2456 2038 2464
rect 2026 2424 2038 2456
rect 2026 2416 2028 2424
rect 2036 2416 2038 2424
rect 2026 2414 2038 2416
rect 2026 2164 2038 2166
rect 2026 2156 2028 2164
rect 2036 2156 2038 2164
rect 2026 2126 2038 2156
rect 2058 2164 2070 2636
rect 2090 2644 2102 2646
rect 2090 2636 2092 2644
rect 2100 2636 2102 2644
rect 2090 2404 2102 2636
rect 2122 2524 2134 2776
rect 2154 2724 2166 2726
rect 2154 2716 2156 2724
rect 2164 2716 2166 2724
rect 2154 2664 2166 2716
rect 2154 2656 2156 2664
rect 2164 2656 2166 2664
rect 2154 2654 2166 2656
rect 2122 2516 2124 2524
rect 2132 2516 2134 2524
rect 2122 2514 2134 2516
rect 2186 2504 2198 2856
rect 2186 2496 2188 2504
rect 2196 2496 2198 2504
rect 2186 2494 2198 2496
rect 2090 2396 2092 2404
rect 2100 2396 2102 2404
rect 2090 2394 2102 2396
rect 2218 2404 2230 2936
rect 2250 2924 2262 3356
rect 2474 3284 2486 3286
rect 2474 3276 2476 3284
rect 2484 3276 2486 3284
rect 2282 3224 2294 3226
rect 2282 3216 2284 3224
rect 2292 3216 2294 3224
rect 2282 3084 2294 3216
rect 2282 3076 2284 3084
rect 2292 3076 2294 3084
rect 2282 3074 2294 3076
rect 2250 2916 2252 2924
rect 2260 2916 2262 2924
rect 2250 2624 2262 2916
rect 2442 2904 2454 2906
rect 2442 2896 2444 2904
rect 2452 2896 2454 2904
rect 2346 2724 2358 2726
rect 2346 2716 2348 2724
rect 2356 2716 2358 2724
rect 2250 2616 2252 2624
rect 2260 2616 2262 2624
rect 2250 2614 2262 2616
rect 2282 2704 2294 2706
rect 2282 2696 2284 2704
rect 2292 2696 2294 2704
rect 2218 2396 2220 2404
rect 2228 2396 2230 2404
rect 2154 2364 2198 2366
rect 2154 2356 2156 2364
rect 2164 2356 2198 2364
rect 2154 2354 2198 2356
rect 2122 2304 2134 2306
rect 2122 2296 2124 2304
rect 2132 2296 2134 2304
rect 2058 2156 2060 2164
rect 2068 2156 2070 2164
rect 2058 2154 2070 2156
rect 2090 2184 2102 2186
rect 2090 2176 2092 2184
rect 2100 2176 2102 2184
rect 2090 2126 2102 2176
rect 2026 2114 2102 2126
rect 1994 2096 1996 2104
rect 2004 2096 2006 2104
rect 1994 2094 2006 2096
rect 1962 1996 1964 2004
rect 1972 1996 1974 2004
rect 1962 1864 1974 1996
rect 2058 2004 2070 2006
rect 2058 1996 2060 2004
rect 2068 1996 2070 2004
rect 1994 1964 2006 1966
rect 1994 1956 1996 1964
rect 2004 1956 2006 1964
rect 1994 1884 2006 1956
rect 1994 1876 1996 1884
rect 2004 1876 2006 1884
rect 1994 1874 2006 1876
rect 1962 1856 1964 1864
rect 1972 1856 1974 1864
rect 1962 1854 1974 1856
rect 1930 1716 1932 1724
rect 1940 1716 1942 1724
rect 1930 1714 1942 1716
rect 1994 1804 2006 1806
rect 1994 1796 1996 1804
rect 2004 1796 2006 1804
rect 1994 1504 2006 1796
rect 2058 1684 2070 1996
rect 2122 1984 2134 2296
rect 2186 2204 2198 2354
rect 2186 2196 2188 2204
rect 2196 2196 2198 2204
rect 2186 2194 2198 2196
rect 2218 2144 2230 2396
rect 2250 2244 2262 2246
rect 2250 2236 2252 2244
rect 2260 2236 2262 2244
rect 2250 2184 2262 2236
rect 2250 2176 2252 2184
rect 2260 2176 2262 2184
rect 2250 2174 2262 2176
rect 2282 2164 2294 2696
rect 2346 2664 2358 2716
rect 2442 2704 2454 2896
rect 2442 2696 2444 2704
rect 2452 2696 2454 2704
rect 2442 2694 2454 2696
rect 2346 2656 2348 2664
rect 2356 2656 2358 2664
rect 2346 2654 2358 2656
rect 2474 2684 2486 3276
rect 2544 3014 2608 3406
rect 2634 3364 2646 3366
rect 2634 3356 2636 3364
rect 2644 3356 2646 3364
rect 2634 3324 2646 3356
rect 2986 3344 2998 3346
rect 2986 3336 2988 3344
rect 2996 3336 2998 3344
rect 2634 3316 2636 3324
rect 2644 3316 2646 3324
rect 2634 3314 2646 3316
rect 2730 3324 2742 3326
rect 2730 3316 2732 3324
rect 2740 3316 2742 3324
rect 2634 3124 2646 3126
rect 2634 3116 2636 3124
rect 2644 3116 2646 3124
rect 2634 3064 2646 3116
rect 2634 3056 2636 3064
rect 2644 3056 2646 3064
rect 2634 3054 2646 3056
rect 2730 3104 2742 3316
rect 2986 3304 2998 3336
rect 2986 3296 2988 3304
rect 2996 3296 2998 3304
rect 2986 3294 2998 3296
rect 2730 3096 2732 3104
rect 2740 3096 2742 3104
rect 2544 3006 2548 3014
rect 2556 3006 2560 3014
rect 2568 3006 2572 3014
rect 2580 3006 2584 3014
rect 2592 3006 2596 3014
rect 2604 3006 2608 3014
rect 2506 2864 2518 2866
rect 2506 2856 2508 2864
rect 2516 2856 2518 2864
rect 2506 2784 2518 2856
rect 2506 2776 2508 2784
rect 2516 2776 2518 2784
rect 2506 2774 2518 2776
rect 2474 2676 2476 2684
rect 2484 2676 2486 2684
rect 2346 2584 2358 2586
rect 2346 2576 2348 2584
rect 2356 2576 2358 2584
rect 2346 2264 2358 2576
rect 2346 2256 2348 2264
rect 2356 2256 2358 2264
rect 2346 2254 2358 2256
rect 2442 2444 2454 2446
rect 2442 2436 2444 2444
rect 2452 2436 2454 2444
rect 2442 2264 2454 2436
rect 2442 2256 2444 2264
rect 2452 2256 2454 2264
rect 2442 2254 2454 2256
rect 2282 2156 2284 2164
rect 2292 2156 2294 2164
rect 2282 2154 2294 2156
rect 2314 2204 2326 2206
rect 2314 2196 2316 2204
rect 2324 2196 2326 2204
rect 2218 2136 2220 2144
rect 2228 2136 2230 2144
rect 2218 2134 2230 2136
rect 2314 2124 2326 2196
rect 2314 2116 2316 2124
rect 2324 2116 2326 2124
rect 2314 2114 2326 2116
rect 2346 2144 2358 2146
rect 2346 2136 2348 2144
rect 2356 2136 2358 2144
rect 2282 2064 2294 2066
rect 2282 2056 2284 2064
rect 2292 2056 2294 2064
rect 2122 1976 2124 1984
rect 2132 1976 2134 1984
rect 2122 1974 2134 1976
rect 2218 2004 2230 2006
rect 2218 1996 2220 2004
rect 2228 1996 2230 2004
rect 2058 1676 2060 1684
rect 2068 1676 2070 1684
rect 2058 1674 2070 1676
rect 2090 1904 2102 1906
rect 2090 1896 2092 1904
rect 2100 1896 2102 1904
rect 1994 1496 1996 1504
rect 2004 1496 2006 1504
rect 1994 1494 2006 1496
rect 2026 1604 2038 1606
rect 2026 1596 2028 1604
rect 2036 1596 2038 1604
rect 2026 1444 2038 1596
rect 2026 1436 2028 1444
rect 2036 1436 2038 1444
rect 2026 1434 2038 1436
rect 2058 1564 2070 1566
rect 2058 1556 2060 1564
rect 2068 1556 2070 1564
rect 2058 1086 2070 1556
rect 2090 1524 2102 1896
rect 2218 1864 2230 1996
rect 2218 1856 2220 1864
rect 2228 1856 2230 1864
rect 2218 1854 2230 1856
rect 2250 1984 2262 1986
rect 2250 1976 2252 1984
rect 2260 1976 2262 1984
rect 2154 1844 2166 1846
rect 2154 1836 2156 1844
rect 2164 1836 2166 1844
rect 2154 1764 2166 1836
rect 2154 1756 2156 1764
rect 2164 1756 2166 1764
rect 2154 1754 2166 1756
rect 2090 1516 2092 1524
rect 2100 1516 2102 1524
rect 2090 1514 2102 1516
rect 2186 1644 2198 1646
rect 2186 1636 2188 1644
rect 2196 1636 2198 1644
rect 2154 1504 2166 1506
rect 2154 1496 2156 1504
rect 2164 1496 2166 1504
rect 1834 1056 1836 1064
rect 1844 1056 1846 1064
rect 1834 1054 1846 1056
rect 1962 1084 1974 1086
rect 1962 1076 1964 1084
rect 1972 1076 1974 1084
rect 1450 936 1452 944
rect 1460 936 1462 944
rect 1162 916 1164 924
rect 1172 916 1174 924
rect 1162 914 1174 916
rect 1226 924 1238 926
rect 1226 916 1228 924
rect 1236 916 1238 924
rect 1040 806 1044 814
rect 1052 806 1056 814
rect 1064 806 1068 814
rect 1076 806 1080 814
rect 1088 806 1092 814
rect 1100 806 1104 814
rect 938 656 940 664
rect 948 656 950 664
rect 938 654 950 656
rect 522 536 524 544
rect 532 536 534 544
rect 522 534 534 536
rect 1040 414 1104 806
rect 1194 784 1206 786
rect 1194 776 1196 784
rect 1204 776 1206 784
rect 1194 584 1206 776
rect 1226 744 1238 916
rect 1226 736 1228 744
rect 1236 736 1238 744
rect 1226 734 1238 736
rect 1194 576 1196 584
rect 1204 576 1206 584
rect 1194 574 1206 576
rect 1290 724 1302 726
rect 1290 716 1292 724
rect 1300 716 1302 724
rect 1040 406 1044 414
rect 1052 406 1056 414
rect 1064 406 1068 414
rect 1076 406 1080 414
rect 1088 406 1092 414
rect 1100 406 1104 414
rect 1040 14 1104 406
rect 1290 304 1302 716
rect 1450 704 1462 936
rect 1610 924 1622 926
rect 1610 916 1612 924
rect 1620 916 1622 924
rect 1610 884 1622 916
rect 1610 876 1612 884
rect 1620 876 1622 884
rect 1610 874 1622 876
rect 1738 924 1750 926
rect 1738 916 1740 924
rect 1748 916 1750 924
rect 1738 844 1750 916
rect 1930 904 1942 906
rect 1930 896 1932 904
rect 1940 896 1942 904
rect 1738 836 1740 844
rect 1748 836 1750 844
rect 1738 834 1750 836
rect 1770 844 1782 846
rect 1770 836 1772 844
rect 1780 836 1782 844
rect 1450 696 1452 704
rect 1460 696 1462 704
rect 1450 694 1462 696
rect 1482 684 1494 686
rect 1482 676 1484 684
rect 1492 676 1494 684
rect 1482 384 1494 676
rect 1546 684 1558 686
rect 1546 676 1548 684
rect 1556 676 1558 684
rect 1546 644 1558 676
rect 1674 684 1686 686
rect 1674 676 1676 684
rect 1684 676 1686 684
rect 1546 636 1548 644
rect 1556 636 1558 644
rect 1546 634 1558 636
rect 1578 644 1590 646
rect 1578 636 1580 644
rect 1588 636 1590 644
rect 1482 376 1484 384
rect 1492 376 1494 384
rect 1482 374 1494 376
rect 1290 296 1292 304
rect 1300 296 1302 304
rect 1290 294 1302 296
rect 1578 144 1590 636
rect 1674 604 1686 676
rect 1770 644 1782 836
rect 1770 636 1772 644
rect 1780 636 1782 644
rect 1770 634 1782 636
rect 1674 596 1676 604
rect 1684 596 1686 604
rect 1674 594 1686 596
rect 1738 564 1750 566
rect 1738 556 1740 564
rect 1748 556 1750 564
rect 1738 484 1750 556
rect 1930 564 1942 896
rect 1930 556 1932 564
rect 1940 556 1942 564
rect 1930 554 1942 556
rect 1962 564 1974 1076
rect 2026 1074 2070 1086
rect 2090 1484 2102 1486
rect 2090 1476 2092 1484
rect 2100 1476 2102 1484
rect 2026 924 2038 1074
rect 2026 916 2028 924
rect 2036 916 2038 924
rect 2026 914 2038 916
rect 2058 1044 2070 1046
rect 2058 1036 2060 1044
rect 2068 1036 2070 1044
rect 2058 804 2070 1036
rect 2058 796 2060 804
rect 2068 796 2070 804
rect 2058 794 2070 796
rect 2090 704 2102 1476
rect 2154 1464 2166 1496
rect 2154 1456 2156 1464
rect 2164 1456 2166 1464
rect 2154 1324 2166 1456
rect 2154 1316 2156 1324
rect 2164 1316 2166 1324
rect 2154 1314 2166 1316
rect 2154 1144 2166 1146
rect 2154 1136 2156 1144
rect 2164 1136 2166 1144
rect 2090 696 2092 704
rect 2100 696 2102 704
rect 2090 694 2102 696
rect 2122 1044 2134 1046
rect 2122 1036 2124 1044
rect 2132 1036 2134 1044
rect 2122 704 2134 1036
rect 2154 884 2166 1136
rect 2186 1084 2198 1636
rect 2218 1604 2230 1606
rect 2218 1596 2220 1604
rect 2228 1596 2230 1604
rect 2218 1224 2230 1596
rect 2250 1344 2262 1976
rect 2282 1704 2294 2056
rect 2346 1724 2358 2136
rect 2346 1716 2348 1724
rect 2356 1716 2358 1724
rect 2346 1714 2358 1716
rect 2378 2104 2390 2106
rect 2378 2096 2380 2104
rect 2388 2096 2390 2104
rect 2282 1696 2284 1704
rect 2292 1696 2294 1704
rect 2282 1694 2294 1696
rect 2378 1664 2390 2096
rect 2442 2104 2454 2106
rect 2442 2096 2444 2104
rect 2452 2096 2454 2104
rect 2410 2084 2422 2086
rect 2410 2076 2412 2084
rect 2420 2076 2422 2084
rect 2410 1924 2422 2076
rect 2442 2004 2454 2096
rect 2442 1996 2444 2004
rect 2452 1996 2454 2004
rect 2442 1994 2454 1996
rect 2410 1916 2412 1924
rect 2420 1916 2422 1924
rect 2410 1914 2422 1916
rect 2378 1656 2380 1664
rect 2388 1656 2390 1664
rect 2378 1654 2390 1656
rect 2410 1864 2422 1866
rect 2410 1856 2412 1864
rect 2420 1856 2422 1864
rect 2282 1564 2294 1566
rect 2282 1556 2284 1564
rect 2292 1556 2294 1564
rect 2282 1404 2294 1556
rect 2378 1564 2390 1566
rect 2378 1556 2380 1564
rect 2388 1556 2390 1564
rect 2282 1396 2284 1404
rect 2292 1396 2294 1404
rect 2282 1394 2294 1396
rect 2346 1464 2358 1466
rect 2346 1456 2348 1464
rect 2356 1456 2358 1464
rect 2250 1336 2252 1344
rect 2260 1336 2262 1344
rect 2250 1334 2262 1336
rect 2218 1216 2220 1224
rect 2228 1216 2230 1224
rect 2218 1214 2230 1216
rect 2186 1076 2188 1084
rect 2196 1076 2198 1084
rect 2186 1074 2198 1076
rect 2250 1144 2262 1146
rect 2250 1136 2252 1144
rect 2260 1136 2262 1144
rect 2154 876 2156 884
rect 2164 876 2166 884
rect 2154 874 2166 876
rect 2122 696 2124 704
rect 2132 696 2134 704
rect 2122 694 2134 696
rect 2154 684 2166 686
rect 2154 676 2156 684
rect 2164 676 2166 684
rect 1962 556 1964 564
rect 1972 556 1974 564
rect 1962 554 1974 556
rect 2090 624 2102 626
rect 2090 616 2092 624
rect 2100 616 2102 624
rect 1738 476 1740 484
rect 1748 476 1750 484
rect 1738 474 1750 476
rect 1578 136 1580 144
rect 1588 136 1590 144
rect 1578 134 1590 136
rect 1802 304 1814 306
rect 1802 296 1804 304
rect 1812 296 1814 304
rect 1802 124 1814 296
rect 2090 204 2102 616
rect 2090 196 2092 204
rect 2100 196 2102 204
rect 2090 194 2102 196
rect 1802 116 1804 124
rect 1812 116 1814 124
rect 1802 114 1814 116
rect 2154 64 2166 676
rect 2186 684 2198 686
rect 2186 676 2188 684
rect 2196 676 2198 684
rect 2186 484 2198 676
rect 2250 544 2262 1136
rect 2346 1124 2358 1456
rect 2378 1284 2390 1556
rect 2410 1384 2422 1856
rect 2474 1724 2486 2676
rect 2506 2644 2518 2646
rect 2506 2636 2508 2644
rect 2516 2636 2518 2644
rect 2506 2364 2518 2636
rect 2506 2356 2508 2364
rect 2516 2356 2518 2364
rect 2506 2354 2518 2356
rect 2544 2614 2608 3006
rect 2544 2606 2548 2614
rect 2556 2606 2560 2614
rect 2568 2606 2572 2614
rect 2580 2606 2584 2614
rect 2592 2606 2596 2614
rect 2604 2606 2608 2614
rect 2506 2244 2518 2246
rect 2506 2236 2508 2244
rect 2516 2236 2518 2244
rect 2506 2144 2518 2236
rect 2506 2136 2508 2144
rect 2516 2136 2518 2144
rect 2506 2134 2518 2136
rect 2544 2214 2608 2606
rect 2666 2964 2678 2966
rect 2666 2956 2668 2964
rect 2676 2956 2678 2964
rect 2666 2604 2678 2956
rect 2666 2596 2668 2604
rect 2676 2596 2678 2604
rect 2666 2594 2678 2596
rect 2666 2524 2694 2526
rect 2666 2516 2684 2524
rect 2692 2516 2694 2524
rect 2666 2514 2694 2516
rect 2666 2446 2678 2514
rect 2634 2444 2678 2446
rect 2634 2436 2636 2444
rect 2644 2436 2678 2444
rect 2634 2434 2678 2436
rect 2666 2324 2678 2326
rect 2666 2316 2668 2324
rect 2676 2316 2678 2324
rect 2544 2206 2548 2214
rect 2556 2206 2560 2214
rect 2568 2206 2572 2214
rect 2580 2206 2584 2214
rect 2592 2206 2596 2214
rect 2604 2206 2608 2214
rect 2474 1716 2476 1724
rect 2484 1716 2486 1724
rect 2410 1376 2412 1384
rect 2420 1376 2422 1384
rect 2410 1374 2422 1376
rect 2442 1604 2454 1606
rect 2442 1596 2444 1604
rect 2452 1596 2454 1604
rect 2442 1304 2454 1596
rect 2474 1504 2486 1716
rect 2474 1496 2476 1504
rect 2484 1496 2486 1504
rect 2474 1494 2486 1496
rect 2544 1814 2608 2206
rect 2634 2304 2646 2306
rect 2634 2296 2636 2304
rect 2644 2296 2646 2304
rect 2634 2204 2646 2296
rect 2634 2196 2636 2204
rect 2644 2196 2646 2204
rect 2634 2194 2646 2196
rect 2666 2284 2678 2316
rect 2666 2276 2668 2284
rect 2676 2276 2678 2284
rect 2666 2064 2678 2276
rect 2666 2056 2668 2064
rect 2676 2056 2678 2064
rect 2666 2054 2678 2056
rect 2698 2124 2710 2126
rect 2698 2116 2700 2124
rect 2708 2116 2710 2124
rect 2698 1984 2710 2116
rect 2730 2124 2742 3096
rect 2890 3244 2902 3246
rect 2890 3236 2892 3244
rect 2900 3236 2902 3244
rect 2890 2904 2902 3236
rect 2890 2896 2892 2904
rect 2900 2896 2902 2904
rect 2890 2894 2902 2896
rect 2922 3184 2934 3186
rect 2922 3176 2924 3184
rect 2932 3176 2934 3184
rect 2762 2884 2774 2886
rect 2762 2876 2764 2884
rect 2772 2876 2774 2884
rect 2762 2844 2774 2876
rect 2762 2836 2764 2844
rect 2772 2836 2774 2844
rect 2762 2834 2774 2836
rect 2794 2884 2806 2886
rect 2794 2876 2796 2884
rect 2804 2876 2806 2884
rect 2794 2764 2806 2876
rect 2794 2756 2796 2764
rect 2804 2756 2806 2764
rect 2794 2754 2806 2756
rect 2922 2724 2934 3176
rect 3722 3144 3734 3146
rect 3722 3136 3724 3144
rect 3732 3136 3734 3144
rect 2922 2716 2924 2724
rect 2932 2716 2934 2724
rect 2922 2714 2934 2716
rect 2986 3104 2998 3106
rect 2986 3096 2988 3104
rect 2996 3096 2998 3104
rect 2986 2644 2998 3096
rect 3082 2964 3094 2966
rect 3082 2956 3084 2964
rect 3092 2956 3094 2964
rect 3082 2864 3094 2956
rect 3082 2856 3084 2864
rect 3092 2856 3094 2864
rect 3082 2854 3094 2856
rect 3338 2864 3350 2866
rect 3338 2856 3340 2864
rect 3348 2856 3350 2864
rect 3274 2844 3286 2846
rect 3274 2836 3276 2844
rect 3284 2836 3286 2844
rect 3274 2724 3286 2836
rect 3274 2716 3276 2724
rect 3284 2716 3286 2724
rect 3274 2714 3286 2716
rect 2986 2636 2988 2644
rect 2996 2636 2998 2644
rect 2986 2634 2998 2636
rect 3050 2664 3062 2666
rect 3050 2656 3052 2664
rect 3060 2656 3062 2664
rect 3050 2646 3062 2656
rect 3050 2644 3158 2646
rect 3050 2636 3148 2644
rect 3156 2636 3158 2644
rect 3050 2634 3158 2636
rect 2730 2116 2732 2124
rect 2740 2116 2742 2124
rect 2730 2114 2742 2116
rect 2762 2604 2774 2606
rect 2762 2596 2764 2604
rect 2772 2596 2774 2604
rect 2762 2444 2774 2596
rect 2762 2436 2764 2444
rect 2772 2436 2774 2444
rect 2762 2344 2774 2436
rect 3018 2604 3030 2606
rect 3018 2596 3020 2604
rect 3028 2596 3030 2604
rect 3018 2424 3030 2596
rect 3018 2416 3020 2424
rect 3028 2416 3030 2424
rect 3018 2414 3030 2416
rect 3050 2524 3062 2526
rect 3050 2516 3052 2524
rect 3060 2516 3062 2524
rect 2762 2336 2764 2344
rect 2772 2336 2774 2344
rect 2762 2284 2774 2336
rect 2890 2404 2902 2406
rect 2890 2396 2892 2404
rect 2900 2396 2902 2404
rect 2762 2276 2764 2284
rect 2772 2276 2774 2284
rect 2698 1976 2700 1984
rect 2708 1976 2710 1984
rect 2698 1974 2710 1976
rect 2762 1964 2774 2276
rect 2826 2324 2838 2326
rect 2826 2316 2828 2324
rect 2836 2316 2838 2324
rect 2826 2284 2838 2316
rect 2826 2276 2828 2284
rect 2836 2276 2838 2284
rect 2826 2274 2838 2276
rect 2858 2244 2870 2246
rect 2858 2236 2860 2244
rect 2868 2236 2870 2244
rect 2762 1956 2764 1964
rect 2772 1956 2774 1964
rect 2762 1954 2774 1956
rect 2826 2004 2838 2006
rect 2826 1996 2828 2004
rect 2836 1996 2838 2004
rect 2544 1806 2548 1814
rect 2556 1806 2560 1814
rect 2568 1806 2572 1814
rect 2580 1806 2584 1814
rect 2592 1806 2596 1814
rect 2604 1806 2608 1814
rect 2442 1296 2444 1304
rect 2452 1296 2454 1304
rect 2442 1294 2454 1296
rect 2544 1414 2608 1806
rect 2794 1864 2806 1866
rect 2794 1856 2796 1864
rect 2804 1856 2806 1864
rect 2762 1764 2774 1766
rect 2762 1756 2764 1764
rect 2772 1756 2774 1764
rect 2544 1406 2548 1414
rect 2556 1406 2560 1414
rect 2568 1406 2572 1414
rect 2580 1406 2584 1414
rect 2592 1406 2596 1414
rect 2604 1406 2608 1414
rect 2378 1276 2380 1284
rect 2388 1276 2390 1284
rect 2378 1274 2390 1276
rect 2346 1116 2348 1124
rect 2356 1116 2358 1124
rect 2346 1114 2358 1116
rect 2442 1244 2454 1246
rect 2442 1236 2444 1244
rect 2452 1236 2454 1244
rect 2442 1184 2454 1236
rect 2442 1176 2444 1184
rect 2452 1176 2454 1184
rect 2410 984 2422 986
rect 2410 976 2412 984
rect 2420 976 2422 984
rect 2346 784 2358 786
rect 2346 776 2348 784
rect 2356 776 2358 784
rect 2346 624 2358 776
rect 2346 616 2348 624
rect 2356 616 2358 624
rect 2346 614 2358 616
rect 2378 764 2390 766
rect 2378 756 2380 764
rect 2388 756 2390 764
rect 2378 704 2390 756
rect 2378 696 2380 704
rect 2388 696 2390 704
rect 2250 536 2252 544
rect 2260 536 2262 544
rect 2250 534 2262 536
rect 2186 476 2188 484
rect 2196 476 2198 484
rect 2186 474 2198 476
rect 2378 144 2390 696
rect 2410 584 2422 976
rect 2442 704 2454 1176
rect 2474 1024 2486 1026
rect 2474 1016 2476 1024
rect 2484 1016 2486 1024
rect 2474 924 2486 1016
rect 2474 916 2476 924
rect 2484 916 2486 924
rect 2474 914 2486 916
rect 2544 1014 2608 1406
rect 2634 1624 2646 1626
rect 2634 1616 2636 1624
rect 2644 1616 2646 1624
rect 2634 1344 2646 1616
rect 2666 1524 2678 1526
rect 2666 1516 2668 1524
rect 2676 1516 2678 1524
rect 2666 1424 2678 1516
rect 2762 1484 2774 1756
rect 2794 1504 2806 1856
rect 2794 1496 2796 1504
rect 2804 1496 2806 1504
rect 2794 1494 2806 1496
rect 2762 1476 2764 1484
rect 2772 1476 2774 1484
rect 2762 1474 2774 1476
rect 2666 1416 2668 1424
rect 2676 1416 2678 1424
rect 2666 1414 2678 1416
rect 2634 1336 2636 1344
rect 2644 1336 2646 1344
rect 2634 1334 2646 1336
rect 2826 1224 2838 1996
rect 2858 1804 2870 2236
rect 2890 2224 2902 2396
rect 2890 2216 2892 2224
rect 2900 2216 2902 2224
rect 2890 2214 2902 2216
rect 2954 2204 2966 2206
rect 2954 2196 2956 2204
rect 2964 2196 2966 2204
rect 2954 1884 2966 2196
rect 3050 2204 3062 2516
rect 3050 2196 3052 2204
rect 3060 2196 3062 2204
rect 3050 2194 3062 2196
rect 3082 2204 3094 2206
rect 3082 2196 3084 2204
rect 3092 2196 3094 2204
rect 3082 2024 3094 2196
rect 3338 2204 3350 2856
rect 3530 2704 3542 2706
rect 3530 2696 3532 2704
rect 3540 2696 3542 2704
rect 3530 2686 3542 2696
rect 3722 2704 3734 3136
rect 3722 2696 3724 2704
rect 3732 2696 3734 2704
rect 3722 2694 3734 2696
rect 3530 2674 3574 2686
rect 3562 2644 3574 2674
rect 3562 2636 3564 2644
rect 3572 2636 3574 2644
rect 3562 2634 3574 2636
rect 3818 2604 3830 2606
rect 3818 2596 3820 2604
rect 3828 2596 3830 2604
rect 3626 2544 3638 2546
rect 3626 2536 3628 2544
rect 3636 2536 3638 2544
rect 3338 2196 3340 2204
rect 3348 2196 3350 2204
rect 3338 2194 3350 2196
rect 3434 2524 3446 2526
rect 3434 2516 3436 2524
rect 3444 2516 3446 2524
rect 3082 2016 3084 2024
rect 3092 2016 3094 2024
rect 3082 2014 3094 2016
rect 3306 1944 3318 1946
rect 3306 1936 3308 1944
rect 3316 1936 3318 1944
rect 2954 1876 2956 1884
rect 2964 1876 2966 1884
rect 2954 1874 2966 1876
rect 2986 1884 2998 1886
rect 2986 1876 2988 1884
rect 2996 1876 2998 1884
rect 2858 1796 2860 1804
rect 2868 1796 2870 1804
rect 2858 1794 2870 1796
rect 2954 1824 2966 1826
rect 2954 1816 2956 1824
rect 2964 1816 2966 1824
rect 2826 1216 2828 1224
rect 2836 1216 2838 1224
rect 2826 1214 2838 1216
rect 2858 1664 2870 1666
rect 2858 1656 2860 1664
rect 2868 1656 2870 1664
rect 2858 1224 2870 1656
rect 2954 1504 2966 1816
rect 2986 1624 2998 1876
rect 3274 1724 3286 1726
rect 3274 1716 3276 1724
rect 3284 1716 3286 1724
rect 2986 1616 2988 1624
rect 2996 1616 2998 1624
rect 2986 1614 2998 1616
rect 3178 1624 3190 1626
rect 3178 1616 3180 1624
rect 3188 1616 3190 1624
rect 2954 1496 2956 1504
rect 2964 1496 2966 1504
rect 2954 1494 2966 1496
rect 3114 1524 3126 1526
rect 3114 1516 3116 1524
rect 3124 1516 3126 1524
rect 3018 1404 3030 1406
rect 3018 1396 3020 1404
rect 3028 1396 3030 1404
rect 2858 1216 2860 1224
rect 2868 1216 2870 1224
rect 2858 1214 2870 1216
rect 2922 1364 2934 1366
rect 2922 1356 2924 1364
rect 2932 1356 2934 1364
rect 2762 1144 2774 1146
rect 2762 1136 2764 1144
rect 2772 1136 2774 1144
rect 2544 1006 2548 1014
rect 2556 1006 2560 1014
rect 2568 1006 2572 1014
rect 2580 1006 2584 1014
rect 2592 1006 2596 1014
rect 2604 1006 2608 1014
rect 2442 696 2444 704
rect 2452 696 2454 704
rect 2442 694 2454 696
rect 2474 824 2486 826
rect 2474 816 2476 824
rect 2484 816 2486 824
rect 2410 576 2412 584
rect 2420 576 2422 584
rect 2410 574 2422 576
rect 2474 584 2486 816
rect 2474 576 2476 584
rect 2484 576 2486 584
rect 2474 574 2486 576
rect 2544 614 2608 1006
rect 2634 1064 2646 1066
rect 2634 1056 2636 1064
rect 2644 1056 2646 1064
rect 2634 924 2646 1056
rect 2762 944 2774 1136
rect 2890 1124 2902 1126
rect 2890 1116 2892 1124
rect 2900 1116 2902 1124
rect 2762 936 2764 944
rect 2772 936 2774 944
rect 2762 934 2774 936
rect 2826 1004 2838 1006
rect 2826 996 2828 1004
rect 2836 996 2838 1004
rect 2634 916 2636 924
rect 2644 916 2646 924
rect 2634 914 2646 916
rect 2826 864 2838 996
rect 2826 856 2828 864
rect 2836 856 2838 864
rect 2826 854 2838 856
rect 2858 1004 2870 1006
rect 2858 996 2860 1004
rect 2868 996 2870 1004
rect 2666 804 2678 806
rect 2666 796 2668 804
rect 2676 796 2678 804
rect 2544 606 2548 614
rect 2556 606 2560 614
rect 2568 606 2572 614
rect 2580 606 2584 614
rect 2592 606 2596 614
rect 2604 606 2608 614
rect 2378 136 2380 144
rect 2388 136 2390 144
rect 2378 134 2390 136
rect 2544 214 2608 606
rect 2634 764 2646 766
rect 2634 756 2636 764
rect 2644 756 2646 764
rect 2634 724 2646 756
rect 2634 716 2636 724
rect 2644 716 2646 724
rect 2634 564 2646 716
rect 2634 556 2636 564
rect 2644 556 2646 564
rect 2634 554 2646 556
rect 2666 444 2678 796
rect 2762 804 2774 806
rect 2762 796 2764 804
rect 2772 796 2774 804
rect 2698 684 2710 686
rect 2698 676 2700 684
rect 2708 676 2710 684
rect 2698 464 2710 676
rect 2698 456 2700 464
rect 2708 456 2710 464
rect 2698 454 2710 456
rect 2730 584 2742 586
rect 2730 576 2732 584
rect 2740 576 2742 584
rect 2666 436 2668 444
rect 2676 436 2678 444
rect 2666 434 2678 436
rect 2730 304 2742 576
rect 2762 524 2774 796
rect 2762 516 2764 524
rect 2772 516 2774 524
rect 2762 514 2774 516
rect 2826 544 2838 546
rect 2826 536 2828 544
rect 2836 536 2838 544
rect 2762 484 2774 486
rect 2762 476 2764 484
rect 2772 476 2774 484
rect 2762 324 2774 476
rect 2762 316 2764 324
rect 2772 316 2774 324
rect 2762 314 2774 316
rect 2730 296 2732 304
rect 2740 296 2742 304
rect 2730 294 2742 296
rect 2544 206 2548 214
rect 2556 206 2560 214
rect 2568 206 2572 214
rect 2580 206 2584 214
rect 2592 206 2596 214
rect 2604 206 2608 214
rect 2154 56 2156 64
rect 2164 56 2166 64
rect 2154 54 2166 56
rect 1040 6 1044 14
rect 1052 6 1056 14
rect 1064 6 1068 14
rect 1076 6 1080 14
rect 1088 6 1092 14
rect 1100 6 1104 14
rect 1040 -10 1104 6
rect 2544 -10 2608 206
rect 2826 164 2838 536
rect 2858 224 2870 996
rect 2890 624 2902 1116
rect 2922 944 2934 1356
rect 2954 1364 2966 1366
rect 2954 1356 2956 1364
rect 2964 1356 2966 1364
rect 2954 1204 2966 1356
rect 3018 1304 3030 1396
rect 3114 1404 3126 1516
rect 3178 1444 3190 1616
rect 3178 1436 3180 1444
rect 3188 1436 3190 1444
rect 3178 1434 3190 1436
rect 3114 1396 3116 1404
rect 3124 1396 3126 1404
rect 3114 1394 3126 1396
rect 3082 1384 3094 1386
rect 3082 1376 3084 1384
rect 3092 1376 3094 1384
rect 3082 1344 3094 1376
rect 3082 1336 3084 1344
rect 3092 1336 3094 1344
rect 3082 1334 3094 1336
rect 3018 1296 3020 1304
rect 3028 1296 3030 1304
rect 3018 1294 3030 1296
rect 2954 1196 2956 1204
rect 2964 1196 2966 1204
rect 2954 1194 2966 1196
rect 3178 1264 3190 1266
rect 3178 1256 3180 1264
rect 3188 1256 3190 1264
rect 2986 1084 2998 1086
rect 2986 1076 2988 1084
rect 2996 1076 2998 1084
rect 2986 1044 2998 1076
rect 2986 1036 2988 1044
rect 2996 1036 2998 1044
rect 2986 1034 2998 1036
rect 3178 964 3190 1256
rect 3178 956 3180 964
rect 3188 956 3190 964
rect 3178 954 3190 956
rect 3210 1204 3222 1206
rect 3210 1196 3212 1204
rect 3220 1196 3222 1204
rect 2922 936 2924 944
rect 2932 936 2934 944
rect 2922 934 2934 936
rect 2954 944 2966 946
rect 2954 936 2956 944
rect 2964 936 2966 944
rect 2922 764 2934 766
rect 2922 756 2924 764
rect 2932 756 2934 764
rect 2922 724 2934 756
rect 2922 716 2924 724
rect 2932 716 2934 724
rect 2922 714 2934 716
rect 2890 616 2892 624
rect 2900 616 2902 624
rect 2890 614 2902 616
rect 2954 664 2966 936
rect 2954 656 2956 664
rect 2964 656 2966 664
rect 2954 564 2966 656
rect 2954 556 2956 564
rect 2964 556 2966 564
rect 2954 554 2966 556
rect 3082 824 3094 826
rect 3082 816 3084 824
rect 3092 816 3094 824
rect 2986 444 2998 446
rect 2986 436 2988 444
rect 2996 436 2998 444
rect 2858 216 2860 224
rect 2868 216 2870 224
rect 2858 214 2870 216
rect 2890 324 2902 326
rect 2890 316 2892 324
rect 2900 316 2902 324
rect 2826 156 2828 164
rect 2836 156 2838 164
rect 2826 154 2838 156
rect 2890 104 2902 316
rect 2986 124 2998 436
rect 3082 324 3094 816
rect 3210 684 3222 1196
rect 3274 1104 3286 1716
rect 3306 1324 3318 1936
rect 3434 1944 3446 2516
rect 3466 2404 3478 2406
rect 3466 2396 3468 2404
rect 3476 2396 3478 2404
rect 3466 2144 3478 2396
rect 3466 2136 3468 2144
rect 3476 2136 3478 2144
rect 3466 2134 3478 2136
rect 3434 1936 3436 1944
rect 3444 1936 3446 1944
rect 3434 1934 3446 1936
rect 3562 2064 3574 2066
rect 3562 2056 3564 2064
rect 3572 2056 3574 2064
rect 3434 1864 3446 1866
rect 3434 1856 3436 1864
rect 3444 1856 3446 1864
rect 3306 1316 3308 1324
rect 3316 1316 3318 1324
rect 3306 1314 3318 1316
rect 3370 1564 3382 1566
rect 3370 1556 3372 1564
rect 3380 1556 3382 1564
rect 3370 1244 3382 1556
rect 3370 1236 3372 1244
rect 3380 1236 3382 1244
rect 3370 1234 3382 1236
rect 3274 1096 3276 1104
rect 3284 1096 3286 1104
rect 3274 1094 3286 1096
rect 3434 1104 3446 1856
rect 3562 1684 3574 2056
rect 3562 1676 3564 1684
rect 3572 1676 3574 1684
rect 3562 1674 3574 1676
rect 3434 1096 3436 1104
rect 3444 1096 3446 1104
rect 3434 1094 3446 1096
rect 3466 1584 3478 1586
rect 3466 1576 3468 1584
rect 3476 1576 3478 1584
rect 3466 1084 3478 1576
rect 3626 1484 3638 2536
rect 3626 1476 3628 1484
rect 3636 1476 3638 1484
rect 3626 1474 3638 1476
rect 3818 2424 3830 2596
rect 3818 2416 3820 2424
rect 3828 2416 3830 2424
rect 3818 1844 3830 2416
rect 3850 2064 3862 3416
rect 3914 3324 3926 3326
rect 3914 3316 3916 3324
rect 3924 3316 3926 3324
rect 3914 2304 3926 3316
rect 3914 2296 3916 2304
rect 3924 2296 3926 2304
rect 3914 2294 3926 2296
rect 4048 3214 4112 3416
rect 4048 3206 4052 3214
rect 4060 3206 4064 3214
rect 4072 3206 4076 3214
rect 4084 3206 4088 3214
rect 4096 3206 4100 3214
rect 4108 3206 4112 3214
rect 4048 2814 4112 3206
rect 4458 3084 4470 3086
rect 4458 3076 4460 3084
rect 4468 3076 4470 3084
rect 4048 2806 4052 2814
rect 4060 2806 4064 2814
rect 4072 2806 4076 2814
rect 4084 2806 4088 2814
rect 4096 2806 4100 2814
rect 4108 2806 4112 2814
rect 4048 2414 4112 2806
rect 4170 2984 4182 2986
rect 4170 2976 4172 2984
rect 4180 2976 4182 2984
rect 4170 2724 4182 2976
rect 4170 2716 4172 2724
rect 4180 2716 4182 2724
rect 4170 2714 4182 2716
rect 4298 2984 4310 2986
rect 4298 2976 4300 2984
rect 4308 2976 4310 2984
rect 4298 2584 4310 2976
rect 4458 2924 4470 3076
rect 4458 2916 4460 2924
rect 4468 2916 4470 2924
rect 4458 2914 4470 2916
rect 4874 2964 4886 2966
rect 4874 2956 4876 2964
rect 4884 2956 4886 2964
rect 4746 2724 4758 2726
rect 4746 2716 4748 2724
rect 4756 2716 4758 2724
rect 4298 2576 4300 2584
rect 4308 2576 4310 2584
rect 4298 2574 4310 2576
rect 4490 2624 4502 2626
rect 4490 2616 4492 2624
rect 4500 2616 4502 2624
rect 4202 2564 4214 2566
rect 4202 2556 4204 2564
rect 4212 2556 4214 2564
rect 4202 2504 4214 2556
rect 4202 2496 4204 2504
rect 4212 2496 4214 2504
rect 4202 2494 4214 2496
rect 4048 2406 4052 2414
rect 4060 2406 4064 2414
rect 4072 2406 4076 2414
rect 4084 2406 4088 2414
rect 4096 2406 4100 2414
rect 4108 2406 4112 2414
rect 3850 2056 3852 2064
rect 3860 2056 3862 2064
rect 3850 2054 3862 2056
rect 3946 2104 3958 2106
rect 3946 2096 3948 2104
rect 3956 2096 3958 2104
rect 3818 1836 3820 1844
rect 3828 1836 3830 1844
rect 3594 1304 3606 1306
rect 3594 1296 3596 1304
rect 3604 1296 3606 1304
rect 3498 1264 3510 1266
rect 3498 1256 3500 1264
rect 3508 1256 3510 1264
rect 3498 1224 3510 1256
rect 3498 1216 3500 1224
rect 3508 1216 3510 1224
rect 3498 1214 3510 1216
rect 3466 1076 3468 1084
rect 3476 1076 3478 1084
rect 3466 1074 3478 1076
rect 3530 1004 3542 1006
rect 3530 996 3532 1004
rect 3540 996 3542 1004
rect 3210 676 3212 684
rect 3220 676 3222 684
rect 3210 674 3222 676
rect 3242 764 3254 766
rect 3242 756 3244 764
rect 3252 756 3254 764
rect 3146 564 3158 566
rect 3146 556 3148 564
rect 3156 556 3158 564
rect 3146 404 3158 556
rect 3242 526 3254 756
rect 3338 584 3350 586
rect 3338 576 3340 584
rect 3348 576 3350 584
rect 3338 566 3350 576
rect 3338 554 3382 566
rect 3370 544 3382 554
rect 3370 536 3372 544
rect 3380 536 3382 544
rect 3370 534 3382 536
rect 3434 564 3446 566
rect 3434 556 3436 564
rect 3444 556 3446 564
rect 3146 396 3148 404
rect 3156 396 3158 404
rect 3082 316 3084 324
rect 3092 316 3094 324
rect 3082 314 3094 316
rect 3114 324 3126 326
rect 3114 316 3116 324
rect 3124 316 3126 324
rect 3114 224 3126 316
rect 3114 216 3116 224
rect 3124 216 3126 224
rect 3114 214 3126 216
rect 3146 224 3158 396
rect 3178 524 3190 526
rect 3178 516 3180 524
rect 3188 516 3190 524
rect 3178 284 3190 516
rect 3178 276 3180 284
rect 3188 276 3190 284
rect 3178 274 3190 276
rect 3210 514 3254 526
rect 3146 216 3148 224
rect 3156 216 3158 224
rect 3146 214 3158 216
rect 3178 144 3190 146
rect 3178 136 3180 144
rect 3188 136 3190 144
rect 3178 126 3190 136
rect 2986 116 2988 124
rect 2996 116 2998 124
rect 2986 114 2998 116
rect 3146 114 3190 126
rect 2890 96 2892 104
rect 2900 96 2902 104
rect 2890 94 2902 96
rect 3146 84 3158 114
rect 3146 76 3148 84
rect 3156 76 3158 84
rect 3146 74 3158 76
rect 3210 64 3222 514
rect 3306 504 3318 506
rect 3306 496 3308 504
rect 3316 496 3318 504
rect 3242 484 3254 486
rect 3242 476 3244 484
rect 3252 476 3254 484
rect 3242 124 3254 476
rect 3306 144 3318 496
rect 3338 284 3350 286
rect 3338 276 3340 284
rect 3348 276 3350 284
rect 3338 224 3350 276
rect 3402 284 3414 286
rect 3402 276 3404 284
rect 3412 276 3414 284
rect 3338 216 3340 224
rect 3348 216 3350 224
rect 3338 214 3350 216
rect 3370 264 3382 266
rect 3370 256 3372 264
rect 3380 256 3382 264
rect 3306 136 3308 144
rect 3316 136 3318 144
rect 3306 134 3318 136
rect 3242 116 3244 124
rect 3252 116 3254 124
rect 3242 114 3254 116
rect 3370 104 3382 256
rect 3402 244 3414 276
rect 3402 236 3404 244
rect 3412 236 3414 244
rect 3402 234 3414 236
rect 3434 144 3446 556
rect 3530 164 3542 996
rect 3594 944 3606 1296
rect 3594 936 3596 944
rect 3604 936 3606 944
rect 3594 934 3606 936
rect 3818 924 3830 1836
rect 3850 1944 3862 1946
rect 3850 1936 3852 1944
rect 3860 1936 3862 1944
rect 3850 1444 3862 1936
rect 3850 1436 3852 1444
rect 3860 1436 3862 1444
rect 3850 1434 3862 1436
rect 3946 1644 3958 2096
rect 3946 1636 3948 1644
rect 3956 1636 3958 1644
rect 3818 916 3820 924
rect 3828 916 3830 924
rect 3818 844 3830 916
rect 3818 836 3820 844
rect 3828 836 3830 844
rect 3818 834 3830 836
rect 3882 864 3894 866
rect 3882 856 3884 864
rect 3892 856 3894 864
rect 3882 524 3894 856
rect 3946 704 3958 1636
rect 4048 2014 4112 2406
rect 4138 2384 4150 2386
rect 4138 2376 4140 2384
rect 4148 2376 4150 2384
rect 4138 2344 4150 2376
rect 4138 2336 4140 2344
rect 4148 2336 4150 2344
rect 4138 2334 4150 2336
rect 4048 2006 4052 2014
rect 4060 2006 4064 2014
rect 4072 2006 4076 2014
rect 4084 2006 4088 2014
rect 4096 2006 4100 2014
rect 4108 2006 4112 2014
rect 4048 1614 4112 2006
rect 4048 1606 4052 1614
rect 4060 1606 4064 1614
rect 4072 1606 4076 1614
rect 4084 1606 4088 1614
rect 4096 1606 4100 1614
rect 4108 1606 4112 1614
rect 3946 696 3948 704
rect 3956 696 3958 704
rect 3946 694 3958 696
rect 3978 1344 3990 1346
rect 3978 1336 3980 1344
rect 3988 1336 3990 1344
rect 3978 684 3990 1336
rect 3978 676 3980 684
rect 3988 676 3990 684
rect 3978 674 3990 676
rect 4048 1214 4112 1606
rect 4138 2144 4150 2146
rect 4138 2136 4140 2144
rect 4148 2136 4150 2144
rect 4138 1804 4150 2136
rect 4490 2144 4502 2616
rect 4746 2304 4758 2716
rect 4746 2296 4748 2304
rect 4756 2296 4758 2304
rect 4746 2294 4758 2296
rect 4778 2684 4790 2686
rect 4778 2676 4780 2684
rect 4788 2676 4790 2684
rect 4490 2136 4492 2144
rect 4500 2136 4502 2144
rect 4490 2134 4502 2136
rect 4138 1796 4140 1804
rect 4148 1796 4150 1804
rect 4138 1424 4150 1796
rect 4522 1844 4534 1846
rect 4522 1836 4524 1844
rect 4532 1836 4534 1844
rect 4138 1416 4140 1424
rect 4148 1416 4150 1424
rect 4138 1414 4150 1416
rect 4234 1784 4246 1786
rect 4234 1776 4236 1784
rect 4244 1776 4246 1784
rect 4048 1206 4052 1214
rect 4060 1206 4064 1214
rect 4072 1206 4076 1214
rect 4084 1206 4088 1214
rect 4096 1206 4100 1214
rect 4108 1206 4112 1214
rect 4048 814 4112 1206
rect 4048 806 4052 814
rect 4060 806 4064 814
rect 4072 806 4076 814
rect 4084 806 4088 814
rect 4096 806 4100 814
rect 4108 806 4112 814
rect 3882 516 3884 524
rect 3892 516 3894 524
rect 3882 514 3894 516
rect 3530 156 3532 164
rect 3540 156 3542 164
rect 3530 154 3542 156
rect 4048 414 4112 806
rect 4234 684 4246 1776
rect 4522 1664 4534 1836
rect 4778 1744 4790 2676
rect 4810 2544 4822 2546
rect 4810 2536 4812 2544
rect 4820 2536 4822 2544
rect 4810 2444 4822 2536
rect 4810 2436 4812 2444
rect 4820 2436 4822 2444
rect 4810 2434 4822 2436
rect 4874 2444 4886 2956
rect 5098 2904 5110 2906
rect 5098 2896 5100 2904
rect 5108 2896 5110 2904
rect 5066 2864 5078 2866
rect 5066 2856 5068 2864
rect 5076 2856 5078 2864
rect 4970 2744 4982 2746
rect 4970 2736 4972 2744
rect 4980 2736 4982 2744
rect 4874 2436 4876 2444
rect 4884 2436 4886 2444
rect 4874 2434 4886 2436
rect 4906 2484 4918 2486
rect 4906 2476 4908 2484
rect 4916 2476 4918 2484
rect 4778 1736 4780 1744
rect 4788 1736 4790 1744
rect 4778 1734 4790 1736
rect 4522 1656 4524 1664
rect 4532 1656 4534 1664
rect 4522 1654 4534 1656
rect 4298 1304 4310 1306
rect 4298 1296 4300 1304
rect 4308 1296 4310 1304
rect 4298 704 4310 1296
rect 4874 1244 4886 1246
rect 4874 1236 4876 1244
rect 4884 1236 4886 1244
rect 4650 1144 4662 1146
rect 4650 1136 4652 1144
rect 4660 1136 4662 1144
rect 4554 1064 4566 1066
rect 4554 1056 4556 1064
rect 4564 1056 4566 1064
rect 4554 724 4566 1056
rect 4554 716 4556 724
rect 4564 716 4566 724
rect 4554 714 4566 716
rect 4618 1004 4630 1006
rect 4618 996 4620 1004
rect 4628 996 4630 1004
rect 4298 696 4300 704
rect 4308 696 4310 704
rect 4298 694 4310 696
rect 4234 676 4236 684
rect 4244 676 4246 684
rect 4234 674 4246 676
rect 4618 624 4630 996
rect 4650 804 4662 1136
rect 4650 796 4652 804
rect 4660 796 4662 804
rect 4650 794 4662 796
rect 4618 616 4620 624
rect 4628 616 4630 624
rect 4618 614 4630 616
rect 4874 524 4886 1236
rect 4906 1224 4918 2476
rect 4970 2484 4982 2736
rect 4970 2476 4972 2484
rect 4980 2476 4982 2484
rect 4970 2474 4982 2476
rect 5034 2604 5046 2606
rect 5034 2596 5036 2604
rect 5044 2596 5046 2604
rect 4938 1904 4950 1906
rect 4938 1896 4940 1904
rect 4948 1896 4950 1904
rect 4938 1764 4950 1896
rect 4938 1756 4940 1764
rect 4948 1756 4950 1764
rect 4938 1754 4950 1756
rect 5034 1344 5046 2596
rect 5066 2544 5078 2856
rect 5066 2536 5068 2544
rect 5076 2536 5078 2544
rect 5066 2534 5078 2536
rect 5066 2504 5078 2506
rect 5066 2496 5068 2504
rect 5076 2496 5078 2504
rect 5066 1944 5078 2496
rect 5066 1936 5068 1944
rect 5076 1936 5078 1944
rect 5066 1934 5078 1936
rect 5098 1964 5110 2896
rect 5098 1956 5100 1964
rect 5108 1956 5110 1964
rect 5066 1884 5078 1886
rect 5066 1876 5068 1884
rect 5076 1876 5078 1884
rect 5066 1704 5078 1876
rect 5066 1696 5068 1704
rect 5076 1696 5078 1704
rect 5066 1694 5078 1696
rect 5034 1336 5036 1344
rect 5044 1336 5046 1344
rect 5034 1334 5046 1336
rect 5066 1364 5078 1366
rect 5066 1356 5068 1364
rect 5076 1356 5078 1364
rect 4906 1216 4908 1224
rect 4916 1216 4918 1224
rect 4906 1214 4918 1216
rect 4938 1124 4950 1126
rect 4938 1116 4940 1124
rect 4948 1116 4950 1124
rect 4938 544 4950 1116
rect 5066 764 5078 1356
rect 5098 1324 5110 1956
rect 5130 1884 5142 1886
rect 5130 1876 5132 1884
rect 5140 1876 5142 1884
rect 5130 1824 5142 1876
rect 5130 1816 5132 1824
rect 5140 1816 5142 1824
rect 5130 1814 5142 1816
rect 5098 1316 5100 1324
rect 5108 1316 5110 1324
rect 5098 1244 5110 1316
rect 5098 1236 5100 1244
rect 5108 1236 5110 1244
rect 5098 1234 5110 1236
rect 5066 756 5068 764
rect 5076 756 5078 764
rect 5066 754 5078 756
rect 4938 536 4940 544
rect 4948 536 4950 544
rect 4938 534 4950 536
rect 4874 516 4876 524
rect 4884 516 4886 524
rect 4874 514 4886 516
rect 4048 406 4052 414
rect 4060 406 4064 414
rect 4072 406 4076 414
rect 4084 406 4088 414
rect 4096 406 4100 414
rect 4108 406 4112 414
rect 3434 136 3436 144
rect 3444 136 3446 144
rect 3434 134 3446 136
rect 3370 96 3372 104
rect 3380 96 3382 104
rect 3370 94 3382 96
rect 3210 56 3212 64
rect 3220 56 3222 64
rect 3210 54 3222 56
rect 4048 14 4112 406
rect 4048 6 4052 14
rect 4060 6 4064 14
rect 4072 6 4076 14
rect 4084 6 4088 14
rect 4096 6 4100 14
rect 4108 6 4112 14
rect 4048 -10 4112 6
use BUFX2  _1426_
timestamp 1591632351
transform -1 0 56 0 -1 210
box -4 -6 52 206
use BUFX2  _1410_
timestamp 1591632351
transform -1 0 104 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1586_
timestamp 1591632351
transform -1 0 296 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _1570_
timestamp 1591632351
transform -1 0 200 0 1 210
box -4 -6 196 206
use DFFPOSX1  _1571_
timestamp 1591632351
transform 1 0 200 0 1 210
box -4 -6 196 206
use OAI21X1  _838_
timestamp 1591632351
transform -1 0 360 0 -1 210
box -4 -6 68 206
use BUFX2  _1427_
timestamp 1591632351
transform -1 0 408 0 -1 210
box -4 -6 52 206
use OAI21X1  _844_
timestamp 1591632351
transform -1 0 472 0 -1 210
box -4 -6 68 206
use OAI21X1  _1367_
timestamp 1591632351
transform -1 0 456 0 1 210
box -4 -6 68 206
use BUFX2  _1407_
timestamp 1591632351
transform -1 0 520 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1583_
timestamp 1591632351
transform -1 0 712 0 -1 210
box -4 -6 196 206
use OAI21X1  _1355_
timestamp 1591632351
transform -1 0 520 0 1 210
box -4 -6 68 206
use OAI21X1  _802_
timestamp 1591632351
transform 1 0 520 0 1 210
box -4 -6 68 206
use OAI21X1  _808_
timestamp 1591632351
transform -1 0 648 0 1 210
box -4 -6 68 206
use OAI21X1  _766_
timestamp 1591632351
transform 1 0 712 0 -1 210
box -4 -6 68 206
use BUFX2  _1411_
timestamp 1591632351
transform -1 0 824 0 -1 210
box -4 -6 52 206
use BUFX2  _1401_
timestamp 1591632351
transform 1 0 648 0 1 210
box -4 -6 52 206
use DFFPOSX1  _1587_
timestamp 1591632351
transform -1 0 888 0 1 210
box -4 -6 196 206
use DFFPOSX1  _1580_
timestamp 1591632351
transform 1 0 824 0 -1 210
box -4 -6 196 206
use OAI21X1  _850_
timestamp 1591632351
transform -1 0 952 0 1 210
box -4 -6 68 206
use OAI21X1  _807_
timestamp 1591632351
transform -1 0 1016 0 1 210
box -4 -6 68 206
use FILL  SFILL10960x2100
timestamp 1591632351
transform 1 0 1096 0 1 210
box -4 -6 20 206
use FILL  SFILL10800x2100
timestamp 1591632351
transform 1 0 1080 0 1 210
box -4 -6 20 206
use FILL  SFILL10640x2100
timestamp 1591632351
transform 1 0 1064 0 1 210
box -4 -6 20 206
use FILL  SFILL10960x100
timestamp 1591632351
transform -1 0 1112 0 -1 210
box -4 -6 20 206
use FILL  SFILL10800x100
timestamp 1591632351
transform -1 0 1096 0 -1 210
box -4 -6 20 206
use FILL  SFILL10640x100
timestamp 1591632351
transform -1 0 1080 0 -1 210
box -4 -6 20 206
use BUFX2  _1408_
timestamp 1591632351
transform -1 0 1064 0 1 210
box -4 -6 52 206
use BUFX2  _1404_
timestamp 1591632351
transform 1 0 1016 0 -1 210
box -4 -6 52 206
use FILL  SFILL11120x2100
timestamp 1591632351
transform 1 0 1112 0 1 210
box -4 -6 20 206
use FILL  SFILL11120x100
timestamp 1591632351
transform -1 0 1128 0 -1 210
box -4 -6 20 206
use OAI21X1  _771_
timestamp 1591632351
transform -1 0 1256 0 -1 210
box -4 -6 68 206
use OAI21X1  _772_
timestamp 1591632351
transform -1 0 1192 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _1584_
timestamp 1591632351
transform -1 0 1320 0 1 210
box -4 -6 196 206
use OAI21X1  _843_
timestamp 1591632351
transform -1 0 1320 0 -1 210
box -4 -6 68 206
use BUFX2  _1403_
timestamp 1591632351
transform -1 0 1368 0 -1 210
box -4 -6 52 206
use BUFX2  _1412_
timestamp 1591632351
transform -1 0 1416 0 -1 210
box -4 -6 52 206
use OAI21X1  _754_
timestamp 1591632351
transform 1 0 1320 0 1 210
box -4 -6 68 206
use DFFPOSX1  _1588_
timestamp 1591632351
transform -1 0 1576 0 1 210
box -4 -6 196 206
use DFFPOSX1  _1579_
timestamp 1591632351
transform -1 0 1608 0 -1 210
box -4 -6 196 206
use BUFX2  _1423_
timestamp 1591632351
transform -1 0 1656 0 -1 210
box -4 -6 52 206
use OAI21X1  _862_
timestamp 1591632351
transform -1 0 1640 0 1 210
box -4 -6 68 206
use DFFPOSX1  _1567_
timestamp 1591632351
transform -1 0 1848 0 -1 210
box -4 -6 196 206
use OAI21X1  _1319_
timestamp 1591632351
transform 1 0 1640 0 1 210
box -4 -6 68 206
use DFFPOSX1  _1572_
timestamp 1591632351
transform 1 0 1704 0 1 210
box -4 -6 196 206
use BUFX2  _1428_
timestamp 1591632351
transform 1 0 1848 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1458_
timestamp 1591632351
transform -1 0 2088 0 -1 210
box -4 -6 196 206
use MUX2X1  _1356_
timestamp 1591632351
transform -1 0 1992 0 1 210
box -4 -6 100 206
use MUX2X1  _839_
timestamp 1591632351
transform -1 0 2088 0 1 210
box -4 -6 100 206
use NAND2X1  _923_
timestamp 1591632351
transform 1 0 2088 0 -1 210
box -4 -6 52 206
use OAI21X1  _924_
timestamp 1591632351
transform -1 0 2200 0 -1 210
box -4 -6 68 206
use OAI22X1  _842_
timestamp 1591632351
transform -1 0 2280 0 -1 210
box -4 -6 84 206
use BUFX2  BUFX2_insert119
timestamp 1591632351
transform 1 0 2088 0 1 210
box -4 -6 52 206
use OAI22X1  _1359_
timestamp 1591632351
transform -1 0 2216 0 1 210
box -4 -6 84 206
use OAI21X1  _841_
timestamp 1591632351
transform -1 0 2344 0 -1 210
box -4 -6 68 206
use NOR2X1  _840_
timestamp 1591632351
transform -1 0 2392 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1501_
timestamp 1591632351
transform 1 0 2392 0 -1 210
box -4 -6 196 206
use OAI21X1  _1358_
timestamp 1591632351
transform -1 0 2280 0 1 210
box -4 -6 68 206
use MUX2X1  _1380_
timestamp 1591632351
transform -1 0 2376 0 1 210
box -4 -6 100 206
use NOR2X1  _1357_
timestamp 1591632351
transform 1 0 2376 0 1 210
box -4 -6 52 206
use MUX2X1  _863_
timestamp 1591632351
transform -1 0 2520 0 1 210
box -4 -6 100 206
use OAI22X1  _1287_
timestamp 1591632351
transform -1 0 2664 0 1 210
box -4 -6 84 206
use FILL  SFILL25840x100
timestamp 1591632351
transform -1 0 2600 0 -1 210
box -4 -6 20 206
use FILL  SFILL26000x100
timestamp 1591632351
transform -1 0 2616 0 -1 210
box -4 -6 20 206
use FILL  SFILL25200x2100
timestamp 1591632351
transform 1 0 2520 0 1 210
box -4 -6 20 206
use FILL  SFILL25360x2100
timestamp 1591632351
transform 1 0 2536 0 1 210
box -4 -6 20 206
use FILL  SFILL25520x2100
timestamp 1591632351
transform 1 0 2552 0 1 210
box -4 -6 20 206
use FILL  SFILL25680x2100
timestamp 1591632351
transform 1 0 2568 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_insert43
timestamp 1591632351
transform -1 0 2696 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1460_
timestamp 1591632351
transform -1 0 2888 0 -1 210
box -4 -6 196 206
use NOR2X1  _1285_
timestamp 1591632351
transform -1 0 2712 0 1 210
box -4 -6 52 206
use OAI21X1  _1286_
timestamp 1591632351
transform -1 0 2776 0 1 210
box -4 -6 68 206
use DFFPOSX1  _1444_
timestamp 1591632351
transform -1 0 2968 0 1 210
box -4 -6 196 206
use FILL  SFILL26160x100
timestamp 1591632351
transform -1 0 2632 0 -1 210
box -4 -6 20 206
use FILL  SFILL26320x100
timestamp 1591632351
transform -1 0 2648 0 -1 210
box -4 -6 20 206
use NAND2X1  _929_
timestamp 1591632351
transform 1 0 2888 0 -1 210
box -4 -6 52 206
use OAI21X1  _930_
timestamp 1591632351
transform -1 0 3000 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _1506_
timestamp 1591632351
transform -1 0 3192 0 -1 210
box -4 -6 196 206
use OAI21X1  _967_
timestamp 1591632351
transform 1 0 2968 0 1 210
box -4 -6 68 206
use NAND2X1  _996_
timestamp 1591632351
transform 1 0 3192 0 -1 210
box -4 -6 52 206
use OAI21X1  _966_
timestamp 1591632351
transform -1 0 3096 0 1 210
box -4 -6 68 206
use MUX2X1  _1320_
timestamp 1591632351
transform -1 0 3192 0 1 210
box -4 -6 100 206
use OAI21X1  _805_
timestamp 1591632351
transform 1 0 3192 0 1 210
box -4 -6 68 206
use OAI21X1  _997_
timestamp 1591632351
transform -1 0 3304 0 -1 210
box -4 -6 68 206
use OAI21X1  _769_
timestamp 1591632351
transform 1 0 3304 0 -1 210
box -4 -6 68 206
use OAI22X1  _770_
timestamp 1591632351
transform -1 0 3448 0 -1 210
box -4 -6 84 206
use OAI22X1  _806_
timestamp 1591632351
transform 1 0 3256 0 1 210
box -4 -6 84 206
use MUX2X1  _1284_
timestamp 1591632351
transform 1 0 3336 0 1 210
box -4 -6 100 206
use NOR2X1  _768_
timestamp 1591632351
transform -1 0 3496 0 -1 210
box -4 -6 52 206
use MUX2X1  _803_
timestamp 1591632351
transform -1 0 3592 0 -1 210
box -4 -6 100 206
use MUX2X1  _767_
timestamp 1591632351
transform 1 0 3592 0 -1 210
box -4 -6 100 206
use DFFPOSX1  _1439_
timestamp 1591632351
transform -1 0 3624 0 1 210
box -4 -6 196 206
use DFFPOSX1  _1436_
timestamp 1591632351
transform -1 0 3880 0 -1 210
box -4 -6 196 206
use OAI21X1  _957_
timestamp 1591632351
transform -1 0 3688 0 1 210
box -4 -6 68 206
use OAI21X1  _950_
timestamp 1591632351
transform 1 0 3688 0 1 210
box -4 -6 68 206
use OAI21X1  _951_
timestamp 1591632351
transform -1 0 3816 0 1 210
box -4 -6 68 206
use DFFPOSX1  _1508_
timestamp 1591632351
transform -1 0 4008 0 1 210
box -4 -6 196 206
use DFFPOSX1  _1452_
timestamp 1591632351
transform -1 0 4072 0 -1 210
box -4 -6 196 206
use NAND2X1  _990_
timestamp 1591632351
transform 1 0 4008 0 1 210
box -4 -6 52 206
use FILL  SFILL41040x2100
timestamp 1591632351
transform 1 0 4104 0 1 210
box -4 -6 20 206
use FILL  SFILL40880x2100
timestamp 1591632351
transform 1 0 4088 0 1 210
box -4 -6 20 206
use FILL  SFILL40720x2100
timestamp 1591632351
transform 1 0 4072 0 1 210
box -4 -6 20 206
use FILL  SFILL40560x2100
timestamp 1591632351
transform 1 0 4056 0 1 210
box -4 -6 20 206
use FILL  SFILL41040x100
timestamp 1591632351
transform -1 0 4120 0 -1 210
box -4 -6 20 206
use FILL  SFILL40880x100
timestamp 1591632351
transform -1 0 4104 0 -1 210
box -4 -6 20 206
use FILL  SFILL40720x100
timestamp 1591632351
transform -1 0 4088 0 -1 210
box -4 -6 20 206
use FILL  SFILL41200x100
timestamp 1591632351
transform -1 0 4136 0 -1 210
box -4 -6 20 206
use OAI21X1  _991_
timestamp 1591632351
transform -1 0 4184 0 1 210
box -4 -6 68 206
use OAI21X1  _906_
timestamp 1591632351
transform -1 0 4248 0 -1 210
box -4 -6 68 206
use NAND2X1  _905_
timestamp 1591632351
transform 1 0 4136 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _1503_
timestamp 1591632351
transform -1 0 4376 0 1 210
box -4 -6 196 206
use DFFPOSX1  _1455_
timestamp 1591632351
transform -1 0 4440 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _1548_
timestamp 1591632351
transform -1 0 4568 0 1 210
box -4 -6 196 206
use OAI21X1  _915_
timestamp 1591632351
transform 1 0 4440 0 -1 210
box -4 -6 68 206
use NAND2X1  _914_
timestamp 1591632351
transform -1 0 4552 0 -1 210
box -4 -6 52 206
use OAI21X1  _985_
timestamp 1591632351
transform 1 0 4552 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _1500_
timestamp 1591632351
transform -1 0 4808 0 -1 210
box -4 -6 196 206
use NAND2X1  _984_
timestamp 1591632351
transform -1 0 4616 0 1 210
box -4 -6 52 206
use INVX1  _1024_
timestamp 1591632351
transform 1 0 4616 0 1 210
box -4 -6 36 206
use DFFPOSX1  _1554_
timestamp 1591632351
transform -1 0 5000 0 -1 210
box -4 -6 196 206
use OAI21X1  _1026_
timestamp 1591632351
transform 1 0 4648 0 1 210
box -4 -6 68 206
use INVX1  _1042_
timestamp 1591632351
transform 1 0 4712 0 1 210
box -4 -6 36 206
use OAI21X1  _1044_
timestamp 1591632351
transform 1 0 4744 0 1 210
box -4 -6 68 206
use INVX1  _1036_
timestamp 1591632351
transform 1 0 4808 0 1 210
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert5
timestamp 1591632351
transform -1 0 5144 0 -1 210
box -4 -6 148 206
use OAI21X1  _1038_
timestamp 1591632351
transform 1 0 4840 0 1 210
box -4 -6 68 206
use DFFPOSX1  _1552_
timestamp 1591632351
transform -1 0 5096 0 1 210
box -4 -6 196 206
use FILL  FILL49040x2100
timestamp 1591632351
transform 1 0 5096 0 1 210
box -4 -6 20 206
use FILL  FILL49200x2100
timestamp 1591632351
transform 1 0 5112 0 1 210
box -4 -6 20 206
use FILL  FILL49360x2100
timestamp 1591632351
transform 1 0 5128 0 1 210
box -4 -6 20 206
use BUFX2  _1420_
timestamp 1591632351
transform -1 0 56 0 -1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert12
timestamp 1591632351
transform 1 0 56 0 -1 610
box -4 -6 148 206
use DFFPOSX1  _1564_
timestamp 1591632351
transform -1 0 392 0 -1 610
box -4 -6 196 206
use OAI21X1  _1283_
timestamp 1591632351
transform -1 0 456 0 -1 610
box -4 -6 68 206
use OAI21X1  _1373_
timestamp 1591632351
transform -1 0 520 0 -1 610
box -4 -6 68 206
use OAI21X1  _1289_
timestamp 1591632351
transform -1 0 584 0 -1 610
box -4 -6 68 206
use OAI21X1  _1361_
timestamp 1591632351
transform -1 0 648 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _1577_
timestamp 1591632351
transform -1 0 840 0 -1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert95
timestamp 1591632351
transform -1 0 888 0 -1 610
box -4 -6 52 206
use OAI21X1  _1288_
timestamp 1591632351
transform -1 0 952 0 -1 610
box -4 -6 68 206
use OAI21X1  _856_
timestamp 1591632351
transform -1 0 1016 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert91
timestamp 1591632351
transform -1 0 1064 0 -1 610
box -4 -6 52 206
use OAI21X1  _855_
timestamp 1591632351
transform -1 0 1192 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert3
timestamp 1591632351
transform -1 0 1240 0 -1 610
box -4 -6 52 206
use FILL  SFILL10640x4100
timestamp 1591632351
transform -1 0 1080 0 -1 610
box -4 -6 20 206
use FILL  SFILL10800x4100
timestamp 1591632351
transform -1 0 1096 0 -1 610
box -4 -6 20 206
use FILL  SFILL10960x4100
timestamp 1591632351
transform -1 0 1112 0 -1 610
box -4 -6 20 206
use FILL  SFILL11120x4100
timestamp 1591632351
transform -1 0 1128 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert0
timestamp 1591632351
transform 1 0 1240 0 -1 610
box -4 -6 52 206
use OAI21X1  _814_
timestamp 1591632351
transform -1 0 1352 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _1526_
timestamp 1591632351
transform -1 0 1544 0 -1 610
box -4 -6 196 206
use OAI21X1  _1360_
timestamp 1591632351
transform -1 0 1608 0 -1 610
box -4 -6 68 206
use OAI21X1  _868_
timestamp 1591632351
transform -1 0 1672 0 -1 610
box -4 -6 68 206
use OAI21X1  _867_
timestamp 1591632351
transform -1 0 1736 0 -1 610
box -4 -6 68 206
use OAI21X1  _820_
timestamp 1591632351
transform -1 0 1800 0 -1 610
box -4 -6 68 206
use OAI21X1  _819_
timestamp 1591632351
transform -1 0 1864 0 -1 610
box -4 -6 68 206
use OAI21X1  _1379_
timestamp 1591632351
transform 1 0 1864 0 -1 610
box -4 -6 68 206
use OAI21X1  _1325_
timestamp 1591632351
transform -1 0 1992 0 -1 610
box -4 -6 68 206
use OAI21X1  _1372_
timestamp 1591632351
transform -1 0 2056 0 -1 610
box -4 -6 68 206
use OAI21X1  _1385_
timestamp 1591632351
transform -1 0 2120 0 -1 610
box -4 -6 68 206
use OAI21X1  _1324_
timestamp 1591632351
transform -1 0 2184 0 -1 610
box -4 -6 68 206
use OAI21X1  _1384_
timestamp 1591632351
transform -1 0 2248 0 -1 610
box -4 -6 68 206
use OAI22X1  _1383_
timestamp 1591632351
transform -1 0 2328 0 -1 610
box -4 -6 84 206
use OAI21X1  _1382_
timestamp 1591632351
transform -1 0 2392 0 -1 610
box -4 -6 68 206
use NOR2X1  _1381_
timestamp 1591632351
transform 1 0 2392 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert121
timestamp 1591632351
transform 1 0 2440 0 -1 610
box -4 -6 52 206
use NAND2X1  _986_
timestamp 1591632351
transform -1 0 2536 0 -1 610
box -4 -6 52 206
use NAND2X1  _998_
timestamp 1591632351
transform 1 0 2600 0 -1 610
box -4 -6 52 206
use FILL  SFILL25360x4100
timestamp 1591632351
transform -1 0 2552 0 -1 610
box -4 -6 20 206
use FILL  SFILL25520x4100
timestamp 1591632351
transform -1 0 2568 0 -1 610
box -4 -6 20 206
use FILL  SFILL25680x4100
timestamp 1591632351
transform -1 0 2584 0 -1 610
box -4 -6 20 206
use FILL  SFILL25840x4100
timestamp 1591632351
transform -1 0 2600 0 -1 610
box -4 -6 20 206
use OAI22X1  _1335_
timestamp 1591632351
transform -1 0 2728 0 -1 610
box -4 -6 84 206
use OAI21X1  _1334_
timestamp 1591632351
transform -1 0 2792 0 -1 610
box -4 -6 68 206
use OAI21X1  _1370_
timestamp 1591632351
transform -1 0 2856 0 -1 610
box -4 -6 68 206
use NOR2X1  _1333_
timestamp 1591632351
transform -1 0 2904 0 -1 610
box -4 -6 52 206
use OAI22X1  _1323_
timestamp 1591632351
transform -1 0 2984 0 -1 610
box -4 -6 84 206
use OAI21X1  _1322_
timestamp 1591632351
transform -1 0 3048 0 -1 610
box -4 -6 68 206
use NOR2X1  _1321_
timestamp 1591632351
transform -1 0 3096 0 -1 610
box -4 -6 52 206
use OAI21X1  _817_
timestamp 1591632351
transform 1 0 3096 0 -1 610
box -4 -6 68 206
use OAI22X1  _818_
timestamp 1591632351
transform 1 0 3160 0 -1 610
box -4 -6 84 206
use NOR2X1  _816_
timestamp 1591632351
transform 1 0 3240 0 -1 610
box -4 -6 52 206
use NOR2X1  _804_
timestamp 1591632351
transform -1 0 3336 0 -1 610
box -4 -6 52 206
use MUX2X1  _1332_
timestamp 1591632351
transform 1 0 3336 0 -1 610
box -4 -6 100 206
use MUX2X1  _815_
timestamp 1591632351
transform -1 0 3528 0 -1 610
box -4 -6 100 206
use OAI21X1  _956_
timestamp 1591632351
transform -1 0 3592 0 -1 610
box -4 -6 68 206
use OAI21X1  _958_
timestamp 1591632351
transform 1 0 3592 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _1440_
timestamp 1591632351
transform -1 0 3848 0 -1 610
box -4 -6 196 206
use OAI21X1  _959_
timestamp 1591632351
transform -1 0 3912 0 -1 610
box -4 -6 68 206
use NAND2X1  _1000_
timestamp 1591632351
transform 1 0 3912 0 -1 610
box -4 -6 52 206
use OAI21X1  _1001_
timestamp 1591632351
transform 1 0 3960 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _1456_
timestamp 1591632351
transform -1 0 4280 0 -1 610
box -4 -6 196 206
use FILL  SFILL40240x4100
timestamp 1591632351
transform -1 0 4040 0 -1 610
box -4 -6 20 206
use FILL  SFILL40400x4100
timestamp 1591632351
transform -1 0 4056 0 -1 610
box -4 -6 20 206
use FILL  SFILL40560x4100
timestamp 1591632351
transform -1 0 4072 0 -1 610
box -4 -6 20 206
use FILL  SFILL40720x4100
timestamp 1591632351
transform -1 0 4088 0 -1 610
box -4 -6 20 206
use NAND2X1  _917_
timestamp 1591632351
transform 1 0 4280 0 -1 610
box -4 -6 52 206
use OAI21X1  _918_
timestamp 1591632351
transform -1 0 4392 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert23
timestamp 1591632351
transform 1 0 4392 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _1555_
timestamp 1591632351
transform -1 0 4632 0 -1 610
box -4 -6 196 206
use INVX2  _904_
timestamp 1591632351
transform -1 0 4664 0 -1 610
box -4 -6 36 206
use NAND3X1  _1025_
timestamp 1591632351
transform -1 0 4728 0 -1 610
box -4 -6 68 206
use INVX2  _922_
timestamp 1591632351
transform -1 0 4760 0 -1 610
box -4 -6 36 206
use NAND3X1  _1043_
timestamp 1591632351
transform 1 0 4760 0 -1 610
box -4 -6 68 206
use INVX2  _916_
timestamp 1591632351
transform -1 0 4856 0 -1 610
box -4 -6 36 206
use NAND3X1  _1037_
timestamp 1591632351
transform -1 0 4920 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _1551_
timestamp 1591632351
transform -1 0 5112 0 -1 610
box -4 -6 196 206
use FILL  FILL49200x4100
timestamp 1591632351
transform -1 0 5128 0 -1 610
box -4 -6 20 206
use FILL  FILL49360x4100
timestamp 1591632351
transform -1 0 5144 0 -1 610
box -4 -6 20 206
use BUFX2  _1405_
timestamp 1591632351
transform -1 0 56 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert100
timestamp 1591632351
transform 1 0 56 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert101
timestamp 1591632351
transform 1 0 104 0 1 610
box -4 -6 52 206
use DFFPOSX1  _1581_
timestamp 1591632351
transform -1 0 344 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert107
timestamp 1591632351
transform 1 0 344 0 1 610
box -4 -6 52 206
use OAI21X1  _778_
timestamp 1591632351
transform -1 0 456 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert105
timestamp 1591632351
transform 1 0 456 0 1 610
box -4 -6 52 206
use OAI21X1  _784_
timestamp 1591632351
transform -1 0 568 0 1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert6
timestamp 1591632351
transform 1 0 568 0 1 610
box -4 -6 148 206
use OAI21X1  _730_
timestamp 1591632351
transform -1 0 776 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert68
timestamp 1591632351
transform 1 0 776 0 1 610
box -4 -6 52 206
use DFFPOSX1  _1494_
timestamp 1591632351
transform 1 0 824 0 1 610
box -4 -6 196 206
use OAI21X1  _973_
timestamp 1591632351
transform 1 0 1016 0 1 610
box -4 -6 68 206
use NAND2X1  _972_
timestamp 1591632351
transform -1 0 1192 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert66
timestamp 1591632351
transform 1 0 1192 0 1 610
box -4 -6 52 206
use FILL  SFILL10800x6100
timestamp 1591632351
transform 1 0 1080 0 1 610
box -4 -6 20 206
use FILL  SFILL10960x6100
timestamp 1591632351
transform 1 0 1096 0 1 610
box -4 -6 20 206
use FILL  SFILL11120x6100
timestamp 1591632351
transform 1 0 1112 0 1 610
box -4 -6 20 206
use FILL  SFILL11280x6100
timestamp 1591632351
transform 1 0 1128 0 1 610
box -4 -6 20 206
use MUX2X1  _1205_
timestamp 1591632351
transform 1 0 1240 0 1 610
box -4 -6 100 206
use MUX2X1  _686_
timestamp 1591632351
transform 1 0 1336 0 1 610
box -4 -6 100 206
use NAND2X1  _1056_
timestamp 1591632351
transform 1 0 1432 0 1 610
box -4 -6 52 206
use OAI21X1  _1057_
timestamp 1591632351
transform -1 0 1544 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert94
timestamp 1591632351
transform 1 0 1544 0 1 610
box -4 -6 52 206
use OAI21X1  _760_
timestamp 1591632351
transform -1 0 1656 0 1 610
box -4 -6 68 206
use OAI21X1  _783_
timestamp 1591632351
transform -1 0 1720 0 1 610
box -4 -6 68 206
use OAI21X1  _1336_
timestamp 1591632351
transform 1 0 1720 0 1 610
box -4 -6 68 206
use OAI21X1  _759_
timestamp 1591632351
transform -1 0 1848 0 1 610
box -4 -6 68 206
use DFFPOSX1  _1442_
timestamp 1591632351
transform -1 0 2040 0 1 610
box -4 -6 196 206
use OAI21X1  _963_
timestamp 1591632351
transform -1 0 2104 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert41
timestamp 1591632351
transform 1 0 2104 0 1 610
box -4 -6 52 206
use OAI22X1  _866_
timestamp 1591632351
transform -1 0 2232 0 1 610
box -4 -6 84 206
use OAI21X1  _865_
timestamp 1591632351
transform -1 0 2296 0 1 610
box -4 -6 68 206
use NOR2X1  _864_
timestamp 1591632351
transform 1 0 2296 0 1 610
box -4 -6 52 206
use OAI22X1  _854_
timestamp 1591632351
transform -1 0 2424 0 1 610
box -4 -6 84 206
use OAI21X1  _987_
timestamp 1591632351
transform 1 0 2424 0 1 610
box -4 -6 68 206
use OAI21X1  _853_
timestamp 1591632351
transform -1 0 2552 0 1 610
box -4 -6 68 206
use FILL  SFILL25520x6100
timestamp 1591632351
transform 1 0 2552 0 1 610
box -4 -6 20 206
use FILL  SFILL25680x6100
timestamp 1591632351
transform 1 0 2568 0 1 610
box -4 -6 20 206
use FILL  SFILL25840x6100
timestamp 1591632351
transform 1 0 2584 0 1 610
box -4 -6 20 206
use FILL  SFILL26000x6100
timestamp 1591632351
transform 1 0 2600 0 1 610
box -4 -6 20 206
use NOR2X1  _852_
timestamp 1591632351
transform -1 0 2664 0 1 610
box -4 -6 52 206
use OAI21X1  _999_
timestamp 1591632351
transform -1 0 2728 0 1 610
box -4 -6 68 206
use OAI22X1  _1371_
timestamp 1591632351
transform -1 0 2808 0 1 610
box -4 -6 84 206
use NOR2X1  _1369_
timestamp 1591632351
transform 1 0 2808 0 1 610
box -4 -6 52 206
use DFFPOSX1  _1507_
timestamp 1591632351
transform 1 0 2856 0 1 610
box -4 -6 196 206
use MUX2X1  _851_
timestamp 1591632351
transform -1 0 3144 0 1 610
box -4 -6 100 206
use MUX2X1  _1368_
timestamp 1591632351
transform -1 0 3240 0 1 610
box -4 -6 100 206
use OAI21X1  _927_
timestamp 1591632351
transform 1 0 3240 0 1 610
box -4 -6 68 206
use NAND2X1  _926_
timestamp 1591632351
transform -1 0 3352 0 1 610
box -4 -6 52 206
use DFFPOSX1  _1459_
timestamp 1591632351
transform -1 0 3544 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert38
timestamp 1591632351
transform 1 0 3544 0 1 610
box -4 -6 52 206
use NAND2X1  _992_
timestamp 1591632351
transform 1 0 3592 0 1 610
box -4 -6 52 206
use DFFPOSX1  _1504_
timestamp 1591632351
transform -1 0 3832 0 1 610
box -4 -6 196 206
use OAI21X1  _993_
timestamp 1591632351
transform -1 0 3896 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert35
timestamp 1591632351
transform -1 0 3944 0 1 610
box -4 -6 52 206
use DFFPOSX1  _1532_
timestamp 1591632351
transform -1 0 4136 0 1 610
box -4 -6 196 206
use NAND2X1  _1068_
timestamp 1591632351
transform 1 0 4200 0 1 610
box -4 -6 52 206
use FILL  SFILL41360x6100
timestamp 1591632351
transform 1 0 4136 0 1 610
box -4 -6 20 206
use FILL  SFILL41520x6100
timestamp 1591632351
transform 1 0 4152 0 1 610
box -4 -6 20 206
use FILL  SFILL41680x6100
timestamp 1591632351
transform 1 0 4168 0 1 610
box -4 -6 20 206
use FILL  SFILL41840x6100
timestamp 1591632351
transform 1 0 4184 0 1 610
box -4 -6 20 206
use OAI21X1  _1069_
timestamp 1591632351
transform -1 0 4312 0 1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert13
timestamp 1591632351
transform -1 0 4456 0 1 610
box -4 -6 148 206
use INVX1  _1045_
timestamp 1591632351
transform 1 0 4456 0 1 610
box -4 -6 36 206
use OAI21X1  _1047_
timestamp 1591632351
transform 1 0 4488 0 1 610
box -4 -6 68 206
use DFFPOSX1  _1510_
timestamp 1591632351
transform -1 0 4744 0 1 610
box -4 -6 196 206
use INVX1  _1088_
timestamp 1591632351
transform 1 0 4744 0 1 610
box -4 -6 36 206
use OAI21X1  _1091_
timestamp 1591632351
transform 1 0 4776 0 1 610
box -4 -6 68 206
use NAND3X1  _1126_
timestamp 1591632351
transform -1 0 4904 0 1 610
box -4 -6 68 206
use INVX1  _1033_
timestamp 1591632351
transform 1 0 4904 0 1 610
box -4 -6 36 206
use OAI21X1  _1035_
timestamp 1591632351
transform 1 0 4936 0 1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert14
timestamp 1591632351
transform -1 0 5144 0 1 610
box -4 -6 148 206
use BUFX2  _1424_
timestamp 1591632351
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use BUFX2  _1414_
timestamp 1591632351
transform -1 0 104 0 -1 1010
box -4 -6 52 206
use OAI21X1  _1331_
timestamp 1591632351
transform -1 0 168 0 -1 1010
box -4 -6 68 206
use OAI21X1  _1337_
timestamp 1591632351
transform -1 0 232 0 -1 1010
box -4 -6 68 206
use OAI21X1  _1211_
timestamp 1591632351
transform 1 0 232 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1558_
timestamp 1591632351
transform -1 0 488 0 -1 1010
box -4 -6 196 206
use OAI21X1  _1217_
timestamp 1591632351
transform -1 0 552 0 -1 1010
box -4 -6 68 206
use NOR2X1  _1210_
timestamp 1591632351
transform 1 0 552 0 -1 1010
box -4 -6 52 206
use NOR2X1  _1282_
timestamp 1591632351
transform 1 0 600 0 -1 1010
box -4 -6 52 206
use NOR2X1  _691_
timestamp 1591632351
transform 1 0 648 0 -1 1010
box -4 -6 52 206
use NOR2X1  _1354_
timestamp 1591632351
transform 1 0 696 0 -1 1010
box -4 -6 52 206
use OAI21X1  _1216_
timestamp 1591632351
transform -1 0 808 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1430_
timestamp 1591632351
transform 1 0 808 0 -1 1010
box -4 -6 196 206
use OAI21X1  _939_
timestamp 1591632351
transform 1 0 1000 0 -1 1010
box -4 -6 68 206
use OAI21X1  _938_
timestamp 1591632351
transform -1 0 1192 0 -1 1010
box -4 -6 68 206
use OAI21X1  _736_
timestamp 1591632351
transform -1 0 1256 0 -1 1010
box -4 -6 68 206
use FILL  SFILL10640x8100
timestamp 1591632351
transform -1 0 1080 0 -1 1010
box -4 -6 20 206
use FILL  SFILL10800x8100
timestamp 1591632351
transform -1 0 1096 0 -1 1010
box -4 -6 20 206
use FILL  SFILL10960x8100
timestamp 1591632351
transform -1 0 1112 0 -1 1010
box -4 -6 20 206
use FILL  SFILL11120x8100
timestamp 1591632351
transform -1 0 1128 0 -1 1010
box -4 -6 20 206
use OAI21X1  _735_
timestamp 1591632351
transform -1 0 1320 0 -1 1010
box -4 -6 68 206
use NOR2X1  _801_
timestamp 1591632351
transform 1 0 1320 0 -1 1010
box -4 -6 52 206
use OAI22X1  _1209_
timestamp 1591632351
transform -1 0 1448 0 -1 1010
box -4 -6 84 206
use OAI21X1  _1208_
timestamp 1591632351
transform -1 0 1512 0 -1 1010
box -4 -6 68 206
use OAI22X1  _690_
timestamp 1591632351
transform -1 0 1592 0 -1 1010
box -4 -6 84 206
use OAI21X1  _689_
timestamp 1591632351
transform -1 0 1656 0 -1 1010
box -4 -6 68 206
use NOR2X1  _837_
timestamp 1591632351
transform 1 0 1656 0 -1 1010
box -4 -6 52 206
use OAI21X1  _835_
timestamp 1591632351
transform -1 0 1768 0 -1 1010
box -4 -6 68 206
use OAI22X1  _836_
timestamp 1591632351
transform 1 0 1768 0 -1 1010
box -4 -6 84 206
use OAI22X1  _1353_
timestamp 1591632351
transform -1 0 1928 0 -1 1010
box -4 -6 84 206
use OAI21X1  _1352_
timestamp 1591632351
transform -1 0 1992 0 -1 1010
box -4 -6 68 206
use OAI21X1  _962_
timestamp 1591632351
transform -1 0 2056 0 -1 1010
box -4 -6 68 206
use MUX2X1  _1350_
timestamp 1591632351
transform 1 0 2056 0 -1 1010
box -4 -6 100 206
use MUX2X1  _833_
timestamp 1591632351
transform -1 0 2248 0 -1 1010
box -4 -6 100 206
use NOR2X1  _765_
timestamp 1591632351
transform 1 0 2248 0 -1 1010
box -4 -6 52 206
use NAND2X1  _1080_
timestamp 1591632351
transform 1 0 2296 0 -1 1010
box -4 -6 52 206
use OAI21X1  _1081_
timestamp 1591632351
transform -1 0 2408 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1538_
timestamp 1591632351
transform -1 0 2600 0 -1 1010
box -4 -6 196 206
use FILL  SFILL26000x8100
timestamp 1591632351
transform -1 0 2616 0 -1 1010
box -4 -6 20 206
use NAND2X1  _908_
timestamp 1591632351
transform -1 0 2712 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert48
timestamp 1591632351
transform -1 0 2760 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert74
timestamp 1591632351
transform -1 0 2808 0 -1 1010
box -4 -6 52 206
use OAI22X1  _782_
timestamp 1591632351
transform -1 0 2888 0 -1 1010
box -4 -6 84 206
use FILL  SFILL26160x8100
timestamp 1591632351
transform -1 0 2632 0 -1 1010
box -4 -6 20 206
use FILL  SFILL26320x8100
timestamp 1591632351
transform -1 0 2648 0 -1 1010
box -4 -6 20 206
use FILL  SFILL26480x8100
timestamp 1591632351
transform -1 0 2664 0 -1 1010
box -4 -6 20 206
use BUFX2  BUFX2_insert81
timestamp 1591632351
transform 1 0 2888 0 -1 1010
box -4 -6 52 206
use OAI21X1  _781_
timestamp 1591632351
transform 1 0 2936 0 -1 1010
box -4 -6 68 206
use OAI22X1  _764_
timestamp 1591632351
transform -1 0 3080 0 -1 1010
box -4 -6 84 206
use OAI21X1  _763_
timestamp 1591632351
transform -1 0 3144 0 -1 1010
box -4 -6 68 206
use NOR2X1  _1279_
timestamp 1591632351
transform -1 0 3192 0 -1 1010
box -4 -6 52 206
use OAI22X1  _1281_
timestamp 1591632351
transform 1 0 3192 0 -1 1010
box -4 -6 84 206
use BUFX2  BUFX2_insert28
timestamp 1591632351
transform 1 0 3272 0 -1 1010
box -4 -6 52 206
use MUX2X1  _1278_
timestamp 1591632351
transform 1 0 3320 0 -1 1010
box -4 -6 100 206
use MUX2X1  _761_
timestamp 1591632351
transform -1 0 3512 0 -1 1010
box -4 -6 100 206
use NOR2X1  _798_
timestamp 1591632351
transform -1 0 3560 0 -1 1010
box -4 -6 52 206
use OAI22X1  _800_
timestamp 1591632351
transform 1 0 3560 0 -1 1010
box -4 -6 84 206
use OAI21X1  _799_
timestamp 1591632351
transform -1 0 3704 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert21
timestamp 1591632351
transform -1 0 3752 0 -1 1010
box -4 -6 52 206
use OAI21X1  _964_
timestamp 1591632351
transform 1 0 3752 0 -1 1010
box -4 -6 68 206
use OAI21X1  _965_
timestamp 1591632351
transform -1 0 3880 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1443_
timestamp 1591632351
transform -1 0 4072 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  _1490_
timestamp 1591632351
transform -1 0 4328 0 -1 1010
box -4 -6 196 206
use FILL  SFILL40720x8100
timestamp 1591632351
transform -1 0 4088 0 -1 1010
box -4 -6 20 206
use FILL  SFILL40880x8100
timestamp 1591632351
transform -1 0 4104 0 -1 1010
box -4 -6 20 206
use FILL  SFILL41040x8100
timestamp 1591632351
transform -1 0 4120 0 -1 1010
box -4 -6 20 206
use FILL  SFILL41200x8100
timestamp 1591632351
transform -1 0 4136 0 -1 1010
box -4 -6 20 206
use OAI21X1  _1163_
timestamp 1591632351
transform -1 0 4392 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1516_
timestamp 1591632351
transform -1 0 4584 0 -1 1010
box -4 -6 196 206
use INVX1  _1107_
timestamp 1591632351
transform 1 0 4584 0 -1 1010
box -4 -6 36 206
use OAI21X1  _1109_
timestamp 1591632351
transform 1 0 4616 0 -1 1010
box -4 -6 68 206
use DFFPOSX1  _1522_
timestamp 1591632351
transform -1 0 4872 0 -1 1010
box -4 -6 196 206
use OAI21X1  _1127_
timestamp 1591632351
transform -1 0 4936 0 -1 1010
box -4 -6 68 206
use INVX1  _1125_
timestamp 1591632351
transform 1 0 4936 0 -1 1010
box -4 -6 36 206
use NAND3X1  _1108_
timestamp 1591632351
transform 1 0 4968 0 -1 1010
box -4 -6 68 206
use NAND3X1  _1090_
timestamp 1591632351
transform -1 0 5096 0 -1 1010
box -4 -6 68 206
use FILL  FILL49040x8100
timestamp 1591632351
transform -1 0 5112 0 -1 1010
box -4 -6 20 206
use FILL  FILL49200x8100
timestamp 1591632351
transform -1 0 5128 0 -1 1010
box -4 -6 20 206
use FILL  FILL49360x8100
timestamp 1591632351
transform -1 0 5144 0 -1 1010
box -4 -6 20 206
use BUFX2  _1398_
timestamp 1591632351
transform -1 0 56 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _1568_
timestamp 1591632351
transform -1 0 248 0 1 1010
box -4 -6 196 206
use OAI21X1  _693_
timestamp 1591632351
transform 1 0 248 0 1 1010
box -4 -6 68 206
use NOR2X1  _698_
timestamp 1591632351
transform -1 0 360 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _1574_
timestamp 1591632351
transform -1 0 552 0 1 1010
box -4 -6 196 206
use OAI21X1  _700_
timestamp 1591632351
transform -1 0 616 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _1446_
timestamp 1591632351
transform 1 0 616 0 1 1010
box -4 -6 196 206
use NAND2X1  _887_
timestamp 1591632351
transform 1 0 808 0 1 1010
box -4 -6 52 206
use OAI21X1  _888_
timestamp 1591632351
transform -1 0 920 0 1 1010
box -4 -6 68 206
use MUX2X1  _1212_
timestamp 1591632351
transform -1 0 1016 0 1 1010
box -4 -6 100 206
use OAI22X1  _1215_
timestamp 1591632351
transform -1 0 1160 0 1 1010
box -4 -6 84 206
use OAI21X1  _1214_
timestamp 1591632351
transform -1 0 1224 0 1 1010
box -4 -6 68 206
use FILL  SFILL10160x10100
timestamp 1591632351
transform 1 0 1016 0 1 1010
box -4 -6 20 206
use FILL  SFILL10320x10100
timestamp 1591632351
transform 1 0 1032 0 1 1010
box -4 -6 20 206
use FILL  SFILL10480x10100
timestamp 1591632351
transform 1 0 1048 0 1 1010
box -4 -6 20 206
use FILL  SFILL10640x10100
timestamp 1591632351
transform 1 0 1064 0 1 1010
box -4 -6 20 206
use MUX2X1  _694_
timestamp 1591632351
transform 1 0 1224 0 1 1010
box -4 -6 100 206
use OAI21X1  _696_
timestamp 1591632351
transform 1 0 1320 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _1478_
timestamp 1591632351
transform -1 0 1576 0 1 1010
box -4 -6 196 206
use NAND2X1  _1138_
timestamp 1591632351
transform 1 0 1576 0 1 1010
box -4 -6 52 206
use OAI21X1  _1139_
timestamp 1591632351
transform -1 0 1688 0 1 1010
box -4 -6 68 206
use NOR2X1  _1207_
timestamp 1591632351
transform -1 0 1736 0 1 1010
box -4 -6 52 206
use NOR2X1  _688_
timestamp 1591632351
transform -1 0 1784 0 1 1010
box -4 -6 52 206
use NOR2X1  _834_
timestamp 1591632351
transform -1 0 1832 0 1 1010
box -4 -6 52 206
use NOR2X1  _1366_
timestamp 1591632351
transform 1 0 1832 0 1 1010
box -4 -6 52 206
use NOR2X1  _1351_
timestamp 1591632351
transform 1 0 1880 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _1474_
timestamp 1591632351
transform -1 0 2120 0 1 1010
box -4 -6 196 206
use OAI21X1  _1197_
timestamp 1591632351
transform -1 0 2184 0 1 1010
box -4 -6 68 206
use NOR2X1  _861_
timestamp 1591632351
transform 1 0 2184 0 1 1010
box -4 -6 52 206
use NOR2X1  _813_
timestamp 1591632351
transform 1 0 2232 0 1 1010
box -4 -6 52 206
use NOR2X1  _849_
timestamp 1591632351
transform 1 0 2280 0 1 1010
box -4 -6 52 206
use NOR2X1  _1378_
timestamp 1591632351
transform -1 0 2376 0 1 1010
box -4 -6 52 206
use NOR2X1  _1318_
timestamp 1591632351
transform 1 0 2376 0 1 1010
box -4 -6 52 206
use OAI21X1  _909_
timestamp 1591632351
transform 1 0 2424 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _1453_
timestamp 1591632351
transform 1 0 2552 0 1 1010
box -4 -6 196 206
use FILL  SFILL24880x10100
timestamp 1591632351
transform 1 0 2488 0 1 1010
box -4 -6 20 206
use FILL  SFILL25040x10100
timestamp 1591632351
transform 1 0 2504 0 1 1010
box -4 -6 20 206
use FILL  SFILL25200x10100
timestamp 1591632351
transform 1 0 2520 0 1 1010
box -4 -6 20 206
use FILL  SFILL25360x10100
timestamp 1591632351
transform 1 0 2536 0 1 1010
box -4 -6 20 206
use BUFX2  BUFX2_insert49
timestamp 1591632351
transform 1 0 2744 0 1 1010
box -4 -6 52 206
use MUX2X1  _779_
timestamp 1591632351
transform -1 0 2888 0 1 1010
box -4 -6 100 206
use MUX2X1  _1296_
timestamp 1591632351
transform 1 0 2888 0 1 1010
box -4 -6 100 206
use OAI22X1  _1299_
timestamp 1591632351
transform -1 0 3064 0 1 1010
box -4 -6 84 206
use OAI21X1  _1298_
timestamp 1591632351
transform 1 0 3064 0 1 1010
box -4 -6 68 206
use NOR2X1  _762_
timestamp 1591632351
transform -1 0 3176 0 1 1010
box -4 -6 52 206
use OAI21X1  _1280_
timestamp 1591632351
transform 1 0 3176 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert30
timestamp 1591632351
transform -1 0 3288 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert42
timestamp 1591632351
transform 1 0 3288 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _1476_
timestamp 1591632351
transform -1 0 3528 0 1 1010
box -4 -6 196 206
use OAI21X1  _1201_
timestamp 1591632351
transform 1 0 3528 0 1 1010
box -4 -6 68 206
use MUX2X1  _797_
timestamp 1591632351
transform 1 0 3592 0 1 1010
box -4 -6 100 206
use MUX2X1  _1314_
timestamp 1591632351
transform 1 0 3688 0 1 1010
box -4 -6 100 206
use DFFPOSX1  _1468_
timestamp 1591632351
transform -1 0 3976 0 1 1010
box -4 -6 196 206
use OAI21X1  _1185_
timestamp 1591632351
transform -1 0 4040 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _1471_
timestamp 1591632351
transform -1 0 4296 0 1 1010
box -4 -6 196 206
use FILL  SFILL40400x10100
timestamp 1591632351
transform 1 0 4040 0 1 1010
box -4 -6 20 206
use FILL  SFILL40560x10100
timestamp 1591632351
transform 1 0 4056 0 1 1010
box -4 -6 20 206
use FILL  SFILL40720x10100
timestamp 1591632351
transform 1 0 4072 0 1 1010
box -4 -6 20 206
use FILL  SFILL40880x10100
timestamp 1591632351
transform 1 0 4088 0 1 1010
box -4 -6 20 206
use NAND2X1  _1162_
timestamp 1591632351
transform 1 0 4296 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _1484_
timestamp 1591632351
transform -1 0 4536 0 1 1010
box -4 -6 196 206
use NAND2X1  _1150_
timestamp 1591632351
transform 1 0 4536 0 1 1010
box -4 -6 52 206
use OAI21X1  _1151_
timestamp 1591632351
transform -1 0 4648 0 1 1010
box -4 -6 68 206
use INVX2  _913_
timestamp 1591632351
transform -1 0 4680 0 1 1010
box -4 -6 36 206
use INVX2  _881_
timestamp 1591632351
transform -1 0 4712 0 1 1010
box -4 -6 36 206
use DFFPOSX1  _1519_
timestamp 1591632351
transform -1 0 4904 0 1 1010
box -4 -6 196 206
use INVX1  _1116_
timestamp 1591632351
transform 1 0 4904 0 1 1010
box -4 -6 36 206
use OAI21X1  _1118_
timestamp 1591632351
transform 1 0 4936 0 1 1010
box -4 -6 68 206
use NAND3X1  _1120_
timestamp 1591632351
transform 1 0 5000 0 1 1010
box -4 -6 68 206
use NAND3X1  _1117_
timestamp 1591632351
transform 1 0 5064 0 1 1010
box -4 -6 68 206
use FILL  FILL49360x10100
timestamp 1591632351
transform 1 0 5128 0 1 1010
box -4 -6 20 206
use BUFX2  _1421_
timestamp 1591632351
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use BUFX2  _1417_
timestamp 1591632351
transform -1 0 104 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _1565_
timestamp 1591632351
transform -1 0 296 0 -1 1410
box -4 -6 196 206
use OAI21X1  _1295_
timestamp 1591632351
transform -1 0 360 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1247_
timestamp 1591632351
transform 1 0 360 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _1561_
timestamp 1591632351
transform -1 0 616 0 -1 1410
box -4 -6 196 206
use OAI21X1  _1301_
timestamp 1591632351
transform -1 0 680 0 -1 1410
box -4 -6 68 206
use INVX4  _685_
timestamp 1591632351
transform 1 0 680 0 -1 1410
box -4 -6 52 206
use OAI21X1  _699_
timestamp 1591632351
transform -1 0 792 0 -1 1410
box -4 -6 68 206
use NOR2X1  _1330_
timestamp 1591632351
transform 1 0 792 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1300_
timestamp 1591632351
transform -1 0 904 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1253_
timestamp 1591632351
transform -1 0 968 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1252_
timestamp 1591632351
transform 1 0 968 0 -1 1410
box -4 -6 68 206
use MUX2X1  _1248_
timestamp 1591632351
transform 1 0 1096 0 -1 1410
box -4 -6 100 206
use OAI22X1  _1251_
timestamp 1591632351
transform -1 0 1272 0 -1 1410
box -4 -6 84 206
use FILL  SFILL10320x12100
timestamp 1591632351
transform -1 0 1048 0 -1 1410
box -4 -6 20 206
use FILL  SFILL10480x12100
timestamp 1591632351
transform -1 0 1064 0 -1 1410
box -4 -6 20 206
use FILL  SFILL10640x12100
timestamp 1591632351
transform -1 0 1080 0 -1 1410
box -4 -6 20 206
use FILL  SFILL10800x12100
timestamp 1591632351
transform -1 0 1096 0 -1 1410
box -4 -6 20 206
use OAI21X1  _1250_
timestamp 1591632351
transform -1 0 1336 0 -1 1410
box -4 -6 68 206
use OAI22X1  _697_
timestamp 1591632351
transform -1 0 1416 0 -1 1410
box -4 -6 84 206
use OAI22X1  _734_
timestamp 1591632351
transform -1 0 1496 0 -1 1410
box -4 -6 84 206
use OAI21X1  _733_
timestamp 1591632351
transform 1 0 1496 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert33
timestamp 1591632351
transform -1 0 1608 0 -1 1410
box -4 -6 52 206
use NOR2X1  _732_
timestamp 1591632351
transform -1 0 1656 0 -1 1410
box -4 -6 52 206
use NOR2X1  _1249_
timestamp 1591632351
transform 1 0 1656 0 -1 1410
box -4 -6 52 206
use NOR2X1  _695_
timestamp 1591632351
transform -1 0 1752 0 -1 1410
box -4 -6 52 206
use NOR2X1  _1213_
timestamp 1591632351
transform -1 0 1800 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert79
timestamp 1591632351
transform -1 0 1848 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert46
timestamp 1591632351
transform -1 0 1896 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert116
timestamp 1591632351
transform -1 0 1944 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert113
timestamp 1591632351
transform -1 0 1992 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1196_
timestamp 1591632351
transform 1 0 1992 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1172_
timestamp 1591632351
transform 1 0 2056 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1173_
timestamp 1591632351
transform -1 0 2184 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _1462_
timestamp 1591632351
transform -1 0 2376 0 -1 1410
box -4 -6 196 206
use BUFX2  BUFX2_insert53
timestamp 1591632351
transform 1 0 2376 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert36
timestamp 1591632351
transform -1 0 2472 0 -1 1410
box -4 -6 52 206
use OAI21X1  _952_
timestamp 1591632351
transform 1 0 2472 0 -1 1410
box -4 -6 68 206
use OAI21X1  _953_
timestamp 1591632351
transform -1 0 2664 0 -1 1410
box -4 -6 68 206
use FILL  SFILL25360x12100
timestamp 1591632351
transform -1 0 2552 0 -1 1410
box -4 -6 20 206
use FILL  SFILL25520x12100
timestamp 1591632351
transform -1 0 2568 0 -1 1410
box -4 -6 20 206
use FILL  SFILL25680x12100
timestamp 1591632351
transform -1 0 2584 0 -1 1410
box -4 -6 20 206
use FILL  SFILL25840x12100
timestamp 1591632351
transform -1 0 2600 0 -1 1410
box -4 -6 20 206
use BUFX2  BUFX2_insert111
timestamp 1591632351
transform 1 0 2664 0 -1 1410
box -4 -6 52 206
use INVX8  _687_
timestamp 1591632351
transform 1 0 2712 0 -1 1410
box -4 -6 84 206
use BUFX2  BUFX2_insert77
timestamp 1591632351
transform 1 0 2792 0 -1 1410
box -4 -6 52 206
use NOR2X1  _780_
timestamp 1591632351
transform -1 0 2888 0 -1 1410
box -4 -6 52 206
use NOR2X1  _1297_
timestamp 1591632351
transform -1 0 2936 0 -1 1410
box -4 -6 52 206
use OAI22X1  _1329_
timestamp 1591632351
transform -1 0 3016 0 -1 1410
box -4 -6 84 206
use NOR2X1  _1327_
timestamp 1591632351
transform -1 0 3064 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1328_
timestamp 1591632351
transform -1 0 3128 0 -1 1410
box -4 -6 68 206
use NOR2X1  _810_
timestamp 1591632351
transform 1 0 3128 0 -1 1410
box -4 -6 52 206
use OAI22X1  _812_
timestamp 1591632351
transform 1 0 3176 0 -1 1410
box -4 -6 84 206
use OAI21X1  _811_
timestamp 1591632351
transform -1 0 3320 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert87
timestamp 1591632351
transform 1 0 3320 0 -1 1410
box -4 -6 52 206
use OAI22X1  _1317_
timestamp 1591632351
transform -1 0 3448 0 -1 1410
box -4 -6 84 206
use NOR2X1  _1315_
timestamp 1591632351
transform -1 0 3496 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1316_
timestamp 1591632351
transform -1 0 3560 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1200_
timestamp 1591632351
transform -1 0 3624 0 -1 1410
box -4 -6 68 206
use MUX2X1  _809_
timestamp 1591632351
transform 1 0 3624 0 -1 1410
box -4 -6 100 206
use MUX2X1  _1326_
timestamp 1591632351
transform 1 0 3720 0 -1 1410
box -4 -6 100 206
use BUFX2  BUFX2_insert52
timestamp 1591632351
transform -1 0 3864 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1184_
timestamp 1591632351
transform -1 0 3928 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1190_
timestamp 1591632351
transform 1 0 3928 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1191_
timestamp 1591632351
transform -1 0 4056 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _1535_
timestamp 1591632351
transform -1 0 4312 0 -1 1410
box -4 -6 196 206
use FILL  SFILL40560x12100
timestamp 1591632351
transform -1 0 4072 0 -1 1410
box -4 -6 20 206
use FILL  SFILL40720x12100
timestamp 1591632351
transform -1 0 4088 0 -1 1410
box -4 -6 20 206
use FILL  SFILL40880x12100
timestamp 1591632351
transform -1 0 4104 0 -1 1410
box -4 -6 20 206
use FILL  SFILL41040x12100
timestamp 1591632351
transform -1 0 4120 0 -1 1410
box -4 -6 20 206
use NAND2X1  _1074_
timestamp 1591632351
transform -1 0 4360 0 -1 1410
box -4 -6 52 206
use OAI21X1  _1075_
timestamp 1591632351
transform -1 0 4424 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1157_
timestamp 1591632351
transform 1 0 4424 0 -1 1410
box -4 -6 68 206
use NAND2X1  _1156_
timestamp 1591632351
transform -1 0 4536 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _1487_
timestamp 1591632351
transform -1 0 4728 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _1520_
timestamp 1591632351
transform -1 0 4920 0 -1 1410
box -4 -6 196 206
use INVX1  _1119_
timestamp 1591632351
transform 1 0 4920 0 -1 1410
box -4 -6 36 206
use OAI21X1  _1121_
timestamp 1591632351
transform 1 0 4952 0 -1 1410
box -4 -6 68 206
use OAI21X1  _1008_
timestamp 1591632351
transform 1 0 5016 0 -1 1410
box -4 -6 68 206
use NAND3X1  _1007_
timestamp 1591632351
transform 1 0 5080 0 -1 1410
box -4 -6 68 206
use BUFX2  _1399_
timestamp 1591632351
transform -1 0 56 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert106
timestamp 1591632351
transform 1 0 56 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert103
timestamp 1591632351
transform 1 0 104 0 1 1410
box -4 -6 52 206
use OAI21X1  _706_
timestamp 1591632351
transform 1 0 152 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _1575_
timestamp 1591632351
transform -1 0 408 0 1 1410
box -4 -6 196 206
use DFFPOSX1  _1481_
timestamp 1591632351
transform 1 0 408 0 1 1410
box -4 -6 196 206
use DFFPOSX1  _1497_
timestamp 1591632351
transform 1 0 600 0 1 1410
box -4 -6 196 206
use BUFX2  BUFX2_insert1
timestamp 1591632351
transform -1 0 840 0 1 1410
box -4 -6 52 206
use NAND2X1  _978_
timestamp 1591632351
transform 1 0 840 0 1 1410
box -4 -6 52 206
use OAI21X1  _979_
timestamp 1591632351
transform -1 0 952 0 1 1410
box -4 -6 68 206
use OAI21X1  _945_
timestamp 1591632351
transform 1 0 952 0 1 1410
box -4 -6 68 206
use OAI21X1  _944_
timestamp 1591632351
transform -1 0 1080 0 1 1410
box -4 -6 68 206
use MUX2X1  _731_
timestamp 1591632351
transform -1 0 1240 0 1 1410
box -4 -6 100 206
use FILL  SFILL10800x14100
timestamp 1591632351
transform 1 0 1080 0 1 1410
box -4 -6 20 206
use FILL  SFILL10960x14100
timestamp 1591632351
transform 1 0 1096 0 1 1410
box -4 -6 20 206
use FILL  SFILL11120x14100
timestamp 1591632351
transform 1 0 1112 0 1 1410
box -4 -6 20 206
use FILL  SFILL11280x14100
timestamp 1591632351
transform 1 0 1128 0 1 1410
box -4 -6 20 206
use NOR2X1  _729_
timestamp 1591632351
transform 1 0 1240 0 1 1410
box -4 -6 52 206
use NOR2X1  _1246_
timestamp 1591632351
transform 1 0 1288 0 1 1410
box -4 -6 52 206
use OAI21X1  _1145_
timestamp 1591632351
transform 1 0 1336 0 1 1410
box -4 -6 68 206
use NAND2X1  _1144_
timestamp 1591632351
transform -1 0 1448 0 1 1410
box -4 -6 52 206
use OAI21X1  _727_
timestamp 1591632351
transform 1 0 1448 0 1 1410
box -4 -6 68 206
use OAI22X1  _728_
timestamp 1591632351
transform 1 0 1512 0 1 1410
box -4 -6 84 206
use NOR2X1  _777_
timestamp 1591632351
transform 1 0 1592 0 1 1410
box -4 -6 52 206
use NOR2X1  _726_
timestamp 1591632351
transform -1 0 1688 0 1 1410
box -4 -6 52 206
use OAI21X1  _1244_
timestamp 1591632351
transform 1 0 1688 0 1 1410
box -4 -6 68 206
use OAI22X1  _1245_
timestamp 1591632351
transform 1 0 1752 0 1 1410
box -4 -6 84 206
use NOR2X1  _1243_
timestamp 1591632351
transform 1 0 1832 0 1 1410
box -4 -6 52 206
use OAI21X1  _1178_
timestamp 1591632351
transform -1 0 1944 0 1 1410
box -4 -6 68 206
use OAI21X1  _1179_
timestamp 1591632351
transform -1 0 2008 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _1465_
timestamp 1591632351
transform -1 0 2200 0 1 1410
box -4 -6 196 206
use BUFX2  BUFX2_insert115
timestamp 1591632351
transform 1 0 2200 0 1 1410
box -4 -6 52 206
use NOR2X1  _1294_
timestamp 1591632351
transform 1 0 2248 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert26
timestamp 1591632351
transform 1 0 2296 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _1437_
timestamp 1591632351
transform 1 0 2344 0 1 1410
box -4 -6 196 206
use BUFX2  BUFX2_insert112
timestamp 1591632351
transform -1 0 2648 0 1 1410
box -4 -6 52 206
use FILL  SFILL25360x14100
timestamp 1591632351
transform 1 0 2536 0 1 1410
box -4 -6 20 206
use FILL  SFILL25520x14100
timestamp 1591632351
transform 1 0 2552 0 1 1410
box -4 -6 20 206
use FILL  SFILL25680x14100
timestamp 1591632351
transform 1 0 2568 0 1 1410
box -4 -6 20 206
use FILL  SFILL25840x14100
timestamp 1591632351
transform 1 0 2584 0 1 1410
box -4 -6 20 206
use OAI21X1  _1186_
timestamp 1591632351
transform 1 0 2648 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert85
timestamp 1591632351
transform -1 0 2760 0 1 1410
box -4 -6 52 206
use OAI21X1  _1187_
timestamp 1591632351
transform -1 0 2824 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert122
timestamp 1591632351
transform 1 0 2824 0 1 1410
box -4 -6 52 206
use NOR2X1  _846_
timestamp 1591632351
transform -1 0 2920 0 1 1410
box -4 -6 52 206
use OAI22X1  _848_
timestamp 1591632351
transform 1 0 2920 0 1 1410
box -4 -6 84 206
use OAI21X1  _847_
timestamp 1591632351
transform -1 0 3064 0 1 1410
box -4 -6 68 206
use OAI21X1  _1364_
timestamp 1591632351
transform -1 0 3128 0 1 1410
box -4 -6 68 206
use OAI22X1  _1365_
timestamp 1591632351
transform 1 0 3128 0 1 1410
box -4 -6 84 206
use NOR2X1  _858_
timestamp 1591632351
transform -1 0 3256 0 1 1410
box -4 -6 52 206
use OAI22X1  _860_
timestamp 1591632351
transform 1 0 3256 0 1 1410
box -4 -6 84 206
use OAI21X1  _859_
timestamp 1591632351
transform -1 0 3400 0 1 1410
box -4 -6 68 206
use NOR2X1  _1375_
timestamp 1591632351
transform 1 0 3400 0 1 1410
box -4 -6 52 206
use OAI22X1  _1377_
timestamp 1591632351
transform 1 0 3448 0 1 1410
box -4 -6 84 206
use OAI21X1  _1376_
timestamp 1591632351
transform -1 0 3592 0 1 1410
box -4 -6 68 206
use OAI21X1  _1192_
timestamp 1591632351
transform 1 0 3592 0 1 1410
box -4 -6 68 206
use NAND2X1  _1166_
timestamp 1591632351
transform 1 0 3656 0 1 1410
box -4 -6 52 206
use OAI21X1  _1167_
timestamp 1591632351
transform -1 0 3768 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _1492_
timestamp 1591632351
transform -1 0 3960 0 1 1410
box -4 -6 196 206
use OAI21X1  _1193_
timestamp 1591632351
transform -1 0 4024 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _1472_
timestamp 1591632351
transform -1 0 4280 0 1 1410
box -4 -6 196 206
use FILL  SFILL40240x14100
timestamp 1591632351
transform 1 0 4024 0 1 1410
box -4 -6 20 206
use FILL  SFILL40400x14100
timestamp 1591632351
transform 1 0 4040 0 1 1410
box -4 -6 20 206
use FILL  SFILL40560x14100
timestamp 1591632351
transform 1 0 4056 0 1 1410
box -4 -6 20 206
use FILL  SFILL40720x14100
timestamp 1591632351
transform 1 0 4072 0 1 1410
box -4 -6 20 206
use DFFPOSX1  _1536_
timestamp 1591632351
transform -1 0 4472 0 1 1410
box -4 -6 196 206
use NAND2X1  _1076_
timestamp 1591632351
transform 1 0 4472 0 1 1410
box -4 -6 52 206
use OAI21X1  _1077_
timestamp 1591632351
transform -1 0 4584 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _1556_
timestamp 1591632351
transform -1 0 4776 0 1 1410
box -4 -6 196 206
use OAI21X1  _1050_
timestamp 1591632351
transform -1 0 4840 0 1 1410
box -4 -6 68 206
use INVX1  _1048_
timestamp 1591632351
transform -1 0 4872 0 1 1410
box -4 -6 36 206
use AND2X2  _1006_
timestamp 1591632351
transform 1 0 4872 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _1542_
timestamp 1591632351
transform -1 0 5128 0 1 1410
box -4 -6 196 206
use FILL  FILL49360x14100
timestamp 1591632351
transform 1 0 5128 0 1 1410
box -4 -6 20 206
use INVX8  _692_
timestamp 1591632351
transform -1 0 88 0 -1 1810
box -4 -6 84 206
use NAND2X1  _884_
timestamp 1591632351
transform -1 0 136 0 -1 1810
box -4 -6 52 206
use AND2X2  _935_
timestamp 1591632351
transform 1 0 136 0 -1 1810
box -4 -6 68 206
use NOR2X1  _885_
timestamp 1591632351
transform -1 0 248 0 -1 1810
box -4 -6 52 206
use NAND2X1  _936_
timestamp 1591632351
transform 1 0 248 0 -1 1810
box -4 -6 52 206
use OAI21X1  _712_
timestamp 1591632351
transform -1 0 360 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  _1433_
timestamp 1591632351
transform 1 0 360 0 -1 1810
box -4 -6 196 206
use DFFPOSX1  _1448_
timestamp 1591632351
transform -1 0 744 0 -1 1810
box -4 -6 196 206
use NAND2X1  _893_
timestamp 1591632351
transform 1 0 744 0 -1 1810
box -4 -6 52 206
use OAI21X1  _894_
timestamp 1591632351
transform -1 0 856 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  _1449_
timestamp 1591632351
transform 1 0 856 0 -1 1810
box -4 -6 196 206
use OAI21X1  _897_
timestamp 1591632351
transform 1 0 1112 0 -1 1810
box -4 -6 68 206
use NAND2X1  _896_
timestamp 1591632351
transform -1 0 1224 0 -1 1810
box -4 -6 52 206
use FILL  SFILL10480x16100
timestamp 1591632351
transform -1 0 1064 0 -1 1810
box -4 -6 20 206
use FILL  SFILL10640x16100
timestamp 1591632351
transform -1 0 1080 0 -1 1810
box -4 -6 20 206
use FILL  SFILL10800x16100
timestamp 1591632351
transform -1 0 1096 0 -1 1810
box -4 -6 20 206
use FILL  SFILL10960x16100
timestamp 1591632351
transform -1 0 1112 0 -1 1810
box -4 -6 20 206
use DFFPOSX1  _1496_
timestamp 1591632351
transform -1 0 1416 0 -1 1810
box -4 -6 196 206
use NAND2X1  _976_
timestamp 1591632351
transform 1 0 1416 0 -1 1810
box -4 -6 52 206
use OAI21X1  _977_
timestamp 1591632351
transform -1 0 1528 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert90
timestamp 1591632351
transform -1 0 1576 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _1464_
timestamp 1591632351
transform -1 0 1768 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_insert51
timestamp 1591632351
transform -1 0 1816 0 -1 1810
box -4 -6 52 206
use MUX2X1  _725_
timestamp 1591632351
transform -1 0 1912 0 -1 1810
box -4 -6 100 206
use MUX2X1  _1242_
timestamp 1591632351
transform -1 0 2008 0 -1 1810
box -4 -6 100 206
use BUFX2  BUFX2_insert22
timestamp 1591632351
transform -1 0 2056 0 -1 1810
box -4 -6 52 206
use INVX8  _1206_
timestamp 1591632351
transform 1 0 2056 0 -1 1810
box -4 -6 84 206
use NAND2X1  _1062_
timestamp 1591632351
transform 1 0 2136 0 -1 1810
box -4 -6 52 206
use OAI21X1  _1063_
timestamp 1591632351
transform -1 0 2248 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  _1529_
timestamp 1591632351
transform -1 0 2440 0 -1 1810
box -4 -6 196 206
use OAI22X1  _1293_
timestamp 1591632351
transform -1 0 2520 0 -1 1810
box -4 -6 84 206
use NOR2X1  _1291_
timestamp 1591632351
transform -1 0 2568 0 -1 1810
box -4 -6 52 206
use FILL  SFILL25680x16100
timestamp 1591632351
transform -1 0 2584 0 -1 1810
box -4 -6 20 206
use FILL  SFILL25840x16100
timestamp 1591632351
transform -1 0 2600 0 -1 1810
box -4 -6 20 206
use FILL  SFILL26000x16100
timestamp 1591632351
transform -1 0 2616 0 -1 1810
box -4 -6 20 206
use NOR2X1  _774_
timestamp 1591632351
transform 1 0 2632 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _1469_
timestamp 1591632351
transform -1 0 2872 0 -1 1810
box -4 -6 196 206
use FILL  SFILL26160x16100
timestamp 1591632351
transform -1 0 2632 0 -1 1810
box -4 -6 20 206
use OAI21X1  _1198_
timestamp 1591632351
transform 1 0 2872 0 -1 1810
box -4 -6 68 206
use OAI21X1  _1199_
timestamp 1591632351
transform -1 0 3000 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  _1475_
timestamp 1591632351
transform 1 0 3000 0 -1 1810
box -4 -6 196 206
use NOR2X1  _1363_
timestamp 1591632351
transform 1 0 3192 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert29
timestamp 1591632351
transform -1 0 3288 0 -1 1810
box -4 -6 52 206
use INVX2  _895_
timestamp 1591632351
transform -1 0 3320 0 -1 1810
box -4 -6 36 206
use MUX2X1  _845_
timestamp 1591632351
transform -1 0 3416 0 -1 1810
box -4 -6 100 206
use MUX2X1  _1362_
timestamp 1591632351
transform -1 0 3512 0 -1 1810
box -4 -6 100 206
use MUX2X1  _857_
timestamp 1591632351
transform -1 0 3608 0 -1 1810
box -4 -6 100 206
use MUX2X1  _1374_
timestamp 1591632351
transform -1 0 3704 0 -1 1810
box -4 -6 100 206
use BUFX2  BUFX2_insert84
timestamp 1591632351
transform 1 0 3704 0 -1 1810
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert8
timestamp 1591632351
transform -1 0 3896 0 -1 1810
box -4 -6 148 206
use NAND2X1  _1158_
timestamp 1591632351
transform -1 0 3944 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _1488_
timestamp 1591632351
transform -1 0 4136 0 -1 1810
box -4 -6 196 206
use OAI21X1  _1159_
timestamp 1591632351
transform -1 0 4264 0 -1 1810
box -4 -6 68 206
use FILL  SFILL41360x16100
timestamp 1591632351
transform -1 0 4152 0 -1 1810
box -4 -6 20 206
use FILL  SFILL41520x16100
timestamp 1591632351
transform -1 0 4168 0 -1 1810
box -4 -6 20 206
use FILL  SFILL41680x16100
timestamp 1591632351
transform -1 0 4184 0 -1 1810
box -4 -6 20 206
use FILL  SFILL41840x16100
timestamp 1591632351
transform -1 0 4200 0 -1 1810
box -4 -6 20 206
use NAND2X1  _934_
timestamp 1591632351
transform -1 0 4312 0 -1 1810
box -4 -6 52 206
use INVX1  _883_
timestamp 1591632351
transform -1 0 4344 0 -1 1810
box -4 -6 36 206
use NAND3X1  _886_
timestamp 1591632351
transform -1 0 4408 0 -1 1810
box -4 -6 68 206
use INVX1  _882_
timestamp 1591632351
transform -1 0 4440 0 -1 1810
box -4 -6 36 206
use NOR2X1  _1054_
timestamp 1591632351
transform -1 0 4488 0 -1 1810
box -4 -6 52 206
use NOR2X1  _970_
timestamp 1591632351
transform -1 0 4536 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert18
timestamp 1591632351
transform 1 0 4536 0 -1 1810
box -4 -6 52 206
use NAND3X1  _1046_
timestamp 1591632351
transform 1 0 4584 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert73
timestamp 1591632351
transform 1 0 4648 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert16
timestamp 1591632351
transform 1 0 4696 0 -1 1810
box -4 -6 52 206
use NAND3X1  _1049_
timestamp 1591632351
transform -1 0 4808 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert97
timestamp 1591632351
transform 1 0 4808 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _1545_
timestamp 1591632351
transform -1 0 5048 0 -1 1810
box -4 -6 196 206
use INVX1  _1015_
timestamp 1591632351
transform 1 0 5048 0 -1 1810
box -4 -6 36 206
use OAI21X1  _1017_
timestamp 1591632351
transform 1 0 5080 0 -1 1810
box -4 -6 68 206
use BUFX2  _1400_
timestamp 1591632351
transform -1 0 56 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert109
timestamp 1591632351
transform 1 0 56 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert104
timestamp 1591632351
transform 1 0 104 0 1 1810
box -4 -6 52 206
use OAI21X1  _718_
timestamp 1591632351
transform 1 0 152 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _1576_
timestamp 1591632351
transform -1 0 408 0 1 1810
box -4 -6 196 206
use BUFX2  BUFX2_insert108
timestamp 1591632351
transform 1 0 408 0 1 1810
box -4 -6 52 206
use OAI21X1  _724_
timestamp 1591632351
transform -1 0 520 0 1 1810
box -4 -6 68 206
use OAI21X1  _723_
timestamp 1591632351
transform -1 0 584 0 1 1810
box -4 -6 68 206
use OAI21X1  _711_
timestamp 1591632351
transform -1 0 648 0 1 1810
box -4 -6 68 206
use NOR2X1  _717_
timestamp 1591632351
transform 1 0 648 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _1432_
timestamp 1591632351
transform 1 0 696 0 1 1810
box -4 -6 196 206
use BUFX2  BUFX2_insert2
timestamp 1591632351
transform 1 0 888 0 1 1810
box -4 -6 52 206
use OAI21X1  _943_
timestamp 1591632351
transform 1 0 936 0 1 1810
box -4 -6 68 206
use OAI21X1  _942_
timestamp 1591632351
transform -1 0 1064 0 1 1810
box -4 -6 68 206
use MUX2X1  _1236_
timestamp 1591632351
transform -1 0 1224 0 1 1810
box -4 -6 100 206
use FILL  SFILL10640x18100
timestamp 1591632351
transform 1 0 1064 0 1 1810
box -4 -6 20 206
use FILL  SFILL10800x18100
timestamp 1591632351
transform 1 0 1080 0 1 1810
box -4 -6 20 206
use FILL  SFILL10960x18100
timestamp 1591632351
transform 1 0 1096 0 1 1810
box -4 -6 20 206
use FILL  SFILL11120x18100
timestamp 1591632351
transform 1 0 1112 0 1 1810
box -4 -6 20 206
use MUX2X1  _719_
timestamp 1591632351
transform 1 0 1224 0 1 1810
box -4 -6 100 206
use OAI22X1  _722_
timestamp 1591632351
transform -1 0 1400 0 1 1810
box -4 -6 84 206
use OAI21X1  _721_
timestamp 1591632351
transform 1 0 1400 0 1 1810
box -4 -6 68 206
use OAI22X1  _716_
timestamp 1591632351
transform -1 0 1544 0 1 1810
box -4 -6 84 206
use OAI21X1  _715_
timestamp 1591632351
transform -1 0 1608 0 1 1810
box -4 -6 68 206
use NOR2X1  _714_
timestamp 1591632351
transform -1 0 1656 0 1 1810
box -4 -6 52 206
use NOR2X1  _705_
timestamp 1591632351
transform 1 0 1656 0 1 1810
box -4 -6 52 206
use OAI21X1  _1177_
timestamp 1591632351
transform -1 0 1768 0 1 1810
box -4 -6 68 206
use OAI21X1  _1176_
timestamp 1591632351
transform -1 0 1832 0 1 1810
box -4 -6 68 206
use OAI21X1  _1220_
timestamp 1591632351
transform 1 0 1832 0 1 1810
box -4 -6 68 206
use OAI22X1  _1221_
timestamp 1591632351
transform 1 0 1896 0 1 1810
box -4 -6 84 206
use NOR2X1  _1219_
timestamp 1591632351
transform -1 0 2024 0 1 1810
box -4 -6 52 206
use OAI21X1  _703_
timestamp 1591632351
transform 1 0 2024 0 1 1810
box -4 -6 68 206
use OAI22X1  _704_
timestamp 1591632351
transform 1 0 2088 0 1 1810
box -4 -6 84 206
use NOR2X1  _702_
timestamp 1591632351
transform 1 0 2168 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert44
timestamp 1591632351
transform 1 0 2216 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert55
timestamp 1591632351
transform -1 0 2312 0 1 1810
box -4 -6 52 206
use OAI22X1  _776_
timestamp 1591632351
transform -1 0 2392 0 1 1810
box -4 -6 84 206
use OAI21X1  _775_
timestamp 1591632351
transform -1 0 2456 0 1 1810
box -4 -6 68 206
use OAI21X1  _1292_
timestamp 1591632351
transform -1 0 2520 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert47
timestamp 1591632351
transform -1 0 2568 0 1 1810
box -4 -6 52 206
use FILL  SFILL25680x18100
timestamp 1591632351
transform 1 0 2568 0 1 1810
box -4 -6 20 206
use FILL  SFILL25840x18100
timestamp 1591632351
transform 1 0 2584 0 1 1810
box -4 -6 20 206
use FILL  SFILL26000x18100
timestamp 1591632351
transform 1 0 2600 0 1 1810
box -4 -6 20 206
use NAND2X1  _1152_
timestamp 1591632351
transform -1 0 2680 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _1485_
timestamp 1591632351
transform -1 0 2872 0 1 1810
box -4 -6 196 206
use FILL  SFILL26160x18100
timestamp 1591632351
transform 1 0 2616 0 1 1810
box -4 -6 20 206
use BUFX2  BUFX2_insert82
timestamp 1591632351
transform -1 0 2920 0 1 1810
box -4 -6 52 206
use OAI21X1  _1153_
timestamp 1591632351
transform -1 0 2984 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert57
timestamp 1591632351
transform -1 0 3032 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert88
timestamp 1591632351
transform -1 0 3080 0 1 1810
box -4 -6 52 206
use NAND2X1  _1164_
timestamp 1591632351
transform 1 0 3080 0 1 1810
box -4 -6 52 206
use OAI21X1  _1165_
timestamp 1591632351
transform -1 0 3192 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _1491_
timestamp 1591632351
transform -1 0 3384 0 1 1810
box -4 -6 196 206
use BUFX2  BUFX2_insert63
timestamp 1591632351
transform 1 0 3384 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert58
timestamp 1591632351
transform 1 0 3432 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert83
timestamp 1591632351
transform 1 0 3480 0 1 1810
box -4 -6 52 206
use NAND2X1  _1082_
timestamp 1591632351
transform 1 0 3528 0 1 1810
box -4 -6 52 206
use OAI21X1  _1083_
timestamp 1591632351
transform -1 0 3640 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _1539_
timestamp 1591632351
transform -1 0 3832 0 1 1810
box -4 -6 196 206
use INVX1  _1027_
timestamp 1591632351
transform 1 0 3832 0 1 1810
box -4 -6 36 206
use DFFPOSX1  _1549_
timestamp 1591632351
transform -1 0 4056 0 1 1810
box -4 -6 196 206
use OAI21X1  _1029_
timestamp 1591632351
transform 1 0 4120 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert62
timestamp 1591632351
transform 1 0 4184 0 1 1810
box -4 -6 52 206
use FILL  SFILL40560x18100
timestamp 1591632351
transform 1 0 4056 0 1 1810
box -4 -6 20 206
use FILL  SFILL40720x18100
timestamp 1591632351
transform 1 0 4072 0 1 1810
box -4 -6 20 206
use FILL  SFILL40880x18100
timestamp 1591632351
transform 1 0 4088 0 1 1810
box -4 -6 20 206
use FILL  SFILL41040x18100
timestamp 1591632351
transform 1 0 4104 0 1 1810
box -4 -6 20 206
use BUFX2  BUFX2_insert60
timestamp 1591632351
transform 1 0 4232 0 1 1810
box -4 -6 52 206
use NAND3X1  _1137_
timestamp 1591632351
transform 1 0 4280 0 1 1810
box -4 -6 68 206
use NAND2X1  _1170_
timestamp 1591632351
transform -1 0 4392 0 1 1810
box -4 -6 52 206
use NAND2X1  _1055_
timestamp 1591632351
transform -1 0 4440 0 1 1810
box -4 -6 52 206
use INVX2  _928_
timestamp 1591632351
transform -1 0 4472 0 1 1810
box -4 -6 36 206
use BUFX2  BUFX2_insert99
timestamp 1591632351
transform 1 0 4472 0 1 1810
box -4 -6 52 206
use INVX2  _925_
timestamp 1591632351
transform -1 0 4552 0 1 1810
box -4 -6 36 206
use NAND3X1  _1129_
timestamp 1591632351
transform -1 0 4616 0 1 1810
box -4 -6 68 206
use NAND3X1  _1099_
timestamp 1591632351
transform -1 0 4680 0 1 1810
box -4 -6 68 206
use NAND3X1  _1132_
timestamp 1591632351
transform -1 0 4744 0 1 1810
box -4 -6 68 206
use INVX1  _1128_
timestamp 1591632351
transform 1 0 4744 0 1 1810
box -4 -6 36 206
use OAI21X1  _1130_
timestamp 1591632351
transform 1 0 4776 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _1523_
timestamp 1591632351
transform -1 0 5032 0 1 1810
box -4 -6 196 206
use NAND3X1  _1016_
timestamp 1591632351
transform -1 0 5096 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert70
timestamp 1591632351
transform -1 0 5144 0 1 1810
box -4 -6 52 206
use BUFX2  _1416_
timestamp 1591632351
transform -1 0 56 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert102
timestamp 1591632351
transform 1 0 56 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1235_
timestamp 1591632351
transform 1 0 104 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _1560_
timestamp 1591632351
transform -1 0 360 0 -1 2210
box -4 -6 196 206
use OAI21X1  _1241_
timestamp 1591632351
transform -1 0 424 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert93
timestamp 1591632351
transform 1 0 424 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1240_
timestamp 1591632351
transform -1 0 536 0 -1 2210
box -4 -6 68 206
use NOR2X1  _1222_
timestamp 1591632351
transform -1 0 584 0 -1 2210
box -4 -6 52 206
use NOR2X1  _1234_
timestamp 1591632351
transform 1 0 584 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert67
timestamp 1591632351
transform -1 0 680 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert92
timestamp 1591632351
transform -1 0 728 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _1528_
timestamp 1591632351
transform 1 0 728 0 -1 2210
box -4 -6 196 206
use NAND2X1  _980_
timestamp 1591632351
transform 1 0 920 0 -1 2210
box -4 -6 52 206
use NAND2X1  _1060_
timestamp 1591632351
transform 1 0 968 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1061_
timestamp 1591632351
transform -1 0 1080 0 -1 2210
box -4 -6 68 206
use OAI22X1  _1239_
timestamp 1591632351
transform -1 0 1224 0 -1 2210
box -4 -6 84 206
use FILL  SFILL10800x20100
timestamp 1591632351
transform -1 0 1096 0 -1 2210
box -4 -6 20 206
use FILL  SFILL10960x20100
timestamp 1591632351
transform -1 0 1112 0 -1 2210
box -4 -6 20 206
use FILL  SFILL11120x20100
timestamp 1591632351
transform -1 0 1128 0 -1 2210
box -4 -6 20 206
use FILL  SFILL11280x20100
timestamp 1591632351
transform -1 0 1144 0 -1 2210
box -4 -6 20 206
use OAI21X1  _1238_
timestamp 1591632351
transform -1 0 1288 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _1480_
timestamp 1591632351
transform 1 0 1288 0 -1 2210
box -4 -6 196 206
use NOR2X1  _720_
timestamp 1591632351
transform -1 0 1528 0 -1 2210
box -4 -6 52 206
use MUX2X1  _713_
timestamp 1591632351
transform -1 0 1624 0 -1 2210
box -4 -6 100 206
use BUFX2  BUFX2_insert40
timestamp 1591632351
transform -1 0 1672 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _1479_
timestamp 1591632351
transform 1 0 1672 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_insert50
timestamp 1591632351
transform -1 0 1912 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert120
timestamp 1591632351
transform 1 0 1912 0 -1 2210
box -4 -6 52 206
use NAND2X1  _1140_
timestamp 1591632351
transform 1 0 1960 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1141_
timestamp 1591632351
transform -1 0 2072 0 -1 2210
box -4 -6 68 206
use NOR2X1  _753_
timestamp 1591632351
transform 1 0 2072 0 -1 2210
box -4 -6 52 206
use NAND2X1  _974_
timestamp 1591632351
transform 1 0 2120 0 -1 2210
box -4 -6 52 206
use OAI21X1  _975_
timestamp 1591632351
transform -1 0 2232 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _1495_
timestamp 1591632351
transform 1 0 2232 0 -1 2210
box -4 -6 196 206
use MUX2X1  _701_
timestamp 1591632351
transform -1 0 2520 0 -1 2210
box -4 -6 100 206
use MUX2X1  _1218_
timestamp 1591632351
transform -1 0 2680 0 -1 2210
box -4 -6 100 206
use FILL  SFILL25200x20100
timestamp 1591632351
transform -1 0 2536 0 -1 2210
box -4 -6 20 206
use FILL  SFILL25360x20100
timestamp 1591632351
transform -1 0 2552 0 -1 2210
box -4 -6 20 206
use FILL  SFILL25520x20100
timestamp 1591632351
transform -1 0 2568 0 -1 2210
box -4 -6 20 206
use FILL  SFILL25680x20100
timestamp 1591632351
transform -1 0 2584 0 -1 2210
box -4 -6 20 206
use BUFX2  BUFX2_insert61
timestamp 1591632351
transform -1 0 2728 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert75
timestamp 1591632351
transform -1 0 2776 0 -1 2210
box -4 -6 52 206
use NAND2X1  _1058_
timestamp 1591632351
transform 1 0 2776 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1059_
timestamp 1591632351
transform -1 0 2888 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _1527_
timestamp 1591632351
transform -1 0 3080 0 -1 2210
box -4 -6 196 206
use MUX2X1  _773_
timestamp 1591632351
transform 1 0 3080 0 -1 2210
box -4 -6 100 206
use MUX2X1  _1290_
timestamp 1591632351
transform 1 0 3176 0 -1 2210
box -4 -6 100 206
use DFFPOSX1  _1463_
timestamp 1591632351
transform -1 0 3464 0 -1 2210
box -4 -6 196 206
use OAI21X1  _1175_
timestamp 1591632351
transform 1 0 3464 0 -1 2210
box -4 -6 68 206
use OAI21X1  _1174_
timestamp 1591632351
transform -1 0 3592 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert56
timestamp 1591632351
transform -1 0 3640 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _1533_
timestamp 1591632351
transform -1 0 3832 0 -1 2210
box -4 -6 196 206
use NAND2X1  _1070_
timestamp 1591632351
transform 1 0 3832 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1071_
timestamp 1591632351
transform -1 0 3944 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert59
timestamp 1591632351
transform 1 0 3944 0 -1 2210
box -4 -6 52 206
use NAND2X1  _1084_
timestamp 1591632351
transform 1 0 3992 0 -1 2210
box -4 -6 52 206
use OAI21X1  _1085_
timestamp 1591632351
transform -1 0 4168 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _1540_
timestamp 1591632351
transform -1 0 4360 0 -1 2210
box -4 -6 196 206
use FILL  SFILL40400x20100
timestamp 1591632351
transform -1 0 4056 0 -1 2210
box -4 -6 20 206
use FILL  SFILL40560x20100
timestamp 1591632351
transform -1 0 4072 0 -1 2210
box -4 -6 20 206
use FILL  SFILL40720x20100
timestamp 1591632351
transform -1 0 4088 0 -1 2210
box -4 -6 20 206
use FILL  SFILL40880x20100
timestamp 1591632351
transform -1 0 4104 0 -1 2210
box -4 -6 20 206
use INVX2  _907_
timestamp 1591632351
transform -1 0 4392 0 -1 2210
box -4 -6 36 206
use NAND2X1  _971_
timestamp 1591632351
transform -1 0 4440 0 -1 2210
box -4 -6 52 206
use NAND3X1  _1028_
timestamp 1591632351
transform 1 0 4440 0 -1 2210
box -4 -6 68 206
use INVX8  _1005_
timestamp 1591632351
transform 1 0 4504 0 -1 2210
box -4 -6 84 206
use DFFPOSX1  _1513_
timestamp 1591632351
transform -1 0 4776 0 -1 2210
box -4 -6 196 206
use OAI21X1  _1100_
timestamp 1591632351
transform -1 0 4840 0 -1 2210
box -4 -6 68 206
use INVX1  _1098_
timestamp 1591632351
transform 1 0 4840 0 -1 2210
box -4 -6 36 206
use OAI21X1  _1133_
timestamp 1591632351
transform 1 0 4872 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _1524_
timestamp 1591632351
transform -1 0 5128 0 -1 2210
box -4 -6 196 206
use FILL  FILL49360x20100
timestamp 1591632351
transform -1 0 5144 0 -1 2210
box -4 -6 20 206
use BUFX2  _1415_
timestamp 1591632351
transform -1 0 56 0 1 2210
box -4 -6 52 206
use BUFX2  _1402_
timestamp 1591632351
transform -1 0 104 0 1 2210
box -4 -6 52 206
use OAI21X1  _1259_
timestamp 1591632351
transform 1 0 104 0 1 2210
box -4 -6 68 206
use OAI21X1  _1223_
timestamp 1591632351
transform 1 0 168 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _1559_
timestamp 1591632351
transform -1 0 424 0 1 2210
box -4 -6 196 206
use OAI21X1  _742_
timestamp 1591632351
transform 1 0 424 0 1 2210
box -4 -6 68 206
use OAI21X1  _1229_
timestamp 1591632351
transform -1 0 552 0 1 2210
box -4 -6 68 206
use OAI21X1  _1228_
timestamp 1591632351
transform -1 0 616 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _1578_
timestamp 1591632351
transform -1 0 808 0 1 2210
box -4 -6 196 206
use OAI21X1  _748_
timestamp 1591632351
transform -1 0 872 0 1 2210
box -4 -6 68 206
use OAI21X1  _747_
timestamp 1591632351
transform -1 0 936 0 1 2210
box -4 -6 68 206
use OAI21X1  _981_
timestamp 1591632351
transform -1 0 1000 0 1 2210
box -4 -6 68 206
use FILL  SFILL10000x22100
timestamp 1591632351
transform 1 0 1000 0 1 2210
box -4 -6 20 206
use DFFPOSX1  _1498_
timestamp 1591632351
transform 1 0 1064 0 1 2210
box -4 -6 196 206
use FILL  SFILL10160x22100
timestamp 1591632351
transform 1 0 1016 0 1 2210
box -4 -6 20 206
use FILL  SFILL10320x22100
timestamp 1591632351
transform 1 0 1032 0 1 2210
box -4 -6 20 206
use FILL  SFILL10480x22100
timestamp 1591632351
transform 1 0 1048 0 1 2210
box -4 -6 20 206
use OAI22X1  _746_
timestamp 1591632351
transform -1 0 1336 0 1 2210
box -4 -6 84 206
use OAI21X1  _745_
timestamp 1591632351
transform -1 0 1400 0 1 2210
box -4 -6 68 206
use OAI21X1  _1262_
timestamp 1591632351
transform 1 0 1400 0 1 2210
box -4 -6 68 206
use NOR2X1  _1237_
timestamp 1591632351
transform -1 0 1512 0 1 2210
box -4 -6 52 206
use NOR2X1  _741_
timestamp 1591632351
transform 1 0 1512 0 1 2210
box -4 -6 52 206
use MUX2X1  _1230_
timestamp 1591632351
transform -1 0 1656 0 1 2210
box -4 -6 100 206
use OAI22X1  _1233_
timestamp 1591632351
transform -1 0 1736 0 1 2210
box -4 -6 84 206
use NOR2X1  _1231_
timestamp 1591632351
transform 1 0 1736 0 1 2210
box -4 -6 52 206
use OAI21X1  _1232_
timestamp 1591632351
transform -1 0 1848 0 1 2210
box -4 -6 68 206
use NAND2X1  _1142_
timestamp 1591632351
transform 1 0 1848 0 1 2210
box -4 -6 52 206
use OAI21X1  _1143_
timestamp 1591632351
transform -1 0 1960 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert114
timestamp 1591632351
transform -1 0 2008 0 1 2210
box -4 -6 52 206
use NOR2X1  _708_
timestamp 1591632351
transform -1 0 2056 0 1 2210
box -4 -6 52 206
use OAI22X1  _710_
timestamp 1591632351
transform -1 0 2136 0 1 2210
box -4 -6 84 206
use OAI21X1  _709_
timestamp 1591632351
transform -1 0 2200 0 1 2210
box -4 -6 68 206
use OAI22X1  _1227_
timestamp 1591632351
transform -1 0 2280 0 1 2210
box -4 -6 84 206
use OAI21X1  _1226_
timestamp 1591632351
transform -1 0 2344 0 1 2210
box -4 -6 68 206
use NOR2X1  _1225_
timestamp 1591632351
transform 1 0 2344 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert34
timestamp 1591632351
transform -1 0 2440 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert64
timestamp 1591632351
transform -1 0 2488 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert110
timestamp 1591632351
transform -1 0 2536 0 1 2210
box -4 -6 52 206
use OAI22X1  _740_
timestamp 1591632351
transform -1 0 2680 0 1 2210
box -4 -6 84 206
use FILL  SFILL25360x22100
timestamp 1591632351
transform 1 0 2536 0 1 2210
box -4 -6 20 206
use FILL  SFILL25520x22100
timestamp 1591632351
transform 1 0 2552 0 1 2210
box -4 -6 20 206
use FILL  SFILL25680x22100
timestamp 1591632351
transform 1 0 2568 0 1 2210
box -4 -6 20 206
use FILL  SFILL25840x22100
timestamp 1591632351
transform 1 0 2584 0 1 2210
box -4 -6 20 206
use OAI21X1  _739_
timestamp 1591632351
transform -1 0 2744 0 1 2210
box -4 -6 68 206
use NOR2X1  _738_
timestamp 1591632351
transform -1 0 2792 0 1 2210
box -4 -6 52 206
use OAI21X1  _1256_
timestamp 1591632351
transform 1 0 2792 0 1 2210
box -4 -6 68 206
use OAI22X1  _1257_
timestamp 1591632351
transform -1 0 2936 0 1 2210
box -4 -6 84 206
use NOR2X1  _1255_
timestamp 1591632351
transform 1 0 2936 0 1 2210
box -4 -6 52 206
use INVX2  _892_
timestamp 1591632351
transform -1 0 3016 0 1 2210
box -4 -6 36 206
use MUX2X1  _737_
timestamp 1591632351
transform 1 0 3016 0 1 2210
box -4 -6 100 206
use MUX2X1  _1254_
timestamp 1591632351
transform 1 0 3112 0 1 2210
box -4 -6 100 206
use BUFX2  BUFX2_insert65
timestamp 1591632351
transform -1 0 3256 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _1466_
timestamp 1591632351
transform -1 0 3448 0 1 2210
box -4 -6 196 206
use OAI21X1  _1181_
timestamp 1591632351
transform 1 0 3448 0 1 2210
box -4 -6 68 206
use OAI21X1  _1180_
timestamp 1591632351
transform -1 0 3576 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert54
timestamp 1591632351
transform 1 0 3576 0 1 2210
box -4 -6 52 206
use DFFPOSX1  _1517_
timestamp 1591632351
transform -1 0 3816 0 1 2210
box -4 -6 196 206
use INVX1  _1110_
timestamp 1591632351
transform 1 0 3816 0 1 2210
box -4 -6 36 206
use OAI21X1  _1112_
timestamp 1591632351
transform 1 0 3848 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert37
timestamp 1591632351
transform -1 0 3960 0 1 2210
box -4 -6 52 206
use NAND2X1  _1064_
timestamp 1591632351
transform 1 0 3960 0 1 2210
box -4 -6 52 206
use OAI21X1  _1065_
timestamp 1591632351
transform -1 0 4072 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _1530_
timestamp 1591632351
transform -1 0 4328 0 1 2210
box -4 -6 196 206
use FILL  SFILL40720x22100
timestamp 1591632351
transform 1 0 4072 0 1 2210
box -4 -6 20 206
use FILL  SFILL40880x22100
timestamp 1591632351
transform 1 0 4088 0 1 2210
box -4 -6 20 206
use FILL  SFILL41040x22100
timestamp 1591632351
transform 1 0 4104 0 1 2210
box -4 -6 20 206
use FILL  SFILL41200x22100
timestamp 1591632351
transform 1 0 4120 0 1 2210
box -4 -6 20 206
use NAND3X1  _1111_
timestamp 1591632351
transform -1 0 4392 0 1 2210
box -4 -6 68 206
use NAND3X1  _1013_
timestamp 1591632351
transform -1 0 4456 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert19
timestamp 1591632351
transform -1 0 4504 0 1 2210
box -4 -6 52 206
use OAI21X1  _1014_
timestamp 1591632351
transform -1 0 4568 0 1 2210
box -4 -6 68 206
use INVX1  _1012_
timestamp 1591632351
transform -1 0 4600 0 1 2210
box -4 -6 36 206
use DFFPOSX1  _1544_
timestamp 1591632351
transform -1 0 4792 0 1 2210
box -4 -6 196 206
use NAND3X1  _1102_
timestamp 1591632351
transform -1 0 4856 0 1 2210
box -4 -6 68 206
use OAI21X1  _1103_
timestamp 1591632351
transform -1 0 4920 0 1 2210
box -4 -6 68 206
use INVX1  _1101_
timestamp 1591632351
transform -1 0 4952 0 1 2210
box -4 -6 36 206
use DFFPOSX1  _1514_
timestamp 1591632351
transform 1 0 4952 0 1 2210
box -4 -6 196 206
use BUFX2  _1406_
timestamp 1591632351
transform -1 0 56 0 -1 2610
box -4 -6 52 206
use BUFX2  _1418_
timestamp 1591632351
transform -1 0 104 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _1562_
timestamp 1591632351
transform -1 0 296 0 -1 2610
box -4 -6 196 206
use OAI21X1  _1265_
timestamp 1591632351
transform -1 0 360 0 -1 2610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert10
timestamp 1591632351
transform -1 0 504 0 -1 2610
box -4 -6 148 206
use OAI21X1  _1264_
timestamp 1591632351
transform -1 0 568 0 -1 2610
box -4 -6 68 206
use OAI21X1  _1276_
timestamp 1591632351
transform -1 0 632 0 -1 2610
box -4 -6 68 206
use NOR2X1  _1258_
timestamp 1591632351
transform 1 0 632 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _1450_
timestamp 1591632351
transform 1 0 680 0 -1 2610
box -4 -6 196 206
use NAND2X1  _899_
timestamp 1591632351
transform 1 0 872 0 -1 2610
box -4 -6 52 206
use OAI21X1  _900_
timestamp 1591632351
transform -1 0 984 0 -1 2610
box -4 -6 68 206
use MUX2X1  _1260_
timestamp 1591632351
transform 1 0 984 0 -1 2610
box -4 -6 100 206
use OAI22X1  _1263_
timestamp 1591632351
transform -1 0 1224 0 -1 2610
box -4 -6 84 206
use FILL  SFILL10800x24100
timestamp 1591632351
transform -1 0 1096 0 -1 2610
box -4 -6 20 206
use FILL  SFILL10960x24100
timestamp 1591632351
transform -1 0 1112 0 -1 2610
box -4 -6 20 206
use FILL  SFILL11120x24100
timestamp 1591632351
transform -1 0 1128 0 -1 2610
box -4 -6 20 206
use FILL  SFILL11280x24100
timestamp 1591632351
transform -1 0 1144 0 -1 2610
box -4 -6 20 206
use MUX2X1  _743_
timestamp 1591632351
transform 1 0 1224 0 -1 2610
box -4 -6 100 206
use NOR2X1  _1261_
timestamp 1591632351
transform 1 0 1320 0 -1 2610
box -4 -6 52 206
use NOR2X1  _744_
timestamp 1591632351
transform -1 0 1416 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _1434_
timestamp 1591632351
transform -1 0 1608 0 -1 2610
box -4 -6 196 206
use OAI21X1  _947_
timestamp 1591632351
transform 1 0 1608 0 -1 2610
box -4 -6 68 206
use OAI21X1  _946_
timestamp 1591632351
transform -1 0 1736 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert31
timestamp 1591632351
transform 1 0 1736 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert45
timestamp 1591632351
transform 1 0 1784 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert89
timestamp 1591632351
transform -1 0 1880 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert118
timestamp 1591632351
transform -1 0 1928 0 -1 2610
box -4 -6 52 206
use OAI21X1  _1182_
timestamp 1591632351
transform -1 0 1992 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert24
timestamp 1591632351
transform 1 0 1992 0 -1 2610
box -4 -6 52 206
use MUX2X1  _707_
timestamp 1591632351
transform -1 0 2136 0 -1 2610
box -4 -6 100 206
use MUX2X1  _1224_
timestamp 1591632351
transform 1 0 2136 0 -1 2610
box -4 -6 100 206
use OAI22X1  _1275_
timestamp 1591632351
transform -1 0 2312 0 -1 2610
box -4 -6 84 206
use OAI21X1  _1274_
timestamp 1591632351
transform -1 0 2376 0 -1 2610
box -4 -6 68 206
use OAI21X1  _757_
timestamp 1591632351
transform 1 0 2376 0 -1 2610
box -4 -6 68 206
use OAI22X1  _758_
timestamp 1591632351
transform -1 0 2520 0 -1 2610
box -4 -6 84 206
use NOR2X1  _756_
timestamp 1591632351
transform -1 0 2568 0 -1 2610
box -4 -6 52 206
use FILL  SFILL25680x24100
timestamp 1591632351
transform -1 0 2584 0 -1 2610
box -4 -6 20 206
use FILL  SFILL25840x24100
timestamp 1591632351
transform -1 0 2600 0 -1 2610
box -4 -6 20 206
use FILL  SFILL26000x24100
timestamp 1591632351
transform -1 0 2616 0 -1 2610
box -4 -6 20 206
use NOR2X1  _1273_
timestamp 1591632351
transform -1 0 2680 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert76
timestamp 1591632351
transform 1 0 2680 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _1482_
timestamp 1591632351
transform -1 0 2920 0 -1 2610
box -4 -6 196 206
use FILL  SFILL26160x24100
timestamp 1591632351
transform -1 0 2632 0 -1 2610
box -4 -6 20 206
use NAND2X1  _1146_
timestamp 1591632351
transform 1 0 2920 0 -1 2610
box -4 -6 52 206
use OAI21X1  _1147_
timestamp 1591632351
transform -1 0 3032 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert117
timestamp 1591632351
transform 1 0 3032 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert39
timestamp 1591632351
transform -1 0 3128 0 -1 2610
box -4 -6 52 206
use DFFPOSX1  _1447_
timestamp 1591632351
transform -1 0 3320 0 -1 2610
box -4 -6 196 206
use NAND2X1  _890_
timestamp 1591632351
transform 1 0 3320 0 -1 2610
box -4 -6 52 206
use OAI21X1  _891_
timestamp 1591632351
transform -1 0 3432 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert86
timestamp 1591632351
transform 1 0 3432 0 -1 2610
box -4 -6 52 206
use OR2X2  _937_
timestamp 1591632351
transform -1 0 3544 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _1486_
timestamp 1591632351
transform -1 0 3736 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  _1531_
timestamp 1591632351
transform -1 0 3928 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  _1499_
timestamp 1591632351
transform -1 0 4120 0 -1 2610
box -4 -6 196 206
use OAI21X1  _983_
timestamp 1591632351
transform -1 0 4248 0 -1 2610
box -4 -6 68 206
use FILL  SFILL41200x24100
timestamp 1591632351
transform -1 0 4136 0 -1 2610
box -4 -6 20 206
use FILL  SFILL41360x24100
timestamp 1591632351
transform -1 0 4152 0 -1 2610
box -4 -6 20 206
use FILL  SFILL41520x24100
timestamp 1591632351
transform -1 0 4168 0 -1 2610
box -4 -6 20 206
use FILL  SFILL41680x24100
timestamp 1591632351
transform -1 0 4184 0 -1 2610
box -4 -6 20 206
use INVX2  _898_
timestamp 1591632351
transform -1 0 4280 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  _1512_
timestamp 1591632351
transform -1 0 4472 0 -1 2610
box -4 -6 196 206
use INVX1  _1095_
timestamp 1591632351
transform 1 0 4472 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  _1547_
timestamp 1591632351
transform -1 0 4696 0 -1 2610
box -4 -6 196 206
use INVX1  _1021_
timestamp 1591632351
transform 1 0 4696 0 -1 2610
box -4 -6 36 206
use OAI21X1  _1023_
timestamp 1591632351
transform 1 0 4728 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _1546_
timestamp 1591632351
transform -1 0 4984 0 -1 2610
box -4 -6 196 206
use NAND3X1  _1019_
timestamp 1591632351
transform -1 0 5048 0 -1 2610
box -4 -6 68 206
use OAI21X1  _1020_
timestamp 1591632351
transform -1 0 5112 0 -1 2610
box -4 -6 68 206
use INVX1  _1018_
timestamp 1591632351
transform -1 0 5144 0 -1 2610
box -4 -6 36 206
use BUFX2  _1419_
timestamp 1591632351
transform -1 0 56 0 1 2610
box -4 -6 52 206
use OAI21X1  _826_
timestamp 1591632351
transform -1 0 120 0 1 2610
box -4 -6 68 206
use OAI21X1  _1271_
timestamp 1591632351
transform 1 0 120 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _1563_
timestamp 1591632351
transform -1 0 376 0 1 2610
box -4 -6 196 206
use OAI21X1  _1277_
timestamp 1591632351
transform -1 0 440 0 1 2610
box -4 -6 68 206
use OAI21X1  _874_
timestamp 1591632351
transform -1 0 504 0 1 2610
box -4 -6 68 206
use OAI21X1  _790_
timestamp 1591632351
transform 1 0 504 0 1 2610
box -4 -6 68 206
use OAI21X1  _832_
timestamp 1591632351
transform -1 0 632 0 1 2610
box -4 -6 68 206
use OAI21X1  _796_
timestamp 1591632351
transform -1 0 696 0 1 2610
box -4 -6 68 206
use OAI21X1  _880_
timestamp 1591632351
transform -1 0 760 0 1 2610
box -4 -6 68 206
use OAI21X1  _795_
timestamp 1591632351
transform -1 0 824 0 1 2610
box -4 -6 68 206
use OAI21X1  _831_
timestamp 1591632351
transform -1 0 888 0 1 2610
box -4 -6 68 206
use OAI21X1  _879_
timestamp 1591632351
transform -1 0 952 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _1509_
timestamp 1591632351
transform 1 0 952 0 1 2610
box -4 -6 196 206
use OAI21X1  _877_
timestamp 1591632351
transform 1 0 1208 0 1 2610
box -4 -6 68 206
use FILL  SFILL11440x26100
timestamp 1591632351
transform 1 0 1144 0 1 2610
box -4 -6 20 206
use FILL  SFILL11600x26100
timestamp 1591632351
transform 1 0 1160 0 1 2610
box -4 -6 20 206
use FILL  SFILL11760x26100
timestamp 1591632351
transform 1 0 1176 0 1 2610
box -4 -6 20 206
use FILL  SFILL11920x26100
timestamp 1591632351
transform 1 0 1192 0 1 2610
box -4 -6 20 206
use OAI22X1  _878_
timestamp 1591632351
transform -1 0 1352 0 1 2610
box -4 -6 84 206
use NOR2X1  _789_
timestamp 1591632351
transform 1 0 1352 0 1 2610
box -4 -6 52 206
use NOR2X1  _873_
timestamp 1591632351
transform 1 0 1400 0 1 2610
box -4 -6 52 206
use NOR2X1  _1270_
timestamp 1591632351
transform 1 0 1448 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert32
timestamp 1591632351
transform -1 0 1544 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _1467_
timestamp 1591632351
transform 1 0 1544 0 1 2610
box -4 -6 196 206
use NOR2X1  _1267_
timestamp 1591632351
transform -1 0 1784 0 1 2610
box -4 -6 52 206
use OAI22X1  _1269_
timestamp 1591632351
transform 1 0 1784 0 1 2610
box -4 -6 84 206
use OAI21X1  _1268_
timestamp 1591632351
transform -1 0 1928 0 1 2610
box -4 -6 68 206
use OAI21X1  _1183_
timestamp 1591632351
transform -1 0 1992 0 1 2610
box -4 -6 68 206
use NOR2X1  _750_
timestamp 1591632351
transform 1 0 1992 0 1 2610
box -4 -6 52 206
use NOR2X1  _825_
timestamp 1591632351
transform 1 0 2040 0 1 2610
box -4 -6 52 206
use OAI21X1  _751_
timestamp 1591632351
transform -1 0 2152 0 1 2610
box -4 -6 68 206
use OAI22X1  _752_
timestamp 1591632351
transform 1 0 2152 0 1 2610
box -4 -6 84 206
use MUX2X1  _1272_
timestamp 1591632351
transform 1 0 2232 0 1 2610
box -4 -6 100 206
use MUX2X1  _1266_
timestamp 1591632351
transform 1 0 2328 0 1 2610
box -4 -6 100 206
use MUX2X1  _749_
timestamp 1591632351
transform 1 0 2424 0 1 2610
box -4 -6 100 206
use BUFX2  BUFX2_insert27
timestamp 1591632351
transform 1 0 2520 0 1 2610
box -4 -6 52 206
use FILL  SFILL25680x26100
timestamp 1591632351
transform 1 0 2568 0 1 2610
box -4 -6 20 206
use FILL  SFILL25840x26100
timestamp 1591632351
transform 1 0 2584 0 1 2610
box -4 -6 20 206
use FILL  SFILL26000x26100
timestamp 1591632351
transform 1 0 2600 0 1 2610
box -4 -6 20 206
use DFFPOSX1  _1489_
timestamp 1591632351
transform -1 0 2824 0 1 2610
box -4 -6 196 206
use FILL  SFILL26160x26100
timestamp 1591632351
transform 1 0 2616 0 1 2610
box -4 -6 20 206
use NAND2X1  _1160_
timestamp 1591632351
transform 1 0 2824 0 1 2610
box -4 -6 52 206
use OAI21X1  _1161_
timestamp 1591632351
transform -1 0 2936 0 1 2610
box -4 -6 68 206
use OAI22X1  _788_
timestamp 1591632351
transform -1 0 3016 0 1 2610
box -4 -6 84 206
use OAI21X1  _787_
timestamp 1591632351
transform 1 0 3016 0 1 2610
box -4 -6 68 206
use NOR2X1  _786_
timestamp 1591632351
transform -1 0 3128 0 1 2610
box -4 -6 52 206
use NOR2X1  _1303_
timestamp 1591632351
transform -1 0 3176 0 1 2610
box -4 -6 52 206
use OAI22X1  _1305_
timestamp 1591632351
transform 1 0 3176 0 1 2610
box -4 -6 84 206
use OAI21X1  _1304_
timestamp 1591632351
transform -1 0 3320 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _1441_
timestamp 1591632351
transform -1 0 3512 0 1 2610
box -4 -6 196 206
use OAI21X1  _960_
timestamp 1591632351
transform -1 0 3576 0 1 2610
box -4 -6 68 206
use OAI21X1  _961_
timestamp 1591632351
transform -1 0 3640 0 1 2610
box -4 -6 68 206
use NAND2X1  _1154_
timestamp 1591632351
transform 1 0 3640 0 1 2610
box -4 -6 52 206
use OAI21X1  _1155_
timestamp 1591632351
transform -1 0 3752 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert25
timestamp 1591632351
transform -1 0 3800 0 1 2610
box -4 -6 52 206
use OR2X2  _1171_
timestamp 1591632351
transform -1 0 3864 0 1 2610
box -4 -6 68 206
use OAI21X1  _1188_
timestamp 1591632351
transform 1 0 3864 0 1 2610
box -4 -6 68 206
use OAI21X1  _1189_
timestamp 1591632351
transform -1 0 3992 0 1 2610
box -4 -6 68 206
use NAND2X1  _1066_
timestamp 1591632351
transform 1 0 3992 0 1 2610
box -4 -6 52 206
use OAI21X1  _1067_
timestamp 1591632351
transform -1 0 4168 0 1 2610
box -4 -6 68 206
use NAND2X1  _982_
timestamp 1591632351
transform 1 0 4168 0 1 2610
box -4 -6 52 206
use OAI21X1  _948_
timestamp 1591632351
transform -1 0 4280 0 1 2610
box -4 -6 68 206
use FILL  SFILL40400x26100
timestamp 1591632351
transform 1 0 4040 0 1 2610
box -4 -6 20 206
use FILL  SFILL40560x26100
timestamp 1591632351
transform 1 0 4056 0 1 2610
box -4 -6 20 206
use FILL  SFILL40720x26100
timestamp 1591632351
transform 1 0 4072 0 1 2610
box -4 -6 20 206
use FILL  SFILL40880x26100
timestamp 1591632351
transform 1 0 4088 0 1 2610
box -4 -6 20 206
use OAI21X1  _954_
timestamp 1591632351
transform -1 0 4344 0 1 2610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert11
timestamp 1591632351
transform -1 0 4488 0 1 2610
box -4 -6 148 206
use OAI21X1  _1097_
timestamp 1591632351
transform 1 0 4488 0 1 2610
box -4 -6 68 206
use NAND3X1  _1096_
timestamp 1591632351
transform 1 0 4552 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert17
timestamp 1591632351
transform -1 0 4664 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert20
timestamp 1591632351
transform 1 0 4664 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _1515_
timestamp 1591632351
transform -1 0 4904 0 1 2610
box -4 -6 196 206
use INVX1  _1104_
timestamp 1591632351
transform 1 0 4904 0 1 2610
box -4 -6 36 206
use OAI21X1  _1106_
timestamp 1591632351
transform 1 0 4936 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert96
timestamp 1591632351
transform -1 0 5048 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert98
timestamp 1591632351
transform 1 0 5048 0 1 2610
box -4 -6 52 206
use FILL  FILL49040x26100
timestamp 1591632351
transform 1 0 5096 0 1 2610
box -4 -6 20 206
use FILL  FILL49200x26100
timestamp 1591632351
transform 1 0 5112 0 1 2610
box -4 -6 20 206
use FILL  FILL49360x26100
timestamp 1591632351
transform 1 0 5128 0 1 2610
box -4 -6 20 206
use DFFPOSX1  _1585_
timestamp 1591632351
transform -1 0 200 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  _1582_
timestamp 1591632351
transform -1 0 392 0 -1 3010
box -4 -6 196 206
use DFFPOSX1  _1589_
timestamp 1591632351
transform -1 0 584 0 -1 3010
box -4 -6 196 206
use INVX4  _1204_
timestamp 1591632351
transform -1 0 632 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1396_
timestamp 1591632351
transform -1 0 696 0 -1 3010
box -4 -6 68 206
use NOR2X1  _1306_
timestamp 1591632351
transform 1 0 696 0 -1 3010
box -4 -6 52 206
use NAND2X1  _1002_
timestamp 1591632351
transform 1 0 744 0 -1 3010
box -4 -6 52 206
use OAI21X1  _1003_
timestamp 1591632351
transform -1 0 856 0 -1 3010
box -4 -6 68 206
use OAI21X1  _1394_
timestamp 1591632351
transform 1 0 856 0 -1 3010
box -4 -6 68 206
use OAI22X1  _1395_
timestamp 1591632351
transform 1 0 920 0 -1 3010
box -4 -6 84 206
use MUX2X1  _1392_
timestamp 1591632351
transform 1 0 1000 0 -1 3010
box -4 -6 100 206
use MUX2X1  _875_
timestamp 1591632351
transform -1 0 1256 0 -1 3010
box -4 -6 100 206
use FILL  SFILL10960x28100
timestamp 1591632351
transform -1 0 1112 0 -1 3010
box -4 -6 20 206
use FILL  SFILL11120x28100
timestamp 1591632351
transform -1 0 1128 0 -1 3010
box -4 -6 20 206
use FILL  SFILL11280x28100
timestamp 1591632351
transform -1 0 1144 0 -1 3010
box -4 -6 20 206
use FILL  SFILL11440x28100
timestamp 1591632351
transform -1 0 1160 0 -1 3010
box -4 -6 20 206
use NOR2X1  _1393_
timestamp 1591632351
transform -1 0 1304 0 -1 3010
box -4 -6 52 206
use NOR2X1  _876_
timestamp 1591632351
transform 1 0 1304 0 -1 3010
box -4 -6 52 206
use MUX2X1  _869_
timestamp 1591632351
transform 1 0 1352 0 -1 3010
box -4 -6 100 206
use OAI22X1  _872_
timestamp 1591632351
transform -1 0 1528 0 -1 3010
box -4 -6 84 206
use OAI21X1  _871_
timestamp 1591632351
transform 1 0 1528 0 -1 3010
box -4 -6 68 206
use NOR2X1  _870_
timestamp 1591632351
transform 1 0 1592 0 -1 3010
box -4 -6 52 206
use OAI21X1  _969_
timestamp 1591632351
transform 1 0 1640 0 -1 3010
box -4 -6 68 206
use OAI21X1  _968_
timestamp 1591632351
transform -1 0 1768 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert80
timestamp 1591632351
transform -1 0 1816 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _1451_
timestamp 1591632351
transform -1 0 2008 0 -1 3010
box -4 -6 196 206
use OAI21X1  _903_
timestamp 1591632351
transform 1 0 2008 0 -1 3010
box -4 -6 68 206
use NAND2X1  _902_
timestamp 1591632351
transform -1 0 2120 0 -1 3010
box -4 -6 52 206
use OAI21X1  _940_
timestamp 1591632351
transform 1 0 2120 0 -1 3010
box -4 -6 68 206
use OAI21X1  _941_
timestamp 1591632351
transform -1 0 2248 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _1431_
timestamp 1591632351
transform -1 0 2440 0 -1 3010
box -4 -6 196 206
use MUX2X1  _755_
timestamp 1591632351
transform 1 0 2440 0 -1 3010
box -4 -6 100 206
use OAI21X1  _1340_
timestamp 1591632351
transform -1 0 2664 0 -1 3010
box -4 -6 68 206
use FILL  SFILL25360x28100
timestamp 1591632351
transform -1 0 2552 0 -1 3010
box -4 -6 20 206
use FILL  SFILL25520x28100
timestamp 1591632351
transform -1 0 2568 0 -1 3010
box -4 -6 20 206
use FILL  SFILL25680x28100
timestamp 1591632351
transform -1 0 2584 0 -1 3010
box -4 -6 20 206
use FILL  SFILL25840x28100
timestamp 1591632351
transform -1 0 2600 0 -1 3010
box -4 -6 20 206
use NOR2X1  _822_
timestamp 1591632351
transform 1 0 2664 0 -1 3010
box -4 -6 52 206
use OAI22X1  _824_
timestamp 1591632351
transform 1 0 2712 0 -1 3010
box -4 -6 84 206
use OAI21X1  _823_
timestamp 1591632351
transform 1 0 2792 0 -1 3010
box -4 -6 68 206
use OAI22X1  _830_
timestamp 1591632351
transform -1 0 2936 0 -1 3010
box -4 -6 84 206
use NOR2X1  _828_
timestamp 1591632351
transform 1 0 2936 0 -1 3010
box -4 -6 52 206
use OAI21X1  _829_
timestamp 1591632351
transform -1 0 3048 0 -1 3010
box -4 -6 68 206
use NOR2X1  _792_
timestamp 1591632351
transform -1 0 3096 0 -1 3010
box -4 -6 52 206
use OAI22X1  _794_
timestamp 1591632351
transform -1 0 3176 0 -1 3010
box -4 -6 84 206
use OAI21X1  _793_
timestamp 1591632351
transform -1 0 3240 0 -1 3010
box -4 -6 68 206
use OAI21X1  _1310_
timestamp 1591632351
transform -1 0 3304 0 -1 3010
box -4 -6 68 206
use MUX2X1  _1302_
timestamp 1591632351
transform 1 0 3304 0 -1 3010
box -4 -6 100 206
use MUX2X1  _785_
timestamp 1591632351
transform 1 0 3400 0 -1 3010
box -4 -6 100 206
use DFFPOSX1  _1505_
timestamp 1591632351
transform -1 0 3688 0 -1 3010
box -4 -6 196 206
use NAND2X1  _994_
timestamp 1591632351
transform 1 0 3688 0 -1 3010
box -4 -6 52 206
use OAI21X1  _995_
timestamp 1591632351
transform -1 0 3800 0 -1 3010
box -4 -6 68 206
use INVX2  _889_
timestamp 1591632351
transform -1 0 3832 0 -1 3010
box -4 -6 36 206
use DFFPOSX1  _1470_
timestamp 1591632351
transform -1 0 4024 0 -1 3010
box -4 -6 196 206
use OAI21X1  _949_
timestamp 1591632351
transform -1 0 4088 0 -1 3010
box -4 -6 68 206
use OAI21X1  _955_
timestamp 1591632351
transform 1 0 4152 0 -1 3010
box -4 -6 68 206
use INVX2  _901_
timestamp 1591632351
transform -1 0 4248 0 -1 3010
box -4 -6 36 206
use FILL  SFILL40880x28100
timestamp 1591632351
transform -1 0 4104 0 -1 3010
box -4 -6 20 206
use FILL  SFILL41040x28100
timestamp 1591632351
transform -1 0 4120 0 -1 3010
box -4 -6 20 206
use FILL  SFILL41200x28100
timestamp 1591632351
transform -1 0 4136 0 -1 3010
box -4 -6 20 206
use FILL  SFILL41360x28100
timestamp 1591632351
transform -1 0 4152 0 -1 3010
box -4 -6 20 206
use OAI21X1  _989_
timestamp 1591632351
transform 1 0 4248 0 -1 3010
box -4 -6 68 206
use NAND2X1  _988_
timestamp 1591632351
transform -1 0 4360 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _1502_
timestamp 1591632351
transform -1 0 4552 0 -1 3010
box -4 -6 196 206
use NAND3X1  _1010_
timestamp 1591632351
transform 1 0 4552 0 -1 3010
box -4 -6 68 206
use INVX1  _1009_
timestamp 1591632351
transform 1 0 4616 0 -1 3010
box -4 -6 36 206
use OAI21X1  _1011_
timestamp 1591632351
transform 1 0 4648 0 -1 3010
box -4 -6 68 206
use DFFPOSX1  _1543_
timestamp 1591632351
transform -1 0 4904 0 -1 3010
box -4 -6 196 206
use NAND3X1  _1022_
timestamp 1591632351
transform 1 0 4904 0 -1 3010
box -4 -6 68 206
use NAND3X1  _1105_
timestamp 1591632351
transform 1 0 4968 0 -1 3010
box -4 -6 68 206
use NAND3X1  _1034_
timestamp 1591632351
transform 1 0 5032 0 -1 3010
box -4 -6 68 206
use FILL  FILL49040x28100
timestamp 1591632351
transform -1 0 5112 0 -1 3010
box -4 -6 20 206
use FILL  FILL49200x28100
timestamp 1591632351
transform -1 0 5128 0 -1 3010
box -4 -6 20 206
use FILL  FILL49360x28100
timestamp 1591632351
transform -1 0 5144 0 -1 3010
box -4 -6 20 206
use BUFX2  _1409_
timestamp 1591632351
transform -1 0 56 0 1 3010
box -4 -6 52 206
use BUFX2  _1429_
timestamp 1591632351
transform -1 0 104 0 1 3010
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert9
timestamp 1591632351
transform -1 0 248 0 1 3010
box -4 -6 148 206
use DFFPOSX1  _1573_
timestamp 1591632351
transform -1 0 440 0 1 3010
box -4 -6 196 206
use OAI21X1  _1391_
timestamp 1591632351
transform -1 0 504 0 1 3010
box -4 -6 68 206
use OAI21X1  _1397_
timestamp 1591632351
transform -1 0 568 0 1 3010
box -4 -6 68 206
use NOR2X1  _1342_
timestamp 1591632351
transform 1 0 568 0 1 3010
box -4 -6 52 206
use OAI21X1  _1348_
timestamp 1591632351
transform -1 0 680 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert69
timestamp 1591632351
transform -1 0 728 0 1 3010
box -4 -6 52 206
use OAI21X1  _1312_
timestamp 1591632351
transform 1 0 728 0 1 3010
box -4 -6 68 206
use NOR2X1  _1390_
timestamp 1591632351
transform 1 0 792 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _1541_
timestamp 1591632351
transform 1 0 840 0 1 3010
box -4 -6 196 206
use NAND2X1  _1086_
timestamp 1591632351
transform 1 0 1096 0 1 3010
box -4 -6 52 206
use OAI21X1  _1087_
timestamp 1591632351
transform -1 0 1208 0 1 3010
box -4 -6 68 206
use OAI22X1  _1389_
timestamp 1591632351
transform -1 0 1288 0 1 3010
box -4 -6 84 206
use FILL  SFILL10320x30100
timestamp 1591632351
transform 1 0 1032 0 1 3010
box -4 -6 20 206
use FILL  SFILL10480x30100
timestamp 1591632351
transform 1 0 1048 0 1 3010
box -4 -6 20 206
use FILL  SFILL10640x30100
timestamp 1591632351
transform 1 0 1064 0 1 3010
box -4 -6 20 206
use FILL  SFILL10800x30100
timestamp 1591632351
transform 1 0 1080 0 1 3010
box -4 -6 20 206
use OAI21X1  _1388_
timestamp 1591632351
transform -1 0 1352 0 1 3010
box -4 -6 68 206
use MUX2X1  _1386_
timestamp 1591632351
transform 1 0 1352 0 1 3010
box -4 -6 100 206
use NOR2X1  _1387_
timestamp 1591632351
transform -1 0 1496 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _1445_
timestamp 1591632351
transform -1 0 1688 0 1 3010
box -4 -6 196 206
use DFFPOSX1  _1525_
timestamp 1591632351
transform -1 0 1880 0 1 3010
box -4 -6 196 206
use INVX1  _1134_
timestamp 1591632351
transform 1 0 1880 0 1 3010
box -4 -6 36 206
use NAND2X1  _1148_
timestamp 1591632351
transform 1 0 1912 0 1 3010
box -4 -6 52 206
use OAI21X1  _1149_
timestamp 1591632351
transform -1 0 2024 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _1483_
timestamp 1591632351
transform 1 0 2024 0 1 3010
box -4 -6 196 206
use OAI21X1  _1136_
timestamp 1591632351
transform 1 0 2216 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert78
timestamp 1591632351
transform 1 0 2280 0 1 3010
box -4 -6 52 206
use NOR2X1  _1339_
timestamp 1591632351
transform 1 0 2328 0 1 3010
box -4 -6 52 206
use OAI22X1  _1341_
timestamp 1591632351
transform 1 0 2376 0 1 3010
box -4 -6 84 206
use OAI22X1  _1347_
timestamp 1591632351
transform -1 0 2536 0 1 3010
box -4 -6 84 206
use NOR2X1  _1345_
timestamp 1591632351
transform -1 0 2648 0 1 3010
box -4 -6 52 206
use FILL  SFILL25360x30100
timestamp 1591632351
transform 1 0 2536 0 1 3010
box -4 -6 20 206
use FILL  SFILL25520x30100
timestamp 1591632351
transform 1 0 2552 0 1 3010
box -4 -6 20 206
use FILL  SFILL25680x30100
timestamp 1591632351
transform 1 0 2568 0 1 3010
box -4 -6 20 206
use FILL  SFILL25840x30100
timestamp 1591632351
transform 1 0 2584 0 1 3010
box -4 -6 20 206
use OAI21X1  _1346_
timestamp 1591632351
transform -1 0 2712 0 1 3010
box -4 -6 68 206
use MUX2X1  _1344_
timestamp 1591632351
transform -1 0 2808 0 1 3010
box -4 -6 100 206
use MUX2X1  _827_
timestamp 1591632351
transform 1 0 2808 0 1 3010
box -4 -6 100 206
use OAI22X1  _1311_
timestamp 1591632351
transform 1 0 2904 0 1 3010
box -4 -6 84 206
use NOR2X1  _1309_
timestamp 1591632351
transform -1 0 3032 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _1457_
timestamp 1591632351
transform -1 0 3224 0 1 3010
box -4 -6 196 206
use NAND2X1  _920_
timestamp 1591632351
transform 1 0 3224 0 1 3010
box -4 -6 52 206
use OAI21X1  _921_
timestamp 1591632351
transform -1 0 3336 0 1 3010
box -4 -6 68 206
use NAND2X1  _911_
timestamp 1591632351
transform 1 0 3336 0 1 3010
box -4 -6 52 206
use OAI21X1  _912_
timestamp 1591632351
transform -1 0 3448 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _1534_
timestamp 1591632351
transform -1 0 3640 0 1 3010
box -4 -6 196 206
use NAND2X1  _1072_
timestamp 1591632351
transform 1 0 3640 0 1 3010
box -4 -6 52 206
use OAI21X1  _1073_
timestamp 1591632351
transform -1 0 3752 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _1435_
timestamp 1591632351
transform -1 0 3944 0 1 3010
box -4 -6 196 206
use NAND3X1  _1093_
timestamp 1591632351
transform 1 0 3944 0 1 3010
box -4 -6 68 206
use FILL  SFILL40080x30100
timestamp 1591632351
transform 1 0 4008 0 1 3010
box -4 -6 20 206
use DFFPOSX1  _1438_
timestamp 1591632351
transform -1 0 4264 0 1 3010
box -4 -6 196 206
use FILL  SFILL40240x30100
timestamp 1591632351
transform 1 0 4024 0 1 3010
box -4 -6 20 206
use FILL  SFILL40400x30100
timestamp 1591632351
transform 1 0 4040 0 1 3010
box -4 -6 20 206
use FILL  SFILL40560x30100
timestamp 1591632351
transform 1 0 4056 0 1 3010
box -4 -6 20 206
use OAI21X1  _1053_
timestamp 1591632351
transform -1 0 4328 0 1 3010
box -4 -6 68 206
use INVX1  _1051_
timestamp 1591632351
transform -1 0 4360 0 1 3010
box -4 -6 36 206
use DFFPOSX1  _1557_
timestamp 1591632351
transform -1 0 4552 0 1 3010
box -4 -6 196 206
use INVX2  _910_
timestamp 1591632351
transform -1 0 4584 0 1 3010
box -4 -6 36 206
use DFFPOSX1  _1518_
timestamp 1591632351
transform -1 0 4776 0 1 3010
box -4 -6 196 206
use OAI21X1  _1115_
timestamp 1591632351
transform -1 0 4840 0 1 3010
box -4 -6 68 206
use INVX1  _1113_
timestamp 1591632351
transform -1 0 4872 0 1 3010
box -4 -6 36 206
use INVX1  _1131_
timestamp 1591632351
transform 1 0 4872 0 1 3010
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert7
timestamp 1591632351
transform -1 0 5048 0 1 3010
box -4 -6 148 206
use BUFX2  BUFX2_insert72
timestamp 1591632351
transform 1 0 5048 0 1 3010
box -4 -6 52 206
use FILL  FILL49040x30100
timestamp 1591632351
transform 1 0 5096 0 1 3010
box -4 -6 20 206
use FILL  FILL49200x30100
timestamp 1591632351
transform 1 0 5112 0 1 3010
box -4 -6 20 206
use FILL  FILL49360x30100
timestamp 1591632351
transform 1 0 5128 0 1 3010
box -4 -6 20 206
use DFFPOSX1  _1569_
timestamp 1591632351
transform -1 0 200 0 -1 3410
box -4 -6 196 206
use BUFX2  _1425_
timestamp 1591632351
transform -1 0 248 0 -1 3410
box -4 -6 52 206
use BUFX2  _1413_
timestamp 1591632351
transform 1 0 248 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1343_
timestamp 1591632351
transform -1 0 360 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1349_
timestamp 1591632351
transform -1 0 424 0 -1 3410
box -4 -6 68 206
use BUFX2  _1422_
timestamp 1591632351
transform -1 0 472 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1307_
timestamp 1591632351
transform 1 0 472 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _1566_
timestamp 1591632351
transform -1 0 728 0 -1 3410
box -4 -6 196 206
use OAI21X1  _1313_
timestamp 1591632351
transform -1 0 792 0 -1 3410
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert15
timestamp 1591632351
transform -1 0 936 0 -1 3410
box -4 -6 148 206
use DFFPOSX1  _1461_
timestamp 1591632351
transform -1 0 1128 0 -1 3410
box -4 -6 196 206
use NAND2X1  _932_
timestamp 1591632351
transform 1 0 1192 0 -1 3410
box -4 -6 52 206
use FILL  SFILL11280x32100
timestamp 1591632351
transform -1 0 1144 0 -1 3410
box -4 -6 20 206
use FILL  SFILL11440x32100
timestamp 1591632351
transform -1 0 1160 0 -1 3410
box -4 -6 20 206
use FILL  SFILL11600x32100
timestamp 1591632351
transform -1 0 1176 0 -1 3410
box -4 -6 20 206
use FILL  SFILL11760x32100
timestamp 1591632351
transform -1 0 1192 0 -1 3410
box -4 -6 20 206
use OAI21X1  _933_
timestamp 1591632351
transform -1 0 1304 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _1493_
timestamp 1591632351
transform -1 0 1496 0 -1 3410
box -4 -6 196 206
use NAND2X1  _1168_
timestamp 1591632351
transform 1 0 1496 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1169_
timestamp 1591632351
transform -1 0 1608 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _1477_
timestamp 1591632351
transform -1 0 1800 0 -1 3410
box -4 -6 196 206
use OAI21X1  _1202_
timestamp 1591632351
transform -1 0 1864 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1203_
timestamp 1591632351
transform -1 0 1928 0 -1 3410
box -4 -6 68 206
use INVX2  _931_
timestamp 1591632351
transform -1 0 1960 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  _1473_
timestamp 1591632351
transform 1 0 1960 0 -1 3410
box -4 -6 196 206
use OAI21X1  _1194_
timestamp 1591632351
transform 1 0 2152 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1195_
timestamp 1591632351
transform -1 0 2280 0 -1 3410
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert4
timestamp 1591632351
transform 1 0 2280 0 -1 3410
box -4 -6 148 206
use DFFPOSX1  _1511_
timestamp 1591632351
transform -1 0 2616 0 -1 3410
box -4 -6 196 206
use INVX1  _1092_
timestamp 1591632351
transform 1 0 2680 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1094_
timestamp 1591632351
transform 1 0 2712 0 -1 3410
box -4 -6 68 206
use MUX2X1  _1338_
timestamp 1591632351
transform -1 0 2872 0 -1 3410
box -4 -6 100 206
use FILL  SFILL26160x32100
timestamp 1591632351
transform -1 0 2632 0 -1 3410
box -4 -6 20 206
use FILL  SFILL26320x32100
timestamp 1591632351
transform -1 0 2648 0 -1 3410
box -4 -6 20 206
use FILL  SFILL26480x32100
timestamp 1591632351
transform -1 0 2664 0 -1 3410
box -4 -6 20 206
use FILL  SFILL26640x32100
timestamp 1591632351
transform -1 0 2680 0 -1 3410
box -4 -6 20 206
use MUX2X1  _821_
timestamp 1591632351
transform -1 0 2968 0 -1 3410
box -4 -6 100 206
use MUX2X1  _1308_
timestamp 1591632351
transform 1 0 2968 0 -1 3410
box -4 -6 100 206
use MUX2X1  _791_
timestamp 1591632351
transform 1 0 3064 0 -1 3410
box -4 -6 100 206
use DFFPOSX1  _1454_
timestamp 1591632351
transform -1 0 3352 0 -1 3410
box -4 -6 196 206
use NAND2X1  _1078_
timestamp 1591632351
transform 1 0 3352 0 -1 3410
box -4 -6 52 206
use OAI21X1  _1079_
timestamp 1591632351
transform -1 0 3464 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _1537_
timestamp 1591632351
transform -1 0 3656 0 -1 3410
box -4 -6 196 206
use INVX2  _919_
timestamp 1591632351
transform -1 0 3688 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  _1521_
timestamp 1591632351
transform -1 0 3880 0 -1 3410
box -4 -6 196 206
use INVX1  _1122_
timestamp 1591632351
transform 1 0 3880 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1124_
timestamp 1591632351
transform 1 0 3912 0 -1 3410
box -4 -6 68 206
use NAND3X1  _1135_
timestamp 1591632351
transform 1 0 3976 0 -1 3410
box -4 -6 68 206
use NAND3X1  _1123_
timestamp 1591632351
transform 1 0 4104 0 -1 3410
box -4 -6 68 206
use NAND3X1  _1052_
timestamp 1591632351
transform 1 0 4168 0 -1 3410
box -4 -6 68 206
use FILL  SFILL40400x32100
timestamp 1591632351
transform -1 0 4056 0 -1 3410
box -4 -6 20 206
use FILL  SFILL40560x32100
timestamp 1591632351
transform -1 0 4072 0 -1 3410
box -4 -6 20 206
use FILL  SFILL40720x32100
timestamp 1591632351
transform -1 0 4088 0 -1 3410
box -4 -6 20 206
use FILL  SFILL40880x32100
timestamp 1591632351
transform -1 0 4104 0 -1 3410
box -4 -6 20 206
use NAND3X1  _1040_
timestamp 1591632351
transform 1 0 4232 0 -1 3410
box -4 -6 68 206
use INVX1  _1039_
timestamp 1591632351
transform 1 0 4296 0 -1 3410
box -4 -6 36 206
use OAI21X1  _1041_
timestamp 1591632351
transform 1 0 4328 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _1553_
timestamp 1591632351
transform -1 0 4584 0 -1 3410
box -4 -6 196 206
use NAND3X1  _1031_
timestamp 1591632351
transform -1 0 4648 0 -1 3410
box -4 -6 68 206
use NAND3X1  _1114_
timestamp 1591632351
transform 1 0 4648 0 -1 3410
box -4 -6 68 206
use OAI21X1  _1032_
timestamp 1591632351
transform -1 0 4776 0 -1 3410
box -4 -6 68 206
use INVX1  _1030_
timestamp 1591632351
transform -1 0 4808 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  _1550_
timestamp 1591632351
transform -1 0 5000 0 -1 3410
box -4 -6 196 206
use INVX1  _1004_
timestamp 1591632351
transform 1 0 5000 0 -1 3410
box -4 -6 36 206
use BUFX2  BUFX2_insert71
timestamp 1591632351
transform -1 0 5080 0 -1 3410
box -4 -6 52 206
use AND2X2  _1089_
timestamp 1591632351
transform 1 0 5080 0 -1 3410
box -4 -6 68 206
<< labels >>
flabel metal4 s 2544 -10 2608 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 1040 -10 1104 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal3 s 5181 137 5187 143 3 FreeSans 24 0 0 0 clock
port 2 nsew
flabel metal2 s 1949 3457 1955 3463 3 FreeSans 24 90 0 0 data_in[15]
port 3 nsew
flabel metal3 s 5181 1757 5187 1763 3 FreeSans 24 0 0 0 data_in[14]
port 4 nsew
flabel metal3 s 5181 1897 5187 1903 3 FreeSans 24 0 0 0 data_in[13]
port 5 nsew
flabel metal3 s 5181 697 5187 703 3 FreeSans 24 0 0 0 data_in[12]
port 6 nsew
flabel metal2 s 3677 3457 3683 3463 3 FreeSans 24 90 0 0 data_in[11]
port 7 nsew
flabel metal3 s 5181 1157 5187 1163 3 FreeSans 24 0 0 0 data_in[10]
port 8 nsew
flabel metal3 s 5181 1197 5187 1203 3 FreeSans 24 0 0 0 data_in[9]
port 9 nsew
flabel metal2 s 4669 3457 4675 3463 3 FreeSans 24 90 0 0 data_in[8]
port 10 nsew
flabel metal3 s 5181 2117 5187 2123 3 FreeSans 24 0 0 0 data_in[7]
port 11 nsew
flabel metal3 s 5181 897 5187 903 3 FreeSans 24 0 0 0 data_in[6]
port 12 nsew
flabel metal3 s 5181 2897 5187 2903 3 FreeSans 24 0 0 0 data_in[5]
port 13 nsew
flabel metal3 s 5181 2497 5187 2503 3 FreeSans 24 0 0 0 data_in[4]
port 14 nsew
flabel metal3 s 5181 1717 5187 1723 3 FreeSans 24 0 0 0 data_in[3]
port 15 nsew
flabel metal2 s 4557 3457 4563 3463 3 FreeSans 24 90 0 0 data_in[2]
port 16 nsew
flabel metal2 s 3949 3457 3955 3463 3 FreeSans 24 90 0 0 data_in[1]
port 17 nsew
flabel metal3 s 5181 1117 5187 1123 3 FreeSans 24 0 0 0 data_in[0]
port 18 nsew
flabel metal3 s -35 1697 -29 1703 7 FreeSans 24 0 0 0 enable
port 19 nsew
flabel metal2 s 1229 -23 1235 -17 7 FreeSans 24 270 0 0 ra_adrs[2]
port 20 nsew
flabel metal2 s 2637 -23 2643 -17 7 FreeSans 24 270 0 0 ra_adrs[1]
port 21 nsew
flabel metal2 s 2253 3457 2259 3463 3 FreeSans 24 90 0 0 ra_adrs[0]
port 22 nsew
flabel metal2 s 269 3457 275 3463 3 FreeSans 24 90 0 0 ra_out[15]
port 23 nsew
flabel metal2 s 1389 -23 1395 -17 7 FreeSans 24 270 0 0 ra_out[14]
port 24 nsew
flabel metal2 s 797 -23 803 -17 7 FreeSans 24 270 0 0 ra_out[13]
port 25 nsew
flabel metal3 s -35 137 -29 143 7 FreeSans 24 0 0 0 ra_out[12]
port 26 nsew
flabel metal3 s -35 3097 -29 3103 7 FreeSans 24 0 0 0 ra_out[11]
port 27 nsew
flabel metal2 s 1133 -23 1139 -17 7 FreeSans 24 270 0 0 ra_out[10]
port 28 nsew
flabel metal2 s 493 -23 499 -17 7 FreeSans 24 270 0 0 ra_out[9]
port 29 nsew
flabel metal3 s -35 2497 -29 2503 7 FreeSans 24 0 0 0 ra_out[8]
port 30 nsew
flabel metal3 s -35 737 -29 743 7 FreeSans 24 0 0 0 ra_out[7]
port 31 nsew
flabel metal2 s 1165 -23 1171 -17 7 FreeSans 24 270 0 0 ra_out[6]
port 32 nsew
flabel metal2 s 1341 -23 1347 -17 7 FreeSans 24 270 0 0 ra_out[5]
port 33 nsew
flabel metal3 s -35 2297 -29 2303 7 FreeSans 24 0 0 0 ra_out[4]
port 34 nsew
flabel metal2 s 669 -23 675 -17 7 FreeSans 24 270 0 0 ra_out[3]
port 35 nsew
flabel metal3 s -35 1897 -29 1903 7 FreeSans 24 0 0 0 ra_out[2]
port 36 nsew
flabel metal3 s -35 1497 -29 1503 7 FreeSans 24 0 0 0 ra_out[1]
port 37 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 ra_out[0]
port 38 nsew
flabel metal2 s 701 3457 707 3463 3 FreeSans 24 90 0 0 rb_adrs[2]
port 39 nsew
flabel metal2 s 2109 -23 2115 -17 7 FreeSans 24 270 0 0 rb_adrs[1]
port 40 nsew
flabel metal2 s 2637 3457 2643 3463 3 FreeSans 24 90 0 0 rb_adrs[0]
port 41 nsew
flabel metal3 s -35 3137 -29 3143 7 FreeSans 24 0 0 0 rb_out[15]
port 42 nsew
flabel metal2 s 1869 -23 1875 -17 7 FreeSans 24 270 0 0 rb_out[14]
port 43 nsew
flabel metal2 s 381 -23 387 -17 7 FreeSans 24 270 0 0 rb_out[13]
port 44 nsew
flabel metal3 s -35 97 -29 103 7 FreeSans 24 0 0 0 rb_out[12]
port 45 nsew
flabel metal2 s 221 3457 227 3463 3 FreeSans 24 90 0 0 rb_out[11]
port 46 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 rb_out[10]
port 47 nsew
flabel metal2 s 1629 -23 1635 -17 7 FreeSans 24 270 0 0 rb_out[9]
port 48 nsew
flabel metal2 s 445 3457 451 3463 3 FreeSans 24 90 0 0 rb_out[8]
port 49 nsew
flabel metal3 s -35 1337 -29 1343 7 FreeSans 24 0 0 0 rb_out[7]
port 50 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 rb_out[6]
port 51 nsew
flabel metal3 s -35 2697 -29 2703 7 FreeSans 24 0 0 0 rb_out[5]
port 52 nsew
flabel metal3 s -35 2537 -29 2543 7 FreeSans 24 0 0 0 rb_out[4]
port 53 nsew
flabel metal3 s -35 1297 -29 1303 7 FreeSans 24 0 0 0 rb_out[3]
port 54 nsew
flabel metal3 s -35 2097 -29 2103 7 FreeSans 24 0 0 0 rb_out[2]
port 55 nsew
flabel metal3 s -35 2337 -29 2343 7 FreeSans 24 0 0 0 rb_out[1]
port 56 nsew
flabel metal3 s -35 937 -29 943 7 FreeSans 24 0 0 0 rb_out[0]
port 57 nsew
flabel metal3 s 5181 1837 5187 1843 3 FreeSans 24 0 0 0 rd_adrs[2]
port 58 nsew
flabel metal3 s 5181 1797 5187 1803 3 FreeSans 24 0 0 0 rd_adrs[1]
port 59 nsew
flabel metal3 s -35 1737 -29 1743 7 FreeSans 24 0 0 0 rd_adrs[0]
port 60 nsew
flabel metal3 s -35 697 -29 703 7 FreeSans 24 0 0 0 wr_en
port 61 nsew
<< end >>
