VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO internal_register
   CLASS BLOCK ;
   FOREIGN internal_register ;
   ORIGIN 3.5000 2.3000 ;
   SIZE 523.8000 BY 348.6000 ;
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.4000 340.4000 514.8000 341.6000 ;
	    RECT 2.8000 336.0000 3.6000 340.4000 ;
	    RECT 8.4000 337.8000 9.2000 340.4000 ;
	    RECT 11.6000 337.8000 12.6000 340.4000 ;
	    RECT 17.2000 335.8000 18.0000 340.4000 ;
	    RECT 22.0000 335.8000 22.8000 340.4000 ;
	    RECT 26.8000 335.8000 27.6000 340.4000 ;
	    RECT 33.2000 336.6000 34.0000 340.4000 ;
	    RECT 39.6000 336.6000 40.4000 340.4000 ;
	    RECT 44.4000 335.8000 45.2000 340.4000 ;
	    RECT 49.2000 336.6000 50.0000 340.4000 ;
	    RECT 55.6000 336.0000 56.4000 340.4000 ;
	    RECT 61.2000 337.8000 62.0000 340.4000 ;
	    RECT 64.4000 337.8000 65.4000 340.4000 ;
	    RECT 70.0000 335.8000 70.8000 340.4000 ;
	    RECT 76.4000 336.6000 77.2000 340.4000 ;
	    RECT 79.6000 335.8000 80.4000 340.4000 ;
	    RECT 82.8000 335.8000 83.6000 340.4000 ;
	    RECT 86.0000 335.8000 86.8000 340.4000 ;
	    RECT 89.2000 335.8000 90.0000 340.4000 ;
	    RECT 92.4000 335.8000 93.2000 340.4000 ;
	    RECT 95.6000 336.0000 96.4000 340.4000 ;
	    RECT 101.2000 337.8000 102.0000 340.4000 ;
	    RECT 104.4000 337.8000 105.4000 340.4000 ;
	    RECT 110.0000 335.8000 110.8000 340.4000 ;
	    RECT 119.6000 335.8000 120.4000 340.4000 ;
	    RECT 127.6000 336.6000 128.4000 340.4000 ;
	    RECT 132.4000 336.0000 133.2000 340.4000 ;
	    RECT 138.0000 337.8000 138.8000 340.4000 ;
	    RECT 141.2000 337.8000 142.2000 340.4000 ;
	    RECT 146.8000 335.8000 147.6000 340.4000 ;
	    RECT 150.0000 335.8000 150.8000 340.4000 ;
	    RECT 158.0000 336.6000 158.8000 340.4000 ;
	    RECT 162.8000 336.0000 163.6000 340.4000 ;
	    RECT 168.4000 337.8000 169.2000 340.4000 ;
	    RECT 171.6000 337.8000 172.6000 340.4000 ;
	    RECT 177.2000 335.8000 178.0000 340.4000 ;
	    RECT 183.6000 336.6000 184.4000 340.4000 ;
	    RECT 190.0000 336.6000 190.8000 340.4000 ;
	    RECT 194.8000 335.8000 195.6000 340.4000 ;
	    RECT 198.0000 335.8000 198.8000 340.4000 ;
	    RECT 203.4000 337.8000 204.4000 340.4000 ;
	    RECT 206.8000 337.8000 207.6000 340.4000 ;
	    RECT 212.4000 336.0000 213.2000 340.4000 ;
	    RECT 217.2000 336.6000 218.0000 340.4000 ;
	    RECT 225.2000 336.6000 226.0000 340.4000 ;
	    RECT 228.4000 335.8000 229.2000 340.4000 ;
	    RECT 231.6000 335.8000 232.4000 340.4000 ;
	    RECT 234.8000 335.8000 235.6000 340.4000 ;
	    RECT 238.0000 335.8000 238.8000 340.4000 ;
	    RECT 241.2000 335.8000 242.0000 340.4000 ;
	    RECT 244.4000 336.0000 245.2000 340.4000 ;
	    RECT 250.0000 337.8000 250.8000 340.4000 ;
	    RECT 253.2000 337.8000 254.2000 340.4000 ;
	    RECT 258.8000 335.8000 259.6000 340.4000 ;
	    RECT 268.4000 337.8000 269.2000 340.4000 ;
	    RECT 273.2000 336.6000 274.0000 340.4000 ;
	    RECT 279.2000 335.0000 280.0000 340.4000 ;
	    RECT 284.4000 335.4000 285.2000 340.4000 ;
	    RECT 288.8000 335.0000 289.6000 340.4000 ;
	    RECT 294.0000 335.4000 294.8000 340.4000 ;
	    RECT 298.8000 335.4000 299.6000 340.4000 ;
	    RECT 304.0000 335.0000 304.8000 340.4000 ;
	    RECT 308.4000 335.4000 309.2000 340.4000 ;
	    RECT 313.6000 335.0000 314.4000 340.4000 ;
	    RECT 318.0000 336.0000 318.8000 340.4000 ;
	    RECT 323.6000 337.8000 324.4000 340.4000 ;
	    RECT 326.8000 337.8000 327.8000 340.4000 ;
	    RECT 332.4000 335.8000 333.2000 340.4000 ;
	    RECT 335.6000 335.8000 336.4000 340.4000 ;
	    RECT 343.6000 336.6000 344.4000 340.4000 ;
	    RECT 348.4000 336.0000 349.2000 340.4000 ;
	    RECT 354.0000 337.8000 354.8000 340.4000 ;
	    RECT 357.2000 337.8000 358.2000 340.4000 ;
	    RECT 362.8000 335.8000 363.6000 340.4000 ;
	    RECT 367.6000 335.8000 368.4000 340.4000 ;
	    RECT 370.8000 336.0000 371.6000 340.4000 ;
	    RECT 376.4000 337.8000 377.2000 340.4000 ;
	    RECT 379.6000 337.8000 380.6000 340.4000 ;
	    RECT 385.2000 335.8000 386.0000 340.4000 ;
	    RECT 388.4000 337.8000 389.2000 340.4000 ;
	    RECT 393.2000 336.6000 394.0000 340.4000 ;
	    RECT 398.0000 333.8000 398.8000 340.4000 ;
	    RECT 410.8000 333.8000 411.6000 340.4000 ;
	    RECT 417.2000 333.8000 418.0000 340.4000 ;
	    RECT 423.6000 333.8000 424.4000 340.4000 ;
	    RECT 430.0000 337.8000 430.8000 340.4000 ;
	    RECT 434.8000 336.6000 435.6000 340.4000 ;
	    RECT 441.2000 336.0000 442.0000 340.4000 ;
	    RECT 446.8000 337.8000 447.6000 340.4000 ;
	    RECT 450.0000 337.8000 451.0000 340.4000 ;
	    RECT 455.6000 335.8000 456.4000 340.4000 ;
	    RECT 463.6000 333.8000 464.4000 340.4000 ;
	    RECT 465.2000 333.8000 466.0000 340.4000 ;
	    RECT 474.8000 336.6000 475.6000 340.4000 ;
	    RECT 479.6000 337.8000 480.4000 340.4000 ;
	    RECT 482.8000 336.0000 483.6000 340.4000 ;
	    RECT 488.4000 337.8000 489.2000 340.4000 ;
	    RECT 491.6000 337.8000 492.6000 340.4000 ;
	    RECT 497.2000 335.8000 498.0000 340.4000 ;
	    RECT 500.4000 337.8000 501.2000 340.4000 ;
	    RECT 505.2000 335.8000 506.0000 340.4000 ;
	    RECT 511.0000 336.0000 511.8000 340.4000 ;
	    RECT 2.8000 301.6000 3.6000 306.2000 ;
	    RECT 7.6000 301.6000 8.4000 306.2000 ;
	    RECT 10.8000 301.6000 11.6000 306.2000 ;
	    RECT 14.0000 301.6000 14.8000 306.2000 ;
	    RECT 17.2000 301.6000 18.0000 306.2000 ;
	    RECT 20.4000 301.6000 21.2000 306.2000 ;
	    RECT 23.6000 301.6000 24.4000 306.2000 ;
	    RECT 26.8000 301.6000 27.6000 306.0000 ;
	    RECT 32.4000 301.6000 33.2000 304.2000 ;
	    RECT 35.6000 301.6000 36.6000 304.2000 ;
	    RECT 41.2000 301.6000 42.0000 306.2000 ;
	    RECT 47.6000 301.6000 48.4000 305.4000 ;
	    RECT 54.0000 301.6000 54.8000 305.4000 ;
	    RECT 57.2000 301.6000 58.0000 304.2000 ;
	    RECT 60.4000 301.6000 61.2000 304.2000 ;
	    RECT 65.2000 301.6000 66.0000 305.4000 ;
	    RECT 70.0000 301.6000 70.8000 306.2000 ;
	    RECT 74.8000 301.6000 75.6000 305.4000 ;
	    RECT 79.6000 301.6000 80.4000 304.2000 ;
	    RECT 82.8000 301.6000 83.6000 304.2000 ;
	    RECT 86.0000 301.6000 86.8000 306.2000 ;
	    RECT 91.4000 301.6000 92.4000 304.2000 ;
	    RECT 94.8000 301.6000 95.6000 304.2000 ;
	    RECT 100.4000 301.6000 101.2000 306.0000 ;
	    RECT 110.0000 301.6000 110.8000 306.2000 ;
	    RECT 118.0000 301.6000 118.8000 305.4000 ;
	    RECT 126.0000 301.6000 126.8000 305.4000 ;
	    RECT 132.4000 301.6000 133.2000 305.4000 ;
	    RECT 137.2000 301.6000 138.0000 306.6000 ;
	    RECT 142.4000 301.6000 143.2000 307.0000 ;
	    RECT 145.2000 301.6000 146.0000 304.2000 ;
	    RECT 148.4000 301.6000 149.2000 304.2000 ;
	    RECT 151.6000 301.6000 152.4000 306.0000 ;
	    RECT 157.2000 301.6000 158.0000 304.2000 ;
	    RECT 160.4000 301.6000 161.4000 304.2000 ;
	    RECT 166.0000 301.6000 166.8000 306.2000 ;
	    RECT 170.8000 301.6000 171.6000 306.0000 ;
	    RECT 176.4000 301.6000 177.2000 304.2000 ;
	    RECT 179.6000 301.6000 180.6000 304.2000 ;
	    RECT 185.2000 301.6000 186.0000 306.2000 ;
	    RECT 188.4000 301.6000 189.2000 304.2000 ;
	    RECT 191.6000 301.6000 192.4000 306.2000 ;
	    RECT 199.6000 301.6000 200.4000 305.4000 ;
	    RECT 204.4000 301.6000 205.2000 306.2000 ;
	    RECT 209.8000 301.6000 210.8000 304.2000 ;
	    RECT 213.2000 301.6000 214.0000 304.2000 ;
	    RECT 218.8000 301.6000 219.6000 306.0000 ;
	    RECT 223.6000 301.6000 224.4000 305.4000 ;
	    RECT 230.0000 301.6000 230.8000 306.2000 ;
	    RECT 233.2000 301.6000 234.0000 304.2000 ;
	    RECT 236.4000 301.6000 237.2000 304.2000 ;
	    RECT 239.6000 301.6000 240.4000 305.4000 ;
	    RECT 250.8000 301.6000 251.6000 305.4000 ;
	    RECT 260.4000 301.6000 261.2000 304.2000 ;
	    RECT 263.6000 301.6000 264.4000 304.2000 ;
	    RECT 268.4000 301.6000 269.2000 305.4000 ;
	    RECT 272.8000 301.6000 273.6000 307.0000 ;
	    RECT 278.0000 301.6000 278.8000 306.6000 ;
	    RECT 282.8000 301.6000 283.6000 306.6000 ;
	    RECT 288.0000 301.6000 288.8000 307.0000 ;
	    RECT 292.4000 301.6000 293.2000 305.4000 ;
	    RECT 298.8000 301.6000 299.6000 304.2000 ;
	    RECT 302.0000 301.6000 302.8000 304.2000 ;
	    RECT 305.2000 301.6000 306.0000 306.0000 ;
	    RECT 310.8000 301.6000 311.6000 304.2000 ;
	    RECT 314.0000 301.6000 315.0000 304.2000 ;
	    RECT 319.6000 301.6000 320.4000 306.2000 ;
	    RECT 322.8000 301.6000 323.6000 306.2000 ;
	    RECT 330.8000 301.6000 331.6000 305.4000 ;
	    RECT 334.0000 301.6000 334.8000 306.2000 ;
	    RECT 342.0000 301.6000 342.8000 305.4000 ;
	    RECT 346.8000 301.6000 347.6000 306.0000 ;
	    RECT 352.4000 301.6000 353.2000 304.2000 ;
	    RECT 355.6000 301.6000 356.6000 304.2000 ;
	    RECT 361.2000 301.6000 362.0000 306.2000 ;
	    RECT 364.4000 301.6000 365.2000 306.2000 ;
	    RECT 372.4000 301.6000 373.2000 305.4000 ;
	    RECT 377.2000 301.6000 378.0000 306.0000 ;
	    RECT 382.8000 301.6000 383.6000 304.2000 ;
	    RECT 386.0000 301.6000 387.0000 304.2000 ;
	    RECT 391.6000 301.6000 392.4000 306.2000 ;
	    RECT 394.8000 301.6000 395.6000 308.2000 ;
	    RECT 409.2000 301.6000 410.0000 306.0000 ;
	    RECT 414.8000 301.6000 415.6000 304.2000 ;
	    RECT 418.0000 301.6000 419.0000 304.2000 ;
	    RECT 423.6000 301.6000 424.4000 306.2000 ;
	    RECT 430.0000 301.6000 430.8000 305.4000 ;
	    RECT 434.8000 301.6000 435.6000 304.2000 ;
	    RECT 438.0000 301.6000 438.8000 306.0000 ;
	    RECT 443.6000 301.6000 444.4000 304.2000 ;
	    RECT 446.8000 301.6000 447.8000 304.2000 ;
	    RECT 452.4000 301.6000 453.2000 306.2000 ;
	    RECT 457.2000 301.6000 458.0000 306.2000 ;
	    RECT 460.4000 301.6000 461.2000 306.0000 ;
	    RECT 466.0000 301.6000 466.8000 304.2000 ;
	    RECT 469.2000 301.6000 470.2000 304.2000 ;
	    RECT 474.8000 301.6000 475.6000 306.2000 ;
	    RECT 481.2000 301.6000 482.0000 305.4000 ;
	    RECT 486.0000 301.6000 486.8000 304.2000 ;
	    RECT 487.6000 301.6000 488.4000 304.2000 ;
	    RECT 490.8000 301.6000 491.6000 306.2000 ;
	    RECT 494.0000 301.6000 494.8000 306.2000 ;
	    RECT 497.2000 301.6000 498.0000 306.2000 ;
	    RECT 500.4000 301.6000 501.2000 306.2000 ;
	    RECT 503.6000 301.6000 504.4000 306.2000 ;
	    RECT 506.8000 301.6000 507.6000 306.2000 ;
	    RECT 0.4000 300.4000 514.8000 301.6000 ;
	    RECT 2.8000 296.0000 3.6000 300.4000 ;
	    RECT 8.4000 297.8000 9.2000 300.4000 ;
	    RECT 11.6000 297.8000 12.6000 300.4000 ;
	    RECT 17.2000 295.8000 18.0000 300.4000 ;
	    RECT 22.0000 296.0000 22.8000 300.4000 ;
	    RECT 27.6000 297.8000 28.4000 300.4000 ;
	    RECT 30.8000 297.8000 31.8000 300.4000 ;
	    RECT 36.4000 295.8000 37.2000 300.4000 ;
	    RECT 41.2000 296.0000 42.0000 300.4000 ;
	    RECT 46.8000 297.8000 47.6000 300.4000 ;
	    RECT 50.0000 297.8000 51.0000 300.4000 ;
	    RECT 55.6000 295.8000 56.4000 300.4000 ;
	    RECT 58.8000 295.8000 59.6000 300.4000 ;
	    RECT 62.0000 295.8000 62.8000 300.4000 ;
	    RECT 66.8000 296.6000 67.6000 300.4000 ;
	    RECT 70.0000 297.8000 70.8000 300.4000 ;
	    RECT 73.2000 297.8000 74.0000 300.4000 ;
	    RECT 74.8000 295.8000 75.6000 300.4000 ;
	    RECT 82.8000 296.6000 83.6000 300.4000 ;
	    RECT 87.6000 296.6000 88.4000 300.4000 ;
	    RECT 94.0000 296.6000 94.8000 300.4000 ;
	    RECT 102.0000 295.4000 102.8000 300.4000 ;
	    RECT 107.2000 295.0000 108.0000 300.4000 ;
	    RECT 117.6000 295.0000 118.4000 300.4000 ;
	    RECT 122.8000 295.4000 123.6000 300.4000 ;
	    RECT 126.0000 297.8000 126.8000 300.4000 ;
	    RECT 129.2000 297.8000 130.0000 300.4000 ;
	    RECT 130.8000 297.8000 131.6000 300.4000 ;
	    RECT 134.0000 297.8000 134.8000 300.4000 ;
	    RECT 137.2000 295.4000 138.0000 300.4000 ;
	    RECT 142.4000 295.0000 143.2000 300.4000 ;
	    RECT 150.0000 296.6000 150.8000 300.4000 ;
	    RECT 154.8000 296.6000 155.6000 300.4000 ;
	    RECT 159.6000 297.8000 160.4000 300.4000 ;
	    RECT 162.8000 297.8000 163.6000 300.4000 ;
	    RECT 166.0000 296.6000 166.8000 300.4000 ;
	    RECT 174.0000 296.6000 174.8000 300.4000 ;
	    RECT 178.8000 295.8000 179.6000 300.4000 ;
	    RECT 183.6000 296.0000 184.4000 300.4000 ;
	    RECT 189.2000 297.8000 190.0000 300.4000 ;
	    RECT 192.4000 297.8000 193.4000 300.4000 ;
	    RECT 198.0000 295.8000 198.8000 300.4000 ;
	    RECT 202.8000 296.6000 203.6000 300.4000 ;
	    RECT 210.8000 295.8000 211.6000 300.4000 ;
	    RECT 214.0000 296.6000 214.8000 300.4000 ;
	    RECT 222.0000 296.6000 222.8000 300.4000 ;
	    RECT 226.8000 296.0000 227.6000 300.4000 ;
	    RECT 232.4000 297.8000 233.2000 300.4000 ;
	    RECT 235.6000 297.8000 236.6000 300.4000 ;
	    RECT 241.2000 295.8000 242.0000 300.4000 ;
	    RECT 246.0000 295.4000 246.8000 300.4000 ;
	    RECT 251.2000 295.0000 252.0000 300.4000 ;
	    RECT 263.6000 296.6000 264.4000 300.4000 ;
	    RECT 266.8000 297.8000 267.6000 300.4000 ;
	    RECT 270.0000 297.8000 270.8000 300.4000 ;
	    RECT 273.2000 296.6000 274.0000 300.4000 ;
	    RECT 281.2000 296.6000 282.0000 300.4000 ;
	    RECT 290.8000 296.6000 291.6000 300.4000 ;
	    RECT 294.0000 297.8000 294.8000 300.4000 ;
	    RECT 297.2000 297.8000 298.0000 300.4000 ;
	    RECT 302.0000 296.6000 302.8000 300.4000 ;
	    RECT 305.2000 297.8000 306.0000 300.4000 ;
	    RECT 308.4000 297.8000 309.2000 300.4000 ;
	    RECT 314.8000 296.6000 315.6000 300.4000 ;
	    RECT 321.2000 296.6000 322.0000 300.4000 ;
	    RECT 327.6000 296.6000 328.4000 300.4000 ;
	    RECT 332.4000 295.4000 333.2000 300.4000 ;
	    RECT 337.6000 295.0000 338.4000 300.4000 ;
	    RECT 342.0000 295.4000 342.8000 300.4000 ;
	    RECT 347.2000 295.0000 348.0000 300.4000 ;
	    RECT 351.6000 296.0000 352.4000 300.4000 ;
	    RECT 357.2000 297.8000 358.0000 300.4000 ;
	    RECT 360.4000 297.8000 361.4000 300.4000 ;
	    RECT 366.0000 295.8000 366.8000 300.4000 ;
	    RECT 369.2000 295.8000 370.0000 300.4000 ;
	    RECT 377.2000 296.6000 378.0000 300.4000 ;
	    RECT 382.0000 295.8000 382.8000 300.4000 ;
	    RECT 385.2000 296.0000 386.0000 300.4000 ;
	    RECT 390.8000 297.8000 391.6000 300.4000 ;
	    RECT 394.0000 297.8000 395.0000 300.4000 ;
	    RECT 399.6000 295.8000 400.4000 300.4000 ;
	    RECT 406.0000 296.6000 406.8000 300.4000 ;
	    RECT 417.2000 296.6000 418.0000 300.4000 ;
	    RECT 423.6000 295.8000 424.4000 300.4000 ;
	    RECT 426.8000 296.6000 427.6000 300.4000 ;
	    RECT 434.8000 295.8000 435.6000 300.4000 ;
	    RECT 438.0000 296.0000 438.8000 300.4000 ;
	    RECT 443.6000 297.8000 444.4000 300.4000 ;
	    RECT 446.8000 297.8000 447.8000 300.4000 ;
	    RECT 452.4000 295.8000 453.2000 300.4000 ;
	    RECT 455.6000 293.8000 456.4000 300.4000 ;
	    RECT 462.0000 297.8000 462.8000 300.4000 ;
	    RECT 466.8000 296.6000 467.6000 300.4000 ;
	    RECT 473.2000 296.0000 474.0000 300.4000 ;
	    RECT 478.8000 297.8000 479.6000 300.4000 ;
	    RECT 482.0000 297.8000 483.0000 300.4000 ;
	    RECT 487.6000 295.8000 488.4000 300.4000 ;
	    RECT 490.8000 293.8000 491.6000 300.4000 ;
	    RECT 497.2000 293.8000 498.0000 300.4000 ;
	    RECT 503.6000 293.8000 504.4000 300.4000 ;
	    RECT 2.8000 261.6000 3.6000 266.2000 ;
	    RECT 9.2000 261.6000 10.0000 265.4000 ;
	    RECT 14.0000 261.6000 14.8000 265.4000 ;
	    RECT 20.4000 261.6000 21.2000 266.0000 ;
	    RECT 26.0000 261.6000 26.8000 264.2000 ;
	    RECT 29.2000 261.6000 30.2000 264.2000 ;
	    RECT 34.8000 261.6000 35.6000 266.2000 ;
	    RECT 41.2000 261.6000 42.0000 265.4000 ;
	    RECT 47.6000 261.6000 48.4000 265.4000 ;
	    RECT 52.4000 261.6000 53.2000 265.4000 ;
	    RECT 60.4000 261.6000 61.2000 265.4000 ;
	    RECT 66.8000 261.6000 67.6000 265.4000 ;
	    RECT 73.2000 261.6000 74.0000 265.4000 ;
	    RECT 79.6000 261.6000 80.4000 265.4000 ;
	    RECT 86.0000 261.6000 86.8000 265.4000 ;
	    RECT 92.4000 261.6000 93.2000 265.4000 ;
	    RECT 97.2000 261.6000 98.0000 266.2000 ;
	    RECT 102.6000 261.6000 103.6000 264.2000 ;
	    RECT 106.0000 261.6000 106.8000 264.2000 ;
	    RECT 111.6000 261.6000 112.4000 266.0000 ;
	    RECT 122.8000 261.6000 123.6000 265.4000 ;
	    RECT 132.4000 261.6000 133.2000 265.4000 ;
	    RECT 135.6000 261.6000 136.4000 264.2000 ;
	    RECT 138.8000 261.6000 139.6000 264.2000 ;
	    RECT 140.4000 261.6000 141.2000 264.2000 ;
	    RECT 143.6000 261.6000 144.4000 264.2000 ;
	    RECT 145.2000 261.6000 146.0000 264.2000 ;
	    RECT 148.4000 261.6000 149.2000 264.2000 ;
	    RECT 151.6000 261.6000 152.4000 266.2000 ;
	    RECT 156.4000 261.6000 157.2000 266.2000 ;
	    RECT 161.8000 261.6000 162.8000 264.2000 ;
	    RECT 165.2000 261.6000 166.0000 264.2000 ;
	    RECT 170.8000 261.6000 171.6000 266.0000 ;
	    RECT 174.0000 261.6000 174.8000 264.2000 ;
	    RECT 177.2000 261.6000 178.0000 264.2000 ;
	    RECT 180.4000 261.6000 181.2000 265.4000 ;
	    RECT 190.0000 261.6000 190.8000 265.4000 ;
	    RECT 196.4000 261.6000 197.2000 265.4000 ;
	    RECT 199.6000 261.6000 200.4000 264.2000 ;
	    RECT 202.8000 261.6000 203.6000 264.2000 ;
	    RECT 204.4000 261.6000 205.2000 264.2000 ;
	    RECT 207.6000 261.6000 208.4000 264.2000 ;
	    RECT 212.4000 261.6000 213.2000 265.4000 ;
	    RECT 217.2000 261.6000 218.0000 265.4000 ;
	    RECT 225.2000 261.6000 226.0000 266.6000 ;
	    RECT 230.4000 261.6000 231.2000 267.0000 ;
	    RECT 234.8000 261.6000 235.6000 266.6000 ;
	    RECT 240.0000 261.6000 240.8000 267.0000 ;
	    RECT 244.4000 261.6000 245.2000 266.6000 ;
	    RECT 249.6000 261.6000 250.4000 267.0000 ;
	    RECT 254.0000 261.6000 254.8000 266.2000 ;
	    RECT 265.2000 261.6000 266.0000 266.0000 ;
	    RECT 270.8000 261.6000 271.6000 264.2000 ;
	    RECT 274.0000 261.6000 275.0000 264.2000 ;
	    RECT 279.6000 261.6000 280.4000 266.2000 ;
	    RECT 282.8000 261.6000 283.6000 266.2000 ;
	    RECT 290.8000 261.6000 291.6000 265.4000 ;
	    RECT 298.8000 261.6000 299.6000 265.4000 ;
	    RECT 303.6000 261.6000 304.4000 265.4000 ;
	    RECT 308.4000 261.6000 309.2000 264.2000 ;
	    RECT 311.6000 261.6000 312.4000 264.2000 ;
	    RECT 313.2000 261.6000 314.0000 264.2000 ;
	    RECT 316.4000 261.6000 317.2000 264.2000 ;
	    RECT 319.6000 261.6000 320.4000 265.4000 ;
	    RECT 329.2000 261.6000 330.0000 265.4000 ;
	    RECT 334.0000 261.6000 334.8000 266.0000 ;
	    RECT 339.6000 261.6000 340.4000 264.2000 ;
	    RECT 342.8000 261.6000 343.8000 264.2000 ;
	    RECT 348.4000 261.6000 349.2000 266.2000 ;
	    RECT 354.8000 261.6000 355.6000 265.4000 ;
	    RECT 361.2000 261.6000 362.0000 265.4000 ;
	    RECT 364.4000 261.6000 365.2000 266.2000 ;
	    RECT 372.4000 261.6000 373.2000 265.4000 ;
	    RECT 377.2000 261.6000 378.0000 266.2000 ;
	    RECT 382.0000 261.6000 382.8000 265.8000 ;
	    RECT 385.2000 261.6000 386.0000 264.2000 ;
	    RECT 388.4000 261.6000 389.2000 265.4000 ;
	    RECT 396.4000 261.6000 397.2000 265.4000 ;
	    RECT 399.6000 261.6000 400.4000 266.2000 ;
	    RECT 414.0000 261.6000 414.8000 265.4000 ;
	    RECT 417.2000 261.6000 418.0000 266.2000 ;
	    RECT 425.2000 261.6000 426.0000 265.4000 ;
	    RECT 431.6000 261.6000 432.4000 265.4000 ;
	    RECT 434.8000 261.6000 435.6000 266.2000 ;
	    RECT 438.0000 261.6000 438.8000 266.2000 ;
	    RECT 441.2000 261.6000 442.0000 266.2000 ;
	    RECT 444.4000 261.6000 445.2000 266.2000 ;
	    RECT 447.6000 261.6000 448.4000 266.2000 ;
	    RECT 450.8000 261.6000 451.6000 265.4000 ;
	    RECT 455.6000 261.6000 456.4000 268.2000 ;
	    RECT 463.6000 261.6000 464.4000 266.2000 ;
	    RECT 468.4000 261.6000 469.2000 266.2000 ;
	    RECT 473.2000 261.6000 474.0000 266.0000 ;
	    RECT 478.8000 261.6000 479.6000 264.2000 ;
	    RECT 482.0000 261.6000 483.0000 264.2000 ;
	    RECT 487.6000 261.6000 488.4000 266.2000 ;
	    RECT 490.8000 261.6000 491.6000 264.2000 ;
	    RECT 495.6000 261.6000 496.4000 265.4000 ;
	    RECT 502.0000 261.6000 502.8000 266.2000 ;
	    RECT 506.8000 261.6000 507.6000 266.2000 ;
	    RECT 0.4000 260.4000 514.8000 261.6000 ;
	    RECT 2.8000 255.8000 3.6000 260.4000 ;
	    RECT 7.6000 255.8000 8.4000 260.4000 ;
	    RECT 12.4000 256.0000 13.2000 260.4000 ;
	    RECT 18.0000 257.8000 18.8000 260.4000 ;
	    RECT 21.2000 257.8000 22.2000 260.4000 ;
	    RECT 26.8000 255.8000 27.6000 260.4000 ;
	    RECT 33.2000 256.6000 34.0000 260.4000 ;
	    RECT 36.4000 255.8000 37.2000 260.4000 ;
	    RECT 39.6000 255.8000 40.4000 260.4000 ;
	    RECT 42.8000 255.8000 43.6000 260.4000 ;
	    RECT 46.0000 255.8000 46.8000 260.4000 ;
	    RECT 49.2000 255.8000 50.0000 260.4000 ;
	    RECT 54.0000 256.6000 54.8000 260.4000 ;
	    RECT 60.4000 256.6000 61.2000 260.4000 ;
	    RECT 63.6000 257.8000 64.4000 260.4000 ;
	    RECT 66.8000 257.8000 67.6000 260.4000 ;
	    RECT 70.0000 255.8000 70.8000 260.4000 ;
	    RECT 75.4000 257.8000 76.4000 260.4000 ;
	    RECT 78.8000 257.8000 79.6000 260.4000 ;
	    RECT 84.4000 256.0000 85.2000 260.4000 ;
	    RECT 87.6000 255.8000 88.4000 260.4000 ;
	    RECT 95.6000 256.6000 96.4000 260.4000 ;
	    RECT 100.4000 255.4000 101.2000 260.4000 ;
	    RECT 105.6000 255.0000 106.4000 260.4000 ;
	    RECT 119.6000 256.6000 120.4000 260.4000 ;
	    RECT 124.4000 255.4000 125.2000 260.4000 ;
	    RECT 129.6000 255.0000 130.4000 260.4000 ;
	    RECT 132.4000 257.8000 133.2000 260.4000 ;
	    RECT 135.6000 257.8000 136.4000 260.4000 ;
	    RECT 137.2000 257.8000 138.0000 260.4000 ;
	    RECT 140.4000 257.8000 141.2000 260.4000 ;
	    RECT 143.6000 256.0000 144.4000 260.4000 ;
	    RECT 149.2000 257.8000 150.0000 260.4000 ;
	    RECT 152.4000 257.8000 153.4000 260.4000 ;
	    RECT 158.0000 255.8000 158.8000 260.4000 ;
	    RECT 162.8000 256.6000 163.6000 260.4000 ;
	    RECT 170.8000 256.6000 171.6000 260.4000 ;
	    RECT 175.6000 255.8000 176.4000 260.4000 ;
	    RECT 180.4000 255.8000 181.2000 260.4000 ;
	    RECT 185.2000 255.8000 186.0000 260.4000 ;
	    RECT 190.0000 255.8000 190.8000 260.4000 ;
	    RECT 196.4000 256.6000 197.2000 260.4000 ;
	    RECT 201.2000 255.8000 202.0000 260.4000 ;
	    RECT 205.6000 255.0000 206.4000 260.4000 ;
	    RECT 210.8000 255.4000 211.6000 260.4000 ;
	    RECT 215.6000 255.4000 216.4000 260.4000 ;
	    RECT 220.8000 255.0000 221.6000 260.4000 ;
	    RECT 228.4000 256.6000 229.2000 260.4000 ;
	    RECT 234.8000 256.6000 235.6000 260.4000 ;
	    RECT 239.6000 256.6000 240.4000 260.4000 ;
	    RECT 249.2000 256.6000 250.0000 260.4000 ;
	    RECT 252.4000 257.8000 253.2000 260.4000 ;
	    RECT 255.6000 257.8000 256.4000 260.4000 ;
	    RECT 263.6000 257.8000 264.4000 260.4000 ;
	    RECT 266.8000 257.8000 267.6000 260.4000 ;
	    RECT 270.0000 255.8000 270.8000 260.4000 ;
	    RECT 274.8000 256.0000 275.6000 260.4000 ;
	    RECT 280.4000 257.8000 281.2000 260.4000 ;
	    RECT 283.6000 257.8000 284.6000 260.4000 ;
	    RECT 289.2000 255.8000 290.0000 260.4000 ;
	    RECT 292.4000 255.8000 293.2000 260.4000 ;
	    RECT 300.4000 256.6000 301.2000 260.4000 ;
	    RECT 305.2000 255.8000 306.0000 260.4000 ;
	    RECT 310.0000 255.8000 310.8000 260.4000 ;
	    RECT 314.8000 256.0000 315.6000 260.4000 ;
	    RECT 320.4000 257.8000 321.2000 260.4000 ;
	    RECT 323.6000 257.8000 324.6000 260.4000 ;
	    RECT 329.2000 255.8000 330.0000 260.4000 ;
	    RECT 332.4000 255.8000 333.2000 260.4000 ;
	    RECT 340.4000 256.6000 341.2000 260.4000 ;
	    RECT 345.2000 255.8000 346.0000 260.4000 ;
	    RECT 350.0000 256.2000 350.8000 260.4000 ;
	    RECT 353.2000 257.8000 354.0000 260.4000 ;
	    RECT 356.4000 256.0000 357.2000 260.4000 ;
	    RECT 362.0000 257.8000 362.8000 260.4000 ;
	    RECT 365.2000 257.8000 366.2000 260.4000 ;
	    RECT 370.8000 255.8000 371.6000 260.4000 ;
	    RECT 375.6000 256.0000 376.4000 260.4000 ;
	    RECT 381.2000 257.8000 382.0000 260.4000 ;
	    RECT 384.4000 257.8000 385.4000 260.4000 ;
	    RECT 390.0000 255.8000 390.8000 260.4000 ;
	    RECT 394.8000 256.0000 395.6000 260.4000 ;
	    RECT 400.4000 257.8000 401.2000 260.4000 ;
	    RECT 403.6000 257.8000 404.6000 260.4000 ;
	    RECT 409.2000 255.8000 410.0000 260.4000 ;
	    RECT 422.0000 256.6000 422.8000 260.4000 ;
	    RECT 426.8000 255.8000 427.6000 260.4000 ;
	    RECT 430.0000 256.0000 430.8000 260.4000 ;
	    RECT 435.6000 257.8000 436.4000 260.4000 ;
	    RECT 438.8000 257.8000 439.8000 260.4000 ;
	    RECT 444.4000 255.8000 445.2000 260.4000 ;
	    RECT 447.6000 257.8000 448.4000 260.4000 ;
	    RECT 452.4000 256.0000 453.2000 260.4000 ;
	    RECT 458.0000 257.8000 458.8000 260.4000 ;
	    RECT 461.2000 257.8000 462.2000 260.4000 ;
	    RECT 466.8000 255.8000 467.6000 260.4000 ;
	    RECT 470.0000 257.8000 470.8000 260.4000 ;
	    RECT 474.8000 256.6000 475.6000 260.4000 ;
	    RECT 481.2000 256.0000 482.0000 260.4000 ;
	    RECT 486.8000 257.8000 487.6000 260.4000 ;
	    RECT 490.0000 257.8000 491.0000 260.4000 ;
	    RECT 495.6000 255.8000 496.4000 260.4000 ;
	    RECT 503.6000 253.8000 504.4000 260.4000 ;
	    RECT 508.4000 256.6000 509.2000 260.4000 ;
	    RECT 513.2000 257.8000 514.0000 260.4000 ;
	    RECT 2.8000 221.6000 3.6000 226.2000 ;
	    RECT 7.6000 221.6000 8.4000 226.2000 ;
	    RECT 12.4000 221.6000 13.2000 225.4000 ;
	    RECT 18.8000 221.6000 19.6000 225.4000 ;
	    RECT 25.2000 221.6000 26.0000 226.0000 ;
	    RECT 30.8000 221.6000 31.6000 224.2000 ;
	    RECT 34.0000 221.6000 35.0000 224.2000 ;
	    RECT 39.6000 221.6000 40.4000 226.2000 ;
	    RECT 44.4000 221.6000 45.2000 225.4000 ;
	    RECT 52.4000 221.6000 53.2000 225.4000 ;
	    RECT 58.8000 221.6000 59.6000 225.4000 ;
	    RECT 63.6000 221.6000 64.4000 226.0000 ;
	    RECT 69.2000 221.6000 70.0000 224.2000 ;
	    RECT 72.4000 221.6000 73.4000 224.2000 ;
	    RECT 78.0000 221.6000 78.8000 226.2000 ;
	    RECT 84.4000 221.6000 85.2000 225.4000 ;
	    RECT 90.8000 221.6000 91.6000 225.4000 ;
	    RECT 97.2000 221.6000 98.0000 225.4000 ;
	    RECT 108.4000 221.6000 109.2000 226.2000 ;
	    RECT 113.8000 221.6000 114.8000 224.2000 ;
	    RECT 117.2000 221.6000 118.0000 224.2000 ;
	    RECT 122.8000 221.6000 123.6000 226.0000 ;
	    RECT 130.8000 221.6000 131.6000 225.4000 ;
	    RECT 137.2000 221.6000 138.0000 225.4000 ;
	    RECT 142.0000 221.6000 142.8000 225.4000 ;
	    RECT 146.8000 221.6000 147.6000 224.2000 ;
	    RECT 150.0000 221.6000 150.8000 224.2000 ;
	    RECT 151.6000 221.6000 152.4000 224.2000 ;
	    RECT 154.8000 221.6000 155.6000 224.2000 ;
	    RECT 157.6000 221.6000 158.4000 227.0000 ;
	    RECT 162.8000 221.6000 163.6000 226.6000 ;
	    RECT 170.8000 221.6000 171.6000 225.4000 ;
	    RECT 174.0000 221.6000 174.8000 224.2000 ;
	    RECT 177.2000 221.6000 178.0000 224.2000 ;
	    RECT 182.0000 221.6000 182.8000 225.4000 ;
	    RECT 185.2000 221.6000 186.0000 226.2000 ;
	    RECT 193.2000 221.6000 194.0000 225.4000 ;
	    RECT 198.0000 221.6000 198.8000 226.2000 ;
	    RECT 201.2000 221.6000 202.0000 224.2000 ;
	    RECT 204.4000 221.6000 205.2000 224.2000 ;
	    RECT 210.8000 221.6000 211.6000 225.4000 ;
	    RECT 217.2000 221.6000 218.0000 225.4000 ;
	    RECT 225.2000 221.6000 226.0000 225.4000 ;
	    RECT 231.6000 221.6000 232.4000 225.4000 ;
	    RECT 234.8000 221.6000 235.6000 224.2000 ;
	    RECT 238.0000 221.6000 238.8000 224.2000 ;
	    RECT 241.2000 221.6000 242.0000 226.2000 ;
	    RECT 246.0000 221.6000 246.8000 226.2000 ;
	    RECT 250.8000 221.6000 251.6000 226.2000 ;
	    RECT 265.2000 221.6000 266.0000 225.4000 ;
	    RECT 271.6000 221.6000 272.4000 225.4000 ;
	    RECT 274.8000 221.6000 275.6000 224.2000 ;
	    RECT 278.0000 221.6000 278.8000 224.2000 ;
	    RECT 281.2000 221.6000 282.0000 225.4000 ;
	    RECT 290.8000 221.6000 291.6000 225.4000 ;
	    RECT 294.0000 221.6000 294.8000 224.2000 ;
	    RECT 297.2000 221.6000 298.0000 224.2000 ;
	    RECT 300.4000 221.6000 301.2000 226.2000 ;
	    RECT 303.6000 221.6000 304.4000 226.6000 ;
	    RECT 308.8000 221.6000 309.6000 227.0000 ;
	    RECT 313.2000 221.6000 314.0000 226.6000 ;
	    RECT 318.4000 221.6000 319.2000 227.0000 ;
	    RECT 322.8000 221.6000 323.6000 226.2000 ;
	    RECT 327.6000 221.6000 328.4000 226.0000 ;
	    RECT 333.2000 221.6000 334.0000 224.2000 ;
	    RECT 336.4000 221.6000 337.4000 224.2000 ;
	    RECT 342.0000 221.6000 342.8000 226.2000 ;
	    RECT 346.8000 221.6000 347.6000 225.4000 ;
	    RECT 354.8000 221.6000 355.6000 225.4000 ;
	    RECT 359.6000 221.6000 360.4000 226.2000 ;
	    RECT 364.4000 221.6000 365.2000 226.0000 ;
	    RECT 370.0000 221.6000 370.8000 224.2000 ;
	    RECT 373.2000 221.6000 374.2000 224.2000 ;
	    RECT 378.8000 221.6000 379.6000 226.2000 ;
	    RECT 382.0000 221.6000 382.8000 224.2000 ;
	    RECT 386.8000 221.6000 387.6000 225.4000 ;
	    RECT 393.2000 221.6000 394.0000 226.2000 ;
	    RECT 396.4000 221.6000 397.2000 226.2000 ;
	    RECT 404.4000 221.6000 405.2000 225.4000 ;
	    RECT 415.6000 221.6000 416.4000 226.0000 ;
	    RECT 421.2000 221.6000 422.0000 224.2000 ;
	    RECT 424.4000 221.6000 425.4000 224.2000 ;
	    RECT 430.0000 221.6000 430.8000 226.2000 ;
	    RECT 438.0000 221.6000 438.8000 228.2000 ;
	    RECT 444.4000 221.6000 445.2000 228.2000 ;
	    RECT 447.6000 221.6000 448.4000 226.2000 ;
	    RECT 454.0000 221.6000 454.8000 225.4000 ;
	    RECT 458.8000 221.6000 459.6000 224.2000 ;
	    RECT 462.0000 221.6000 462.8000 226.0000 ;
	    RECT 467.6000 221.6000 468.4000 224.2000 ;
	    RECT 470.8000 221.6000 471.8000 224.2000 ;
	    RECT 476.4000 221.6000 477.2000 226.2000 ;
	    RECT 484.4000 221.6000 485.2000 228.2000 ;
	    RECT 489.2000 221.6000 490.0000 225.4000 ;
	    RECT 494.0000 221.6000 494.8000 224.2000 ;
	    RECT 497.2000 221.6000 498.0000 226.2000 ;
	    RECT 502.6000 221.6000 503.6000 224.2000 ;
	    RECT 506.0000 221.6000 506.8000 224.2000 ;
	    RECT 511.6000 221.6000 512.4000 226.0000 ;
	    RECT 0.4000 220.4000 514.8000 221.6000 ;
	    RECT 2.8000 215.8000 3.6000 220.4000 ;
	    RECT 7.6000 215.8000 8.4000 220.4000 ;
	    RECT 12.4000 216.6000 13.2000 220.4000 ;
	    RECT 18.8000 216.0000 19.6000 220.4000 ;
	    RECT 24.4000 217.8000 25.2000 220.4000 ;
	    RECT 27.6000 217.8000 28.6000 220.4000 ;
	    RECT 33.2000 215.8000 34.0000 220.4000 ;
	    RECT 39.6000 216.6000 40.4000 220.4000 ;
	    RECT 44.4000 215.8000 45.2000 220.4000 ;
	    RECT 50.8000 216.6000 51.6000 220.4000 ;
	    RECT 54.0000 217.8000 54.8000 220.4000 ;
	    RECT 57.2000 217.8000 58.0000 220.4000 ;
	    RECT 58.8000 217.8000 59.6000 220.4000 ;
	    RECT 62.0000 217.8000 62.8000 220.4000 ;
	    RECT 65.2000 215.8000 66.0000 220.4000 ;
	    RECT 70.0000 215.8000 70.8000 220.4000 ;
	    RECT 74.8000 215.8000 75.6000 220.4000 ;
	    RECT 80.2000 217.8000 81.2000 220.4000 ;
	    RECT 83.6000 217.8000 84.4000 220.4000 ;
	    RECT 89.2000 216.0000 90.0000 220.4000 ;
	    RECT 92.4000 215.8000 93.2000 220.4000 ;
	    RECT 97.2000 215.8000 98.0000 220.4000 ;
	    RECT 105.2000 216.6000 106.0000 220.4000 ;
	    RECT 119.6000 216.6000 120.4000 220.4000 ;
	    RECT 126.0000 216.6000 126.8000 220.4000 ;
	    RECT 130.8000 215.8000 131.6000 220.4000 ;
	    RECT 136.2000 217.8000 137.2000 220.4000 ;
	    RECT 139.6000 217.8000 140.4000 220.4000 ;
	    RECT 145.2000 216.0000 146.0000 220.4000 ;
	    RECT 148.4000 217.8000 149.2000 220.4000 ;
	    RECT 151.6000 217.8000 152.4000 220.4000 ;
	    RECT 154.4000 215.0000 155.2000 220.4000 ;
	    RECT 159.6000 215.4000 160.4000 220.4000 ;
	    RECT 164.4000 215.8000 165.2000 220.4000 ;
	    RECT 169.2000 215.8000 170.0000 220.4000 ;
	    RECT 174.6000 217.8000 175.6000 220.4000 ;
	    RECT 178.0000 217.8000 178.8000 220.4000 ;
	    RECT 183.6000 216.0000 184.4000 220.4000 ;
	    RECT 188.4000 215.8000 189.2000 220.4000 ;
	    RECT 193.2000 215.8000 194.0000 220.4000 ;
	    RECT 196.4000 215.8000 197.2000 220.4000 ;
	    RECT 204.4000 216.6000 205.2000 220.4000 ;
	    RECT 207.6000 217.8000 208.4000 220.4000 ;
	    RECT 210.8000 217.8000 211.6000 220.4000 ;
	    RECT 212.4000 215.8000 213.2000 220.4000 ;
	    RECT 220.4000 216.6000 221.2000 220.4000 ;
	    RECT 225.2000 215.8000 226.0000 220.4000 ;
	    RECT 230.6000 217.8000 231.6000 220.4000 ;
	    RECT 234.0000 217.8000 234.8000 220.4000 ;
	    RECT 239.6000 216.0000 240.4000 220.4000 ;
	    RECT 244.0000 215.0000 244.8000 220.4000 ;
	    RECT 249.2000 215.4000 250.0000 220.4000 ;
	    RECT 260.0000 215.0000 260.8000 220.4000 ;
	    RECT 265.2000 215.4000 266.0000 220.4000 ;
	    RECT 270.0000 215.8000 270.8000 220.4000 ;
	    RECT 274.8000 215.8000 275.6000 220.4000 ;
	    RECT 278.0000 215.8000 278.8000 220.4000 ;
	    RECT 286.0000 216.6000 286.8000 220.4000 ;
	    RECT 290.8000 216.0000 291.6000 220.4000 ;
	    RECT 296.4000 217.8000 297.2000 220.4000 ;
	    RECT 299.6000 217.8000 300.6000 220.4000 ;
	    RECT 305.2000 215.8000 306.0000 220.4000 ;
	    RECT 310.0000 215.4000 310.8000 220.4000 ;
	    RECT 315.2000 215.0000 316.0000 220.4000 ;
	    RECT 319.6000 215.4000 320.4000 220.4000 ;
	    RECT 324.8000 215.0000 325.6000 220.4000 ;
	    RECT 329.2000 216.0000 330.0000 220.4000 ;
	    RECT 334.8000 217.8000 335.6000 220.4000 ;
	    RECT 338.0000 217.8000 339.0000 220.4000 ;
	    RECT 343.6000 215.8000 344.4000 220.4000 ;
	    RECT 348.4000 216.6000 349.2000 220.4000 ;
	    RECT 356.4000 216.6000 357.2000 220.4000 ;
	    RECT 361.2000 215.8000 362.0000 220.4000 ;
	    RECT 366.0000 216.0000 366.8000 220.4000 ;
	    RECT 371.6000 217.8000 372.4000 220.4000 ;
	    RECT 374.8000 217.8000 375.8000 220.4000 ;
	    RECT 380.4000 215.8000 381.2000 220.4000 ;
	    RECT 383.6000 215.8000 384.4000 220.4000 ;
	    RECT 391.6000 216.6000 392.4000 220.4000 ;
	    RECT 396.4000 215.8000 397.2000 220.4000 ;
	    RECT 399.6000 215.8000 400.4000 220.4000 ;
	    RECT 414.0000 216.6000 414.8000 220.4000 ;
	    RECT 418.8000 216.0000 419.6000 220.4000 ;
	    RECT 424.4000 217.8000 425.2000 220.4000 ;
	    RECT 427.6000 217.8000 428.6000 220.4000 ;
	    RECT 433.2000 215.8000 434.0000 220.4000 ;
	    RECT 438.0000 215.8000 438.8000 220.4000 ;
	    RECT 442.8000 215.8000 443.6000 220.4000 ;
	    RECT 444.4000 213.8000 445.2000 220.4000 ;
	    RECT 450.8000 215.8000 451.6000 220.4000 ;
	    RECT 454.0000 215.8000 454.8000 220.4000 ;
	    RECT 457.2000 215.8000 458.0000 220.4000 ;
	    RECT 460.4000 216.0000 461.2000 220.4000 ;
	    RECT 466.0000 217.8000 466.8000 220.4000 ;
	    RECT 469.2000 217.8000 470.2000 220.4000 ;
	    RECT 474.8000 215.8000 475.6000 220.4000 ;
	    RECT 481.2000 216.6000 482.0000 220.4000 ;
	    RECT 484.4000 217.8000 485.2000 220.4000 ;
	    RECT 489.2000 216.6000 490.0000 220.4000 ;
	    RECT 495.6000 216.0000 496.4000 220.4000 ;
	    RECT 501.2000 217.8000 502.0000 220.4000 ;
	    RECT 504.4000 217.8000 505.4000 220.4000 ;
	    RECT 510.0000 215.8000 510.8000 220.4000 ;
	    RECT 2.8000 181.6000 3.6000 186.2000 ;
	    RECT 7.6000 181.6000 8.4000 186.2000 ;
	    RECT 12.4000 181.6000 13.2000 186.2000 ;
	    RECT 17.2000 181.6000 18.0000 185.4000 ;
	    RECT 23.6000 181.6000 24.4000 186.0000 ;
	    RECT 29.2000 181.6000 30.0000 184.2000 ;
	    RECT 32.4000 181.6000 33.4000 184.2000 ;
	    RECT 38.0000 181.6000 38.8000 186.2000 ;
	    RECT 42.8000 181.6000 43.6000 186.2000 ;
	    RECT 49.2000 181.6000 50.0000 185.4000 ;
	    RECT 55.6000 181.6000 56.4000 185.4000 ;
	    RECT 62.0000 181.6000 62.8000 185.4000 ;
	    RECT 65.2000 181.6000 66.0000 184.2000 ;
	    RECT 68.4000 181.6000 69.2000 184.2000 ;
	    RECT 71.6000 181.6000 72.4000 186.2000 ;
	    RECT 77.0000 181.6000 78.0000 184.2000 ;
	    RECT 80.4000 181.6000 81.2000 184.2000 ;
	    RECT 86.0000 181.6000 86.8000 186.0000 ;
	    RECT 90.8000 181.6000 91.6000 186.2000 ;
	    RECT 95.6000 181.6000 96.4000 185.4000 ;
	    RECT 103.6000 181.6000 104.4000 185.4000 ;
	    RECT 114.4000 181.6000 115.2000 187.0000 ;
	    RECT 119.6000 181.6000 120.4000 186.6000 ;
	    RECT 124.4000 181.6000 125.2000 186.6000 ;
	    RECT 129.6000 181.6000 130.4000 187.0000 ;
	    RECT 137.2000 181.6000 138.0000 185.4000 ;
	    RECT 142.0000 181.6000 142.8000 185.4000 ;
	    RECT 151.6000 181.6000 152.4000 185.4000 ;
	    RECT 158.0000 181.6000 158.8000 185.4000 ;
	    RECT 161.2000 181.6000 162.0000 184.2000 ;
	    RECT 164.4000 181.6000 165.2000 184.2000 ;
	    RECT 166.0000 181.6000 166.8000 184.2000 ;
	    RECT 169.2000 181.6000 170.0000 184.2000 ;
	    RECT 174.0000 181.6000 174.8000 185.4000 ;
	    RECT 180.4000 181.6000 181.2000 185.4000 ;
	    RECT 185.2000 181.6000 186.0000 185.4000 ;
	    RECT 191.6000 181.6000 192.4000 185.4000 ;
	    RECT 198.0000 181.6000 198.8000 184.2000 ;
	    RECT 201.2000 181.6000 202.0000 184.2000 ;
	    RECT 204.4000 181.6000 205.2000 185.4000 ;
	    RECT 210.8000 181.6000 211.6000 185.4000 ;
	    RECT 217.2000 181.6000 218.0000 184.2000 ;
	    RECT 220.4000 181.6000 221.2000 184.2000 ;
	    RECT 223.6000 181.6000 224.4000 186.2000 ;
	    RECT 228.4000 181.6000 229.2000 186.2000 ;
	    RECT 236.4000 181.6000 237.2000 185.4000 ;
	    RECT 242.8000 181.6000 243.6000 185.4000 ;
	    RECT 249.2000 181.6000 250.0000 185.4000 ;
	    RECT 254.0000 181.6000 254.8000 186.2000 ;
	    RECT 266.8000 181.6000 267.6000 186.2000 ;
	    RECT 270.0000 181.6000 270.8000 186.0000 ;
	    RECT 275.6000 181.6000 276.4000 184.2000 ;
	    RECT 278.8000 181.6000 279.8000 184.2000 ;
	    RECT 284.4000 181.6000 285.2000 186.2000 ;
	    RECT 289.2000 181.6000 290.0000 186.2000 ;
	    RECT 295.6000 181.6000 296.4000 185.4000 ;
	    RECT 300.4000 181.6000 301.2000 186.2000 ;
	    RECT 305.2000 181.6000 306.0000 186.2000 ;
	    RECT 308.4000 181.6000 309.2000 186.2000 ;
	    RECT 316.4000 181.6000 317.2000 185.4000 ;
	    RECT 321.2000 181.6000 322.0000 186.0000 ;
	    RECT 326.8000 181.6000 327.6000 184.2000 ;
	    RECT 330.0000 181.6000 331.0000 184.2000 ;
	    RECT 335.6000 181.6000 336.4000 186.2000 ;
	    RECT 340.4000 181.6000 341.2000 186.2000 ;
	    RECT 345.2000 181.6000 346.0000 186.2000 ;
	    RECT 350.0000 181.6000 350.8000 186.2000 ;
	    RECT 353.2000 181.6000 354.0000 186.2000 ;
	    RECT 361.2000 181.6000 362.0000 185.4000 ;
	    RECT 366.0000 181.6000 366.8000 186.0000 ;
	    RECT 371.6000 181.6000 372.4000 184.2000 ;
	    RECT 374.8000 181.6000 375.8000 184.2000 ;
	    RECT 380.4000 181.6000 381.2000 186.2000 ;
	    RECT 383.6000 181.6000 384.4000 184.2000 ;
	    RECT 388.4000 181.6000 389.2000 186.0000 ;
	    RECT 394.0000 181.6000 394.8000 184.2000 ;
	    RECT 397.2000 181.6000 398.2000 184.2000 ;
	    RECT 402.8000 181.6000 403.6000 186.2000 ;
	    RECT 414.0000 181.6000 414.8000 185.4000 ;
	    RECT 420.4000 181.6000 421.2000 186.2000 ;
	    RECT 425.2000 181.6000 426.0000 186.2000 ;
	    RECT 428.4000 181.6000 429.2000 188.2000 ;
	    RECT 438.0000 181.6000 438.8000 186.2000 ;
	    RECT 442.8000 181.6000 443.6000 186.2000 ;
	    RECT 446.0000 181.6000 446.8000 186.2000 ;
	    RECT 449.2000 181.6000 450.0000 186.2000 ;
	    RECT 454.0000 181.6000 454.8000 186.2000 ;
	    RECT 460.4000 181.6000 461.2000 188.2000 ;
	    RECT 466.8000 181.6000 467.6000 188.2000 ;
	    RECT 473.2000 181.6000 474.0000 188.2000 ;
	    RECT 474.8000 181.6000 475.6000 184.2000 ;
	    RECT 479.6000 181.6000 480.4000 185.4000 ;
	    RECT 486.0000 181.6000 486.8000 186.0000 ;
	    RECT 491.6000 181.6000 492.4000 184.2000 ;
	    RECT 494.8000 181.6000 495.8000 184.2000 ;
	    RECT 500.4000 181.6000 501.2000 186.2000 ;
	    RECT 508.4000 181.6000 509.2000 188.2000 ;
	    RECT 511.6000 181.6000 512.4000 186.2000 ;
	    RECT 0.4000 180.4000 514.8000 181.6000 ;
	    RECT 1.2000 175.8000 2.0000 180.4000 ;
	    RECT 4.4000 175.8000 5.2000 180.4000 ;
	    RECT 7.6000 175.8000 8.4000 180.4000 ;
	    RECT 12.4000 175.8000 13.2000 180.4000 ;
	    RECT 16.6000 176.0000 17.4000 180.4000 ;
	    RECT 20.4000 177.8000 21.2000 180.4000 ;
	    RECT 23.6000 177.8000 24.4000 180.4000 ;
	    RECT 25.2000 175.8000 26.0000 180.4000 ;
	    RECT 33.2000 176.6000 34.0000 180.4000 ;
	    RECT 38.0000 175.8000 38.8000 180.4000 ;
	    RECT 43.4000 177.8000 44.4000 180.4000 ;
	    RECT 46.8000 177.8000 47.6000 180.4000 ;
	    RECT 52.4000 176.0000 53.2000 180.4000 ;
	    RECT 57.2000 176.0000 58.0000 180.4000 ;
	    RECT 62.8000 177.8000 63.6000 180.4000 ;
	    RECT 66.0000 177.8000 67.0000 180.4000 ;
	    RECT 71.6000 175.8000 72.4000 180.4000 ;
	    RECT 74.8000 175.8000 75.6000 180.4000 ;
	    RECT 82.8000 176.6000 83.6000 180.4000 ;
	    RECT 87.6000 175.8000 88.4000 180.4000 ;
	    RECT 93.0000 177.8000 94.0000 180.4000 ;
	    RECT 96.4000 177.8000 97.2000 180.4000 ;
	    RECT 102.0000 176.0000 102.8000 180.4000 ;
	    RECT 113.2000 176.6000 114.0000 180.4000 ;
	    RECT 121.2000 175.8000 122.0000 180.4000 ;
	    RECT 124.4000 176.0000 125.2000 180.4000 ;
	    RECT 130.0000 177.8000 130.8000 180.4000 ;
	    RECT 133.2000 177.8000 134.2000 180.4000 ;
	    RECT 138.8000 175.8000 139.6000 180.4000 ;
	    RECT 142.0000 175.8000 142.8000 180.4000 ;
	    RECT 150.0000 176.6000 150.8000 180.4000 ;
	    RECT 154.8000 175.8000 155.6000 180.4000 ;
	    RECT 159.6000 176.0000 160.4000 180.4000 ;
	    RECT 165.2000 177.8000 166.0000 180.4000 ;
	    RECT 168.4000 177.8000 169.4000 180.4000 ;
	    RECT 174.0000 175.8000 174.8000 180.4000 ;
	    RECT 178.8000 175.8000 179.6000 180.4000 ;
	    RECT 183.2000 175.0000 184.0000 180.4000 ;
	    RECT 188.4000 175.4000 189.2000 180.4000 ;
	    RECT 192.8000 175.0000 193.6000 180.4000 ;
	    RECT 198.0000 175.4000 198.8000 180.4000 ;
	    RECT 202.8000 175.8000 203.6000 180.4000 ;
	    RECT 206.0000 175.8000 206.8000 180.4000 ;
	    RECT 209.2000 175.8000 210.0000 180.4000 ;
	    RECT 212.4000 175.8000 213.2000 180.4000 ;
	    RECT 214.0000 175.8000 214.8000 180.4000 ;
	    RECT 222.0000 176.6000 222.8000 180.4000 ;
	    RECT 226.8000 176.0000 227.6000 180.4000 ;
	    RECT 232.4000 177.8000 233.2000 180.4000 ;
	    RECT 235.6000 177.8000 236.6000 180.4000 ;
	    RECT 241.2000 175.8000 242.0000 180.4000 ;
	    RECT 249.2000 176.6000 250.0000 180.4000 ;
	    RECT 252.4000 177.8000 253.2000 180.4000 ;
	    RECT 255.6000 177.8000 256.4000 180.4000 ;
	    RECT 263.6000 177.8000 264.4000 180.4000 ;
	    RECT 266.8000 177.8000 267.6000 180.4000 ;
	    RECT 270.0000 176.0000 270.8000 180.4000 ;
	    RECT 275.6000 177.8000 276.4000 180.4000 ;
	    RECT 278.8000 177.8000 279.8000 180.4000 ;
	    RECT 284.4000 175.8000 285.2000 180.4000 ;
	    RECT 289.2000 176.6000 290.0000 180.4000 ;
	    RECT 297.2000 176.6000 298.0000 180.4000 ;
	    RECT 302.0000 175.8000 302.8000 180.4000 ;
	    RECT 307.4000 177.8000 308.4000 180.4000 ;
	    RECT 310.8000 177.8000 311.6000 180.4000 ;
	    RECT 316.4000 176.0000 317.2000 180.4000 ;
	    RECT 319.6000 177.8000 320.4000 180.4000 ;
	    RECT 322.8000 177.8000 323.6000 180.4000 ;
	    RECT 326.0000 175.8000 326.8000 180.4000 ;
	    RECT 330.8000 175.8000 331.6000 180.4000 ;
	    RECT 333.6000 175.0000 334.4000 180.4000 ;
	    RECT 338.8000 175.4000 339.6000 180.4000 ;
	    RECT 343.2000 175.0000 344.0000 180.4000 ;
	    RECT 348.4000 175.4000 349.2000 180.4000 ;
	    RECT 352.8000 175.0000 353.6000 180.4000 ;
	    RECT 358.0000 175.4000 358.8000 180.4000 ;
	    RECT 362.4000 175.0000 363.2000 180.4000 ;
	    RECT 367.6000 175.4000 368.4000 180.4000 ;
	    RECT 372.4000 175.8000 373.2000 180.4000 ;
	    RECT 375.6000 175.8000 376.4000 180.4000 ;
	    RECT 378.8000 175.8000 379.6000 180.4000 ;
	    RECT 382.0000 175.8000 382.8000 180.4000 ;
	    RECT 385.2000 175.8000 386.0000 180.4000 ;
	    RECT 388.4000 175.8000 389.2000 180.4000 ;
	    RECT 393.2000 175.8000 394.0000 180.4000 ;
	    RECT 396.4000 176.0000 397.2000 180.4000 ;
	    RECT 402.0000 177.8000 402.8000 180.4000 ;
	    RECT 405.2000 177.8000 406.2000 180.4000 ;
	    RECT 410.8000 175.8000 411.6000 180.4000 ;
	    RECT 423.6000 176.6000 424.4000 180.4000 ;
	    RECT 430.0000 175.8000 430.8000 180.4000 ;
	    RECT 433.2000 177.8000 434.0000 180.4000 ;
	    RECT 439.6000 173.8000 440.4000 180.4000 ;
	    RECT 442.8000 177.8000 443.6000 180.4000 ;
	    RECT 444.4000 177.8000 445.2000 180.4000 ;
	    RECT 447.6000 177.8000 448.4000 180.4000 ;
	    RECT 449.2000 177.8000 450.0000 180.4000 ;
	    RECT 452.4000 177.8000 453.2000 180.4000 ;
	    RECT 455.6000 175.8000 456.4000 180.4000 ;
	    RECT 458.8000 173.8000 459.6000 180.4000 ;
	    RECT 466.8000 175.8000 467.6000 180.4000 ;
	    RECT 471.6000 175.8000 472.4000 180.4000 ;
	    RECT 479.6000 173.8000 480.4000 180.4000 ;
	    RECT 482.8000 175.8000 483.6000 180.4000 ;
	    RECT 487.6000 176.0000 488.4000 180.4000 ;
	    RECT 493.2000 177.8000 494.0000 180.4000 ;
	    RECT 496.4000 177.8000 497.4000 180.4000 ;
	    RECT 502.0000 175.8000 502.8000 180.4000 ;
	    RECT 505.2000 177.8000 506.0000 180.4000 ;
	    RECT 510.0000 176.6000 510.8000 180.4000 ;
	    RECT 2.8000 141.6000 3.6000 146.2000 ;
	    RECT 7.6000 141.6000 8.4000 146.2000 ;
	    RECT 12.4000 141.6000 13.2000 146.2000 ;
	    RECT 17.2000 141.6000 18.0000 145.4000 ;
	    RECT 23.6000 141.6000 24.4000 146.0000 ;
	    RECT 29.2000 141.6000 30.0000 144.2000 ;
	    RECT 32.4000 141.6000 33.4000 144.2000 ;
	    RECT 38.0000 141.6000 38.8000 146.2000 ;
	    RECT 42.8000 141.6000 43.6000 146.2000 ;
	    RECT 48.2000 141.6000 49.2000 144.2000 ;
	    RECT 51.6000 141.6000 52.4000 144.2000 ;
	    RECT 57.2000 141.6000 58.0000 146.0000 ;
	    RECT 62.0000 141.6000 62.8000 146.2000 ;
	    RECT 67.4000 141.6000 68.4000 144.2000 ;
	    RECT 70.8000 141.6000 71.6000 144.2000 ;
	    RECT 76.4000 141.6000 77.2000 146.0000 ;
	    RECT 81.2000 141.6000 82.0000 146.2000 ;
	    RECT 84.4000 141.6000 85.2000 146.2000 ;
	    RECT 92.4000 141.6000 93.2000 145.4000 ;
	    RECT 97.2000 141.6000 98.0000 145.4000 ;
	    RECT 105.2000 141.6000 106.0000 145.4000 ;
	    RECT 116.0000 141.6000 116.8000 147.0000 ;
	    RECT 121.2000 141.6000 122.0000 146.6000 ;
	    RECT 124.4000 141.6000 125.2000 144.2000 ;
	    RECT 127.6000 141.6000 128.4000 144.2000 ;
	    RECT 129.2000 141.6000 130.0000 144.2000 ;
	    RECT 132.4000 141.6000 133.2000 144.2000 ;
	    RECT 135.6000 141.6000 136.4000 145.4000 ;
	    RECT 143.6000 141.6000 144.4000 146.2000 ;
	    RECT 146.8000 141.6000 147.6000 145.4000 ;
	    RECT 153.2000 141.6000 154.0000 145.4000 ;
	    RECT 159.6000 141.6000 160.4000 144.2000 ;
	    RECT 162.8000 141.6000 163.6000 144.2000 ;
	    RECT 164.4000 141.6000 165.2000 144.2000 ;
	    RECT 167.6000 141.6000 168.4000 144.2000 ;
	    RECT 170.8000 141.6000 171.6000 145.4000 ;
	    RECT 177.2000 141.6000 178.0000 145.4000 ;
	    RECT 183.6000 141.6000 184.4000 144.2000 ;
	    RECT 186.8000 141.6000 187.6000 144.2000 ;
	    RECT 191.6000 141.6000 192.4000 145.4000 ;
	    RECT 198.0000 141.6000 198.8000 145.4000 ;
	    RECT 202.8000 141.6000 203.6000 146.0000 ;
	    RECT 208.4000 141.6000 209.2000 144.2000 ;
	    RECT 211.6000 141.6000 212.6000 144.2000 ;
	    RECT 217.2000 141.6000 218.0000 146.2000 ;
	    RECT 222.0000 141.6000 222.8000 146.2000 ;
	    RECT 225.2000 141.6000 226.0000 144.2000 ;
	    RECT 228.4000 141.6000 229.2000 144.2000 ;
	    RECT 231.6000 141.6000 232.4000 146.2000 ;
	    RECT 236.4000 141.6000 237.2000 146.2000 ;
	    RECT 241.8000 141.6000 242.8000 144.2000 ;
	    RECT 245.2000 141.6000 246.0000 144.2000 ;
	    RECT 250.8000 141.6000 251.6000 146.0000 ;
	    RECT 262.0000 141.6000 262.8000 146.2000 ;
	    RECT 266.8000 141.6000 267.6000 145.4000 ;
	    RECT 273.2000 141.6000 274.0000 146.2000 ;
	    RECT 279.6000 141.6000 280.4000 145.4000 ;
	    RECT 284.4000 141.6000 285.2000 146.2000 ;
	    RECT 287.6000 141.6000 288.4000 144.2000 ;
	    RECT 290.8000 141.6000 291.6000 144.2000 ;
	    RECT 294.0000 141.6000 294.8000 145.4000 ;
	    RECT 303.6000 141.6000 304.4000 145.4000 ;
	    RECT 310.0000 141.6000 310.8000 145.4000 ;
	    RECT 314.8000 141.6000 315.6000 145.4000 ;
	    RECT 321.2000 141.6000 322.0000 144.2000 ;
	    RECT 324.4000 141.6000 325.2000 144.2000 ;
	    RECT 327.6000 141.6000 328.4000 145.4000 ;
	    RECT 337.2000 141.6000 338.0000 145.4000 ;
	    RECT 340.4000 141.6000 341.2000 144.2000 ;
	    RECT 343.6000 141.6000 344.4000 144.2000 ;
	    RECT 346.8000 141.6000 347.6000 145.4000 ;
	    RECT 356.4000 141.6000 357.2000 145.4000 ;
	    RECT 361.2000 141.6000 362.0000 145.4000 ;
	    RECT 366.0000 141.6000 366.8000 146.2000 ;
	    RECT 374.0000 141.6000 374.8000 145.4000 ;
	    RECT 378.8000 141.6000 379.6000 146.0000 ;
	    RECT 384.4000 141.6000 385.2000 144.2000 ;
	    RECT 387.6000 141.6000 388.6000 144.2000 ;
	    RECT 393.2000 141.6000 394.0000 146.2000 ;
	    RECT 399.6000 141.6000 400.4000 145.4000 ;
	    RECT 410.8000 141.6000 411.6000 146.0000 ;
	    RECT 416.4000 141.6000 417.2000 144.2000 ;
	    RECT 419.6000 141.6000 420.6000 144.2000 ;
	    RECT 425.2000 141.6000 426.0000 146.2000 ;
	    RECT 430.0000 141.6000 430.8000 146.0000 ;
	    RECT 435.6000 141.6000 436.4000 144.2000 ;
	    RECT 438.8000 141.6000 439.8000 144.2000 ;
	    RECT 444.4000 141.6000 445.2000 146.2000 ;
	    RECT 447.6000 141.6000 448.4000 146.2000 ;
	    RECT 455.6000 141.6000 456.4000 145.4000 ;
	    RECT 460.4000 141.6000 461.2000 146.0000 ;
	    RECT 466.0000 141.6000 466.8000 144.2000 ;
	    RECT 469.2000 141.6000 470.2000 144.2000 ;
	    RECT 474.8000 141.6000 475.6000 146.2000 ;
	    RECT 481.2000 141.6000 482.0000 145.4000 ;
	    RECT 486.0000 141.6000 486.8000 144.2000 ;
	    RECT 490.2000 141.6000 491.0000 146.0000 ;
	    RECT 495.6000 141.6000 496.4000 146.0000 ;
	    RECT 501.2000 141.6000 502.0000 144.2000 ;
	    RECT 504.4000 141.6000 505.4000 144.2000 ;
	    RECT 510.0000 141.6000 510.8000 146.2000 ;
	    RECT 0.4000 140.4000 514.8000 141.6000 ;
	    RECT 2.8000 135.8000 3.6000 140.4000 ;
	    RECT 7.6000 135.8000 8.4000 140.4000 ;
	    RECT 12.4000 136.0000 13.2000 140.4000 ;
	    RECT 18.0000 137.8000 18.8000 140.4000 ;
	    RECT 21.2000 137.8000 22.2000 140.4000 ;
	    RECT 26.8000 135.8000 27.6000 140.4000 ;
	    RECT 33.2000 136.6000 34.0000 140.4000 ;
	    RECT 38.0000 136.6000 38.8000 140.4000 ;
	    RECT 44.4000 136.0000 45.2000 140.4000 ;
	    RECT 50.0000 137.8000 50.8000 140.4000 ;
	    RECT 53.2000 137.8000 54.2000 140.4000 ;
	    RECT 58.8000 135.8000 59.6000 140.4000 ;
	    RECT 65.2000 136.6000 66.0000 140.4000 ;
	    RECT 68.4000 135.8000 69.2000 140.4000 ;
	    RECT 71.6000 135.8000 72.4000 140.4000 ;
	    RECT 76.4000 136.6000 77.2000 140.4000 ;
	    RECT 79.6000 137.8000 80.4000 140.4000 ;
	    RECT 82.8000 137.8000 83.6000 140.4000 ;
	    RECT 87.6000 136.6000 88.4000 140.4000 ;
	    RECT 94.0000 136.6000 94.8000 140.4000 ;
	    RECT 98.8000 136.6000 99.6000 140.4000 ;
	    RECT 111.6000 135.4000 112.4000 140.4000 ;
	    RECT 116.8000 135.0000 117.6000 140.4000 ;
	    RECT 124.4000 136.6000 125.2000 140.4000 ;
	    RECT 130.8000 136.6000 131.6000 140.4000 ;
	    RECT 138.8000 136.6000 139.6000 140.4000 ;
	    RECT 146.8000 136.6000 147.6000 140.4000 ;
	    RECT 151.6000 136.6000 152.4000 140.4000 ;
	    RECT 158.0000 135.8000 158.8000 140.4000 ;
	    RECT 161.2000 137.8000 162.0000 140.4000 ;
	    RECT 164.4000 137.8000 165.2000 140.4000 ;
	    RECT 166.0000 137.8000 166.8000 140.4000 ;
	    RECT 169.2000 137.8000 170.0000 140.4000 ;
	    RECT 170.8000 137.8000 171.6000 140.4000 ;
	    RECT 174.0000 137.8000 174.8000 140.4000 ;
	    RECT 175.6000 137.8000 176.4000 140.4000 ;
	    RECT 178.8000 137.8000 179.6000 140.4000 ;
	    RECT 182.0000 135.8000 182.8000 140.4000 ;
	    RECT 186.8000 135.8000 187.6000 140.4000 ;
	    RECT 191.6000 135.8000 192.4000 140.4000 ;
	    RECT 196.4000 135.8000 197.2000 140.4000 ;
	    RECT 201.2000 136.6000 202.0000 140.4000 ;
	    RECT 207.6000 136.6000 208.4000 140.4000 ;
	    RECT 215.6000 136.6000 216.4000 140.4000 ;
	    RECT 220.4000 136.0000 221.2000 140.4000 ;
	    RECT 226.0000 137.8000 226.8000 140.4000 ;
	    RECT 229.2000 137.8000 230.2000 140.4000 ;
	    RECT 234.8000 135.8000 235.6000 140.4000 ;
	    RECT 239.6000 135.8000 240.4000 140.4000 ;
	    RECT 244.4000 135.8000 245.2000 140.4000 ;
	    RECT 249.2000 136.6000 250.0000 140.4000 ;
	    RECT 263.6000 136.6000 264.4000 140.4000 ;
	    RECT 268.4000 135.8000 269.2000 140.4000 ;
	    RECT 271.6000 135.8000 272.4000 140.4000 ;
	    RECT 274.8000 135.8000 275.6000 140.4000 ;
	    RECT 278.0000 135.8000 278.8000 140.4000 ;
	    RECT 281.2000 135.8000 282.0000 140.4000 ;
	    RECT 284.4000 137.8000 285.2000 140.4000 ;
	    RECT 287.6000 137.8000 288.4000 140.4000 ;
	    RECT 289.2000 137.8000 290.0000 140.4000 ;
	    RECT 292.4000 137.8000 293.2000 140.4000 ;
	    RECT 298.8000 136.6000 299.6000 140.4000 ;
	    RECT 302.0000 137.8000 302.8000 140.4000 ;
	    RECT 305.2000 137.8000 306.0000 140.4000 ;
	    RECT 310.0000 136.6000 310.8000 140.4000 ;
	    RECT 313.2000 137.8000 314.0000 140.4000 ;
	    RECT 316.4000 137.8000 317.2000 140.4000 ;
	    RECT 319.6000 136.6000 320.4000 140.4000 ;
	    RECT 329.2000 136.6000 330.0000 140.4000 ;
	    RECT 334.0000 135.8000 334.8000 140.4000 ;
	    RECT 342.0000 136.6000 342.8000 140.4000 ;
	    RECT 345.2000 137.8000 346.0000 140.4000 ;
	    RECT 348.4000 137.8000 349.2000 140.4000 ;
	    RECT 353.2000 136.6000 354.0000 140.4000 ;
	    RECT 359.6000 136.6000 360.4000 140.4000 ;
	    RECT 364.4000 135.4000 365.2000 140.4000 ;
	    RECT 369.6000 135.0000 370.4000 140.4000 ;
	    RECT 374.0000 135.4000 374.8000 140.4000 ;
	    RECT 379.2000 135.0000 380.0000 140.4000 ;
	    RECT 383.6000 135.8000 384.4000 140.4000 ;
	    RECT 390.0000 136.6000 390.8000 140.4000 ;
	    RECT 394.8000 136.6000 395.6000 140.4000 ;
	    RECT 402.8000 136.6000 403.6000 140.4000 ;
	    RECT 414.0000 136.0000 414.8000 140.4000 ;
	    RECT 419.6000 137.8000 420.4000 140.4000 ;
	    RECT 422.8000 137.8000 423.8000 140.4000 ;
	    RECT 428.4000 135.8000 429.2000 140.4000 ;
	    RECT 434.8000 135.8000 435.6000 140.4000 ;
	    RECT 439.6000 136.6000 440.4000 140.4000 ;
	    RECT 444.4000 136.6000 445.2000 140.4000 ;
	    RECT 452.4000 135.8000 453.2000 140.4000 ;
	    RECT 455.6000 136.0000 456.4000 140.4000 ;
	    RECT 461.2000 137.8000 462.0000 140.4000 ;
	    RECT 464.4000 137.8000 465.4000 140.4000 ;
	    RECT 470.0000 135.8000 470.8000 140.4000 ;
	    RECT 474.8000 136.0000 475.6000 140.4000 ;
	    RECT 480.4000 137.8000 481.2000 140.4000 ;
	    RECT 483.6000 137.8000 484.6000 140.4000 ;
	    RECT 489.2000 135.8000 490.0000 140.4000 ;
	    RECT 492.4000 137.8000 493.2000 140.4000 ;
	    RECT 497.2000 136.6000 498.0000 140.4000 ;
	    RECT 503.6000 136.6000 504.4000 140.4000 ;
	    RECT 508.4000 133.8000 509.2000 140.4000 ;
	    RECT 2.8000 101.6000 3.6000 106.2000 ;
	    RECT 7.6000 101.6000 8.4000 106.0000 ;
	    RECT 13.2000 101.6000 14.0000 104.2000 ;
	    RECT 16.4000 101.6000 17.4000 104.2000 ;
	    RECT 22.0000 101.6000 22.8000 106.2000 ;
	    RECT 26.8000 101.6000 27.6000 105.4000 ;
	    RECT 31.6000 101.6000 32.4000 104.2000 ;
	    RECT 34.8000 101.6000 35.6000 104.2000 ;
	    RECT 38.0000 101.6000 38.8000 106.0000 ;
	    RECT 43.6000 101.6000 44.4000 104.2000 ;
	    RECT 46.8000 101.6000 47.8000 104.2000 ;
	    RECT 52.4000 101.6000 53.2000 106.2000 ;
	    RECT 58.8000 101.6000 59.6000 105.4000 ;
	    RECT 63.6000 101.6000 64.4000 106.2000 ;
	    RECT 69.0000 101.6000 70.0000 104.2000 ;
	    RECT 72.4000 101.6000 73.2000 104.2000 ;
	    RECT 78.0000 101.6000 78.8000 106.0000 ;
	    RECT 81.2000 101.6000 82.0000 106.2000 ;
	    RECT 89.2000 101.6000 90.0000 105.4000 ;
	    RECT 93.6000 101.6000 94.4000 107.0000 ;
	    RECT 98.8000 101.6000 99.6000 106.6000 ;
	    RECT 113.2000 101.6000 114.0000 105.4000 ;
	    RECT 119.6000 101.6000 120.4000 105.4000 ;
	    RECT 124.4000 101.6000 125.2000 106.6000 ;
	    RECT 129.6000 101.6000 130.4000 107.0000 ;
	    RECT 134.0000 101.6000 134.8000 105.4000 ;
	    RECT 140.4000 101.6000 141.2000 106.0000 ;
	    RECT 146.0000 101.6000 146.8000 104.2000 ;
	    RECT 149.2000 101.6000 150.2000 104.2000 ;
	    RECT 154.8000 101.6000 155.6000 106.2000 ;
	    RECT 158.0000 101.6000 158.8000 106.2000 ;
	    RECT 166.0000 101.6000 166.8000 105.4000 ;
	    RECT 169.2000 101.6000 170.0000 104.2000 ;
	    RECT 172.4000 101.6000 173.2000 104.2000 ;
	    RECT 174.0000 101.6000 174.8000 104.2000 ;
	    RECT 177.2000 101.6000 178.0000 104.2000 ;
	    RECT 178.8000 101.6000 179.6000 104.2000 ;
	    RECT 182.0000 101.6000 182.8000 104.2000 ;
	    RECT 183.6000 101.6000 184.4000 104.2000 ;
	    RECT 186.8000 101.6000 187.6000 104.2000 ;
	    RECT 188.4000 101.6000 189.2000 104.2000 ;
	    RECT 191.6000 101.6000 192.4000 104.2000 ;
	    RECT 194.8000 101.6000 195.6000 106.0000 ;
	    RECT 200.4000 101.6000 201.2000 104.2000 ;
	    RECT 203.6000 101.6000 204.6000 104.2000 ;
	    RECT 209.2000 101.6000 210.0000 106.2000 ;
	    RECT 215.6000 101.6000 216.4000 105.4000 ;
	    RECT 218.8000 101.6000 219.6000 104.2000 ;
	    RECT 222.0000 101.6000 222.8000 104.2000 ;
	    RECT 223.6000 101.6000 224.4000 104.2000 ;
	    RECT 226.8000 101.6000 227.6000 104.2000 ;
	    RECT 228.4000 101.6000 229.2000 104.2000 ;
	    RECT 231.6000 101.6000 232.4000 104.2000 ;
	    RECT 233.2000 101.6000 234.0000 104.2000 ;
	    RECT 236.4000 101.6000 237.2000 104.2000 ;
	    RECT 238.0000 101.6000 238.8000 104.2000 ;
	    RECT 241.2000 101.6000 242.0000 104.2000 ;
	    RECT 244.4000 101.6000 245.2000 105.4000 ;
	    RECT 257.2000 101.6000 258.0000 106.2000 ;
	    RECT 262.6000 101.6000 263.6000 104.2000 ;
	    RECT 266.0000 101.6000 266.8000 104.2000 ;
	    RECT 271.6000 101.6000 272.4000 106.0000 ;
	    RECT 276.4000 101.6000 277.2000 106.2000 ;
	    RECT 280.8000 101.6000 281.6000 107.0000 ;
	    RECT 286.0000 101.6000 286.8000 106.6000 ;
	    RECT 290.8000 101.6000 291.6000 106.6000 ;
	    RECT 296.0000 101.6000 296.8000 107.0000 ;
	    RECT 303.6000 101.6000 304.4000 105.4000 ;
	    RECT 308.4000 101.6000 309.2000 105.4000 ;
	    RECT 313.2000 101.6000 314.0000 104.2000 ;
	    RECT 316.4000 101.6000 317.2000 104.2000 ;
	    RECT 319.6000 101.6000 320.4000 105.4000 ;
	    RECT 326.0000 101.6000 326.8000 106.2000 ;
	    RECT 330.8000 101.6000 331.6000 106.2000 ;
	    RECT 335.6000 101.6000 336.4000 106.0000 ;
	    RECT 341.2000 101.6000 342.0000 104.2000 ;
	    RECT 344.4000 101.6000 345.4000 104.2000 ;
	    RECT 350.0000 101.6000 350.8000 106.2000 ;
	    RECT 354.8000 101.6000 355.6000 105.4000 ;
	    RECT 361.2000 101.6000 362.0000 106.6000 ;
	    RECT 366.4000 101.6000 367.2000 107.0000 ;
	    RECT 370.8000 101.6000 371.6000 106.6000 ;
	    RECT 376.0000 101.6000 376.8000 107.0000 ;
	    RECT 380.4000 101.6000 381.2000 106.0000 ;
	    RECT 386.0000 101.6000 386.8000 104.2000 ;
	    RECT 389.2000 101.6000 390.2000 104.2000 ;
	    RECT 394.8000 101.6000 395.6000 106.2000 ;
	    RECT 401.2000 101.6000 402.0000 105.4000 ;
	    RECT 412.4000 101.6000 413.2000 106.0000 ;
	    RECT 418.0000 101.6000 418.8000 104.2000 ;
	    RECT 421.2000 101.6000 422.2000 104.2000 ;
	    RECT 426.8000 101.6000 427.6000 106.2000 ;
	    RECT 430.0000 101.6000 430.8000 106.2000 ;
	    RECT 436.4000 101.6000 437.2000 106.0000 ;
	    RECT 442.0000 101.6000 442.8000 104.2000 ;
	    RECT 445.2000 101.6000 446.2000 104.2000 ;
	    RECT 450.8000 101.6000 451.6000 106.2000 ;
	    RECT 454.0000 101.6000 454.8000 106.2000 ;
	    RECT 462.0000 101.6000 462.8000 105.4000 ;
	    RECT 466.8000 101.6000 467.6000 106.2000 ;
	    RECT 470.0000 101.6000 470.8000 106.2000 ;
	    RECT 473.2000 101.6000 474.0000 106.0000 ;
	    RECT 478.8000 101.6000 479.6000 104.2000 ;
	    RECT 482.0000 101.6000 483.0000 104.2000 ;
	    RECT 487.6000 101.6000 488.4000 106.2000 ;
	    RECT 490.8000 101.6000 491.6000 104.2000 ;
	    RECT 495.6000 101.6000 496.4000 105.4000 ;
	    RECT 500.4000 101.6000 501.2000 108.2000 ;
	    RECT 506.8000 101.6000 507.6000 108.2000 ;
	    RECT 0.4000 100.4000 514.8000 101.6000 ;
	    RECT 2.8000 95.8000 3.6000 100.4000 ;
	    RECT 7.6000 95.8000 8.4000 100.4000 ;
	    RECT 14.0000 96.6000 14.8000 100.4000 ;
	    RECT 20.4000 96.6000 21.2000 100.4000 ;
	    RECT 25.2000 96.6000 26.0000 100.4000 ;
	    RECT 31.6000 96.0000 32.4000 100.4000 ;
	    RECT 37.2000 97.8000 38.0000 100.4000 ;
	    RECT 40.4000 97.8000 41.4000 100.4000 ;
	    RECT 46.0000 95.8000 46.8000 100.4000 ;
	    RECT 52.4000 96.6000 53.2000 100.4000 ;
	    RECT 55.6000 97.8000 56.4000 100.4000 ;
	    RECT 58.8000 97.8000 59.6000 100.4000 ;
	    RECT 60.4000 97.8000 61.2000 100.4000 ;
	    RECT 63.6000 97.8000 64.4000 100.4000 ;
	    RECT 65.2000 97.8000 66.0000 100.4000 ;
	    RECT 68.4000 97.8000 69.2000 100.4000 ;
	    RECT 70.0000 97.8000 70.8000 100.4000 ;
	    RECT 73.2000 97.8000 74.0000 100.4000 ;
	    RECT 78.0000 96.6000 78.8000 100.4000 ;
	    RECT 82.8000 95.8000 83.6000 100.4000 ;
	    RECT 88.2000 97.8000 89.2000 100.4000 ;
	    RECT 91.6000 97.8000 92.4000 100.4000 ;
	    RECT 97.2000 96.0000 98.0000 100.4000 ;
	    RECT 102.0000 96.6000 102.8000 100.4000 ;
	    RECT 116.4000 96.6000 117.2000 100.4000 ;
	    RECT 122.8000 96.6000 123.6000 100.4000 ;
	    RECT 129.2000 96.6000 130.0000 100.4000 ;
	    RECT 132.4000 97.8000 133.2000 100.4000 ;
	    RECT 135.6000 97.8000 136.4000 100.4000 ;
	    RECT 142.0000 96.6000 142.8000 100.4000 ;
	    RECT 148.4000 96.6000 149.2000 100.4000 ;
	    RECT 156.4000 96.6000 157.2000 100.4000 ;
	    RECT 162.8000 96.6000 163.6000 100.4000 ;
	    RECT 166.0000 97.8000 166.8000 100.4000 ;
	    RECT 169.2000 97.8000 170.0000 100.4000 ;
	    RECT 174.0000 96.6000 174.8000 100.4000 ;
	    RECT 178.8000 96.6000 179.6000 100.4000 ;
	    RECT 190.0000 96.6000 190.8000 100.4000 ;
	    RECT 196.4000 96.6000 197.2000 100.4000 ;
	    RECT 202.8000 96.6000 203.6000 100.4000 ;
	    RECT 207.6000 95.4000 208.4000 100.4000 ;
	    RECT 212.8000 95.0000 213.6000 100.4000 ;
	    RECT 216.8000 95.0000 217.6000 100.4000 ;
	    RECT 222.0000 95.4000 222.8000 100.4000 ;
	    RECT 225.2000 97.8000 226.0000 100.4000 ;
	    RECT 228.4000 97.8000 229.2000 100.4000 ;
	    RECT 230.0000 95.8000 230.8000 100.4000 ;
	    RECT 238.0000 96.6000 238.8000 100.4000 ;
	    RECT 242.8000 96.0000 243.6000 100.4000 ;
	    RECT 248.4000 97.8000 249.2000 100.4000 ;
	    RECT 251.6000 97.8000 252.6000 100.4000 ;
	    RECT 257.2000 95.8000 258.0000 100.4000 ;
	    RECT 270.0000 95.8000 270.8000 100.4000 ;
	    RECT 273.2000 95.8000 274.0000 100.4000 ;
	    RECT 278.0000 95.8000 278.8000 100.4000 ;
	    RECT 286.0000 96.6000 286.8000 100.4000 ;
	    RECT 290.8000 95.8000 291.6000 100.4000 ;
	    RECT 295.6000 96.6000 296.4000 100.4000 ;
	    RECT 305.2000 96.6000 306.0000 100.4000 ;
	    RECT 311.6000 96.6000 312.4000 100.4000 ;
	    RECT 314.8000 97.8000 315.6000 100.4000 ;
	    RECT 318.0000 97.8000 318.8000 100.4000 ;
	    RECT 321.2000 96.6000 322.0000 100.4000 ;
	    RECT 329.2000 95.8000 330.0000 100.4000 ;
	    RECT 334.0000 95.4000 334.8000 100.4000 ;
	    RECT 339.2000 95.0000 340.0000 100.4000 ;
	    RECT 343.2000 95.0000 344.0000 100.4000 ;
	    RECT 348.4000 95.4000 349.2000 100.4000 ;
	    RECT 351.6000 97.8000 352.4000 100.4000 ;
	    RECT 354.8000 97.8000 355.6000 100.4000 ;
	    RECT 358.0000 96.6000 358.8000 100.4000 ;
	    RECT 367.6000 96.6000 368.4000 100.4000 ;
	    RECT 372.4000 95.8000 373.2000 100.4000 ;
	    RECT 377.2000 96.6000 378.0000 100.4000 ;
	    RECT 385.2000 96.6000 386.0000 100.4000 ;
	    RECT 390.0000 96.0000 390.8000 100.4000 ;
	    RECT 395.6000 97.8000 396.4000 100.4000 ;
	    RECT 398.8000 97.8000 399.8000 100.4000 ;
	    RECT 404.4000 95.8000 405.2000 100.4000 ;
	    RECT 415.6000 96.0000 416.4000 100.4000 ;
	    RECT 421.2000 97.8000 422.0000 100.4000 ;
	    RECT 424.4000 97.8000 425.4000 100.4000 ;
	    RECT 430.0000 95.8000 430.8000 100.4000 ;
	    RECT 436.4000 96.6000 437.2000 100.4000 ;
	    RECT 441.2000 96.0000 442.0000 100.4000 ;
	    RECT 446.8000 97.8000 447.6000 100.4000 ;
	    RECT 450.0000 97.8000 451.0000 100.4000 ;
	    RECT 455.6000 95.8000 456.4000 100.4000 ;
	    RECT 458.8000 97.8000 459.6000 100.4000 ;
	    RECT 463.6000 96.6000 464.4000 100.4000 ;
	    RECT 470.0000 96.0000 470.8000 100.4000 ;
	    RECT 475.6000 97.8000 476.4000 100.4000 ;
	    RECT 478.8000 97.8000 479.8000 100.4000 ;
	    RECT 484.4000 95.8000 485.2000 100.4000 ;
	    RECT 490.8000 96.6000 491.6000 100.4000 ;
	    RECT 494.0000 97.8000 494.8000 100.4000 ;
	    RECT 497.2000 93.8000 498.0000 100.4000 ;
	    RECT 508.4000 93.8000 509.2000 100.4000 ;
	    RECT 2.8000 61.6000 3.6000 66.2000 ;
	    RECT 7.6000 61.6000 8.4000 66.2000 ;
	    RECT 12.4000 61.6000 13.2000 66.2000 ;
	    RECT 17.2000 61.6000 18.0000 66.0000 ;
	    RECT 22.8000 61.6000 23.6000 64.2000 ;
	    RECT 26.0000 61.6000 27.0000 64.2000 ;
	    RECT 31.6000 61.6000 32.4000 66.2000 ;
	    RECT 36.4000 61.6000 37.2000 66.2000 ;
	    RECT 42.8000 61.6000 43.6000 65.4000 ;
	    RECT 47.6000 61.6000 48.4000 66.2000 ;
	    RECT 54.0000 61.6000 54.8000 65.4000 ;
	    RECT 57.2000 61.6000 58.0000 66.2000 ;
	    RECT 60.4000 61.6000 61.2000 66.2000 ;
	    RECT 63.6000 61.6000 64.4000 66.2000 ;
	    RECT 66.8000 61.6000 67.6000 66.2000 ;
	    RECT 70.0000 61.6000 70.8000 66.2000 ;
	    RECT 74.8000 61.6000 75.6000 65.4000 ;
	    RECT 79.6000 61.6000 80.4000 66.2000 ;
	    RECT 84.4000 61.6000 85.2000 66.2000 ;
	    RECT 89.8000 61.6000 90.8000 64.2000 ;
	    RECT 93.2000 61.6000 94.0000 64.2000 ;
	    RECT 98.8000 61.6000 99.6000 66.0000 ;
	    RECT 103.6000 61.6000 104.4000 65.4000 ;
	    RECT 118.0000 61.6000 118.8000 66.2000 ;
	    RECT 121.2000 61.6000 122.0000 66.2000 ;
	    RECT 126.0000 61.6000 126.8000 66.6000 ;
	    RECT 131.2000 61.6000 132.0000 67.0000 ;
	    RECT 135.6000 61.6000 136.4000 66.6000 ;
	    RECT 140.8000 61.6000 141.6000 67.0000 ;
	    RECT 143.6000 61.6000 144.4000 66.2000 ;
	    RECT 151.6000 61.6000 152.4000 65.4000 ;
	    RECT 156.4000 61.6000 157.2000 66.2000 ;
	    RECT 162.8000 61.6000 163.6000 65.4000 ;
	    RECT 169.2000 61.6000 170.0000 65.4000 ;
	    RECT 174.0000 61.6000 174.8000 65.4000 ;
	    RECT 182.0000 61.6000 182.8000 65.4000 ;
	    RECT 186.8000 61.6000 187.6000 66.0000 ;
	    RECT 192.4000 61.6000 193.2000 64.2000 ;
	    RECT 195.6000 61.6000 196.6000 64.2000 ;
	    RECT 201.2000 61.6000 202.0000 66.2000 ;
	    RECT 207.6000 61.6000 208.4000 65.4000 ;
	    RECT 212.4000 61.6000 213.2000 66.2000 ;
	    RECT 220.4000 61.6000 221.2000 65.4000 ;
	    RECT 226.8000 61.6000 227.6000 65.4000 ;
	    RECT 230.0000 61.6000 230.8000 64.2000 ;
	    RECT 233.2000 61.6000 234.0000 64.2000 ;
	    RECT 239.6000 61.6000 240.4000 65.4000 ;
	    RECT 244.4000 61.6000 245.2000 65.4000 ;
	    RECT 252.4000 61.6000 253.2000 65.4000 ;
	    RECT 262.0000 61.6000 262.8000 64.2000 ;
	    RECT 265.2000 61.6000 266.0000 64.2000 ;
	    RECT 270.0000 61.6000 270.8000 65.4000 ;
	    RECT 278.0000 61.6000 278.8000 65.4000 ;
	    RECT 281.2000 61.6000 282.0000 64.2000 ;
	    RECT 284.4000 61.6000 285.2000 64.2000 ;
	    RECT 287.6000 61.6000 288.4000 66.2000 ;
	    RECT 293.0000 61.6000 294.0000 64.2000 ;
	    RECT 296.4000 61.6000 297.2000 64.2000 ;
	    RECT 302.0000 61.6000 302.8000 66.0000 ;
	    RECT 306.4000 61.6000 307.2000 67.0000 ;
	    RECT 311.6000 61.6000 312.4000 66.6000 ;
	    RECT 316.0000 61.6000 316.8000 67.0000 ;
	    RECT 321.2000 61.6000 322.0000 66.6000 ;
	    RECT 326.0000 61.6000 326.8000 65.4000 ;
	    RECT 334.0000 61.6000 334.8000 66.2000 ;
	    RECT 337.2000 61.6000 338.0000 66.0000 ;
	    RECT 342.8000 61.6000 343.6000 64.2000 ;
	    RECT 346.0000 61.6000 347.0000 64.2000 ;
	    RECT 351.6000 61.6000 352.4000 66.2000 ;
	    RECT 356.4000 61.6000 357.2000 66.2000 ;
	    RECT 359.6000 61.6000 360.4000 66.2000 ;
	    RECT 366.0000 61.6000 366.8000 66.0000 ;
	    RECT 371.6000 61.6000 372.4000 64.2000 ;
	    RECT 374.8000 61.6000 375.8000 64.2000 ;
	    RECT 380.4000 61.6000 381.2000 66.2000 ;
	    RECT 386.8000 61.6000 387.6000 65.4000 ;
	    RECT 391.6000 61.6000 392.4000 66.2000 ;
	    RECT 396.4000 61.6000 397.2000 66.0000 ;
	    RECT 402.0000 61.6000 402.8000 64.2000 ;
	    RECT 405.2000 61.6000 406.2000 64.2000 ;
	    RECT 410.8000 61.6000 411.6000 66.2000 ;
	    RECT 420.4000 61.6000 421.2000 66.2000 ;
	    RECT 428.4000 61.6000 429.2000 65.4000 ;
	    RECT 431.6000 61.6000 432.4000 66.2000 ;
	    RECT 434.8000 61.6000 435.6000 66.2000 ;
	    RECT 438.0000 61.6000 438.8000 66.2000 ;
	    RECT 441.2000 61.6000 442.0000 66.2000 ;
	    RECT 444.4000 61.6000 445.2000 66.2000 ;
	    RECT 446.0000 61.6000 446.8000 64.2000 ;
	    RECT 450.8000 61.6000 451.6000 65.4000 ;
	    RECT 457.2000 61.6000 458.0000 66.0000 ;
	    RECT 462.8000 61.6000 463.6000 64.2000 ;
	    RECT 466.0000 61.6000 467.0000 64.2000 ;
	    RECT 471.6000 61.6000 472.4000 66.2000 ;
	    RECT 474.8000 61.6000 475.6000 64.2000 ;
	    RECT 479.6000 61.6000 480.4000 65.4000 ;
	    RECT 489.2000 61.6000 490.0000 68.2000 ;
	    RECT 490.8000 61.6000 491.6000 64.2000 ;
	    RECT 495.6000 61.6000 496.4000 65.4000 ;
	    RECT 500.4000 61.6000 501.2000 66.2000 ;
	    RECT 503.6000 61.6000 504.4000 66.2000 ;
	    RECT 506.8000 61.6000 507.6000 66.2000 ;
	    RECT 510.0000 61.6000 510.8000 66.2000 ;
	    RECT 513.2000 61.6000 514.0000 66.2000 ;
	    RECT 0.4000 60.4000 514.8000 61.6000 ;
	    RECT 2.8000 55.8000 3.6000 60.4000 ;
	    RECT 6.0000 55.8000 6.8000 60.4000 ;
	    RECT 9.2000 55.8000 10.0000 60.4000 ;
	    RECT 12.4000 55.8000 13.2000 60.4000 ;
	    RECT 15.6000 55.8000 16.4000 60.4000 ;
	    RECT 18.8000 55.8000 19.6000 60.4000 ;
	    RECT 22.0000 56.0000 22.8000 60.4000 ;
	    RECT 27.6000 57.8000 28.4000 60.4000 ;
	    RECT 30.8000 57.8000 31.8000 60.4000 ;
	    RECT 36.4000 55.8000 37.2000 60.4000 ;
	    RECT 42.8000 56.6000 43.6000 60.4000 ;
	    RECT 49.2000 56.6000 50.0000 60.4000 ;
	    RECT 55.6000 56.6000 56.4000 60.4000 ;
	    RECT 62.0000 56.6000 62.8000 60.4000 ;
	    RECT 66.8000 56.0000 67.6000 60.4000 ;
	    RECT 72.4000 57.8000 73.2000 60.4000 ;
	    RECT 75.6000 57.8000 76.6000 60.4000 ;
	    RECT 81.2000 55.8000 82.0000 60.4000 ;
	    RECT 86.0000 55.8000 86.8000 60.4000 ;
	    RECT 92.4000 56.6000 93.2000 60.4000 ;
	    RECT 98.8000 56.6000 99.6000 60.4000 ;
	    RECT 103.6000 55.8000 104.4000 60.4000 ;
	    RECT 116.4000 56.6000 117.2000 60.4000 ;
	    RECT 121.2000 55.8000 122.0000 60.4000 ;
	    RECT 126.0000 55.8000 126.8000 60.4000 ;
	    RECT 132.4000 56.6000 133.2000 60.4000 ;
	    RECT 137.2000 56.0000 138.0000 60.4000 ;
	    RECT 142.8000 57.8000 143.6000 60.4000 ;
	    RECT 146.0000 57.8000 147.0000 60.4000 ;
	    RECT 151.6000 55.8000 152.4000 60.4000 ;
	    RECT 158.0000 56.6000 158.8000 60.4000 ;
	    RECT 164.4000 56.6000 165.2000 60.4000 ;
	    RECT 170.8000 56.6000 171.6000 60.4000 ;
	    RECT 177.2000 56.6000 178.0000 60.4000 ;
	    RECT 183.6000 56.6000 184.4000 60.4000 ;
	    RECT 188.4000 56.6000 189.2000 60.4000 ;
	    RECT 196.4000 56.6000 197.2000 60.4000 ;
	    RECT 202.8000 56.6000 203.6000 60.4000 ;
	    RECT 209.2000 56.6000 210.0000 60.4000 ;
	    RECT 215.6000 56.6000 216.4000 60.4000 ;
	    RECT 222.0000 56.6000 222.8000 60.4000 ;
	    RECT 230.0000 56.6000 230.8000 60.4000 ;
	    RECT 236.4000 56.6000 237.2000 60.4000 ;
	    RECT 239.6000 57.8000 240.4000 60.4000 ;
	    RECT 242.8000 57.8000 243.6000 60.4000 ;
	    RECT 246.0000 55.8000 246.8000 60.4000 ;
	    RECT 252.4000 55.8000 253.2000 60.4000 ;
	    RECT 260.4000 55.8000 261.2000 60.4000 ;
	    RECT 270.0000 56.6000 270.8000 60.4000 ;
	    RECT 276.4000 56.6000 277.2000 60.4000 ;
	    RECT 282.8000 56.6000 283.6000 60.4000 ;
	    RECT 286.0000 57.8000 286.8000 60.4000 ;
	    RECT 289.2000 57.8000 290.0000 60.4000 ;
	    RECT 295.6000 56.6000 296.4000 60.4000 ;
	    RECT 302.0000 56.6000 302.8000 60.4000 ;
	    RECT 305.2000 57.8000 306.0000 60.4000 ;
	    RECT 308.4000 57.8000 309.2000 60.4000 ;
	    RECT 311.6000 56.6000 312.4000 60.4000 ;
	    RECT 318.0000 56.6000 318.8000 60.4000 ;
	    RECT 324.4000 57.8000 325.2000 60.4000 ;
	    RECT 327.6000 57.8000 328.4000 60.4000 ;
	    RECT 329.2000 57.8000 330.0000 60.4000 ;
	    RECT 332.4000 57.8000 333.2000 60.4000 ;
	    RECT 335.6000 55.4000 336.4000 60.4000 ;
	    RECT 340.8000 55.0000 341.6000 60.4000 ;
	    RECT 344.8000 55.0000 345.6000 60.4000 ;
	    RECT 350.0000 55.4000 350.8000 60.4000 ;
	    RECT 356.4000 56.6000 357.2000 60.4000 ;
	    RECT 361.2000 56.6000 362.0000 60.4000 ;
	    RECT 367.6000 56.0000 368.4000 60.4000 ;
	    RECT 373.2000 57.8000 374.0000 60.4000 ;
	    RECT 376.4000 57.8000 377.4000 60.4000 ;
	    RECT 382.0000 55.8000 382.8000 60.4000 ;
	    RECT 388.4000 56.6000 389.2000 60.4000 ;
	    RECT 391.6000 55.8000 392.4000 60.4000 ;
	    RECT 398.0000 56.6000 398.8000 60.4000 ;
	    RECT 410.8000 56.0000 411.6000 60.4000 ;
	    RECT 416.4000 57.8000 417.2000 60.4000 ;
	    RECT 419.6000 57.8000 420.6000 60.4000 ;
	    RECT 425.2000 55.8000 426.0000 60.4000 ;
	    RECT 428.4000 55.8000 429.2000 60.4000 ;
	    RECT 436.4000 56.6000 437.2000 60.4000 ;
	    RECT 441.2000 55.8000 442.0000 60.4000 ;
	    RECT 446.0000 56.0000 446.8000 60.4000 ;
	    RECT 451.6000 57.8000 452.4000 60.4000 ;
	    RECT 454.8000 57.8000 455.8000 60.4000 ;
	    RECT 460.4000 55.8000 461.2000 60.4000 ;
	    RECT 465.2000 55.8000 466.0000 60.4000 ;
	    RECT 471.6000 53.8000 472.4000 60.4000 ;
	    RECT 474.8000 55.8000 475.6000 60.4000 ;
	    RECT 476.4000 53.8000 477.2000 60.4000 ;
	    RECT 484.4000 55.8000 485.2000 60.4000 ;
	    RECT 490.8000 53.8000 491.6000 60.4000 ;
	    RECT 494.0000 56.0000 494.8000 60.4000 ;
	    RECT 499.6000 57.8000 500.4000 60.4000 ;
	    RECT 502.8000 57.8000 503.8000 60.4000 ;
	    RECT 508.4000 55.8000 509.2000 60.4000 ;
	    RECT 2.8000 21.6000 3.6000 26.0000 ;
	    RECT 8.4000 21.6000 9.2000 24.2000 ;
	    RECT 11.6000 21.6000 12.6000 24.2000 ;
	    RECT 17.2000 21.6000 18.0000 26.2000 ;
	    RECT 22.0000 21.6000 22.8000 26.2000 ;
	    RECT 27.4000 21.6000 28.4000 24.2000 ;
	    RECT 30.8000 21.6000 31.6000 24.2000 ;
	    RECT 36.4000 21.6000 37.2000 26.0000 ;
	    RECT 42.8000 21.6000 43.6000 25.4000 ;
	    RECT 49.2000 21.6000 50.0000 25.4000 ;
	    RECT 54.0000 21.6000 54.8000 25.4000 ;
	    RECT 62.0000 21.6000 62.8000 25.4000 ;
	    RECT 66.8000 21.6000 67.6000 26.2000 ;
	    RECT 71.6000 21.6000 72.4000 26.0000 ;
	    RECT 77.2000 21.6000 78.0000 24.2000 ;
	    RECT 80.4000 21.6000 81.4000 24.2000 ;
	    RECT 86.0000 21.6000 86.8000 26.2000 ;
	    RECT 92.4000 21.6000 93.2000 25.4000 ;
	    RECT 98.8000 21.6000 99.6000 25.4000 ;
	    RECT 103.6000 21.6000 104.4000 26.2000 ;
	    RECT 114.8000 21.6000 115.6000 26.0000 ;
	    RECT 120.4000 21.6000 121.2000 24.2000 ;
	    RECT 123.6000 21.6000 124.6000 24.2000 ;
	    RECT 129.2000 21.6000 130.0000 26.2000 ;
	    RECT 134.0000 21.6000 134.8000 25.4000 ;
	    RECT 140.4000 21.6000 141.2000 26.0000 ;
	    RECT 146.0000 21.6000 146.8000 24.2000 ;
	    RECT 149.2000 21.6000 150.2000 24.2000 ;
	    RECT 154.8000 21.6000 155.6000 26.2000 ;
	    RECT 161.2000 21.6000 162.0000 25.4000 ;
	    RECT 166.0000 21.6000 166.8000 25.4000 ;
	    RECT 172.4000 21.6000 173.2000 26.2000 ;
	    RECT 177.8000 21.6000 178.8000 24.2000 ;
	    RECT 181.2000 21.6000 182.0000 24.2000 ;
	    RECT 186.8000 21.6000 187.6000 26.0000 ;
	    RECT 191.2000 21.6000 192.0000 27.0000 ;
	    RECT 196.4000 21.6000 197.2000 26.6000 ;
	    RECT 200.8000 21.6000 201.6000 27.0000 ;
	    RECT 206.0000 21.6000 206.8000 26.6000 ;
	    RECT 210.8000 21.6000 211.6000 26.2000 ;
	    RECT 218.8000 21.6000 219.6000 25.4000 ;
	    RECT 225.2000 21.6000 226.0000 25.4000 ;
	    RECT 229.6000 21.6000 230.4000 27.0000 ;
	    RECT 234.8000 21.6000 235.6000 26.6000 ;
	    RECT 238.0000 21.6000 238.8000 24.2000 ;
	    RECT 241.2000 21.6000 242.0000 24.2000 ;
	    RECT 244.0000 21.6000 244.8000 27.0000 ;
	    RECT 249.2000 21.6000 250.0000 26.6000 ;
	    RECT 263.6000 21.6000 264.4000 25.4000 ;
	    RECT 266.8000 21.6000 267.6000 24.2000 ;
	    RECT 270.0000 21.6000 270.8000 24.2000 ;
	    RECT 274.8000 21.6000 275.6000 25.4000 ;
	    RECT 279.6000 21.6000 280.4000 26.0000 ;
	    RECT 285.2000 21.6000 286.0000 24.2000 ;
	    RECT 288.4000 21.6000 289.4000 24.2000 ;
	    RECT 294.0000 21.6000 294.8000 26.2000 ;
	    RECT 298.8000 21.6000 299.6000 25.4000 ;
	    RECT 306.8000 21.6000 307.6000 25.4000 ;
	    RECT 311.2000 21.6000 312.0000 27.0000 ;
	    RECT 316.4000 21.6000 317.2000 26.6000 ;
	    RECT 321.2000 21.6000 322.0000 25.4000 ;
	    RECT 327.6000 21.6000 328.4000 25.4000 ;
	    RECT 335.6000 21.6000 336.4000 26.6000 ;
	    RECT 340.8000 21.6000 341.6000 27.0000 ;
	    RECT 345.2000 21.6000 346.0000 26.0000 ;
	    RECT 350.8000 21.6000 351.6000 24.2000 ;
	    RECT 354.0000 21.6000 355.0000 24.2000 ;
	    RECT 359.6000 21.6000 360.4000 26.2000 ;
	    RECT 366.0000 21.6000 366.8000 25.4000 ;
	    RECT 370.8000 21.6000 371.6000 25.4000 ;
	    RECT 378.8000 21.6000 379.6000 25.4000 ;
	    RECT 383.6000 21.6000 384.4000 26.0000 ;
	    RECT 389.2000 21.6000 390.0000 24.2000 ;
	    RECT 392.4000 21.6000 393.4000 24.2000 ;
	    RECT 398.0000 21.6000 398.8000 26.2000 ;
	    RECT 401.2000 21.6000 402.0000 26.2000 ;
	    RECT 415.6000 21.6000 416.4000 25.4000 ;
	    RECT 420.4000 21.6000 421.2000 26.0000 ;
	    RECT 426.0000 21.6000 426.8000 24.2000 ;
	    RECT 429.2000 21.6000 430.2000 24.2000 ;
	    RECT 434.8000 21.6000 435.6000 26.2000 ;
	    RECT 439.6000 21.6000 440.4000 26.0000 ;
	    RECT 445.2000 21.6000 446.0000 24.2000 ;
	    RECT 448.4000 21.6000 449.4000 24.2000 ;
	    RECT 454.0000 21.6000 454.8000 26.2000 ;
	    RECT 460.4000 21.6000 461.2000 26.2000 ;
	    RECT 462.0000 21.6000 462.8000 24.2000 ;
	    RECT 466.8000 21.6000 467.6000 25.4000 ;
	    RECT 471.6000 21.6000 472.4000 24.2000 ;
	    RECT 476.4000 21.6000 477.2000 25.4000 ;
	    RECT 481.2000 21.6000 482.0000 24.2000 ;
	    RECT 486.0000 21.6000 486.8000 25.4000 ;
	    RECT 492.4000 21.6000 493.2000 26.0000 ;
	    RECT 498.0000 21.6000 498.8000 24.2000 ;
	    RECT 501.2000 21.6000 502.2000 24.2000 ;
	    RECT 506.8000 21.6000 507.6000 26.2000 ;
	    RECT 0.4000 20.4000 514.8000 21.6000 ;
	    RECT 2.8000 15.8000 3.6000 20.4000 ;
	    RECT 7.6000 15.8000 8.4000 20.4000 ;
	    RECT 12.4000 16.0000 13.2000 20.4000 ;
	    RECT 18.0000 17.8000 18.8000 20.4000 ;
	    RECT 21.2000 17.8000 22.2000 20.4000 ;
	    RECT 26.8000 15.8000 27.6000 20.4000 ;
	    RECT 33.2000 16.6000 34.0000 20.4000 ;
	    RECT 38.0000 15.8000 38.8000 20.4000 ;
	    RECT 44.4000 16.6000 45.2000 20.4000 ;
	    RECT 49.2000 15.8000 50.0000 20.4000 ;
	    RECT 54.0000 16.0000 54.8000 20.4000 ;
	    RECT 59.6000 17.8000 60.4000 20.4000 ;
	    RECT 62.8000 17.8000 63.8000 20.4000 ;
	    RECT 68.4000 15.8000 69.2000 20.4000 ;
	    RECT 73.2000 16.6000 74.0000 20.4000 ;
	    RECT 79.6000 15.8000 80.4000 20.4000 ;
	    RECT 84.4000 15.8000 85.2000 20.4000 ;
	    RECT 89.8000 17.8000 90.8000 20.4000 ;
	    RECT 93.2000 17.8000 94.0000 20.4000 ;
	    RECT 98.8000 16.0000 99.6000 20.4000 ;
	    RECT 103.6000 15.8000 104.4000 20.4000 ;
	    RECT 116.4000 16.6000 117.2000 20.4000 ;
	    RECT 122.8000 16.6000 123.6000 20.4000 ;
	    RECT 129.2000 16.6000 130.0000 20.4000 ;
	    RECT 134.0000 15.8000 134.8000 20.4000 ;
	    RECT 138.8000 15.8000 139.6000 20.4000 ;
	    RECT 143.6000 16.0000 144.4000 20.4000 ;
	    RECT 149.2000 17.8000 150.0000 20.4000 ;
	    RECT 152.4000 17.8000 153.4000 20.4000 ;
	    RECT 158.0000 15.8000 158.8000 20.4000 ;
	    RECT 162.8000 15.8000 163.6000 20.4000 ;
	    RECT 167.6000 16.0000 168.4000 20.4000 ;
	    RECT 173.2000 17.8000 174.0000 20.4000 ;
	    RECT 176.4000 17.8000 177.4000 20.4000 ;
	    RECT 182.0000 15.8000 182.8000 20.4000 ;
	    RECT 186.8000 15.8000 187.6000 20.4000 ;
	    RECT 191.6000 16.0000 192.4000 20.4000 ;
	    RECT 197.2000 17.8000 198.0000 20.4000 ;
	    RECT 200.4000 17.8000 201.4000 20.4000 ;
	    RECT 206.0000 15.8000 206.8000 20.4000 ;
	    RECT 209.2000 15.8000 210.0000 20.4000 ;
	    RECT 217.2000 16.6000 218.0000 20.4000 ;
	    RECT 225.2000 16.6000 226.0000 20.4000 ;
	    RECT 231.6000 16.6000 232.4000 20.4000 ;
	    RECT 234.8000 17.8000 235.6000 20.4000 ;
	    RECT 238.0000 17.8000 238.8000 20.4000 ;
	    RECT 241.2000 15.8000 242.0000 20.4000 ;
	    RECT 246.6000 17.8000 247.6000 20.4000 ;
	    RECT 250.0000 17.8000 250.8000 20.4000 ;
	    RECT 255.6000 16.0000 256.4000 20.4000 ;
	    RECT 266.8000 15.8000 267.6000 20.4000 ;
	    RECT 271.6000 16.0000 272.4000 20.4000 ;
	    RECT 277.2000 17.8000 278.0000 20.4000 ;
	    RECT 280.4000 17.8000 281.4000 20.4000 ;
	    RECT 286.0000 15.8000 286.8000 20.4000 ;
	    RECT 289.2000 15.8000 290.0000 20.4000 ;
	    RECT 297.2000 16.6000 298.0000 20.4000 ;
	    RECT 302.0000 16.0000 302.8000 20.4000 ;
	    RECT 307.6000 17.8000 308.4000 20.4000 ;
	    RECT 310.8000 17.8000 311.8000 20.4000 ;
	    RECT 316.4000 15.8000 317.2000 20.4000 ;
	    RECT 319.6000 15.8000 320.4000 20.4000 ;
	    RECT 327.6000 16.6000 328.4000 20.4000 ;
	    RECT 332.4000 16.6000 333.2000 20.4000 ;
	    RECT 342.0000 16.6000 342.8000 20.4000 ;
	    RECT 345.2000 17.8000 346.0000 20.4000 ;
	    RECT 348.4000 17.8000 349.2000 20.4000 ;
	    RECT 351.2000 15.0000 352.0000 20.4000 ;
	    RECT 356.4000 15.4000 357.2000 20.4000 ;
	    RECT 361.2000 15.4000 362.0000 20.4000 ;
	    RECT 366.4000 15.0000 367.2000 20.4000 ;
	    RECT 370.8000 16.0000 371.6000 20.4000 ;
	    RECT 376.4000 17.8000 377.2000 20.4000 ;
	    RECT 379.6000 17.8000 380.6000 20.4000 ;
	    RECT 385.2000 15.8000 386.0000 20.4000 ;
	    RECT 390.0000 16.0000 390.8000 20.4000 ;
	    RECT 395.6000 17.8000 396.4000 20.4000 ;
	    RECT 398.8000 17.8000 399.8000 20.4000 ;
	    RECT 404.4000 15.8000 405.2000 20.4000 ;
	    RECT 414.0000 15.8000 414.8000 20.4000 ;
	    RECT 422.0000 16.6000 422.8000 20.4000 ;
	    RECT 426.8000 16.0000 427.6000 20.4000 ;
	    RECT 432.4000 17.8000 433.2000 20.4000 ;
	    RECT 435.6000 17.8000 436.6000 20.4000 ;
	    RECT 441.2000 15.8000 442.0000 20.4000 ;
	    RECT 446.0000 16.6000 446.8000 20.4000 ;
	    RECT 454.0000 15.8000 454.8000 20.4000 ;
	    RECT 457.2000 16.6000 458.0000 20.4000 ;
	    RECT 463.6000 16.0000 464.4000 20.4000 ;
	    RECT 469.2000 17.8000 470.0000 20.4000 ;
	    RECT 472.4000 17.8000 473.4000 20.4000 ;
	    RECT 478.0000 15.8000 478.8000 20.4000 ;
	    RECT 482.8000 16.0000 483.6000 20.4000 ;
	    RECT 488.4000 17.8000 489.2000 20.4000 ;
	    RECT 491.6000 17.8000 492.6000 20.4000 ;
	    RECT 497.2000 15.8000 498.0000 20.4000 ;
	    RECT 500.4000 15.8000 501.2000 20.4000 ;
	    RECT 503.6000 15.8000 504.4000 20.4000 ;
	    RECT 506.8000 15.8000 507.6000 20.4000 ;
	    RECT 510.0000 15.8000 510.8000 20.4000 ;
	    RECT 513.2000 15.8000 514.0000 20.4000 ;
         LAYER metal2 ;
	    RECT 257.0000 341.4000 258.2000 341.6000 ;
	    RECT 254.7000 340.6000 260.5000 341.4000 ;
	    RECT 257.0000 340.4000 258.2000 340.6000 ;
	    RECT 257.0000 301.4000 258.2000 301.6000 ;
	    RECT 254.7000 300.6000 260.5000 301.4000 ;
	    RECT 257.0000 300.4000 258.2000 300.6000 ;
	    RECT 257.0000 261.4000 258.2000 261.6000 ;
	    RECT 254.7000 260.6000 260.5000 261.4000 ;
	    RECT 257.0000 260.4000 258.2000 260.6000 ;
	    RECT 257.0000 221.4000 258.2000 221.6000 ;
	    RECT 254.7000 220.6000 260.5000 221.4000 ;
	    RECT 257.0000 220.4000 258.2000 220.6000 ;
	    RECT 257.0000 181.4000 258.2000 181.6000 ;
	    RECT 254.7000 180.6000 260.5000 181.4000 ;
	    RECT 257.0000 180.4000 258.2000 180.6000 ;
	    RECT 257.0000 141.4000 258.2000 141.6000 ;
	    RECT 254.7000 140.6000 260.5000 141.4000 ;
	    RECT 257.0000 140.4000 258.2000 140.6000 ;
	    RECT 257.0000 101.4000 258.2000 101.6000 ;
	    RECT 254.7000 100.6000 260.5000 101.4000 ;
	    RECT 257.0000 100.4000 258.2000 100.6000 ;
	    RECT 257.0000 61.4000 258.2000 61.6000 ;
	    RECT 254.7000 60.6000 260.5000 61.4000 ;
	    RECT 257.0000 60.4000 258.2000 60.6000 ;
	    RECT 257.0000 21.4000 258.2000 21.6000 ;
	    RECT 254.7000 20.6000 260.5000 21.4000 ;
	    RECT 257.0000 20.4000 258.2000 20.6000 ;
         LAYER metal3 ;
	    RECT 254.6000 340.4000 260.6000 341.6000 ;
	    RECT 254.6000 300.4000 260.6000 301.6000 ;
	    RECT 254.6000 260.4000 260.6000 261.6000 ;
	    RECT 254.6000 220.4000 260.6000 221.6000 ;
	    RECT 254.6000 180.4000 260.6000 181.6000 ;
	    RECT 254.6000 140.4000 260.6000 141.6000 ;
	    RECT 254.6000 100.4000 260.6000 101.6000 ;
	    RECT 254.6000 60.4000 260.6000 61.6000 ;
	    RECT 254.6000 20.4000 260.6000 21.6000 ;
         LAYER metal4 ;
	    RECT 254.4000 -1.0000 260.8000 341.6000 ;
      END
   END gnd
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 2.8000 321.6000 3.6000 330.2000 ;
	    RECT 8.4000 321.6000 9.2000 326.2000 ;
	    RECT 11.6000 321.6000 12.4000 326.2000 ;
	    RECT 17.2000 321.6000 18.0000 330.0000 ;
	    RECT 22.0000 321.6000 22.8000 329.0000 ;
	    RECT 26.8000 321.6000 27.6000 329.0000 ;
	    RECT 30.6000 321.6000 31.4000 326.2000 ;
	    RECT 34.8000 321.6000 35.6000 330.2000 ;
	    RECT 37.0000 321.6000 37.8000 326.2000 ;
	    RECT 41.2000 321.6000 42.0000 330.2000 ;
	    RECT 44.4000 321.6000 45.2000 329.0000 ;
	    RECT 47.6000 321.6000 48.4000 330.2000 ;
	    RECT 51.8000 321.6000 52.6000 326.2000 ;
	    RECT 55.6000 321.6000 56.4000 330.2000 ;
	    RECT 61.2000 321.6000 62.0000 326.2000 ;
	    RECT 64.4000 321.6000 65.2000 326.2000 ;
	    RECT 70.0000 321.6000 70.8000 330.0000 ;
	    RECT 73.8000 321.6000 74.6000 326.2000 ;
	    RECT 78.0000 321.6000 78.8000 330.2000 ;
	    RECT 79.6000 321.6000 80.4000 330.2000 ;
	    RECT 82.8000 321.6000 83.6000 330.2000 ;
	    RECT 86.0000 321.6000 86.8000 330.2000 ;
	    RECT 89.2000 321.6000 90.0000 330.2000 ;
	    RECT 92.4000 321.6000 93.2000 330.2000 ;
	    RECT 95.6000 321.6000 96.4000 330.2000 ;
	    RECT 101.2000 321.6000 102.0000 326.2000 ;
	    RECT 104.4000 321.6000 105.2000 326.2000 ;
	    RECT 110.0000 321.6000 110.8000 330.0000 ;
	    RECT 119.6000 321.6000 120.4000 326.2000 ;
	    RECT 122.8000 321.6000 123.6000 326.2000 ;
	    RECT 125.0000 321.6000 125.8000 326.2000 ;
	    RECT 129.2000 321.6000 130.0000 330.2000 ;
	    RECT 132.4000 321.6000 133.2000 330.2000 ;
	    RECT 138.0000 321.6000 138.8000 326.2000 ;
	    RECT 141.2000 321.6000 142.0000 326.2000 ;
	    RECT 146.8000 321.6000 147.6000 330.0000 ;
	    RECT 150.0000 321.6000 150.8000 326.2000 ;
	    RECT 153.2000 321.6000 154.0000 326.2000 ;
	    RECT 155.4000 321.6000 156.2000 326.2000 ;
	    RECT 159.6000 321.6000 160.4000 330.2000 ;
	    RECT 162.8000 321.6000 163.6000 330.2000 ;
	    RECT 168.4000 321.6000 169.2000 326.2000 ;
	    RECT 171.6000 321.6000 172.4000 326.2000 ;
	    RECT 177.2000 321.6000 178.0000 330.0000 ;
	    RECT 181.0000 321.6000 181.8000 326.2000 ;
	    RECT 185.2000 321.6000 186.0000 330.2000 ;
	    RECT 187.4000 321.6000 188.2000 326.2000 ;
	    RECT 191.6000 321.6000 192.4000 330.2000 ;
	    RECT 194.8000 321.6000 195.6000 330.2000 ;
	    RECT 198.0000 321.6000 198.8000 330.0000 ;
	    RECT 203.6000 321.6000 204.4000 326.2000 ;
	    RECT 206.8000 321.6000 207.6000 326.2000 ;
	    RECT 212.4000 321.6000 213.2000 330.2000 ;
	    RECT 215.6000 321.6000 216.4000 330.2000 ;
	    RECT 219.8000 321.6000 220.6000 326.2000 ;
	    RECT 222.6000 321.6000 223.4000 326.2000 ;
	    RECT 226.8000 321.6000 227.6000 330.2000 ;
	    RECT 228.4000 321.6000 229.2000 330.2000 ;
	    RECT 231.6000 321.6000 232.4000 330.2000 ;
	    RECT 234.8000 321.6000 235.6000 330.2000 ;
	    RECT 238.0000 321.6000 238.8000 330.2000 ;
	    RECT 241.2000 321.6000 242.0000 330.2000 ;
	    RECT 244.4000 321.6000 245.2000 330.2000 ;
	    RECT 250.0000 321.6000 250.8000 326.2000 ;
	    RECT 253.2000 321.6000 254.0000 326.2000 ;
	    RECT 258.8000 321.6000 259.6000 330.0000 ;
	    RECT 268.4000 321.6000 269.2000 326.2000 ;
	    RECT 271.6000 321.6000 272.4000 330.2000 ;
	    RECT 275.8000 321.6000 276.6000 326.2000 ;
	    RECT 279.2000 321.6000 280.0000 330.2000 ;
	    RECT 284.4000 321.6000 285.2000 329.8000 ;
	    RECT 288.8000 321.6000 289.6000 330.2000 ;
	    RECT 294.0000 321.6000 294.8000 329.8000 ;
	    RECT 298.8000 321.6000 299.6000 329.8000 ;
	    RECT 304.0000 321.6000 304.8000 330.2000 ;
	    RECT 308.4000 321.6000 309.2000 329.8000 ;
	    RECT 313.6000 321.6000 314.4000 330.2000 ;
	    RECT 318.0000 321.6000 318.8000 330.2000 ;
	    RECT 323.6000 321.6000 324.4000 326.2000 ;
	    RECT 326.8000 321.6000 327.6000 326.2000 ;
	    RECT 332.4000 321.6000 333.2000 330.0000 ;
	    RECT 335.6000 321.6000 336.4000 326.2000 ;
	    RECT 338.8000 321.6000 339.6000 326.2000 ;
	    RECT 341.0000 321.6000 341.8000 326.2000 ;
	    RECT 345.2000 321.6000 346.0000 330.2000 ;
	    RECT 348.4000 321.6000 349.2000 330.2000 ;
	    RECT 354.0000 321.6000 354.8000 326.2000 ;
	    RECT 357.2000 321.6000 358.0000 326.2000 ;
	    RECT 362.8000 321.6000 363.6000 330.0000 ;
	    RECT 367.6000 321.6000 368.4000 330.2000 ;
	    RECT 370.8000 321.6000 371.6000 330.2000 ;
	    RECT 376.4000 321.6000 377.2000 326.2000 ;
	    RECT 379.6000 321.6000 380.4000 326.2000 ;
	    RECT 385.2000 321.6000 386.0000 330.0000 ;
	    RECT 388.4000 321.6000 389.2000 326.2000 ;
	    RECT 391.6000 321.6000 392.4000 330.2000 ;
	    RECT 395.8000 321.6000 396.6000 326.2000 ;
	    RECT 398.0000 321.6000 398.8000 326.2000 ;
	    RECT 401.2000 321.6000 402.0000 325.8000 ;
	    RECT 410.8000 321.6000 411.6000 326.2000 ;
	    RECT 414.0000 321.6000 414.8000 325.8000 ;
	    RECT 417.2000 321.6000 418.0000 326.2000 ;
	    RECT 420.4000 321.6000 421.2000 325.8000 ;
	    RECT 423.6000 321.6000 424.4000 326.2000 ;
	    RECT 426.8000 321.6000 427.6000 325.8000 ;
	    RECT 430.0000 321.6000 430.8000 326.2000 ;
	    RECT 433.2000 321.6000 434.0000 330.2000 ;
	    RECT 437.4000 321.6000 438.2000 326.2000 ;
	    RECT 441.2000 321.6000 442.0000 330.2000 ;
	    RECT 446.8000 321.6000 447.6000 326.2000 ;
	    RECT 450.0000 321.6000 450.8000 326.2000 ;
	    RECT 455.6000 321.6000 456.4000 330.0000 ;
	    RECT 460.4000 321.6000 461.2000 325.8000 ;
	    RECT 463.6000 321.6000 464.4000 326.2000 ;
	    RECT 465.2000 321.6000 466.0000 326.2000 ;
	    RECT 468.4000 321.6000 469.2000 325.8000 ;
	    RECT 472.2000 321.6000 473.0000 326.2000 ;
	    RECT 476.4000 321.6000 477.2000 330.2000 ;
	    RECT 479.6000 321.6000 480.4000 326.2000 ;
	    RECT 482.8000 321.6000 483.6000 330.2000 ;
	    RECT 488.4000 321.6000 489.2000 326.2000 ;
	    RECT 491.6000 321.6000 492.4000 326.2000 ;
	    RECT 497.2000 321.6000 498.0000 330.0000 ;
	    RECT 500.4000 321.6000 501.2000 326.2000 ;
	    RECT 505.2000 321.6000 506.0000 329.0000 ;
	    RECT 508.4000 321.6000 509.2000 326.2000 ;
	    RECT 511.6000 321.6000 512.4000 329.8000 ;
	    RECT 0.4000 320.4000 514.8000 321.6000 ;
	    RECT 2.8000 313.0000 3.6000 320.4000 ;
	    RECT 7.6000 313.0000 8.4000 320.4000 ;
	    RECT 10.8000 311.8000 11.6000 320.4000 ;
	    RECT 14.0000 311.8000 14.8000 320.4000 ;
	    RECT 17.2000 311.8000 18.0000 320.4000 ;
	    RECT 20.4000 311.8000 21.2000 320.4000 ;
	    RECT 23.6000 311.8000 24.4000 320.4000 ;
	    RECT 26.8000 311.8000 27.6000 320.4000 ;
	    RECT 32.4000 315.8000 33.2000 320.4000 ;
	    RECT 35.6000 315.8000 36.4000 320.4000 ;
	    RECT 41.2000 312.0000 42.0000 320.4000 ;
	    RECT 45.0000 315.8000 45.8000 320.4000 ;
	    RECT 49.2000 311.8000 50.0000 320.4000 ;
	    RECT 51.4000 315.8000 52.2000 320.4000 ;
	    RECT 55.6000 311.8000 56.4000 320.4000 ;
	    RECT 57.2000 311.8000 58.0000 320.4000 ;
	    RECT 62.6000 315.8000 63.4000 320.4000 ;
	    RECT 66.8000 311.8000 67.6000 320.4000 ;
	    RECT 70.0000 313.0000 70.8000 320.4000 ;
	    RECT 73.2000 311.8000 74.0000 320.4000 ;
	    RECT 77.4000 315.8000 78.2000 320.4000 ;
	    RECT 79.6000 311.8000 80.4000 320.4000 ;
	    RECT 86.0000 312.0000 86.8000 320.4000 ;
	    RECT 91.6000 315.8000 92.4000 320.4000 ;
	    RECT 94.8000 315.8000 95.6000 320.4000 ;
	    RECT 100.4000 311.8000 101.2000 320.4000 ;
	    RECT 110.0000 315.8000 110.8000 320.4000 ;
	    RECT 113.2000 315.8000 114.0000 320.4000 ;
	    RECT 115.4000 315.8000 116.2000 320.4000 ;
	    RECT 119.6000 311.8000 120.4000 320.4000 ;
	    RECT 121.2000 311.8000 122.0000 320.4000 ;
	    RECT 127.6000 311.8000 128.4000 320.4000 ;
	    RECT 129.8000 315.8000 130.6000 320.4000 ;
	    RECT 134.0000 311.8000 134.8000 320.4000 ;
	    RECT 137.2000 312.2000 138.0000 320.4000 ;
	    RECT 142.4000 311.8000 143.2000 320.4000 ;
	    RECT 148.4000 311.8000 149.2000 320.4000 ;
	    RECT 151.6000 311.8000 152.4000 320.4000 ;
	    RECT 157.2000 315.8000 158.0000 320.4000 ;
	    RECT 160.4000 315.8000 161.2000 320.4000 ;
	    RECT 166.0000 312.0000 166.8000 320.4000 ;
	    RECT 170.8000 311.8000 171.6000 320.4000 ;
	    RECT 176.4000 315.8000 177.2000 320.4000 ;
	    RECT 179.6000 315.8000 180.4000 320.4000 ;
	    RECT 185.2000 312.0000 186.0000 320.4000 ;
	    RECT 188.4000 315.8000 189.2000 320.4000 ;
	    RECT 191.6000 315.8000 192.4000 320.4000 ;
	    RECT 194.8000 315.8000 195.6000 320.4000 ;
	    RECT 197.0000 315.8000 197.8000 320.4000 ;
	    RECT 201.2000 311.8000 202.0000 320.4000 ;
	    RECT 204.4000 312.0000 205.2000 320.4000 ;
	    RECT 210.0000 315.8000 210.8000 320.4000 ;
	    RECT 213.2000 315.8000 214.0000 320.4000 ;
	    RECT 218.8000 311.8000 219.6000 320.4000 ;
	    RECT 222.0000 311.8000 222.8000 320.4000 ;
	    RECT 226.2000 315.8000 227.0000 320.4000 ;
	    RECT 230.0000 313.0000 230.8000 320.4000 ;
	    RECT 233.2000 311.8000 234.0000 320.4000 ;
	    RECT 238.0000 311.8000 238.8000 320.4000 ;
	    RECT 244.4000 311.8000 245.2000 320.4000 ;
	    RECT 246.0000 311.8000 246.8000 320.4000 ;
	    RECT 252.4000 311.8000 253.2000 320.4000 ;
	    RECT 263.6000 311.8000 264.4000 320.4000 ;
	    RECT 265.8000 315.8000 266.6000 320.4000 ;
	    RECT 270.0000 311.8000 270.8000 320.4000 ;
	    RECT 272.8000 311.8000 273.6000 320.4000 ;
	    RECT 278.0000 312.2000 278.8000 320.4000 ;
	    RECT 282.8000 312.2000 283.6000 320.4000 ;
	    RECT 288.0000 311.8000 288.8000 320.4000 ;
	    RECT 290.8000 311.8000 291.6000 320.4000 ;
	    RECT 297.2000 311.8000 298.0000 320.4000 ;
	    RECT 302.0000 311.8000 302.8000 320.4000 ;
	    RECT 305.2000 311.8000 306.0000 320.4000 ;
	    RECT 310.8000 315.8000 311.6000 320.4000 ;
	    RECT 314.0000 315.8000 314.8000 320.4000 ;
	    RECT 319.6000 312.0000 320.4000 320.4000 ;
	    RECT 322.8000 315.8000 323.6000 320.4000 ;
	    RECT 326.0000 315.8000 326.8000 320.4000 ;
	    RECT 328.2000 315.8000 329.0000 320.4000 ;
	    RECT 332.4000 311.8000 333.2000 320.4000 ;
	    RECT 334.0000 315.8000 334.8000 320.4000 ;
	    RECT 337.2000 315.8000 338.0000 320.4000 ;
	    RECT 339.4000 315.8000 340.2000 320.4000 ;
	    RECT 343.6000 311.8000 344.4000 320.4000 ;
	    RECT 346.8000 311.8000 347.6000 320.4000 ;
	    RECT 352.4000 315.8000 353.2000 320.4000 ;
	    RECT 355.6000 315.8000 356.4000 320.4000 ;
	    RECT 361.2000 312.0000 362.0000 320.4000 ;
	    RECT 364.4000 315.8000 365.2000 320.4000 ;
	    RECT 367.6000 315.8000 368.4000 320.4000 ;
	    RECT 369.8000 315.8000 370.6000 320.4000 ;
	    RECT 374.0000 311.8000 374.8000 320.4000 ;
	    RECT 377.2000 311.8000 378.0000 320.4000 ;
	    RECT 382.8000 315.8000 383.6000 320.4000 ;
	    RECT 386.0000 315.8000 386.8000 320.4000 ;
	    RECT 391.6000 312.0000 392.4000 320.4000 ;
	    RECT 394.8000 315.8000 395.6000 320.4000 ;
	    RECT 398.0000 316.2000 398.8000 320.4000 ;
	    RECT 409.2000 311.8000 410.0000 320.4000 ;
	    RECT 414.8000 315.8000 415.6000 320.4000 ;
	    RECT 418.0000 315.8000 418.8000 320.4000 ;
	    RECT 423.6000 312.0000 424.4000 320.4000 ;
	    RECT 427.4000 315.8000 428.2000 320.4000 ;
	    RECT 431.6000 311.8000 432.4000 320.4000 ;
	    RECT 434.8000 315.8000 435.6000 320.4000 ;
	    RECT 438.0000 311.8000 438.8000 320.4000 ;
	    RECT 443.6000 315.8000 444.4000 320.4000 ;
	    RECT 446.8000 315.8000 447.6000 320.4000 ;
	    RECT 452.4000 312.0000 453.2000 320.4000 ;
	    RECT 457.2000 311.8000 458.0000 320.4000 ;
	    RECT 460.4000 311.8000 461.2000 320.4000 ;
	    RECT 466.0000 315.8000 466.8000 320.4000 ;
	    RECT 469.2000 315.8000 470.0000 320.4000 ;
	    RECT 474.8000 312.0000 475.6000 320.4000 ;
	    RECT 478.6000 315.8000 479.4000 320.4000 ;
	    RECT 482.8000 311.8000 483.6000 320.4000 ;
	    RECT 486.0000 315.8000 486.8000 320.4000 ;
	    RECT 487.6000 315.8000 488.4000 320.4000 ;
	    RECT 490.8000 311.8000 491.6000 320.4000 ;
	    RECT 494.0000 311.8000 494.8000 320.4000 ;
	    RECT 497.2000 311.8000 498.0000 320.4000 ;
	    RECT 500.4000 311.8000 501.2000 320.4000 ;
	    RECT 503.6000 311.8000 504.4000 320.4000 ;
	    RECT 506.8000 313.0000 507.6000 320.4000 ;
	    RECT 2.8000 281.6000 3.6000 290.2000 ;
	    RECT 8.4000 281.6000 9.2000 286.2000 ;
	    RECT 11.6000 281.6000 12.4000 286.2000 ;
	    RECT 17.2000 281.6000 18.0000 290.0000 ;
	    RECT 22.0000 281.6000 22.8000 290.2000 ;
	    RECT 27.6000 281.6000 28.4000 286.2000 ;
	    RECT 30.8000 281.6000 31.6000 286.2000 ;
	    RECT 36.4000 281.6000 37.2000 290.0000 ;
	    RECT 41.2000 281.6000 42.0000 290.2000 ;
	    RECT 46.8000 281.6000 47.6000 286.2000 ;
	    RECT 50.0000 281.6000 50.8000 286.2000 ;
	    RECT 55.6000 281.6000 56.4000 290.0000 ;
	    RECT 58.8000 281.6000 59.6000 290.2000 ;
	    RECT 62.0000 281.6000 62.8000 290.2000 ;
	    RECT 64.2000 281.6000 65.0000 286.2000 ;
	    RECT 68.4000 281.6000 69.2000 290.2000 ;
	    RECT 70.0000 281.6000 70.8000 290.2000 ;
	    RECT 74.8000 281.6000 75.6000 286.2000 ;
	    RECT 78.0000 281.6000 78.8000 286.2000 ;
	    RECT 80.2000 281.6000 81.0000 286.2000 ;
	    RECT 84.4000 281.6000 85.2000 290.2000 ;
	    RECT 86.0000 281.6000 86.8000 290.2000 ;
	    RECT 90.2000 281.6000 91.0000 286.2000 ;
	    RECT 92.4000 281.6000 93.2000 290.2000 ;
	    RECT 98.8000 281.6000 99.6000 290.2000 ;
	    RECT 102.0000 281.6000 102.8000 289.8000 ;
	    RECT 107.2000 281.6000 108.0000 290.2000 ;
	    RECT 117.6000 281.6000 118.4000 290.2000 ;
	    RECT 122.8000 281.6000 123.6000 289.8000 ;
	    RECT 129.2000 281.6000 130.0000 290.2000 ;
	    RECT 130.8000 281.6000 131.6000 290.2000 ;
	    RECT 137.2000 281.6000 138.0000 289.8000 ;
	    RECT 142.4000 281.6000 143.2000 290.2000 ;
	    RECT 145.2000 281.6000 146.0000 290.2000 ;
	    RECT 151.6000 281.6000 152.4000 290.2000 ;
	    RECT 153.2000 281.6000 154.0000 290.2000 ;
	    RECT 157.4000 281.6000 158.2000 286.2000 ;
	    RECT 159.6000 281.6000 160.4000 290.2000 ;
	    RECT 164.4000 281.6000 165.2000 290.2000 ;
	    RECT 168.6000 281.6000 169.4000 286.2000 ;
	    RECT 171.4000 281.6000 172.2000 286.2000 ;
	    RECT 175.6000 281.6000 176.4000 290.2000 ;
	    RECT 178.8000 281.6000 179.6000 289.0000 ;
	    RECT 183.6000 281.6000 184.4000 290.2000 ;
	    RECT 189.2000 281.6000 190.0000 286.2000 ;
	    RECT 192.4000 281.6000 193.2000 286.2000 ;
	    RECT 198.0000 281.6000 198.8000 290.0000 ;
	    RECT 201.2000 281.6000 202.0000 290.2000 ;
	    RECT 205.4000 281.6000 206.2000 286.2000 ;
	    RECT 207.6000 281.6000 208.4000 286.2000 ;
	    RECT 210.8000 281.6000 211.6000 286.2000 ;
	    RECT 212.4000 281.6000 213.2000 290.2000 ;
	    RECT 216.6000 281.6000 217.4000 286.2000 ;
	    RECT 219.4000 281.6000 220.2000 286.2000 ;
	    RECT 223.6000 281.6000 224.4000 290.2000 ;
	    RECT 226.8000 281.6000 227.6000 290.2000 ;
	    RECT 232.4000 281.6000 233.2000 286.2000 ;
	    RECT 235.6000 281.6000 236.4000 286.2000 ;
	    RECT 241.2000 281.6000 242.0000 290.0000 ;
	    RECT 246.0000 281.6000 246.8000 289.8000 ;
	    RECT 251.2000 281.6000 252.0000 290.2000 ;
	    RECT 261.0000 281.6000 261.8000 286.2000 ;
	    RECT 265.2000 281.6000 266.0000 290.2000 ;
	    RECT 266.8000 281.6000 267.6000 290.2000 ;
	    RECT 271.6000 281.6000 272.4000 290.2000 ;
	    RECT 278.0000 281.6000 278.8000 290.2000 ;
	    RECT 279.6000 281.6000 280.4000 290.2000 ;
	    RECT 283.8000 281.6000 284.6000 286.2000 ;
	    RECT 286.0000 281.6000 286.8000 290.2000 ;
	    RECT 292.4000 281.6000 293.2000 290.2000 ;
	    RECT 294.0000 281.6000 294.8000 290.2000 ;
	    RECT 299.4000 281.6000 300.2000 286.2000 ;
	    RECT 303.6000 281.6000 304.4000 290.2000 ;
	    RECT 308.4000 281.6000 309.2000 290.2000 ;
	    RECT 310.0000 281.6000 310.8000 290.2000 ;
	    RECT 316.4000 281.6000 317.2000 290.2000 ;
	    RECT 318.6000 281.6000 319.4000 286.2000 ;
	    RECT 322.8000 281.6000 323.6000 290.2000 ;
	    RECT 325.0000 281.6000 325.8000 286.2000 ;
	    RECT 329.2000 281.6000 330.0000 290.2000 ;
	    RECT 332.4000 281.6000 333.2000 289.8000 ;
	    RECT 337.6000 281.6000 338.4000 290.2000 ;
	    RECT 342.0000 281.6000 342.8000 289.8000 ;
	    RECT 347.2000 281.6000 348.0000 290.2000 ;
	    RECT 351.6000 281.6000 352.4000 290.2000 ;
	    RECT 357.2000 281.6000 358.0000 286.2000 ;
	    RECT 360.4000 281.6000 361.2000 286.2000 ;
	    RECT 366.0000 281.6000 366.8000 290.0000 ;
	    RECT 369.2000 281.6000 370.0000 286.2000 ;
	    RECT 372.4000 281.6000 373.2000 286.2000 ;
	    RECT 374.6000 281.6000 375.4000 286.2000 ;
	    RECT 378.8000 281.6000 379.6000 290.2000 ;
	    RECT 382.0000 281.6000 382.8000 290.2000 ;
	    RECT 385.2000 281.6000 386.0000 290.2000 ;
	    RECT 390.8000 281.6000 391.6000 286.2000 ;
	    RECT 394.0000 281.6000 394.8000 286.2000 ;
	    RECT 399.6000 281.6000 400.4000 290.0000 ;
	    RECT 403.4000 281.6000 404.2000 286.2000 ;
	    RECT 407.6000 281.6000 408.4000 290.2000 ;
	    RECT 415.6000 281.6000 416.4000 290.2000 ;
	    RECT 419.8000 281.6000 420.6000 286.2000 ;
	    RECT 423.6000 281.6000 424.4000 290.2000 ;
	    RECT 425.2000 281.6000 426.0000 290.2000 ;
	    RECT 429.4000 281.6000 430.2000 286.2000 ;
	    RECT 431.6000 281.6000 432.4000 286.2000 ;
	    RECT 434.8000 281.6000 435.6000 286.2000 ;
	    RECT 438.0000 281.6000 438.8000 290.2000 ;
	    RECT 443.6000 281.6000 444.4000 286.2000 ;
	    RECT 446.8000 281.6000 447.6000 286.2000 ;
	    RECT 452.4000 281.6000 453.2000 290.0000 ;
	    RECT 455.6000 281.6000 456.4000 286.2000 ;
	    RECT 458.8000 281.6000 459.6000 285.8000 ;
	    RECT 462.0000 281.6000 462.8000 286.2000 ;
	    RECT 465.2000 281.6000 466.0000 290.2000 ;
	    RECT 469.4000 281.6000 470.2000 286.2000 ;
	    RECT 473.2000 281.6000 474.0000 290.2000 ;
	    RECT 478.8000 281.6000 479.6000 286.2000 ;
	    RECT 482.0000 281.6000 482.8000 286.2000 ;
	    RECT 487.6000 281.6000 488.4000 290.0000 ;
	    RECT 490.8000 281.6000 491.6000 286.2000 ;
	    RECT 494.0000 281.6000 494.8000 285.8000 ;
	    RECT 497.2000 281.6000 498.0000 286.2000 ;
	    RECT 500.4000 281.6000 501.2000 285.8000 ;
	    RECT 503.6000 281.6000 504.4000 286.2000 ;
	    RECT 506.8000 281.6000 507.6000 285.8000 ;
	    RECT 0.4000 280.4000 514.8000 281.6000 ;
	    RECT 2.8000 273.0000 3.6000 280.4000 ;
	    RECT 6.6000 275.8000 7.4000 280.4000 ;
	    RECT 10.8000 271.8000 11.6000 280.4000 ;
	    RECT 12.4000 271.8000 13.2000 280.4000 ;
	    RECT 16.6000 275.8000 17.4000 280.4000 ;
	    RECT 20.4000 271.8000 21.2000 280.4000 ;
	    RECT 26.0000 275.8000 26.8000 280.4000 ;
	    RECT 29.2000 275.8000 30.0000 280.4000 ;
	    RECT 34.8000 272.0000 35.6000 280.4000 ;
	    RECT 38.6000 275.8000 39.4000 280.4000 ;
	    RECT 42.8000 271.8000 43.6000 280.4000 ;
	    RECT 45.0000 275.8000 45.8000 280.4000 ;
	    RECT 49.2000 271.8000 50.0000 280.4000 ;
	    RECT 50.8000 271.8000 51.6000 280.4000 ;
	    RECT 55.0000 275.8000 55.8000 280.4000 ;
	    RECT 57.8000 275.8000 58.6000 280.4000 ;
	    RECT 62.0000 271.8000 62.8000 280.4000 ;
	    RECT 64.2000 275.8000 65.0000 280.4000 ;
	    RECT 68.4000 271.8000 69.2000 280.4000 ;
	    RECT 70.6000 275.8000 71.4000 280.4000 ;
	    RECT 74.8000 271.8000 75.6000 280.4000 ;
	    RECT 77.0000 275.8000 77.8000 280.4000 ;
	    RECT 81.2000 271.8000 82.0000 280.4000 ;
	    RECT 83.4000 275.8000 84.2000 280.4000 ;
	    RECT 87.6000 271.8000 88.4000 280.4000 ;
	    RECT 89.8000 275.8000 90.6000 280.4000 ;
	    RECT 94.0000 271.8000 94.8000 280.4000 ;
	    RECT 97.2000 272.0000 98.0000 280.4000 ;
	    RECT 102.8000 275.8000 103.6000 280.4000 ;
	    RECT 106.0000 275.8000 106.8000 280.4000 ;
	    RECT 111.6000 271.8000 112.4000 280.4000 ;
	    RECT 121.2000 271.8000 122.0000 280.4000 ;
	    RECT 125.4000 275.8000 126.2000 280.4000 ;
	    RECT 127.6000 271.8000 128.4000 280.4000 ;
	    RECT 134.0000 271.8000 134.8000 280.4000 ;
	    RECT 135.6000 271.8000 136.4000 280.4000 ;
	    RECT 140.4000 271.8000 141.2000 280.4000 ;
	    RECT 145.2000 271.8000 146.0000 280.4000 ;
	    RECT 151.6000 273.0000 152.4000 280.4000 ;
	    RECT 156.4000 272.0000 157.2000 280.4000 ;
	    RECT 162.0000 275.8000 162.8000 280.4000 ;
	    RECT 165.2000 275.8000 166.0000 280.4000 ;
	    RECT 170.8000 271.8000 171.6000 280.4000 ;
	    RECT 177.2000 271.8000 178.0000 280.4000 ;
	    RECT 178.8000 271.8000 179.6000 280.4000 ;
	    RECT 185.2000 271.8000 186.0000 280.4000 ;
	    RECT 187.4000 275.8000 188.2000 280.4000 ;
	    RECT 191.6000 271.8000 192.4000 280.4000 ;
	    RECT 193.8000 275.8000 194.6000 280.4000 ;
	    RECT 198.0000 271.8000 198.8000 280.4000 ;
	    RECT 199.6000 271.8000 200.4000 280.4000 ;
	    RECT 204.4000 271.8000 205.2000 280.4000 ;
	    RECT 209.8000 275.8000 210.6000 280.4000 ;
	    RECT 214.0000 271.8000 214.8000 280.4000 ;
	    RECT 215.6000 271.8000 216.4000 280.4000 ;
	    RECT 222.0000 271.8000 222.8000 280.4000 ;
	    RECT 225.2000 272.2000 226.0000 280.4000 ;
	    RECT 230.4000 271.8000 231.2000 280.4000 ;
	    RECT 234.8000 272.2000 235.6000 280.4000 ;
	    RECT 240.0000 271.8000 240.8000 280.4000 ;
	    RECT 244.4000 272.2000 245.2000 280.4000 ;
	    RECT 249.6000 271.8000 250.4000 280.4000 ;
	    RECT 254.0000 273.0000 254.8000 280.4000 ;
	    RECT 265.2000 271.8000 266.0000 280.4000 ;
	    RECT 270.8000 275.8000 271.6000 280.4000 ;
	    RECT 274.0000 275.8000 274.8000 280.4000 ;
	    RECT 279.6000 272.0000 280.4000 280.4000 ;
	    RECT 282.8000 275.8000 283.6000 280.4000 ;
	    RECT 286.0000 275.8000 286.8000 280.4000 ;
	    RECT 288.2000 275.8000 289.0000 280.4000 ;
	    RECT 292.4000 271.8000 293.2000 280.4000 ;
	    RECT 294.0000 271.8000 294.8000 280.4000 ;
	    RECT 300.4000 271.8000 301.2000 280.4000 ;
	    RECT 302.0000 271.8000 302.8000 280.4000 ;
	    RECT 306.2000 275.8000 307.0000 280.4000 ;
	    RECT 311.6000 271.8000 312.4000 280.4000 ;
	    RECT 316.4000 271.8000 317.2000 280.4000 ;
	    RECT 318.0000 271.8000 318.8000 280.4000 ;
	    RECT 324.4000 271.8000 325.2000 280.4000 ;
	    RECT 326.6000 275.8000 327.4000 280.4000 ;
	    RECT 330.8000 271.8000 331.6000 280.4000 ;
	    RECT 334.0000 271.8000 334.8000 280.4000 ;
	    RECT 339.6000 275.8000 340.4000 280.4000 ;
	    RECT 342.8000 275.8000 343.6000 280.4000 ;
	    RECT 348.4000 272.0000 349.2000 280.4000 ;
	    RECT 352.2000 275.8000 353.0000 280.4000 ;
	    RECT 356.4000 271.8000 357.2000 280.4000 ;
	    RECT 358.6000 275.8000 359.4000 280.4000 ;
	    RECT 362.8000 271.8000 363.6000 280.4000 ;
	    RECT 364.4000 275.8000 365.2000 280.4000 ;
	    RECT 367.6000 275.8000 368.4000 280.4000 ;
	    RECT 369.8000 275.8000 370.6000 280.4000 ;
	    RECT 374.0000 271.8000 374.8000 280.4000 ;
	    RECT 377.2000 273.0000 378.0000 280.4000 ;
	    RECT 382.6000 271.8000 383.4000 280.4000 ;
	    RECT 386.8000 271.8000 387.6000 280.4000 ;
	    RECT 391.0000 275.8000 391.8000 280.4000 ;
	    RECT 393.8000 275.8000 394.6000 280.4000 ;
	    RECT 398.0000 271.8000 398.8000 280.4000 ;
	    RECT 399.6000 275.8000 400.4000 280.4000 ;
	    RECT 402.8000 275.8000 403.6000 280.4000 ;
	    RECT 411.4000 275.8000 412.2000 280.4000 ;
	    RECT 415.6000 271.8000 416.4000 280.4000 ;
	    RECT 417.2000 275.8000 418.0000 280.4000 ;
	    RECT 420.4000 275.8000 421.2000 280.4000 ;
	    RECT 422.6000 275.8000 423.4000 280.4000 ;
	    RECT 426.8000 271.8000 427.6000 280.4000 ;
	    RECT 429.0000 275.8000 429.8000 280.4000 ;
	    RECT 433.2000 271.8000 434.0000 280.4000 ;
	    RECT 434.8000 271.8000 435.6000 280.4000 ;
	    RECT 438.0000 271.8000 438.8000 280.4000 ;
	    RECT 441.2000 271.8000 442.0000 280.4000 ;
	    RECT 444.4000 271.8000 445.2000 280.4000 ;
	    RECT 447.6000 271.8000 448.4000 280.4000 ;
	    RECT 449.2000 271.8000 450.0000 280.4000 ;
	    RECT 453.4000 275.8000 454.2000 280.4000 ;
	    RECT 455.6000 275.8000 456.4000 280.4000 ;
	    RECT 458.8000 276.2000 459.6000 280.4000 ;
	    RECT 463.6000 273.0000 464.4000 280.4000 ;
	    RECT 468.4000 273.0000 469.2000 280.4000 ;
	    RECT 473.2000 271.8000 474.0000 280.4000 ;
	    RECT 478.8000 275.8000 479.6000 280.4000 ;
	    RECT 482.0000 275.8000 482.8000 280.4000 ;
	    RECT 487.6000 272.0000 488.4000 280.4000 ;
	    RECT 490.8000 275.8000 491.6000 280.4000 ;
	    RECT 494.0000 271.8000 494.8000 280.4000 ;
	    RECT 498.2000 275.8000 499.0000 280.4000 ;
	    RECT 502.0000 273.0000 502.8000 280.4000 ;
	    RECT 506.8000 273.0000 507.6000 280.4000 ;
	    RECT 2.8000 241.6000 3.6000 249.0000 ;
	    RECT 7.6000 241.6000 8.4000 249.0000 ;
	    RECT 12.4000 241.6000 13.2000 250.2000 ;
	    RECT 18.0000 241.6000 18.8000 246.2000 ;
	    RECT 21.2000 241.6000 22.0000 246.2000 ;
	    RECT 26.8000 241.6000 27.6000 250.0000 ;
	    RECT 30.6000 241.6000 31.4000 246.2000 ;
	    RECT 34.8000 241.6000 35.6000 250.2000 ;
	    RECT 36.4000 241.6000 37.2000 250.2000 ;
	    RECT 39.6000 241.6000 40.4000 250.2000 ;
	    RECT 42.8000 241.6000 43.6000 250.2000 ;
	    RECT 46.0000 241.6000 46.8000 250.2000 ;
	    RECT 49.2000 241.6000 50.0000 250.2000 ;
	    RECT 51.4000 241.6000 52.2000 246.2000 ;
	    RECT 55.6000 241.6000 56.4000 250.2000 ;
	    RECT 57.8000 241.6000 58.6000 246.2000 ;
	    RECT 62.0000 241.6000 62.8000 250.2000 ;
	    RECT 63.6000 241.6000 64.4000 250.2000 ;
	    RECT 70.0000 241.6000 70.8000 250.0000 ;
	    RECT 75.6000 241.6000 76.4000 246.2000 ;
	    RECT 78.8000 241.6000 79.6000 246.2000 ;
	    RECT 84.4000 241.6000 85.2000 250.2000 ;
	    RECT 87.6000 241.6000 88.4000 246.2000 ;
	    RECT 90.8000 241.6000 91.6000 246.2000 ;
	    RECT 93.0000 241.6000 93.8000 246.2000 ;
	    RECT 97.2000 241.6000 98.0000 250.2000 ;
	    RECT 100.4000 241.6000 101.2000 249.8000 ;
	    RECT 105.6000 241.6000 106.4000 250.2000 ;
	    RECT 114.8000 241.6000 115.6000 250.2000 ;
	    RECT 121.2000 241.6000 122.0000 250.2000 ;
	    RECT 124.4000 241.6000 125.2000 249.8000 ;
	    RECT 129.6000 241.6000 130.4000 250.2000 ;
	    RECT 132.4000 241.6000 133.2000 250.2000 ;
	    RECT 140.4000 241.6000 141.2000 250.2000 ;
	    RECT 143.6000 241.6000 144.4000 250.2000 ;
	    RECT 149.2000 241.6000 150.0000 246.2000 ;
	    RECT 152.4000 241.6000 153.2000 246.2000 ;
	    RECT 158.0000 241.6000 158.8000 250.0000 ;
	    RECT 161.2000 241.6000 162.0000 250.2000 ;
	    RECT 165.4000 241.6000 166.2000 246.2000 ;
	    RECT 168.2000 241.6000 169.0000 246.2000 ;
	    RECT 172.4000 241.6000 173.2000 250.2000 ;
	    RECT 175.6000 241.6000 176.4000 249.0000 ;
	    RECT 180.4000 241.6000 181.2000 249.0000 ;
	    RECT 185.2000 241.6000 186.0000 249.0000 ;
	    RECT 190.0000 241.6000 190.8000 249.0000 ;
	    RECT 193.8000 241.6000 194.6000 246.2000 ;
	    RECT 198.0000 241.6000 198.8000 250.2000 ;
	    RECT 201.2000 241.6000 202.0000 249.0000 ;
	    RECT 205.6000 241.6000 206.4000 250.2000 ;
	    RECT 210.8000 241.6000 211.6000 249.8000 ;
	    RECT 215.6000 241.6000 216.4000 249.8000 ;
	    RECT 220.8000 241.6000 221.6000 250.2000 ;
	    RECT 223.6000 241.6000 224.4000 250.2000 ;
	    RECT 230.0000 241.6000 230.8000 250.2000 ;
	    RECT 232.2000 241.6000 233.0000 246.2000 ;
	    RECT 236.4000 241.6000 237.2000 250.2000 ;
	    RECT 238.0000 241.6000 238.8000 250.2000 ;
	    RECT 242.2000 241.6000 243.0000 246.2000 ;
	    RECT 244.4000 241.6000 245.2000 250.2000 ;
	    RECT 250.8000 241.6000 251.6000 250.2000 ;
	    RECT 255.6000 241.6000 256.4000 250.2000 ;
	    RECT 266.8000 241.6000 267.6000 250.2000 ;
	    RECT 270.0000 241.6000 270.8000 249.0000 ;
	    RECT 274.8000 241.6000 275.6000 250.2000 ;
	    RECT 280.4000 241.6000 281.2000 246.2000 ;
	    RECT 283.6000 241.6000 284.4000 246.2000 ;
	    RECT 289.2000 241.6000 290.0000 250.0000 ;
	    RECT 292.4000 241.6000 293.2000 246.2000 ;
	    RECT 295.6000 241.6000 296.4000 246.2000 ;
	    RECT 297.8000 241.6000 298.6000 246.2000 ;
	    RECT 302.0000 241.6000 302.8000 250.2000 ;
	    RECT 305.2000 241.6000 306.0000 249.0000 ;
	    RECT 310.0000 241.6000 310.8000 249.0000 ;
	    RECT 314.8000 241.6000 315.6000 250.2000 ;
	    RECT 320.4000 241.6000 321.2000 246.2000 ;
	    RECT 323.6000 241.6000 324.4000 246.2000 ;
	    RECT 329.2000 241.6000 330.0000 250.0000 ;
	    RECT 332.4000 241.6000 333.2000 246.2000 ;
	    RECT 335.6000 241.6000 336.4000 246.2000 ;
	    RECT 337.8000 241.6000 338.6000 246.2000 ;
	    RECT 342.0000 241.6000 342.8000 250.2000 ;
	    RECT 345.2000 241.6000 346.0000 249.0000 ;
	    RECT 350.6000 241.6000 351.4000 250.2000 ;
	    RECT 356.4000 241.6000 357.2000 250.2000 ;
	    RECT 362.0000 241.6000 362.8000 246.2000 ;
	    RECT 365.2000 241.6000 366.0000 246.2000 ;
	    RECT 370.8000 241.6000 371.6000 250.0000 ;
	    RECT 375.6000 241.6000 376.4000 250.2000 ;
	    RECT 381.2000 241.6000 382.0000 246.2000 ;
	    RECT 384.4000 241.6000 385.2000 246.2000 ;
	    RECT 390.0000 241.6000 390.8000 250.0000 ;
	    RECT 394.8000 241.6000 395.6000 250.2000 ;
	    RECT 400.4000 241.6000 401.2000 246.2000 ;
	    RECT 403.6000 241.6000 404.4000 246.2000 ;
	    RECT 409.2000 241.6000 410.0000 250.0000 ;
	    RECT 419.4000 241.6000 420.2000 246.2000 ;
	    RECT 423.6000 241.6000 424.4000 250.2000 ;
	    RECT 426.8000 241.6000 427.6000 250.2000 ;
	    RECT 430.0000 241.6000 430.8000 250.2000 ;
	    RECT 435.6000 241.6000 436.4000 246.2000 ;
	    RECT 438.8000 241.6000 439.6000 246.2000 ;
	    RECT 444.4000 241.6000 445.2000 250.0000 ;
	    RECT 447.6000 241.6000 448.4000 246.2000 ;
	    RECT 452.4000 241.6000 453.2000 250.2000 ;
	    RECT 458.0000 241.6000 458.8000 246.2000 ;
	    RECT 461.2000 241.6000 462.0000 246.2000 ;
	    RECT 466.8000 241.6000 467.6000 250.0000 ;
	    RECT 470.0000 241.6000 470.8000 246.2000 ;
	    RECT 473.2000 241.6000 474.0000 250.2000 ;
	    RECT 477.4000 241.6000 478.2000 246.2000 ;
	    RECT 481.2000 241.6000 482.0000 250.2000 ;
	    RECT 486.8000 241.6000 487.6000 246.2000 ;
	    RECT 490.0000 241.6000 490.8000 246.2000 ;
	    RECT 495.6000 241.6000 496.4000 250.0000 ;
	    RECT 500.4000 241.6000 501.2000 245.8000 ;
	    RECT 503.6000 241.6000 504.4000 246.2000 ;
	    RECT 505.8000 241.6000 506.6000 246.2000 ;
	    RECT 510.0000 241.6000 510.8000 250.2000 ;
	    RECT 513.2000 241.6000 514.0000 246.2000 ;
	    RECT 0.4000 240.4000 514.8000 241.6000 ;
	    RECT 2.8000 233.0000 3.6000 240.4000 ;
	    RECT 7.6000 233.0000 8.4000 240.4000 ;
	    RECT 10.8000 231.8000 11.6000 240.4000 ;
	    RECT 15.0000 235.8000 15.8000 240.4000 ;
	    RECT 17.2000 231.8000 18.0000 240.4000 ;
	    RECT 21.4000 235.8000 22.2000 240.4000 ;
	    RECT 25.2000 231.8000 26.0000 240.4000 ;
	    RECT 30.8000 235.8000 31.6000 240.4000 ;
	    RECT 34.0000 235.8000 34.8000 240.4000 ;
	    RECT 39.6000 232.0000 40.4000 240.4000 ;
	    RECT 42.8000 231.8000 43.6000 240.4000 ;
	    RECT 47.0000 235.8000 47.8000 240.4000 ;
	    RECT 49.8000 235.8000 50.6000 240.4000 ;
	    RECT 54.0000 231.8000 54.8000 240.4000 ;
	    RECT 56.2000 235.8000 57.0000 240.4000 ;
	    RECT 60.4000 231.8000 61.2000 240.4000 ;
	    RECT 63.6000 231.8000 64.4000 240.4000 ;
	    RECT 69.2000 235.8000 70.0000 240.4000 ;
	    RECT 72.4000 235.8000 73.2000 240.4000 ;
	    RECT 78.0000 232.0000 78.8000 240.4000 ;
	    RECT 81.8000 235.8000 82.6000 240.4000 ;
	    RECT 86.0000 231.8000 86.8000 240.4000 ;
	    RECT 88.2000 235.8000 89.0000 240.4000 ;
	    RECT 92.4000 231.8000 93.2000 240.4000 ;
	    RECT 94.6000 235.8000 95.4000 240.4000 ;
	    RECT 98.8000 231.8000 99.6000 240.4000 ;
	    RECT 108.4000 232.0000 109.2000 240.4000 ;
	    RECT 114.0000 235.8000 114.8000 240.4000 ;
	    RECT 117.2000 235.8000 118.0000 240.4000 ;
	    RECT 122.8000 231.8000 123.6000 240.4000 ;
	    RECT 126.0000 231.8000 126.8000 240.4000 ;
	    RECT 132.4000 231.8000 133.2000 240.4000 ;
	    RECT 134.6000 235.8000 135.4000 240.4000 ;
	    RECT 138.8000 231.8000 139.6000 240.4000 ;
	    RECT 140.4000 231.8000 141.2000 240.4000 ;
	    RECT 144.6000 235.8000 145.4000 240.4000 ;
	    RECT 150.0000 231.8000 150.8000 240.4000 ;
	    RECT 151.6000 231.8000 152.4000 240.4000 ;
	    RECT 157.6000 231.8000 158.4000 240.4000 ;
	    RECT 162.8000 232.2000 163.6000 240.4000 ;
	    RECT 166.0000 231.8000 166.8000 240.4000 ;
	    RECT 172.4000 231.8000 173.2000 240.4000 ;
	    RECT 174.0000 231.8000 174.8000 240.4000 ;
	    RECT 179.4000 235.8000 180.2000 240.4000 ;
	    RECT 183.6000 231.8000 184.4000 240.4000 ;
	    RECT 185.2000 235.8000 186.0000 240.4000 ;
	    RECT 188.4000 235.8000 189.2000 240.4000 ;
	    RECT 190.6000 235.8000 191.4000 240.4000 ;
	    RECT 194.8000 231.8000 195.6000 240.4000 ;
	    RECT 198.0000 233.0000 198.8000 240.4000 ;
	    RECT 204.4000 231.8000 205.2000 240.4000 ;
	    RECT 206.0000 231.8000 206.8000 240.4000 ;
	    RECT 212.4000 231.8000 213.2000 240.4000 ;
	    RECT 214.6000 235.8000 215.4000 240.4000 ;
	    RECT 218.8000 231.8000 219.6000 240.4000 ;
	    RECT 220.4000 231.8000 221.2000 240.4000 ;
	    RECT 226.8000 231.8000 227.6000 240.4000 ;
	    RECT 229.0000 235.8000 229.8000 240.4000 ;
	    RECT 233.2000 231.8000 234.0000 240.4000 ;
	    RECT 234.8000 231.8000 235.6000 240.4000 ;
	    RECT 241.2000 233.0000 242.0000 240.4000 ;
	    RECT 246.0000 233.0000 246.8000 240.4000 ;
	    RECT 250.8000 233.0000 251.6000 240.4000 ;
	    RECT 260.4000 231.8000 261.2000 240.4000 ;
	    RECT 266.8000 231.8000 267.6000 240.4000 ;
	    RECT 269.0000 235.8000 269.8000 240.4000 ;
	    RECT 273.2000 231.8000 274.0000 240.4000 ;
	    RECT 278.0000 231.8000 278.8000 240.4000 ;
	    RECT 279.6000 231.8000 280.4000 240.4000 ;
	    RECT 283.8000 235.8000 284.6000 240.4000 ;
	    RECT 286.0000 231.8000 286.8000 240.4000 ;
	    RECT 292.4000 231.8000 293.2000 240.4000 ;
	    RECT 294.0000 231.8000 294.8000 240.4000 ;
	    RECT 300.4000 231.8000 301.2000 240.4000 ;
	    RECT 303.6000 232.2000 304.4000 240.4000 ;
	    RECT 308.8000 231.8000 309.6000 240.4000 ;
	    RECT 313.2000 232.2000 314.0000 240.4000 ;
	    RECT 318.4000 231.8000 319.2000 240.4000 ;
	    RECT 322.8000 233.0000 323.6000 240.4000 ;
	    RECT 327.6000 231.8000 328.4000 240.4000 ;
	    RECT 333.2000 235.8000 334.0000 240.4000 ;
	    RECT 336.4000 235.8000 337.2000 240.4000 ;
	    RECT 342.0000 232.0000 342.8000 240.4000 ;
	    RECT 345.2000 231.8000 346.0000 240.4000 ;
	    RECT 349.4000 235.8000 350.2000 240.4000 ;
	    RECT 352.2000 235.8000 353.0000 240.4000 ;
	    RECT 356.4000 231.8000 357.2000 240.4000 ;
	    RECT 359.6000 233.0000 360.4000 240.4000 ;
	    RECT 364.4000 231.8000 365.2000 240.4000 ;
	    RECT 370.0000 235.8000 370.8000 240.4000 ;
	    RECT 373.2000 235.8000 374.0000 240.4000 ;
	    RECT 378.8000 232.0000 379.6000 240.4000 ;
	    RECT 382.0000 235.8000 382.8000 240.4000 ;
	    RECT 385.2000 231.8000 386.0000 240.4000 ;
	    RECT 389.4000 235.8000 390.2000 240.4000 ;
	    RECT 393.2000 233.0000 394.0000 240.4000 ;
	    RECT 396.4000 235.8000 397.2000 240.4000 ;
	    RECT 399.6000 235.8000 400.4000 240.4000 ;
	    RECT 401.8000 235.8000 402.6000 240.4000 ;
	    RECT 406.0000 231.8000 406.8000 240.4000 ;
	    RECT 415.6000 231.8000 416.4000 240.4000 ;
	    RECT 421.2000 235.8000 422.0000 240.4000 ;
	    RECT 424.4000 235.8000 425.2000 240.4000 ;
	    RECT 430.0000 232.0000 430.8000 240.4000 ;
	    RECT 434.8000 236.2000 435.6000 240.4000 ;
	    RECT 438.0000 235.8000 438.8000 240.4000 ;
	    RECT 441.2000 236.2000 442.0000 240.4000 ;
	    RECT 444.4000 235.8000 445.2000 240.4000 ;
	    RECT 447.6000 233.0000 448.4000 240.4000 ;
	    RECT 451.4000 235.8000 452.2000 240.4000 ;
	    RECT 455.6000 231.8000 456.4000 240.4000 ;
	    RECT 458.8000 235.8000 459.6000 240.4000 ;
	    RECT 462.0000 231.8000 462.8000 240.4000 ;
	    RECT 467.6000 235.8000 468.4000 240.4000 ;
	    RECT 470.8000 235.8000 471.6000 240.4000 ;
	    RECT 476.4000 232.0000 477.2000 240.4000 ;
	    RECT 481.2000 236.2000 482.0000 240.4000 ;
	    RECT 484.4000 235.8000 485.2000 240.4000 ;
	    RECT 486.6000 235.8000 487.4000 240.4000 ;
	    RECT 490.8000 231.8000 491.6000 240.4000 ;
	    RECT 494.0000 235.8000 494.8000 240.4000 ;
	    RECT 497.2000 232.0000 498.0000 240.4000 ;
	    RECT 502.8000 235.8000 503.6000 240.4000 ;
	    RECT 506.0000 235.8000 506.8000 240.4000 ;
	    RECT 511.6000 231.8000 512.4000 240.4000 ;
	    RECT 2.8000 201.6000 3.6000 209.0000 ;
	    RECT 7.6000 201.6000 8.4000 209.0000 ;
	    RECT 10.8000 201.6000 11.6000 210.2000 ;
	    RECT 15.0000 201.6000 15.8000 206.2000 ;
	    RECT 18.8000 201.6000 19.6000 210.2000 ;
	    RECT 24.4000 201.6000 25.2000 206.2000 ;
	    RECT 27.6000 201.6000 28.4000 206.2000 ;
	    RECT 33.2000 201.6000 34.0000 210.0000 ;
	    RECT 37.0000 201.6000 37.8000 206.2000 ;
	    RECT 41.2000 201.6000 42.0000 210.2000 ;
	    RECT 44.4000 201.6000 45.2000 209.0000 ;
	    RECT 48.2000 201.6000 49.0000 206.2000 ;
	    RECT 52.4000 201.6000 53.2000 210.2000 ;
	    RECT 57.2000 201.6000 58.0000 210.2000 ;
	    RECT 58.8000 201.6000 59.6000 210.2000 ;
	    RECT 65.2000 201.6000 66.0000 209.0000 ;
	    RECT 70.0000 201.6000 70.8000 209.0000 ;
	    RECT 74.8000 201.6000 75.6000 210.0000 ;
	    RECT 80.4000 201.6000 81.2000 206.2000 ;
	    RECT 83.6000 201.6000 84.4000 206.2000 ;
	    RECT 89.2000 201.6000 90.0000 210.2000 ;
	    RECT 92.4000 201.6000 93.2000 206.2000 ;
	    RECT 95.6000 201.6000 96.4000 206.2000 ;
	    RECT 97.2000 201.6000 98.0000 206.2000 ;
	    RECT 100.4000 201.6000 101.2000 206.2000 ;
	    RECT 102.6000 201.6000 103.4000 206.2000 ;
	    RECT 106.8000 201.6000 107.6000 210.2000 ;
	    RECT 114.8000 201.6000 115.6000 210.2000 ;
	    RECT 121.2000 201.6000 122.0000 210.2000 ;
	    RECT 123.4000 201.6000 124.2000 206.2000 ;
	    RECT 127.6000 201.6000 128.4000 210.2000 ;
	    RECT 130.8000 201.6000 131.6000 210.0000 ;
	    RECT 136.4000 201.6000 137.2000 206.2000 ;
	    RECT 139.6000 201.6000 140.4000 206.2000 ;
	    RECT 145.2000 201.6000 146.0000 210.2000 ;
	    RECT 151.6000 201.6000 152.4000 210.2000 ;
	    RECT 154.4000 201.6000 155.2000 210.2000 ;
	    RECT 159.6000 201.6000 160.4000 209.8000 ;
	    RECT 164.4000 201.6000 165.2000 209.0000 ;
	    RECT 169.2000 201.6000 170.0000 210.0000 ;
	    RECT 174.8000 201.6000 175.6000 206.2000 ;
	    RECT 178.0000 201.6000 178.8000 206.2000 ;
	    RECT 183.6000 201.6000 184.4000 210.2000 ;
	    RECT 188.4000 201.6000 189.2000 209.0000 ;
	    RECT 193.2000 201.6000 194.0000 209.0000 ;
	    RECT 196.4000 201.6000 197.2000 206.2000 ;
	    RECT 199.6000 201.6000 200.4000 206.2000 ;
	    RECT 201.8000 201.6000 202.6000 206.2000 ;
	    RECT 206.0000 201.6000 206.8000 210.2000 ;
	    RECT 207.6000 201.6000 208.4000 210.2000 ;
	    RECT 212.4000 201.6000 213.2000 206.2000 ;
	    RECT 215.6000 201.6000 216.4000 206.2000 ;
	    RECT 217.8000 201.6000 218.6000 206.2000 ;
	    RECT 222.0000 201.6000 222.8000 210.2000 ;
	    RECT 225.2000 201.6000 226.0000 210.0000 ;
	    RECT 230.8000 201.6000 231.6000 206.2000 ;
	    RECT 234.0000 201.6000 234.8000 206.2000 ;
	    RECT 239.6000 201.6000 240.4000 210.2000 ;
	    RECT 244.0000 201.6000 244.8000 210.2000 ;
	    RECT 249.2000 201.6000 250.0000 209.8000 ;
	    RECT 260.0000 201.6000 260.8000 210.2000 ;
	    RECT 265.2000 201.6000 266.0000 209.8000 ;
	    RECT 270.0000 201.6000 270.8000 209.0000 ;
	    RECT 274.8000 201.6000 275.6000 209.0000 ;
	    RECT 278.0000 201.6000 278.8000 206.2000 ;
	    RECT 281.2000 201.6000 282.0000 206.2000 ;
	    RECT 283.4000 201.6000 284.2000 206.2000 ;
	    RECT 287.6000 201.6000 288.4000 210.2000 ;
	    RECT 290.8000 201.6000 291.6000 210.2000 ;
	    RECT 296.4000 201.6000 297.2000 206.2000 ;
	    RECT 299.6000 201.6000 300.4000 206.2000 ;
	    RECT 305.2000 201.6000 306.0000 210.0000 ;
	    RECT 310.0000 201.6000 310.8000 209.8000 ;
	    RECT 315.2000 201.6000 316.0000 210.2000 ;
	    RECT 319.6000 201.6000 320.4000 209.8000 ;
	    RECT 324.8000 201.6000 325.6000 210.2000 ;
	    RECT 329.2000 201.6000 330.0000 210.2000 ;
	    RECT 334.8000 201.6000 335.6000 206.2000 ;
	    RECT 338.0000 201.6000 338.8000 206.2000 ;
	    RECT 343.6000 201.6000 344.4000 210.0000 ;
	    RECT 346.8000 201.6000 347.6000 210.2000 ;
	    RECT 351.0000 201.6000 351.8000 206.2000 ;
	    RECT 353.8000 201.6000 354.6000 206.2000 ;
	    RECT 358.0000 201.6000 358.8000 210.2000 ;
	    RECT 361.2000 201.6000 362.0000 209.0000 ;
	    RECT 366.0000 201.6000 366.8000 210.2000 ;
	    RECT 371.6000 201.6000 372.4000 206.2000 ;
	    RECT 374.8000 201.6000 375.6000 206.2000 ;
	    RECT 380.4000 201.6000 381.2000 210.0000 ;
	    RECT 383.6000 201.6000 384.4000 206.2000 ;
	    RECT 386.8000 201.6000 387.6000 206.2000 ;
	    RECT 389.0000 201.6000 389.8000 206.2000 ;
	    RECT 393.2000 201.6000 394.0000 210.2000 ;
	    RECT 396.4000 201.6000 397.2000 209.0000 ;
	    RECT 399.6000 201.6000 400.4000 206.2000 ;
	    RECT 402.8000 201.6000 403.6000 206.2000 ;
	    RECT 411.4000 201.6000 412.2000 206.2000 ;
	    RECT 415.6000 201.6000 416.4000 210.2000 ;
	    RECT 418.8000 201.6000 419.6000 210.2000 ;
	    RECT 424.4000 201.6000 425.2000 206.2000 ;
	    RECT 427.6000 201.6000 428.4000 206.2000 ;
	    RECT 433.2000 201.6000 434.0000 210.0000 ;
	    RECT 438.0000 201.6000 438.8000 210.2000 ;
	    RECT 439.6000 201.6000 440.4000 206.2000 ;
	    RECT 442.8000 201.6000 443.6000 206.2000 ;
	    RECT 444.4000 201.6000 445.2000 206.2000 ;
	    RECT 447.6000 201.6000 448.4000 205.8000 ;
	    RECT 450.8000 201.6000 451.6000 210.2000 ;
	    RECT 454.0000 201.6000 454.8000 210.2000 ;
	    RECT 457.2000 201.6000 458.0000 210.2000 ;
	    RECT 460.4000 201.6000 461.2000 210.2000 ;
	    RECT 466.0000 201.6000 466.8000 206.2000 ;
	    RECT 469.2000 201.6000 470.0000 206.2000 ;
	    RECT 474.8000 201.6000 475.6000 210.0000 ;
	    RECT 478.6000 201.6000 479.4000 206.2000 ;
	    RECT 482.8000 201.6000 483.6000 210.2000 ;
	    RECT 484.4000 201.6000 485.2000 206.2000 ;
	    RECT 487.6000 201.6000 488.4000 210.2000 ;
	    RECT 491.8000 201.6000 492.6000 206.2000 ;
	    RECT 495.6000 201.6000 496.4000 210.2000 ;
	    RECT 501.2000 201.6000 502.0000 206.2000 ;
	    RECT 504.4000 201.6000 505.2000 206.2000 ;
	    RECT 510.0000 201.6000 510.8000 210.0000 ;
	    RECT 0.4000 200.4000 514.8000 201.6000 ;
	    RECT 2.8000 193.0000 3.6000 200.4000 ;
	    RECT 7.6000 193.0000 8.4000 200.4000 ;
	    RECT 12.4000 193.0000 13.2000 200.4000 ;
	    RECT 15.6000 191.8000 16.4000 200.4000 ;
	    RECT 19.8000 195.8000 20.6000 200.4000 ;
	    RECT 23.6000 191.8000 24.4000 200.4000 ;
	    RECT 29.2000 195.8000 30.0000 200.4000 ;
	    RECT 32.4000 195.8000 33.2000 200.4000 ;
	    RECT 38.0000 192.0000 38.8000 200.4000 ;
	    RECT 42.8000 193.0000 43.6000 200.4000 ;
	    RECT 46.6000 195.8000 47.4000 200.4000 ;
	    RECT 50.8000 191.8000 51.6000 200.4000 ;
	    RECT 53.0000 195.8000 53.8000 200.4000 ;
	    RECT 57.2000 191.8000 58.0000 200.4000 ;
	    RECT 59.4000 195.8000 60.2000 200.4000 ;
	    RECT 63.6000 191.8000 64.4000 200.4000 ;
	    RECT 65.2000 191.8000 66.0000 200.4000 ;
	    RECT 71.6000 192.0000 72.4000 200.4000 ;
	    RECT 77.2000 195.8000 78.0000 200.4000 ;
	    RECT 80.4000 195.8000 81.2000 200.4000 ;
	    RECT 86.0000 191.8000 86.8000 200.4000 ;
	    RECT 90.8000 193.0000 91.6000 200.4000 ;
	    RECT 94.0000 191.8000 94.8000 200.4000 ;
	    RECT 98.2000 195.8000 99.0000 200.4000 ;
	    RECT 101.0000 195.8000 101.8000 200.4000 ;
	    RECT 105.2000 191.8000 106.0000 200.4000 ;
	    RECT 114.4000 191.8000 115.2000 200.4000 ;
	    RECT 119.6000 192.2000 120.4000 200.4000 ;
	    RECT 124.4000 192.2000 125.2000 200.4000 ;
	    RECT 129.6000 191.8000 130.4000 200.4000 ;
	    RECT 132.4000 191.8000 133.2000 200.4000 ;
	    RECT 138.8000 191.8000 139.6000 200.4000 ;
	    RECT 140.4000 191.8000 141.2000 200.4000 ;
	    RECT 144.6000 195.8000 145.4000 200.4000 ;
	    RECT 146.8000 191.8000 147.6000 200.4000 ;
	    RECT 153.2000 191.8000 154.0000 200.4000 ;
	    RECT 155.4000 195.8000 156.2000 200.4000 ;
	    RECT 159.6000 191.8000 160.4000 200.4000 ;
	    RECT 164.4000 191.8000 165.2000 200.4000 ;
	    RECT 166.0000 191.8000 166.8000 200.4000 ;
	    RECT 171.4000 195.8000 172.2000 200.4000 ;
	    RECT 175.6000 191.8000 176.4000 200.4000 ;
	    RECT 177.8000 195.8000 178.6000 200.4000 ;
	    RECT 182.0000 191.8000 182.8000 200.4000 ;
	    RECT 183.6000 191.8000 184.4000 200.4000 ;
	    RECT 187.8000 195.8000 188.6000 200.4000 ;
	    RECT 190.0000 191.8000 190.8000 200.4000 ;
	    RECT 196.4000 191.8000 197.2000 200.4000 ;
	    RECT 201.2000 191.8000 202.0000 200.4000 ;
	    RECT 202.8000 191.8000 203.6000 200.4000 ;
	    RECT 207.0000 195.8000 207.8000 200.4000 ;
	    RECT 209.2000 191.8000 210.0000 200.4000 ;
	    RECT 215.6000 191.8000 216.4000 200.4000 ;
	    RECT 217.2000 191.8000 218.0000 200.4000 ;
	    RECT 223.6000 193.0000 224.4000 200.4000 ;
	    RECT 228.4000 193.0000 229.2000 200.4000 ;
	    RECT 231.6000 191.8000 232.4000 200.4000 ;
	    RECT 238.0000 191.8000 238.8000 200.4000 ;
	    RECT 240.2000 195.8000 241.0000 200.4000 ;
	    RECT 244.4000 191.8000 245.2000 200.4000 ;
	    RECT 246.6000 195.8000 247.4000 200.4000 ;
	    RECT 250.8000 191.8000 251.6000 200.4000 ;
	    RECT 254.0000 193.0000 254.8000 200.4000 ;
	    RECT 263.6000 195.8000 264.4000 200.4000 ;
	    RECT 266.8000 195.8000 267.6000 200.4000 ;
	    RECT 270.0000 191.8000 270.8000 200.4000 ;
	    RECT 275.6000 195.8000 276.4000 200.4000 ;
	    RECT 278.8000 195.8000 279.6000 200.4000 ;
	    RECT 284.4000 192.0000 285.2000 200.4000 ;
	    RECT 289.2000 193.0000 290.0000 200.4000 ;
	    RECT 293.0000 195.8000 293.8000 200.4000 ;
	    RECT 297.2000 191.8000 298.0000 200.4000 ;
	    RECT 300.4000 193.0000 301.2000 200.4000 ;
	    RECT 305.2000 193.0000 306.0000 200.4000 ;
	    RECT 308.4000 195.8000 309.2000 200.4000 ;
	    RECT 311.6000 195.8000 312.4000 200.4000 ;
	    RECT 313.8000 195.8000 314.6000 200.4000 ;
	    RECT 318.0000 191.8000 318.8000 200.4000 ;
	    RECT 321.2000 191.8000 322.0000 200.4000 ;
	    RECT 326.8000 195.8000 327.6000 200.4000 ;
	    RECT 330.0000 195.8000 330.8000 200.4000 ;
	    RECT 335.6000 192.0000 336.4000 200.4000 ;
	    RECT 340.4000 193.0000 341.2000 200.4000 ;
	    RECT 345.2000 193.0000 346.0000 200.4000 ;
	    RECT 350.0000 193.0000 350.8000 200.4000 ;
	    RECT 353.2000 195.8000 354.0000 200.4000 ;
	    RECT 356.4000 195.8000 357.2000 200.4000 ;
	    RECT 358.6000 195.8000 359.4000 200.4000 ;
	    RECT 362.8000 191.8000 363.6000 200.4000 ;
	    RECT 366.0000 191.8000 366.8000 200.4000 ;
	    RECT 371.6000 195.8000 372.4000 200.4000 ;
	    RECT 374.8000 195.8000 375.6000 200.4000 ;
	    RECT 380.4000 192.0000 381.2000 200.4000 ;
	    RECT 383.6000 195.8000 384.4000 200.4000 ;
	    RECT 388.4000 191.8000 389.2000 200.4000 ;
	    RECT 394.0000 195.8000 394.8000 200.4000 ;
	    RECT 397.2000 195.8000 398.0000 200.4000 ;
	    RECT 402.8000 192.0000 403.6000 200.4000 ;
	    RECT 412.4000 191.8000 413.2000 200.4000 ;
	    RECT 416.6000 195.8000 417.4000 200.4000 ;
	    RECT 420.4000 193.0000 421.2000 200.4000 ;
	    RECT 425.2000 193.0000 426.0000 200.4000 ;
	    RECT 428.4000 195.8000 429.2000 200.4000 ;
	    RECT 431.6000 196.2000 432.4000 200.4000 ;
	    RECT 434.8000 195.8000 435.6000 200.4000 ;
	    RECT 438.0000 195.8000 438.8000 200.4000 ;
	    RECT 439.6000 195.8000 440.4000 200.4000 ;
	    RECT 442.8000 195.8000 443.6000 200.4000 ;
	    RECT 446.0000 191.8000 446.8000 200.4000 ;
	    RECT 449.2000 193.0000 450.0000 200.4000 ;
	    RECT 454.0000 191.8000 454.8000 200.4000 ;
	    RECT 457.2000 196.2000 458.0000 200.4000 ;
	    RECT 460.4000 195.8000 461.2000 200.4000 ;
	    RECT 463.6000 196.2000 464.4000 200.4000 ;
	    RECT 466.8000 195.8000 467.6000 200.4000 ;
	    RECT 470.0000 196.2000 470.8000 200.4000 ;
	    RECT 473.2000 195.8000 474.0000 200.4000 ;
	    RECT 474.8000 195.8000 475.6000 200.4000 ;
	    RECT 478.0000 191.8000 478.8000 200.4000 ;
	    RECT 482.2000 195.8000 483.0000 200.4000 ;
	    RECT 486.0000 191.8000 486.8000 200.4000 ;
	    RECT 491.6000 195.8000 492.4000 200.4000 ;
	    RECT 494.8000 195.8000 495.6000 200.4000 ;
	    RECT 500.4000 192.0000 501.2000 200.4000 ;
	    RECT 505.2000 196.2000 506.0000 200.4000 ;
	    RECT 508.4000 195.8000 509.2000 200.4000 ;
	    RECT 511.6000 193.0000 512.4000 200.4000 ;
	    RECT 1.2000 161.6000 2.0000 170.2000 ;
	    RECT 4.4000 161.6000 5.2000 170.2000 ;
	    RECT 7.6000 161.6000 8.4000 170.2000 ;
	    RECT 9.2000 161.6000 10.0000 166.2000 ;
	    RECT 12.4000 161.6000 13.2000 166.2000 ;
	    RECT 14.0000 161.6000 14.8000 166.2000 ;
	    RECT 17.2000 161.6000 18.0000 169.8000 ;
	    RECT 23.6000 161.6000 24.4000 170.2000 ;
	    RECT 25.2000 161.6000 26.0000 166.2000 ;
	    RECT 28.4000 161.6000 29.2000 166.2000 ;
	    RECT 30.6000 161.6000 31.4000 166.2000 ;
	    RECT 34.8000 161.6000 35.6000 170.2000 ;
	    RECT 38.0000 161.6000 38.8000 170.0000 ;
	    RECT 43.6000 161.6000 44.4000 166.2000 ;
	    RECT 46.8000 161.6000 47.6000 166.2000 ;
	    RECT 52.4000 161.6000 53.2000 170.2000 ;
	    RECT 57.2000 161.6000 58.0000 170.2000 ;
	    RECT 62.8000 161.6000 63.6000 166.2000 ;
	    RECT 66.0000 161.6000 66.8000 166.2000 ;
	    RECT 71.6000 161.6000 72.4000 170.0000 ;
	    RECT 74.8000 161.6000 75.6000 166.2000 ;
	    RECT 78.0000 161.6000 78.8000 166.2000 ;
	    RECT 80.2000 161.6000 81.0000 166.2000 ;
	    RECT 84.4000 161.6000 85.2000 170.2000 ;
	    RECT 87.6000 161.6000 88.4000 170.0000 ;
	    RECT 93.2000 161.6000 94.0000 166.2000 ;
	    RECT 96.4000 161.6000 97.2000 166.2000 ;
	    RECT 102.0000 161.6000 102.8000 170.2000 ;
	    RECT 111.6000 161.6000 112.4000 170.2000 ;
	    RECT 115.8000 161.6000 116.6000 166.2000 ;
	    RECT 118.0000 161.6000 118.8000 166.2000 ;
	    RECT 121.2000 161.6000 122.0000 166.2000 ;
	    RECT 124.4000 161.6000 125.2000 170.2000 ;
	    RECT 130.0000 161.6000 130.8000 166.2000 ;
	    RECT 133.2000 161.6000 134.0000 166.2000 ;
	    RECT 138.8000 161.6000 139.6000 170.0000 ;
	    RECT 142.0000 161.6000 142.8000 166.2000 ;
	    RECT 145.2000 161.6000 146.0000 166.2000 ;
	    RECT 147.4000 161.6000 148.2000 166.2000 ;
	    RECT 151.6000 161.6000 152.4000 170.2000 ;
	    RECT 154.8000 161.6000 155.6000 169.0000 ;
	    RECT 159.6000 161.6000 160.4000 170.2000 ;
	    RECT 165.2000 161.6000 166.0000 166.2000 ;
	    RECT 168.4000 161.6000 169.2000 166.2000 ;
	    RECT 174.0000 161.6000 174.8000 170.0000 ;
	    RECT 178.8000 161.6000 179.6000 169.0000 ;
	    RECT 183.2000 161.6000 184.0000 170.2000 ;
	    RECT 188.4000 161.6000 189.2000 169.8000 ;
	    RECT 192.8000 161.6000 193.6000 170.2000 ;
	    RECT 198.0000 161.6000 198.8000 169.8000 ;
	    RECT 202.8000 161.6000 203.6000 169.0000 ;
	    RECT 206.0000 161.6000 206.8000 170.2000 ;
	    RECT 209.2000 161.6000 210.0000 170.2000 ;
	    RECT 212.4000 161.6000 213.2000 170.2000 ;
	    RECT 214.0000 161.6000 214.8000 166.2000 ;
	    RECT 217.2000 161.6000 218.0000 166.2000 ;
	    RECT 219.4000 161.6000 220.2000 166.2000 ;
	    RECT 223.6000 161.6000 224.4000 170.2000 ;
	    RECT 226.8000 161.6000 227.6000 170.2000 ;
	    RECT 232.4000 161.6000 233.2000 166.2000 ;
	    RECT 235.6000 161.6000 236.4000 166.2000 ;
	    RECT 241.2000 161.6000 242.0000 170.0000 ;
	    RECT 244.4000 161.6000 245.2000 170.2000 ;
	    RECT 250.8000 161.6000 251.6000 170.2000 ;
	    RECT 255.6000 161.6000 256.4000 170.2000 ;
	    RECT 263.6000 161.6000 264.4000 170.2000 ;
	    RECT 270.0000 161.6000 270.8000 170.2000 ;
	    RECT 275.6000 161.6000 276.4000 166.2000 ;
	    RECT 278.8000 161.6000 279.6000 166.2000 ;
	    RECT 284.4000 161.6000 285.2000 170.0000 ;
	    RECT 287.6000 161.6000 288.4000 170.2000 ;
	    RECT 291.8000 161.6000 292.6000 166.2000 ;
	    RECT 294.6000 161.6000 295.4000 166.2000 ;
	    RECT 298.8000 161.6000 299.6000 170.2000 ;
	    RECT 302.0000 161.6000 302.8000 170.0000 ;
	    RECT 307.6000 161.6000 308.4000 166.2000 ;
	    RECT 310.8000 161.6000 311.6000 166.2000 ;
	    RECT 316.4000 161.6000 317.2000 170.2000 ;
	    RECT 319.6000 161.6000 320.4000 170.2000 ;
	    RECT 326.0000 161.6000 326.8000 169.0000 ;
	    RECT 330.8000 161.6000 331.6000 170.2000 ;
	    RECT 333.6000 161.6000 334.4000 170.2000 ;
	    RECT 338.8000 161.6000 339.6000 169.8000 ;
	    RECT 343.2000 161.6000 344.0000 170.2000 ;
	    RECT 348.4000 161.6000 349.2000 169.8000 ;
	    RECT 352.8000 161.6000 353.6000 170.2000 ;
	    RECT 358.0000 161.6000 358.8000 169.8000 ;
	    RECT 362.4000 161.6000 363.2000 170.2000 ;
	    RECT 367.6000 161.6000 368.4000 169.8000 ;
	    RECT 372.4000 161.6000 373.2000 169.0000 ;
	    RECT 375.6000 161.6000 376.4000 170.2000 ;
	    RECT 378.8000 161.6000 379.6000 170.2000 ;
	    RECT 382.0000 161.6000 382.8000 170.2000 ;
	    RECT 385.2000 161.6000 386.0000 170.2000 ;
	    RECT 388.4000 161.6000 389.2000 170.2000 ;
	    RECT 390.0000 161.6000 390.8000 166.2000 ;
	    RECT 393.2000 161.6000 394.0000 166.2000 ;
	    RECT 396.4000 161.6000 397.2000 170.2000 ;
	    RECT 402.0000 161.6000 402.8000 166.2000 ;
	    RECT 405.2000 161.6000 406.0000 166.2000 ;
	    RECT 410.8000 161.6000 411.6000 170.0000 ;
	    RECT 421.0000 161.6000 421.8000 166.2000 ;
	    RECT 425.2000 161.6000 426.0000 170.2000 ;
	    RECT 426.8000 161.6000 427.6000 166.2000 ;
	    RECT 430.0000 161.6000 430.8000 166.2000 ;
	    RECT 433.2000 161.6000 434.0000 166.2000 ;
	    RECT 436.4000 161.6000 437.2000 165.8000 ;
	    RECT 439.6000 161.6000 440.4000 166.2000 ;
	    RECT 442.8000 161.6000 443.6000 166.2000 ;
	    RECT 447.6000 161.6000 448.4000 170.2000 ;
	    RECT 452.4000 161.6000 453.2000 170.2000 ;
	    RECT 455.6000 161.6000 456.4000 169.0000 ;
	    RECT 458.8000 161.6000 459.6000 166.2000 ;
	    RECT 462.0000 161.6000 462.8000 165.8000 ;
	    RECT 466.8000 161.6000 467.6000 169.0000 ;
	    RECT 471.6000 161.6000 472.4000 169.0000 ;
	    RECT 476.4000 161.6000 477.2000 165.8000 ;
	    RECT 479.6000 161.6000 480.4000 166.2000 ;
	    RECT 482.8000 161.6000 483.6000 169.0000 ;
	    RECT 487.6000 161.6000 488.4000 170.2000 ;
	    RECT 493.2000 161.6000 494.0000 166.2000 ;
	    RECT 496.4000 161.6000 497.2000 166.2000 ;
	    RECT 502.0000 161.6000 502.8000 170.0000 ;
	    RECT 505.2000 161.6000 506.0000 166.2000 ;
	    RECT 508.4000 161.6000 509.2000 170.2000 ;
	    RECT 512.6000 161.6000 513.4000 166.2000 ;
	    RECT 0.4000 160.4000 514.8000 161.6000 ;
	    RECT 2.8000 153.0000 3.6000 160.4000 ;
	    RECT 7.6000 153.0000 8.4000 160.4000 ;
	    RECT 12.4000 153.0000 13.2000 160.4000 ;
	    RECT 15.6000 151.8000 16.4000 160.4000 ;
	    RECT 19.8000 155.8000 20.6000 160.4000 ;
	    RECT 23.6000 151.8000 24.4000 160.4000 ;
	    RECT 29.2000 155.8000 30.0000 160.4000 ;
	    RECT 32.4000 155.8000 33.2000 160.4000 ;
	    RECT 38.0000 152.0000 38.8000 160.4000 ;
	    RECT 42.8000 152.0000 43.6000 160.4000 ;
	    RECT 48.4000 155.8000 49.2000 160.4000 ;
	    RECT 51.6000 155.8000 52.4000 160.4000 ;
	    RECT 57.2000 151.8000 58.0000 160.4000 ;
	    RECT 62.0000 152.0000 62.8000 160.4000 ;
	    RECT 67.6000 155.8000 68.4000 160.4000 ;
	    RECT 70.8000 155.8000 71.6000 160.4000 ;
	    RECT 76.4000 151.8000 77.2000 160.4000 ;
	    RECT 81.2000 153.0000 82.0000 160.4000 ;
	    RECT 84.4000 155.8000 85.2000 160.4000 ;
	    RECT 87.6000 155.8000 88.4000 160.4000 ;
	    RECT 89.8000 155.8000 90.6000 160.4000 ;
	    RECT 94.0000 151.8000 94.8000 160.4000 ;
	    RECT 95.6000 151.8000 96.4000 160.4000 ;
	    RECT 99.8000 155.8000 100.6000 160.4000 ;
	    RECT 102.6000 155.8000 103.4000 160.4000 ;
	    RECT 106.8000 151.8000 107.6000 160.4000 ;
	    RECT 116.0000 151.8000 116.8000 160.4000 ;
	    RECT 121.2000 152.2000 122.0000 160.4000 ;
	    RECT 124.4000 151.8000 125.2000 160.4000 ;
	    RECT 129.2000 151.8000 130.0000 160.4000 ;
	    RECT 134.0000 151.8000 134.8000 160.4000 ;
	    RECT 138.2000 155.8000 139.0000 160.4000 ;
	    RECT 140.4000 155.8000 141.2000 160.4000 ;
	    RECT 143.6000 155.8000 144.4000 160.4000 ;
	    RECT 145.2000 151.8000 146.0000 160.4000 ;
	    RECT 149.4000 155.8000 150.2000 160.4000 ;
	    RECT 151.6000 151.8000 152.4000 160.4000 ;
	    RECT 158.0000 151.8000 158.8000 160.4000 ;
	    RECT 159.6000 151.8000 160.4000 160.4000 ;
	    RECT 167.6000 151.8000 168.4000 160.4000 ;
	    RECT 169.2000 151.8000 170.0000 160.4000 ;
	    RECT 173.4000 155.8000 174.2000 160.4000 ;
	    RECT 175.6000 151.8000 176.4000 160.4000 ;
	    RECT 182.0000 151.8000 182.8000 160.4000 ;
	    RECT 183.6000 151.8000 184.4000 160.4000 ;
	    RECT 189.0000 155.8000 189.8000 160.4000 ;
	    RECT 193.2000 151.8000 194.0000 160.4000 ;
	    RECT 195.4000 155.8000 196.2000 160.4000 ;
	    RECT 199.6000 151.8000 200.4000 160.4000 ;
	    RECT 202.8000 151.8000 203.6000 160.4000 ;
	    RECT 208.4000 155.8000 209.2000 160.4000 ;
	    RECT 211.6000 155.8000 212.4000 160.4000 ;
	    RECT 217.2000 152.0000 218.0000 160.4000 ;
	    RECT 222.0000 153.0000 222.8000 160.4000 ;
	    RECT 225.2000 151.8000 226.0000 160.4000 ;
	    RECT 231.6000 153.0000 232.4000 160.4000 ;
	    RECT 236.4000 152.0000 237.2000 160.4000 ;
	    RECT 242.0000 155.8000 242.8000 160.4000 ;
	    RECT 245.2000 155.8000 246.0000 160.4000 ;
	    RECT 250.8000 151.8000 251.6000 160.4000 ;
	    RECT 262.0000 153.0000 262.8000 160.4000 ;
	    RECT 265.2000 151.8000 266.0000 160.4000 ;
	    RECT 269.4000 155.8000 270.2000 160.4000 ;
	    RECT 273.2000 153.0000 274.0000 160.4000 ;
	    RECT 277.0000 155.8000 277.8000 160.4000 ;
	    RECT 281.2000 151.8000 282.0000 160.4000 ;
	    RECT 284.4000 153.0000 285.2000 160.4000 ;
	    RECT 290.8000 151.8000 291.6000 160.4000 ;
	    RECT 292.4000 151.8000 293.2000 160.4000 ;
	    RECT 298.8000 151.8000 299.6000 160.4000 ;
	    RECT 301.0000 155.8000 301.8000 160.4000 ;
	    RECT 305.2000 151.8000 306.0000 160.4000 ;
	    RECT 307.4000 155.8000 308.2000 160.4000 ;
	    RECT 311.6000 151.8000 312.4000 160.4000 ;
	    RECT 313.2000 151.8000 314.0000 160.4000 ;
	    RECT 319.6000 151.8000 320.4000 160.4000 ;
	    RECT 324.4000 151.8000 325.2000 160.4000 ;
	    RECT 326.0000 151.8000 326.8000 160.4000 ;
	    RECT 332.4000 151.8000 333.2000 160.4000 ;
	    RECT 334.6000 155.8000 335.4000 160.4000 ;
	    RECT 338.8000 151.8000 339.6000 160.4000 ;
	    RECT 340.4000 151.8000 341.2000 160.4000 ;
	    RECT 345.2000 151.8000 346.0000 160.4000 ;
	    RECT 351.6000 151.8000 352.4000 160.4000 ;
	    RECT 353.8000 155.8000 354.6000 160.4000 ;
	    RECT 358.0000 151.8000 358.8000 160.4000 ;
	    RECT 359.6000 151.8000 360.4000 160.4000 ;
	    RECT 363.8000 155.8000 364.6000 160.4000 ;
	    RECT 366.0000 155.8000 366.8000 160.4000 ;
	    RECT 369.2000 155.8000 370.0000 160.4000 ;
	    RECT 371.4000 155.8000 372.2000 160.4000 ;
	    RECT 375.6000 151.8000 376.4000 160.4000 ;
	    RECT 378.8000 151.8000 379.6000 160.4000 ;
	    RECT 384.4000 155.8000 385.2000 160.4000 ;
	    RECT 387.6000 155.8000 388.4000 160.4000 ;
	    RECT 393.2000 152.0000 394.0000 160.4000 ;
	    RECT 397.0000 155.8000 397.8000 160.4000 ;
	    RECT 401.2000 151.8000 402.0000 160.4000 ;
	    RECT 410.8000 151.8000 411.6000 160.4000 ;
	    RECT 416.4000 155.8000 417.2000 160.4000 ;
	    RECT 419.6000 155.8000 420.4000 160.4000 ;
	    RECT 425.2000 152.0000 426.0000 160.4000 ;
	    RECT 430.0000 151.8000 430.8000 160.4000 ;
	    RECT 435.6000 155.8000 436.4000 160.4000 ;
	    RECT 438.8000 155.8000 439.6000 160.4000 ;
	    RECT 444.4000 152.0000 445.2000 160.4000 ;
	    RECT 447.6000 155.8000 448.4000 160.4000 ;
	    RECT 450.8000 155.8000 451.6000 160.4000 ;
	    RECT 453.0000 155.8000 453.8000 160.4000 ;
	    RECT 457.2000 151.8000 458.0000 160.4000 ;
	    RECT 460.4000 151.8000 461.2000 160.4000 ;
	    RECT 466.0000 155.8000 466.8000 160.4000 ;
	    RECT 469.2000 155.8000 470.0000 160.4000 ;
	    RECT 474.8000 152.0000 475.6000 160.4000 ;
	    RECT 478.6000 155.8000 479.4000 160.4000 ;
	    RECT 482.8000 151.8000 483.6000 160.4000 ;
	    RECT 486.0000 155.8000 486.8000 160.4000 ;
	    RECT 487.6000 155.8000 488.4000 160.4000 ;
	    RECT 490.8000 152.2000 491.6000 160.4000 ;
	    RECT 495.6000 151.8000 496.4000 160.4000 ;
	    RECT 501.2000 155.8000 502.0000 160.4000 ;
	    RECT 504.4000 155.8000 505.2000 160.4000 ;
	    RECT 510.0000 152.0000 510.8000 160.4000 ;
	    RECT 2.8000 121.6000 3.6000 129.0000 ;
	    RECT 7.6000 121.6000 8.4000 129.0000 ;
	    RECT 12.4000 121.6000 13.2000 130.2000 ;
	    RECT 18.0000 121.6000 18.8000 126.2000 ;
	    RECT 21.2000 121.6000 22.0000 126.2000 ;
	    RECT 26.8000 121.6000 27.6000 130.0000 ;
	    RECT 30.6000 121.6000 31.4000 126.2000 ;
	    RECT 34.8000 121.6000 35.6000 130.2000 ;
	    RECT 36.4000 121.6000 37.2000 130.2000 ;
	    RECT 40.6000 121.6000 41.4000 126.2000 ;
	    RECT 44.4000 121.6000 45.2000 130.2000 ;
	    RECT 50.0000 121.6000 50.8000 126.2000 ;
	    RECT 53.2000 121.6000 54.0000 126.2000 ;
	    RECT 58.8000 121.6000 59.6000 130.0000 ;
	    RECT 62.6000 121.6000 63.4000 126.2000 ;
	    RECT 66.8000 121.6000 67.6000 130.2000 ;
	    RECT 68.4000 121.6000 69.2000 130.2000 ;
	    RECT 71.6000 121.6000 72.4000 130.2000 ;
	    RECT 73.8000 121.6000 74.6000 126.2000 ;
	    RECT 78.0000 121.6000 78.8000 130.2000 ;
	    RECT 79.6000 121.6000 80.4000 130.2000 ;
	    RECT 85.0000 121.6000 85.8000 126.2000 ;
	    RECT 89.2000 121.6000 90.0000 130.2000 ;
	    RECT 91.4000 121.6000 92.2000 126.2000 ;
	    RECT 95.6000 121.6000 96.4000 130.2000 ;
	    RECT 97.2000 121.6000 98.0000 130.2000 ;
	    RECT 101.4000 121.6000 102.2000 126.2000 ;
	    RECT 111.6000 121.6000 112.4000 129.8000 ;
	    RECT 116.8000 121.6000 117.6000 130.2000 ;
	    RECT 119.6000 121.6000 120.4000 130.2000 ;
	    RECT 126.0000 121.6000 126.8000 130.2000 ;
	    RECT 128.2000 121.6000 129.0000 126.2000 ;
	    RECT 132.4000 121.6000 133.2000 130.2000 ;
	    RECT 134.0000 121.6000 134.8000 130.2000 ;
	    RECT 140.4000 121.6000 141.2000 130.2000 ;
	    RECT 142.0000 121.6000 142.8000 130.2000 ;
	    RECT 148.4000 121.6000 149.2000 130.2000 ;
	    RECT 150.0000 121.6000 150.8000 130.2000 ;
	    RECT 154.2000 121.6000 155.0000 126.2000 ;
	    RECT 158.0000 121.6000 158.8000 129.0000 ;
	    RECT 164.4000 121.6000 165.2000 130.2000 ;
	    RECT 166.0000 121.6000 166.8000 130.2000 ;
	    RECT 174.0000 121.6000 174.8000 130.2000 ;
	    RECT 178.8000 121.6000 179.6000 130.2000 ;
	    RECT 182.0000 121.6000 182.8000 129.0000 ;
	    RECT 186.8000 121.6000 187.6000 129.0000 ;
	    RECT 191.6000 121.6000 192.4000 129.0000 ;
	    RECT 196.4000 121.6000 197.2000 129.0000 ;
	    RECT 199.6000 121.6000 200.4000 130.2000 ;
	    RECT 203.8000 121.6000 204.6000 126.2000 ;
	    RECT 206.0000 121.6000 206.8000 130.2000 ;
	    RECT 210.2000 121.6000 211.0000 126.2000 ;
	    RECT 213.0000 121.6000 213.8000 126.2000 ;
	    RECT 217.2000 121.6000 218.0000 130.2000 ;
	    RECT 220.4000 121.6000 221.2000 130.2000 ;
	    RECT 226.0000 121.6000 226.8000 126.2000 ;
	    RECT 229.2000 121.6000 230.0000 126.2000 ;
	    RECT 234.8000 121.6000 235.6000 130.0000 ;
	    RECT 239.6000 121.6000 240.4000 129.0000 ;
	    RECT 244.4000 121.6000 245.2000 129.0000 ;
	    RECT 247.6000 121.6000 248.4000 130.2000 ;
	    RECT 251.8000 121.6000 252.6000 126.2000 ;
	    RECT 261.0000 121.6000 261.8000 126.2000 ;
	    RECT 265.2000 121.6000 266.0000 130.2000 ;
	    RECT 268.4000 121.6000 269.2000 129.0000 ;
	    RECT 271.6000 121.6000 272.4000 130.2000 ;
	    RECT 274.8000 121.6000 275.6000 130.2000 ;
	    RECT 278.0000 121.6000 278.8000 130.2000 ;
	    RECT 281.2000 121.6000 282.0000 129.0000 ;
	    RECT 287.6000 121.6000 288.4000 130.2000 ;
	    RECT 292.4000 121.6000 293.2000 130.2000 ;
	    RECT 294.0000 121.6000 294.8000 130.2000 ;
	    RECT 300.4000 121.6000 301.2000 130.2000 ;
	    RECT 305.2000 121.6000 306.0000 130.2000 ;
	    RECT 307.4000 121.6000 308.2000 126.2000 ;
	    RECT 311.6000 121.6000 312.4000 130.2000 ;
	    RECT 313.2000 121.6000 314.0000 130.2000 ;
	    RECT 318.0000 121.6000 318.8000 130.2000 ;
	    RECT 324.4000 121.6000 325.2000 130.2000 ;
	    RECT 326.6000 121.6000 327.4000 126.2000 ;
	    RECT 330.8000 121.6000 331.6000 130.2000 ;
	    RECT 334.0000 121.6000 334.8000 129.0000 ;
	    RECT 337.2000 121.6000 338.0000 130.2000 ;
	    RECT 343.6000 121.6000 344.4000 130.2000 ;
	    RECT 348.4000 121.6000 349.2000 130.2000 ;
	    RECT 350.6000 121.6000 351.4000 126.2000 ;
	    RECT 354.8000 121.6000 355.6000 130.2000 ;
	    RECT 357.0000 121.6000 357.8000 126.2000 ;
	    RECT 361.2000 121.6000 362.0000 130.2000 ;
	    RECT 364.4000 121.6000 365.2000 129.8000 ;
	    RECT 369.6000 121.6000 370.4000 130.2000 ;
	    RECT 374.0000 121.6000 374.8000 129.8000 ;
	    RECT 379.2000 121.6000 380.0000 130.2000 ;
	    RECT 383.6000 121.6000 384.4000 129.0000 ;
	    RECT 387.4000 121.6000 388.2000 126.2000 ;
	    RECT 391.6000 121.6000 392.4000 130.2000 ;
	    RECT 393.2000 121.6000 394.0000 130.2000 ;
	    RECT 397.4000 121.6000 398.2000 126.2000 ;
	    RECT 400.2000 121.6000 401.0000 126.2000 ;
	    RECT 404.4000 121.6000 405.2000 130.2000 ;
	    RECT 414.0000 121.6000 414.8000 130.2000 ;
	    RECT 419.6000 121.6000 420.4000 126.2000 ;
	    RECT 422.8000 121.6000 423.6000 126.2000 ;
	    RECT 428.4000 121.6000 429.2000 130.0000 ;
	    RECT 431.6000 121.6000 432.4000 126.2000 ;
	    RECT 434.8000 121.6000 435.6000 126.2000 ;
	    RECT 437.0000 121.6000 437.8000 126.2000 ;
	    RECT 441.2000 121.6000 442.0000 130.2000 ;
	    RECT 442.8000 121.6000 443.6000 130.2000 ;
	    RECT 447.0000 121.6000 447.8000 126.2000 ;
	    RECT 449.2000 121.6000 450.0000 126.2000 ;
	    RECT 452.4000 121.6000 453.2000 126.2000 ;
	    RECT 455.6000 121.6000 456.4000 130.2000 ;
	    RECT 461.2000 121.6000 462.0000 126.2000 ;
	    RECT 464.4000 121.6000 465.2000 126.2000 ;
	    RECT 470.0000 121.6000 470.8000 130.0000 ;
	    RECT 474.8000 121.6000 475.6000 130.2000 ;
	    RECT 480.4000 121.6000 481.2000 126.2000 ;
	    RECT 483.6000 121.6000 484.4000 126.2000 ;
	    RECT 489.2000 121.6000 490.0000 130.0000 ;
	    RECT 492.4000 121.6000 493.2000 126.2000 ;
	    RECT 495.6000 121.6000 496.4000 130.2000 ;
	    RECT 499.8000 121.6000 500.6000 126.2000 ;
	    RECT 502.0000 121.6000 502.8000 130.2000 ;
	    RECT 506.2000 121.6000 507.0000 126.2000 ;
	    RECT 508.4000 121.6000 509.2000 126.2000 ;
	    RECT 511.6000 121.6000 512.4000 125.8000 ;
	    RECT 0.4000 120.4000 514.8000 121.6000 ;
	    RECT 2.8000 113.0000 3.6000 120.4000 ;
	    RECT 7.6000 111.8000 8.4000 120.4000 ;
	    RECT 13.2000 115.8000 14.0000 120.4000 ;
	    RECT 16.4000 115.8000 17.2000 120.4000 ;
	    RECT 22.0000 112.0000 22.8000 120.4000 ;
	    RECT 25.2000 111.8000 26.0000 120.4000 ;
	    RECT 29.4000 115.8000 30.2000 120.4000 ;
	    RECT 34.8000 111.8000 35.6000 120.4000 ;
	    RECT 38.0000 111.8000 38.8000 120.4000 ;
	    RECT 43.6000 115.8000 44.4000 120.4000 ;
	    RECT 46.8000 115.8000 47.6000 120.4000 ;
	    RECT 52.4000 112.0000 53.2000 120.4000 ;
	    RECT 56.2000 115.8000 57.0000 120.4000 ;
	    RECT 60.4000 111.8000 61.2000 120.4000 ;
	    RECT 63.6000 112.0000 64.4000 120.4000 ;
	    RECT 69.2000 115.8000 70.0000 120.4000 ;
	    RECT 72.4000 115.8000 73.2000 120.4000 ;
	    RECT 78.0000 111.8000 78.8000 120.4000 ;
	    RECT 81.2000 115.8000 82.0000 120.4000 ;
	    RECT 84.4000 115.8000 85.2000 120.4000 ;
	    RECT 86.6000 115.8000 87.4000 120.4000 ;
	    RECT 90.8000 111.8000 91.6000 120.4000 ;
	    RECT 93.6000 111.8000 94.4000 120.4000 ;
	    RECT 98.8000 112.2000 99.6000 120.4000 ;
	    RECT 108.4000 111.8000 109.2000 120.4000 ;
	    RECT 114.8000 111.8000 115.6000 120.4000 ;
	    RECT 117.0000 115.8000 117.8000 120.4000 ;
	    RECT 121.2000 111.8000 122.0000 120.4000 ;
	    RECT 124.4000 112.2000 125.2000 120.4000 ;
	    RECT 129.6000 111.8000 130.4000 120.4000 ;
	    RECT 132.4000 111.8000 133.2000 120.4000 ;
	    RECT 136.6000 115.8000 137.4000 120.4000 ;
	    RECT 140.4000 111.8000 141.2000 120.4000 ;
	    RECT 146.0000 115.8000 146.8000 120.4000 ;
	    RECT 149.2000 115.8000 150.0000 120.4000 ;
	    RECT 154.8000 112.0000 155.6000 120.4000 ;
	    RECT 158.0000 115.8000 158.8000 120.4000 ;
	    RECT 161.2000 115.8000 162.0000 120.4000 ;
	    RECT 163.4000 115.8000 164.2000 120.4000 ;
	    RECT 167.6000 111.8000 168.4000 120.4000 ;
	    RECT 172.4000 111.8000 173.2000 120.4000 ;
	    RECT 177.2000 111.8000 178.0000 120.4000 ;
	    RECT 182.0000 111.8000 182.8000 120.4000 ;
	    RECT 183.6000 111.8000 184.4000 120.4000 ;
	    RECT 188.4000 111.8000 189.2000 120.4000 ;
	    RECT 194.8000 111.8000 195.6000 120.4000 ;
	    RECT 200.4000 115.8000 201.2000 120.4000 ;
	    RECT 203.6000 115.8000 204.4000 120.4000 ;
	    RECT 209.2000 112.0000 210.0000 120.4000 ;
	    RECT 213.0000 115.8000 213.8000 120.4000 ;
	    RECT 217.2000 111.8000 218.0000 120.4000 ;
	    RECT 218.8000 111.8000 219.6000 120.4000 ;
	    RECT 223.6000 111.8000 224.4000 120.4000 ;
	    RECT 228.4000 111.8000 229.2000 120.4000 ;
	    RECT 236.4000 111.8000 237.2000 120.4000 ;
	    RECT 238.0000 111.8000 238.8000 120.4000 ;
	    RECT 242.8000 111.8000 243.6000 120.4000 ;
	    RECT 247.0000 115.8000 247.8000 120.4000 ;
	    RECT 257.2000 112.0000 258.0000 120.4000 ;
	    RECT 262.8000 115.8000 263.6000 120.4000 ;
	    RECT 266.0000 115.8000 266.8000 120.4000 ;
	    RECT 271.6000 111.8000 272.4000 120.4000 ;
	    RECT 276.4000 113.0000 277.2000 120.4000 ;
	    RECT 280.8000 111.8000 281.6000 120.4000 ;
	    RECT 286.0000 112.2000 286.8000 120.4000 ;
	    RECT 290.8000 112.2000 291.6000 120.4000 ;
	    RECT 296.0000 111.8000 296.8000 120.4000 ;
	    RECT 298.8000 111.8000 299.6000 120.4000 ;
	    RECT 305.2000 111.8000 306.0000 120.4000 ;
	    RECT 306.8000 111.8000 307.6000 120.4000 ;
	    RECT 311.0000 115.8000 311.8000 120.4000 ;
	    RECT 316.4000 111.8000 317.2000 120.4000 ;
	    RECT 318.0000 111.8000 318.8000 120.4000 ;
	    RECT 322.2000 115.8000 323.0000 120.4000 ;
	    RECT 326.0000 113.0000 326.8000 120.4000 ;
	    RECT 330.8000 113.0000 331.6000 120.4000 ;
	    RECT 335.6000 111.8000 336.4000 120.4000 ;
	    RECT 341.2000 115.8000 342.0000 120.4000 ;
	    RECT 344.4000 115.8000 345.2000 120.4000 ;
	    RECT 350.0000 112.0000 350.8000 120.4000 ;
	    RECT 353.2000 111.8000 354.0000 120.4000 ;
	    RECT 357.4000 115.8000 358.2000 120.4000 ;
	    RECT 361.2000 112.2000 362.0000 120.4000 ;
	    RECT 366.4000 111.8000 367.2000 120.4000 ;
	    RECT 370.8000 112.2000 371.6000 120.4000 ;
	    RECT 376.0000 111.8000 376.8000 120.4000 ;
	    RECT 380.4000 111.8000 381.2000 120.4000 ;
	    RECT 386.0000 115.8000 386.8000 120.4000 ;
	    RECT 389.2000 115.8000 390.0000 120.4000 ;
	    RECT 394.8000 112.0000 395.6000 120.4000 ;
	    RECT 398.6000 115.8000 399.4000 120.4000 ;
	    RECT 402.8000 111.8000 403.6000 120.4000 ;
	    RECT 412.4000 111.8000 413.2000 120.4000 ;
	    RECT 418.0000 115.8000 418.8000 120.4000 ;
	    RECT 421.2000 115.8000 422.0000 120.4000 ;
	    RECT 426.8000 112.0000 427.6000 120.4000 ;
	    RECT 430.0000 115.8000 430.8000 120.4000 ;
	    RECT 433.2000 115.8000 434.0000 120.4000 ;
	    RECT 436.4000 111.8000 437.2000 120.4000 ;
	    RECT 442.0000 115.8000 442.8000 120.4000 ;
	    RECT 445.2000 115.8000 446.0000 120.4000 ;
	    RECT 450.8000 112.0000 451.6000 120.4000 ;
	    RECT 454.0000 115.8000 454.8000 120.4000 ;
	    RECT 457.2000 115.8000 458.0000 120.4000 ;
	    RECT 459.4000 115.8000 460.2000 120.4000 ;
	    RECT 463.6000 111.8000 464.4000 120.4000 ;
	    RECT 466.8000 111.8000 467.6000 120.4000 ;
	    RECT 470.0000 111.8000 470.8000 120.4000 ;
	    RECT 473.2000 111.8000 474.0000 120.4000 ;
	    RECT 478.8000 115.8000 479.6000 120.4000 ;
	    RECT 482.0000 115.8000 482.8000 120.4000 ;
	    RECT 487.6000 112.0000 488.4000 120.4000 ;
	    RECT 490.8000 115.8000 491.6000 120.4000 ;
	    RECT 494.0000 111.8000 494.8000 120.4000 ;
	    RECT 498.2000 115.8000 499.0000 120.4000 ;
	    RECT 500.4000 115.8000 501.2000 120.4000 ;
	    RECT 503.6000 116.2000 504.4000 120.4000 ;
	    RECT 506.8000 115.8000 507.6000 120.4000 ;
	    RECT 510.0000 116.2000 510.8000 120.4000 ;
	    RECT 2.8000 81.6000 3.6000 89.0000 ;
	    RECT 7.6000 81.6000 8.4000 89.0000 ;
	    RECT 11.4000 81.6000 12.2000 86.2000 ;
	    RECT 15.6000 81.6000 16.4000 90.2000 ;
	    RECT 17.8000 81.6000 18.6000 86.2000 ;
	    RECT 22.0000 81.6000 22.8000 90.2000 ;
	    RECT 23.6000 81.6000 24.4000 90.2000 ;
	    RECT 27.8000 81.6000 28.6000 86.2000 ;
	    RECT 31.6000 81.6000 32.4000 90.2000 ;
	    RECT 37.2000 81.6000 38.0000 86.2000 ;
	    RECT 40.4000 81.6000 41.2000 86.2000 ;
	    RECT 46.0000 81.6000 46.8000 90.0000 ;
	    RECT 49.8000 81.6000 50.6000 86.2000 ;
	    RECT 54.0000 81.6000 54.8000 90.2000 ;
	    RECT 55.6000 81.6000 56.4000 90.2000 ;
	    RECT 60.4000 81.6000 61.2000 90.2000 ;
	    RECT 65.2000 81.6000 66.0000 90.2000 ;
	    RECT 70.0000 81.6000 70.8000 90.2000 ;
	    RECT 75.4000 81.6000 76.2000 86.2000 ;
	    RECT 79.6000 81.6000 80.4000 90.2000 ;
	    RECT 82.8000 81.6000 83.6000 90.0000 ;
	    RECT 88.4000 81.6000 89.2000 86.2000 ;
	    RECT 91.6000 81.6000 92.4000 86.2000 ;
	    RECT 97.2000 81.6000 98.0000 90.2000 ;
	    RECT 100.4000 81.6000 101.2000 90.2000 ;
	    RECT 104.6000 81.6000 105.4000 86.2000 ;
	    RECT 113.8000 81.6000 114.6000 86.2000 ;
	    RECT 118.0000 81.6000 118.8000 90.2000 ;
	    RECT 120.2000 81.6000 121.0000 86.2000 ;
	    RECT 124.4000 81.6000 125.2000 90.2000 ;
	    RECT 126.6000 81.6000 127.4000 86.2000 ;
	    RECT 130.8000 81.6000 131.6000 90.2000 ;
	    RECT 132.4000 81.6000 133.2000 90.2000 ;
	    RECT 137.2000 81.6000 138.0000 90.2000 ;
	    RECT 143.6000 81.6000 144.4000 90.2000 ;
	    RECT 145.8000 81.6000 146.6000 86.2000 ;
	    RECT 150.0000 81.6000 150.8000 90.2000 ;
	    RECT 151.6000 81.6000 152.4000 90.2000 ;
	    RECT 158.0000 81.6000 158.8000 90.2000 ;
	    RECT 160.2000 81.6000 161.0000 86.2000 ;
	    RECT 164.4000 81.6000 165.2000 90.2000 ;
	    RECT 166.0000 81.6000 166.8000 90.2000 ;
	    RECT 171.4000 81.6000 172.2000 86.2000 ;
	    RECT 175.6000 81.6000 176.4000 90.2000 ;
	    RECT 177.2000 81.6000 178.0000 90.2000 ;
	    RECT 183.6000 81.6000 184.4000 90.2000 ;
	    RECT 185.2000 81.6000 186.0000 90.2000 ;
	    RECT 191.6000 81.6000 192.4000 90.2000 ;
	    RECT 193.8000 81.6000 194.6000 86.2000 ;
	    RECT 198.0000 81.6000 198.8000 90.2000 ;
	    RECT 200.2000 81.6000 201.0000 86.2000 ;
	    RECT 204.4000 81.6000 205.2000 90.2000 ;
	    RECT 207.6000 81.6000 208.4000 89.8000 ;
	    RECT 212.8000 81.6000 213.6000 90.2000 ;
	    RECT 216.8000 81.6000 217.6000 90.2000 ;
	    RECT 222.0000 81.6000 222.8000 89.8000 ;
	    RECT 225.2000 81.6000 226.0000 90.2000 ;
	    RECT 230.0000 81.6000 230.8000 86.2000 ;
	    RECT 233.2000 81.6000 234.0000 86.2000 ;
	    RECT 235.4000 81.6000 236.2000 86.2000 ;
	    RECT 239.6000 81.6000 240.4000 90.2000 ;
	    RECT 242.8000 81.6000 243.6000 90.2000 ;
	    RECT 248.4000 81.6000 249.2000 86.2000 ;
	    RECT 251.6000 81.6000 252.4000 86.2000 ;
	    RECT 257.2000 81.6000 258.0000 90.0000 ;
	    RECT 266.8000 81.6000 267.6000 86.2000 ;
	    RECT 270.0000 81.6000 270.8000 86.2000 ;
	    RECT 273.2000 81.6000 274.0000 89.0000 ;
	    RECT 278.0000 81.6000 278.8000 89.0000 ;
	    RECT 281.2000 81.6000 282.0000 90.2000 ;
	    RECT 287.6000 81.6000 288.4000 90.2000 ;
	    RECT 290.8000 81.6000 291.6000 89.0000 ;
	    RECT 294.0000 81.6000 294.8000 90.2000 ;
	    RECT 298.2000 81.6000 299.0000 86.2000 ;
	    RECT 300.4000 81.6000 301.2000 90.2000 ;
	    RECT 306.8000 81.6000 307.6000 90.2000 ;
	    RECT 309.0000 81.6000 309.8000 86.2000 ;
	    RECT 313.2000 81.6000 314.0000 90.2000 ;
	    RECT 318.0000 81.6000 318.8000 90.2000 ;
	    RECT 319.6000 81.6000 320.4000 90.2000 ;
	    RECT 326.0000 81.6000 326.8000 90.2000 ;
	    RECT 329.2000 81.6000 330.0000 89.0000 ;
	    RECT 334.0000 81.6000 334.8000 89.8000 ;
	    RECT 339.2000 81.6000 340.0000 90.2000 ;
	    RECT 343.2000 81.6000 344.0000 90.2000 ;
	    RECT 348.4000 81.6000 349.2000 89.8000 ;
	    RECT 354.8000 81.6000 355.6000 90.2000 ;
	    RECT 356.4000 81.6000 357.2000 90.2000 ;
	    RECT 362.8000 81.6000 363.6000 90.2000 ;
	    RECT 365.0000 81.6000 365.8000 86.2000 ;
	    RECT 369.2000 81.6000 370.0000 90.2000 ;
	    RECT 372.4000 81.6000 373.2000 89.0000 ;
	    RECT 375.6000 81.6000 376.4000 90.2000 ;
	    RECT 379.8000 81.6000 380.6000 86.2000 ;
	    RECT 382.6000 81.6000 383.4000 86.2000 ;
	    RECT 386.8000 81.6000 387.6000 90.2000 ;
	    RECT 390.0000 81.6000 390.8000 90.2000 ;
	    RECT 395.6000 81.6000 396.4000 86.2000 ;
	    RECT 398.8000 81.6000 399.6000 86.2000 ;
	    RECT 404.4000 81.6000 405.2000 90.0000 ;
	    RECT 415.6000 81.6000 416.4000 90.2000 ;
	    RECT 421.2000 81.6000 422.0000 86.2000 ;
	    RECT 424.4000 81.6000 425.2000 86.2000 ;
	    RECT 430.0000 81.6000 430.8000 90.0000 ;
	    RECT 433.8000 81.6000 434.6000 86.2000 ;
	    RECT 438.0000 81.6000 438.8000 90.2000 ;
	    RECT 441.2000 81.6000 442.0000 90.2000 ;
	    RECT 446.8000 81.6000 447.6000 86.2000 ;
	    RECT 450.0000 81.6000 450.8000 86.2000 ;
	    RECT 455.6000 81.6000 456.4000 90.0000 ;
	    RECT 458.8000 81.6000 459.6000 86.2000 ;
	    RECT 462.0000 81.6000 462.8000 90.2000 ;
	    RECT 466.2000 81.6000 467.0000 86.2000 ;
	    RECT 470.0000 81.6000 470.8000 90.2000 ;
	    RECT 475.6000 81.6000 476.4000 86.2000 ;
	    RECT 478.8000 81.6000 479.6000 86.2000 ;
	    RECT 484.4000 81.6000 485.2000 90.0000 ;
	    RECT 488.2000 81.6000 489.0000 86.2000 ;
	    RECT 492.4000 81.6000 493.2000 90.2000 ;
	    RECT 494.0000 81.6000 494.8000 86.2000 ;
	    RECT 497.2000 81.6000 498.0000 86.2000 ;
	    RECT 500.4000 81.6000 501.2000 85.8000 ;
	    RECT 505.2000 81.6000 506.0000 85.8000 ;
	    RECT 508.4000 81.6000 509.2000 86.2000 ;
	    RECT 0.4000 80.4000 514.8000 81.6000 ;
	    RECT 2.8000 73.0000 3.6000 80.4000 ;
	    RECT 7.6000 73.0000 8.4000 80.4000 ;
	    RECT 12.4000 73.0000 13.2000 80.4000 ;
	    RECT 17.2000 71.8000 18.0000 80.4000 ;
	    RECT 22.8000 75.8000 23.6000 80.4000 ;
	    RECT 26.0000 75.8000 26.8000 80.4000 ;
	    RECT 31.6000 72.0000 32.4000 80.4000 ;
	    RECT 36.4000 73.0000 37.2000 80.4000 ;
	    RECT 40.2000 75.8000 41.0000 80.4000 ;
	    RECT 44.4000 71.8000 45.2000 80.4000 ;
	    RECT 47.6000 73.0000 48.4000 80.4000 ;
	    RECT 51.4000 75.8000 52.2000 80.4000 ;
	    RECT 55.6000 71.8000 56.4000 80.4000 ;
	    RECT 57.2000 71.8000 58.0000 80.4000 ;
	    RECT 60.4000 71.8000 61.2000 80.4000 ;
	    RECT 63.6000 71.8000 64.4000 80.4000 ;
	    RECT 66.8000 71.8000 67.6000 80.4000 ;
	    RECT 70.0000 71.8000 70.8000 80.4000 ;
	    RECT 72.2000 75.8000 73.0000 80.4000 ;
	    RECT 76.4000 71.8000 77.2000 80.4000 ;
	    RECT 79.6000 73.0000 80.4000 80.4000 ;
	    RECT 84.4000 72.0000 85.2000 80.4000 ;
	    RECT 90.0000 75.8000 90.8000 80.4000 ;
	    RECT 93.2000 75.8000 94.0000 80.4000 ;
	    RECT 98.8000 71.8000 99.6000 80.4000 ;
	    RECT 102.0000 71.8000 102.8000 80.4000 ;
	    RECT 106.2000 75.8000 107.0000 80.4000 ;
	    RECT 114.8000 75.8000 115.6000 80.4000 ;
	    RECT 118.0000 75.8000 118.8000 80.4000 ;
	    RECT 121.2000 73.0000 122.0000 80.4000 ;
	    RECT 126.0000 72.2000 126.8000 80.4000 ;
	    RECT 131.2000 71.8000 132.0000 80.4000 ;
	    RECT 135.6000 72.2000 136.4000 80.4000 ;
	    RECT 140.8000 71.8000 141.6000 80.4000 ;
	    RECT 143.6000 75.8000 144.4000 80.4000 ;
	    RECT 146.8000 75.8000 147.6000 80.4000 ;
	    RECT 149.0000 75.8000 149.8000 80.4000 ;
	    RECT 153.2000 71.8000 154.0000 80.4000 ;
	    RECT 156.4000 73.0000 157.2000 80.4000 ;
	    RECT 160.2000 75.8000 161.0000 80.4000 ;
	    RECT 164.4000 71.8000 165.2000 80.4000 ;
	    RECT 166.6000 75.8000 167.4000 80.4000 ;
	    RECT 170.8000 71.8000 171.6000 80.4000 ;
	    RECT 172.4000 71.8000 173.2000 80.4000 ;
	    RECT 176.6000 75.8000 177.4000 80.4000 ;
	    RECT 179.4000 75.8000 180.2000 80.4000 ;
	    RECT 183.6000 71.8000 184.4000 80.4000 ;
	    RECT 186.8000 71.8000 187.6000 80.4000 ;
	    RECT 192.4000 75.8000 193.2000 80.4000 ;
	    RECT 195.6000 75.8000 196.4000 80.4000 ;
	    RECT 201.2000 72.0000 202.0000 80.4000 ;
	    RECT 205.0000 75.8000 205.8000 80.4000 ;
	    RECT 209.2000 71.8000 210.0000 80.4000 ;
	    RECT 212.4000 73.0000 213.2000 80.4000 ;
	    RECT 215.6000 71.8000 216.4000 80.4000 ;
	    RECT 222.0000 71.8000 222.8000 80.4000 ;
	    RECT 224.2000 75.8000 225.0000 80.4000 ;
	    RECT 228.4000 71.8000 229.2000 80.4000 ;
	    RECT 230.0000 71.8000 230.8000 80.4000 ;
	    RECT 234.8000 71.8000 235.6000 80.4000 ;
	    RECT 241.2000 71.8000 242.0000 80.4000 ;
	    RECT 242.8000 71.8000 243.6000 80.4000 ;
	    RECT 247.0000 75.8000 247.8000 80.4000 ;
	    RECT 249.8000 75.8000 250.6000 80.4000 ;
	    RECT 254.0000 71.8000 254.8000 80.4000 ;
	    RECT 265.2000 71.8000 266.0000 80.4000 ;
	    RECT 267.4000 75.8000 268.2000 80.4000 ;
	    RECT 271.6000 71.8000 272.4000 80.4000 ;
	    RECT 273.2000 71.8000 274.0000 80.4000 ;
	    RECT 279.6000 71.8000 280.4000 80.4000 ;
	    RECT 281.2000 71.8000 282.0000 80.4000 ;
	    RECT 287.6000 72.0000 288.4000 80.4000 ;
	    RECT 293.2000 75.8000 294.0000 80.4000 ;
	    RECT 296.4000 75.8000 297.2000 80.4000 ;
	    RECT 302.0000 71.8000 302.8000 80.4000 ;
	    RECT 306.4000 71.8000 307.2000 80.4000 ;
	    RECT 311.6000 72.2000 312.4000 80.4000 ;
	    RECT 316.0000 71.8000 316.8000 80.4000 ;
	    RECT 321.2000 72.2000 322.0000 80.4000 ;
	    RECT 324.4000 71.8000 325.2000 80.4000 ;
	    RECT 328.6000 75.8000 329.4000 80.4000 ;
	    RECT 330.8000 75.8000 331.6000 80.4000 ;
	    RECT 334.0000 75.8000 334.8000 80.4000 ;
	    RECT 337.2000 71.8000 338.0000 80.4000 ;
	    RECT 342.8000 75.8000 343.6000 80.4000 ;
	    RECT 346.0000 75.8000 346.8000 80.4000 ;
	    RECT 351.6000 72.0000 352.4000 80.4000 ;
	    RECT 356.4000 73.0000 357.2000 80.4000 ;
	    RECT 359.6000 75.8000 360.4000 80.4000 ;
	    RECT 362.8000 75.8000 363.6000 80.4000 ;
	    RECT 366.0000 71.8000 366.8000 80.4000 ;
	    RECT 371.6000 75.8000 372.4000 80.4000 ;
	    RECT 374.8000 75.8000 375.6000 80.4000 ;
	    RECT 380.4000 72.0000 381.2000 80.4000 ;
	    RECT 384.2000 75.8000 385.0000 80.4000 ;
	    RECT 388.4000 71.8000 389.2000 80.4000 ;
	    RECT 391.6000 73.0000 392.4000 80.4000 ;
	    RECT 396.4000 71.8000 397.2000 80.4000 ;
	    RECT 402.0000 75.8000 402.8000 80.4000 ;
	    RECT 405.2000 75.8000 406.0000 80.4000 ;
	    RECT 410.8000 72.0000 411.6000 80.4000 ;
	    RECT 420.4000 75.8000 421.2000 80.4000 ;
	    RECT 423.6000 75.8000 424.4000 80.4000 ;
	    RECT 425.8000 75.8000 426.6000 80.4000 ;
	    RECT 430.0000 71.8000 430.8000 80.4000 ;
	    RECT 431.6000 71.8000 432.4000 80.4000 ;
	    RECT 434.8000 71.8000 435.6000 80.4000 ;
	    RECT 438.0000 71.8000 438.8000 80.4000 ;
	    RECT 441.2000 71.8000 442.0000 80.4000 ;
	    RECT 444.4000 71.8000 445.2000 80.4000 ;
	    RECT 446.0000 75.8000 446.8000 80.4000 ;
	    RECT 449.2000 71.8000 450.0000 80.4000 ;
	    RECT 453.4000 75.8000 454.2000 80.4000 ;
	    RECT 457.2000 71.8000 458.0000 80.4000 ;
	    RECT 462.8000 75.8000 463.6000 80.4000 ;
	    RECT 466.0000 75.8000 466.8000 80.4000 ;
	    RECT 471.6000 72.0000 472.4000 80.4000 ;
	    RECT 474.8000 75.8000 475.6000 80.4000 ;
	    RECT 478.0000 71.8000 478.8000 80.4000 ;
	    RECT 482.2000 75.8000 483.0000 80.4000 ;
	    RECT 486.0000 76.2000 486.8000 80.4000 ;
	    RECT 489.2000 75.8000 490.0000 80.4000 ;
	    RECT 490.8000 75.8000 491.6000 80.4000 ;
	    RECT 494.0000 71.8000 494.8000 80.4000 ;
	    RECT 498.2000 75.8000 499.0000 80.4000 ;
	    RECT 500.4000 71.8000 501.2000 80.4000 ;
	    RECT 503.6000 71.8000 504.4000 80.4000 ;
	    RECT 506.8000 71.8000 507.6000 80.4000 ;
	    RECT 510.0000 71.8000 510.8000 80.4000 ;
	    RECT 513.2000 71.8000 514.0000 80.4000 ;
	    RECT 2.8000 41.6000 3.6000 49.0000 ;
	    RECT 6.0000 41.6000 6.8000 50.2000 ;
	    RECT 9.2000 41.6000 10.0000 50.2000 ;
	    RECT 12.4000 41.6000 13.2000 50.2000 ;
	    RECT 15.6000 41.6000 16.4000 50.2000 ;
	    RECT 18.8000 41.6000 19.6000 50.2000 ;
	    RECT 22.0000 41.6000 22.8000 50.2000 ;
	    RECT 27.6000 41.6000 28.4000 46.2000 ;
	    RECT 30.8000 41.6000 31.6000 46.2000 ;
	    RECT 36.4000 41.6000 37.2000 50.0000 ;
	    RECT 40.2000 41.6000 41.0000 46.2000 ;
	    RECT 44.4000 41.6000 45.2000 50.2000 ;
	    RECT 46.6000 41.6000 47.4000 46.2000 ;
	    RECT 50.8000 41.6000 51.6000 50.2000 ;
	    RECT 53.0000 41.6000 53.8000 46.2000 ;
	    RECT 57.2000 41.6000 58.0000 50.2000 ;
	    RECT 59.4000 41.6000 60.2000 46.2000 ;
	    RECT 63.6000 41.6000 64.4000 50.2000 ;
	    RECT 66.8000 41.6000 67.6000 50.2000 ;
	    RECT 72.4000 41.6000 73.2000 46.2000 ;
	    RECT 75.6000 41.6000 76.4000 46.2000 ;
	    RECT 81.2000 41.6000 82.0000 50.0000 ;
	    RECT 86.0000 41.6000 86.8000 49.0000 ;
	    RECT 89.8000 41.6000 90.6000 46.2000 ;
	    RECT 94.0000 41.6000 94.8000 50.2000 ;
	    RECT 96.2000 41.6000 97.0000 46.2000 ;
	    RECT 100.4000 41.6000 101.2000 50.2000 ;
	    RECT 103.6000 41.6000 104.4000 49.0000 ;
	    RECT 113.8000 41.6000 114.6000 46.2000 ;
	    RECT 118.0000 41.6000 118.8000 50.2000 ;
	    RECT 121.2000 41.6000 122.0000 49.0000 ;
	    RECT 126.0000 41.6000 126.8000 49.0000 ;
	    RECT 129.8000 41.6000 130.6000 46.2000 ;
	    RECT 134.0000 41.6000 134.8000 50.2000 ;
	    RECT 137.2000 41.6000 138.0000 50.2000 ;
	    RECT 142.8000 41.6000 143.6000 46.2000 ;
	    RECT 146.0000 41.6000 146.8000 46.2000 ;
	    RECT 151.6000 41.6000 152.4000 50.0000 ;
	    RECT 155.4000 41.6000 156.2000 46.2000 ;
	    RECT 159.6000 41.6000 160.4000 50.2000 ;
	    RECT 161.8000 41.6000 162.6000 46.2000 ;
	    RECT 166.0000 41.6000 166.8000 50.2000 ;
	    RECT 168.2000 41.6000 169.0000 46.2000 ;
	    RECT 172.4000 41.6000 173.2000 50.2000 ;
	    RECT 174.6000 41.6000 175.4000 46.2000 ;
	    RECT 178.8000 41.6000 179.6000 50.2000 ;
	    RECT 181.0000 41.6000 181.8000 46.2000 ;
	    RECT 185.2000 41.6000 186.0000 50.2000 ;
	    RECT 186.8000 41.6000 187.6000 50.2000 ;
	    RECT 191.0000 41.6000 191.8000 46.2000 ;
	    RECT 193.8000 41.6000 194.6000 46.2000 ;
	    RECT 198.0000 41.6000 198.8000 50.2000 ;
	    RECT 200.2000 41.6000 201.0000 46.2000 ;
	    RECT 204.4000 41.6000 205.2000 50.2000 ;
	    RECT 206.6000 41.6000 207.4000 46.2000 ;
	    RECT 210.8000 41.6000 211.6000 50.2000 ;
	    RECT 213.0000 41.6000 213.8000 46.2000 ;
	    RECT 217.2000 41.6000 218.0000 50.2000 ;
	    RECT 219.4000 41.6000 220.2000 46.2000 ;
	    RECT 223.6000 41.6000 224.4000 50.2000 ;
	    RECT 225.2000 41.6000 226.0000 50.2000 ;
	    RECT 231.6000 41.6000 232.4000 50.2000 ;
	    RECT 233.8000 41.6000 234.6000 46.2000 ;
	    RECT 238.0000 41.6000 238.8000 50.2000 ;
	    RECT 239.6000 41.6000 240.4000 50.2000 ;
	    RECT 246.0000 41.6000 246.8000 49.0000 ;
	    RECT 249.2000 41.6000 250.0000 46.2000 ;
	    RECT 252.4000 41.6000 253.2000 46.2000 ;
	    RECT 260.4000 41.6000 261.2000 46.2000 ;
	    RECT 263.6000 41.6000 264.4000 46.2000 ;
	    RECT 265.2000 41.6000 266.0000 50.2000 ;
	    RECT 271.6000 41.6000 272.4000 50.2000 ;
	    RECT 273.8000 41.6000 274.6000 46.2000 ;
	    RECT 278.0000 41.6000 278.8000 50.2000 ;
	    RECT 280.2000 41.6000 281.0000 46.2000 ;
	    RECT 284.4000 41.6000 285.2000 50.2000 ;
	    RECT 289.2000 41.6000 290.0000 50.2000 ;
	    RECT 290.8000 41.6000 291.6000 50.2000 ;
	    RECT 297.2000 41.6000 298.0000 50.2000 ;
	    RECT 299.4000 41.6000 300.2000 46.2000 ;
	    RECT 303.6000 41.6000 304.4000 50.2000 ;
	    RECT 308.4000 41.6000 309.2000 50.2000 ;
	    RECT 310.0000 41.6000 310.8000 50.2000 ;
	    RECT 314.2000 41.6000 315.0000 46.2000 ;
	    RECT 316.4000 41.6000 317.2000 50.2000 ;
	    RECT 322.8000 41.6000 323.6000 50.2000 ;
	    RECT 324.4000 41.6000 325.2000 50.2000 ;
	    RECT 332.4000 41.6000 333.2000 50.2000 ;
	    RECT 335.6000 41.6000 336.4000 49.8000 ;
	    RECT 340.8000 41.6000 341.6000 50.2000 ;
	    RECT 344.8000 41.6000 345.6000 50.2000 ;
	    RECT 350.0000 41.6000 350.8000 49.8000 ;
	    RECT 353.8000 41.6000 354.6000 46.2000 ;
	    RECT 358.0000 41.6000 358.8000 50.2000 ;
	    RECT 359.6000 41.6000 360.4000 50.2000 ;
	    RECT 363.8000 41.6000 364.6000 46.2000 ;
	    RECT 367.6000 41.6000 368.4000 50.2000 ;
	    RECT 373.2000 41.6000 374.0000 46.2000 ;
	    RECT 376.4000 41.6000 377.2000 46.2000 ;
	    RECT 382.0000 41.6000 382.8000 50.0000 ;
	    RECT 385.8000 41.6000 386.6000 46.2000 ;
	    RECT 390.0000 41.6000 390.8000 50.2000 ;
	    RECT 391.6000 41.6000 392.4000 46.2000 ;
	    RECT 394.8000 41.6000 395.6000 46.2000 ;
	    RECT 396.4000 41.6000 397.2000 50.2000 ;
	    RECT 400.6000 41.6000 401.4000 46.2000 ;
	    RECT 410.8000 41.6000 411.6000 50.2000 ;
	    RECT 416.4000 41.6000 417.2000 46.2000 ;
	    RECT 419.6000 41.6000 420.4000 46.2000 ;
	    RECT 425.2000 41.6000 426.0000 50.0000 ;
	    RECT 428.4000 41.6000 429.2000 46.2000 ;
	    RECT 431.6000 41.6000 432.4000 46.2000 ;
	    RECT 433.8000 41.6000 434.6000 46.2000 ;
	    RECT 438.0000 41.6000 438.8000 50.2000 ;
	    RECT 441.2000 41.6000 442.0000 49.0000 ;
	    RECT 446.0000 41.6000 446.8000 50.2000 ;
	    RECT 451.6000 41.6000 452.4000 46.2000 ;
	    RECT 454.8000 41.6000 455.6000 46.2000 ;
	    RECT 460.4000 41.6000 461.2000 50.0000 ;
	    RECT 465.2000 41.6000 466.0000 50.2000 ;
	    RECT 468.4000 41.6000 469.2000 45.8000 ;
	    RECT 471.6000 41.6000 472.4000 46.2000 ;
	    RECT 474.8000 41.6000 475.6000 50.2000 ;
	    RECT 476.4000 41.6000 477.2000 46.2000 ;
	    RECT 479.6000 41.6000 480.4000 45.8000 ;
	    RECT 484.4000 41.6000 485.2000 50.2000 ;
	    RECT 487.6000 41.6000 488.4000 45.8000 ;
	    RECT 490.8000 41.6000 491.6000 46.2000 ;
	    RECT 494.0000 41.6000 494.8000 50.2000 ;
	    RECT 499.6000 41.6000 500.4000 46.2000 ;
	    RECT 502.8000 41.6000 503.6000 46.2000 ;
	    RECT 508.4000 41.6000 509.2000 50.0000 ;
	    RECT 0.4000 40.4000 514.8000 41.6000 ;
	    RECT 2.8000 31.8000 3.6000 40.4000 ;
	    RECT 8.4000 35.8000 9.2000 40.4000 ;
	    RECT 11.6000 35.8000 12.4000 40.4000 ;
	    RECT 17.2000 32.0000 18.0000 40.4000 ;
	    RECT 22.0000 32.0000 22.8000 40.4000 ;
	    RECT 27.6000 35.8000 28.4000 40.4000 ;
	    RECT 30.8000 35.8000 31.6000 40.4000 ;
	    RECT 36.4000 31.8000 37.2000 40.4000 ;
	    RECT 40.2000 35.8000 41.0000 40.4000 ;
	    RECT 44.4000 31.8000 45.2000 40.4000 ;
	    RECT 46.6000 35.8000 47.4000 40.4000 ;
	    RECT 50.8000 31.8000 51.6000 40.4000 ;
	    RECT 52.4000 31.8000 53.2000 40.4000 ;
	    RECT 56.6000 35.8000 57.4000 40.4000 ;
	    RECT 59.4000 35.8000 60.2000 40.4000 ;
	    RECT 63.6000 31.8000 64.4000 40.4000 ;
	    RECT 66.8000 33.0000 67.6000 40.4000 ;
	    RECT 71.6000 31.8000 72.4000 40.4000 ;
	    RECT 77.2000 35.8000 78.0000 40.4000 ;
	    RECT 80.4000 35.8000 81.2000 40.4000 ;
	    RECT 86.0000 32.0000 86.8000 40.4000 ;
	    RECT 89.8000 35.8000 90.6000 40.4000 ;
	    RECT 94.0000 31.8000 94.8000 40.4000 ;
	    RECT 96.2000 35.8000 97.0000 40.4000 ;
	    RECT 100.4000 31.8000 101.2000 40.4000 ;
	    RECT 103.6000 33.0000 104.4000 40.4000 ;
	    RECT 114.8000 31.8000 115.6000 40.4000 ;
	    RECT 120.4000 35.8000 121.2000 40.4000 ;
	    RECT 123.6000 35.8000 124.4000 40.4000 ;
	    RECT 129.2000 32.0000 130.0000 40.4000 ;
	    RECT 132.4000 31.8000 133.2000 40.4000 ;
	    RECT 136.6000 35.8000 137.4000 40.4000 ;
	    RECT 140.4000 31.8000 141.2000 40.4000 ;
	    RECT 146.0000 35.8000 146.8000 40.4000 ;
	    RECT 149.2000 35.8000 150.0000 40.4000 ;
	    RECT 154.8000 32.0000 155.6000 40.4000 ;
	    RECT 158.6000 35.8000 159.4000 40.4000 ;
	    RECT 162.8000 31.8000 163.6000 40.4000 ;
	    RECT 164.4000 31.8000 165.2000 40.4000 ;
	    RECT 168.6000 35.8000 169.4000 40.4000 ;
	    RECT 172.4000 32.0000 173.2000 40.4000 ;
	    RECT 178.0000 35.8000 178.8000 40.4000 ;
	    RECT 181.2000 35.8000 182.0000 40.4000 ;
	    RECT 186.8000 31.8000 187.6000 40.4000 ;
	    RECT 191.2000 31.8000 192.0000 40.4000 ;
	    RECT 196.4000 32.2000 197.2000 40.4000 ;
	    RECT 200.8000 31.8000 201.6000 40.4000 ;
	    RECT 206.0000 32.2000 206.8000 40.4000 ;
	    RECT 210.8000 33.0000 211.6000 40.4000 ;
	    RECT 214.0000 31.8000 214.8000 40.4000 ;
	    RECT 220.4000 31.8000 221.2000 40.4000 ;
	    RECT 222.6000 35.8000 223.4000 40.4000 ;
	    RECT 226.8000 31.8000 227.6000 40.4000 ;
	    RECT 229.6000 31.8000 230.4000 40.4000 ;
	    RECT 234.8000 32.2000 235.6000 40.4000 ;
	    RECT 238.0000 31.8000 238.8000 40.4000 ;
	    RECT 244.0000 31.8000 244.8000 40.4000 ;
	    RECT 249.2000 32.2000 250.0000 40.4000 ;
	    RECT 258.8000 31.8000 259.6000 40.4000 ;
	    RECT 265.2000 31.8000 266.0000 40.4000 ;
	    RECT 270.0000 31.8000 270.8000 40.4000 ;
	    RECT 272.2000 35.8000 273.0000 40.4000 ;
	    RECT 276.4000 31.8000 277.2000 40.4000 ;
	    RECT 279.6000 31.8000 280.4000 40.4000 ;
	    RECT 285.2000 35.8000 286.0000 40.4000 ;
	    RECT 288.4000 35.8000 289.2000 40.4000 ;
	    RECT 294.0000 32.0000 294.8000 40.4000 ;
	    RECT 297.2000 31.8000 298.0000 40.4000 ;
	    RECT 301.4000 35.8000 302.2000 40.4000 ;
	    RECT 304.2000 35.8000 305.0000 40.4000 ;
	    RECT 308.4000 31.8000 309.2000 40.4000 ;
	    RECT 311.2000 31.8000 312.0000 40.4000 ;
	    RECT 316.4000 32.2000 317.2000 40.4000 ;
	    RECT 319.6000 31.8000 320.4000 40.4000 ;
	    RECT 323.8000 35.8000 324.6000 40.4000 ;
	    RECT 326.0000 31.8000 326.8000 40.4000 ;
	    RECT 332.4000 31.8000 333.2000 40.4000 ;
	    RECT 335.6000 32.2000 336.4000 40.4000 ;
	    RECT 340.8000 31.8000 341.6000 40.4000 ;
	    RECT 345.2000 31.8000 346.0000 40.4000 ;
	    RECT 350.8000 35.8000 351.6000 40.4000 ;
	    RECT 354.0000 35.8000 354.8000 40.4000 ;
	    RECT 359.6000 32.0000 360.4000 40.4000 ;
	    RECT 363.4000 35.8000 364.2000 40.4000 ;
	    RECT 367.6000 31.8000 368.4000 40.4000 ;
	    RECT 369.2000 31.8000 370.0000 40.4000 ;
	    RECT 373.4000 35.8000 374.2000 40.4000 ;
	    RECT 376.2000 35.8000 377.0000 40.4000 ;
	    RECT 380.4000 31.8000 381.2000 40.4000 ;
	    RECT 383.6000 31.8000 384.4000 40.4000 ;
	    RECT 389.2000 35.8000 390.0000 40.4000 ;
	    RECT 392.4000 35.8000 393.2000 40.4000 ;
	    RECT 398.0000 32.0000 398.8000 40.4000 ;
	    RECT 401.2000 35.8000 402.0000 40.4000 ;
	    RECT 404.4000 35.8000 405.2000 40.4000 ;
	    RECT 413.0000 35.8000 413.8000 40.4000 ;
	    RECT 417.2000 31.8000 418.0000 40.4000 ;
	    RECT 420.4000 31.8000 421.2000 40.4000 ;
	    RECT 426.0000 35.8000 426.8000 40.4000 ;
	    RECT 429.2000 35.8000 430.0000 40.4000 ;
	    RECT 434.8000 32.0000 435.6000 40.4000 ;
	    RECT 439.6000 31.8000 440.4000 40.4000 ;
	    RECT 445.2000 35.8000 446.0000 40.4000 ;
	    RECT 448.4000 35.8000 449.2000 40.4000 ;
	    RECT 454.0000 32.0000 454.8000 40.4000 ;
	    RECT 457.2000 35.8000 458.0000 40.4000 ;
	    RECT 460.4000 35.8000 461.2000 40.4000 ;
	    RECT 462.0000 35.8000 462.8000 40.4000 ;
	    RECT 465.2000 31.8000 466.0000 40.4000 ;
	    RECT 469.4000 35.8000 470.2000 40.4000 ;
	    RECT 471.6000 35.8000 472.4000 40.4000 ;
	    RECT 474.8000 31.8000 475.6000 40.4000 ;
	    RECT 479.0000 35.8000 479.8000 40.4000 ;
	    RECT 481.2000 35.8000 482.0000 40.4000 ;
	    RECT 484.4000 31.8000 485.2000 40.4000 ;
	    RECT 488.6000 35.8000 489.4000 40.4000 ;
	    RECT 492.4000 31.8000 493.2000 40.4000 ;
	    RECT 498.0000 35.8000 498.8000 40.4000 ;
	    RECT 501.2000 35.8000 502.0000 40.4000 ;
	    RECT 506.8000 32.0000 507.6000 40.4000 ;
	    RECT 2.8000 1.6000 3.6000 9.0000 ;
	    RECT 7.6000 1.6000 8.4000 9.0000 ;
	    RECT 12.4000 1.6000 13.2000 10.2000 ;
	    RECT 18.0000 1.6000 18.8000 6.2000 ;
	    RECT 21.2000 1.6000 22.0000 6.2000 ;
	    RECT 26.8000 1.6000 27.6000 10.0000 ;
	    RECT 30.6000 1.6000 31.4000 6.2000 ;
	    RECT 34.8000 1.6000 35.6000 10.2000 ;
	    RECT 38.0000 1.6000 38.8000 9.0000 ;
	    RECT 41.8000 1.6000 42.6000 6.2000 ;
	    RECT 46.0000 1.6000 46.8000 10.2000 ;
	    RECT 49.2000 1.6000 50.0000 9.0000 ;
	    RECT 54.0000 1.6000 54.8000 10.2000 ;
	    RECT 59.6000 1.6000 60.4000 6.2000 ;
	    RECT 62.8000 1.6000 63.6000 6.2000 ;
	    RECT 68.4000 1.6000 69.2000 10.0000 ;
	    RECT 71.6000 1.6000 72.4000 10.2000 ;
	    RECT 75.8000 1.6000 76.6000 6.2000 ;
	    RECT 79.6000 1.6000 80.4000 9.0000 ;
	    RECT 84.4000 1.6000 85.2000 10.0000 ;
	    RECT 90.0000 1.6000 90.8000 6.2000 ;
	    RECT 93.2000 1.6000 94.0000 6.2000 ;
	    RECT 98.8000 1.6000 99.6000 10.2000 ;
	    RECT 103.6000 1.6000 104.4000 9.0000 ;
	    RECT 113.8000 1.6000 114.6000 6.2000 ;
	    RECT 118.0000 1.6000 118.8000 10.2000 ;
	    RECT 120.2000 1.6000 121.0000 6.2000 ;
	    RECT 124.4000 1.6000 125.2000 10.2000 ;
	    RECT 126.6000 1.6000 127.4000 6.2000 ;
	    RECT 130.8000 1.6000 131.6000 10.2000 ;
	    RECT 134.0000 1.6000 134.8000 9.0000 ;
	    RECT 138.8000 1.6000 139.6000 9.0000 ;
	    RECT 143.6000 1.6000 144.4000 10.2000 ;
	    RECT 149.2000 1.6000 150.0000 6.2000 ;
	    RECT 152.4000 1.6000 153.2000 6.2000 ;
	    RECT 158.0000 1.6000 158.8000 10.0000 ;
	    RECT 162.8000 1.6000 163.6000 9.0000 ;
	    RECT 167.6000 1.6000 168.4000 10.2000 ;
	    RECT 173.2000 1.6000 174.0000 6.2000 ;
	    RECT 176.4000 1.6000 177.2000 6.2000 ;
	    RECT 182.0000 1.6000 182.8000 10.0000 ;
	    RECT 186.8000 1.6000 187.6000 9.0000 ;
	    RECT 191.6000 1.6000 192.4000 10.2000 ;
	    RECT 197.2000 1.6000 198.0000 6.2000 ;
	    RECT 200.4000 1.6000 201.2000 6.2000 ;
	    RECT 206.0000 1.6000 206.8000 10.0000 ;
	    RECT 209.2000 1.6000 210.0000 6.2000 ;
	    RECT 212.4000 1.6000 213.2000 6.2000 ;
	    RECT 214.6000 1.6000 215.4000 6.2000 ;
	    RECT 218.8000 1.6000 219.6000 10.2000 ;
	    RECT 220.4000 1.6000 221.2000 10.2000 ;
	    RECT 226.8000 1.6000 227.6000 10.2000 ;
	    RECT 229.0000 1.6000 229.8000 6.2000 ;
	    RECT 233.2000 1.6000 234.0000 10.2000 ;
	    RECT 238.0000 1.6000 238.8000 10.2000 ;
	    RECT 241.2000 1.6000 242.0000 10.0000 ;
	    RECT 246.8000 1.6000 247.6000 6.2000 ;
	    RECT 250.0000 1.6000 250.8000 6.2000 ;
	    RECT 255.6000 1.6000 256.4000 10.2000 ;
	    RECT 266.8000 1.6000 267.6000 9.0000 ;
	    RECT 271.6000 1.6000 272.4000 10.2000 ;
	    RECT 277.2000 1.6000 278.0000 6.2000 ;
	    RECT 280.4000 1.6000 281.2000 6.2000 ;
	    RECT 286.0000 1.6000 286.8000 10.0000 ;
	    RECT 289.2000 1.6000 290.0000 6.2000 ;
	    RECT 292.4000 1.6000 293.2000 6.2000 ;
	    RECT 294.6000 1.6000 295.4000 6.2000 ;
	    RECT 298.8000 1.6000 299.6000 10.2000 ;
	    RECT 302.0000 1.6000 302.8000 10.2000 ;
	    RECT 307.6000 1.6000 308.4000 6.2000 ;
	    RECT 310.8000 1.6000 311.6000 6.2000 ;
	    RECT 316.4000 1.6000 317.2000 10.0000 ;
	    RECT 319.6000 1.6000 320.4000 6.2000 ;
	    RECT 322.8000 1.6000 323.6000 6.2000 ;
	    RECT 325.0000 1.6000 325.8000 6.2000 ;
	    RECT 329.2000 1.6000 330.0000 10.2000 ;
	    RECT 330.8000 1.6000 331.6000 10.2000 ;
	    RECT 335.0000 1.6000 335.8000 6.2000 ;
	    RECT 337.2000 1.6000 338.0000 10.2000 ;
	    RECT 343.6000 1.6000 344.4000 10.2000 ;
	    RECT 348.4000 1.6000 349.2000 10.2000 ;
	    RECT 351.2000 1.6000 352.0000 10.2000 ;
	    RECT 356.4000 1.6000 357.2000 9.8000 ;
	    RECT 361.2000 1.6000 362.0000 9.8000 ;
	    RECT 366.4000 1.6000 367.2000 10.2000 ;
	    RECT 370.8000 1.6000 371.6000 10.2000 ;
	    RECT 376.4000 1.6000 377.2000 6.2000 ;
	    RECT 379.6000 1.6000 380.4000 6.2000 ;
	    RECT 385.2000 1.6000 386.0000 10.0000 ;
	    RECT 390.0000 1.6000 390.8000 10.2000 ;
	    RECT 395.6000 1.6000 396.4000 6.2000 ;
	    RECT 398.8000 1.6000 399.6000 6.2000 ;
	    RECT 404.4000 1.6000 405.2000 10.0000 ;
	    RECT 414.0000 1.6000 414.8000 6.2000 ;
	    RECT 417.2000 1.6000 418.0000 6.2000 ;
	    RECT 419.4000 1.6000 420.2000 6.2000 ;
	    RECT 423.6000 1.6000 424.4000 10.2000 ;
	    RECT 426.8000 1.6000 427.6000 10.2000 ;
	    RECT 432.4000 1.6000 433.2000 6.2000 ;
	    RECT 435.6000 1.6000 436.4000 6.2000 ;
	    RECT 441.2000 1.6000 442.0000 10.0000 ;
	    RECT 444.4000 1.6000 445.2000 10.2000 ;
	    RECT 448.6000 1.6000 449.4000 6.2000 ;
	    RECT 450.8000 1.6000 451.6000 6.2000 ;
	    RECT 454.0000 1.6000 454.8000 6.2000 ;
	    RECT 455.6000 1.6000 456.4000 10.2000 ;
	    RECT 459.8000 1.6000 460.6000 6.2000 ;
	    RECT 463.6000 1.6000 464.4000 10.2000 ;
	    RECT 469.2000 1.6000 470.0000 6.2000 ;
	    RECT 472.4000 1.6000 473.2000 6.2000 ;
	    RECT 478.0000 1.6000 478.8000 10.0000 ;
	    RECT 482.8000 1.6000 483.6000 10.2000 ;
	    RECT 488.4000 1.6000 489.2000 6.2000 ;
	    RECT 491.6000 1.6000 492.4000 6.2000 ;
	    RECT 497.2000 1.6000 498.0000 10.0000 ;
	    RECT 500.4000 1.6000 501.2000 10.2000 ;
	    RECT 503.6000 1.6000 504.4000 10.2000 ;
	    RECT 506.8000 1.6000 507.6000 10.2000 ;
	    RECT 510.0000 1.6000 510.8000 10.2000 ;
	    RECT 513.2000 1.6000 514.0000 10.2000 ;
	    RECT 0.4000 0.4000 514.8000 1.6000 ;
         LAYER metal2 ;
	    RECT 106.6000 321.4000 107.8000 321.6000 ;
	    RECT 407.4000 321.4000 408.6000 321.6000 ;
	    RECT 104.3000 320.6000 110.1000 321.4000 ;
	    RECT 405.1000 320.6000 410.9000 321.4000 ;
	    RECT 106.6000 320.4000 107.8000 320.6000 ;
	    RECT 407.4000 320.4000 408.6000 320.6000 ;
	    RECT 106.6000 281.4000 107.8000 281.6000 ;
	    RECT 407.4000 281.4000 408.6000 281.6000 ;
	    RECT 104.3000 280.6000 110.1000 281.4000 ;
	    RECT 405.1000 280.6000 410.9000 281.4000 ;
	    RECT 106.6000 280.4000 107.8000 280.6000 ;
	    RECT 407.4000 280.4000 408.6000 280.6000 ;
	    RECT 106.6000 241.4000 107.8000 241.6000 ;
	    RECT 407.4000 241.4000 408.6000 241.6000 ;
	    RECT 104.3000 240.6000 110.1000 241.4000 ;
	    RECT 405.1000 240.6000 410.9000 241.4000 ;
	    RECT 106.6000 240.4000 107.8000 240.6000 ;
	    RECT 407.4000 240.4000 408.6000 240.6000 ;
	    RECT 106.6000 201.4000 107.8000 201.6000 ;
	    RECT 407.4000 201.4000 408.6000 201.6000 ;
	    RECT 104.3000 200.6000 110.1000 201.4000 ;
	    RECT 405.1000 200.6000 410.9000 201.4000 ;
	    RECT 106.6000 200.4000 107.8000 200.6000 ;
	    RECT 407.4000 200.4000 408.6000 200.6000 ;
	    RECT 106.6000 161.4000 107.8000 161.6000 ;
	    RECT 407.4000 161.4000 408.6000 161.6000 ;
	    RECT 104.3000 160.6000 110.1000 161.4000 ;
	    RECT 405.1000 160.6000 410.9000 161.4000 ;
	    RECT 106.6000 160.4000 107.8000 160.6000 ;
	    RECT 407.4000 160.4000 408.6000 160.6000 ;
	    RECT 106.6000 121.4000 107.8000 121.6000 ;
	    RECT 407.4000 121.4000 408.6000 121.6000 ;
	    RECT 104.3000 120.6000 110.1000 121.4000 ;
	    RECT 405.1000 120.6000 410.9000 121.4000 ;
	    RECT 106.6000 120.4000 107.8000 120.6000 ;
	    RECT 407.4000 120.4000 408.6000 120.6000 ;
	    RECT 106.6000 81.4000 107.8000 81.6000 ;
	    RECT 407.4000 81.4000 408.6000 81.6000 ;
	    RECT 104.3000 80.6000 110.1000 81.4000 ;
	    RECT 405.1000 80.6000 410.9000 81.4000 ;
	    RECT 106.6000 80.4000 107.8000 80.6000 ;
	    RECT 407.4000 80.4000 408.6000 80.6000 ;
	    RECT 106.6000 41.4000 107.8000 41.6000 ;
	    RECT 407.4000 41.4000 408.6000 41.6000 ;
	    RECT 104.3000 40.6000 110.1000 41.4000 ;
	    RECT 405.1000 40.6000 410.9000 41.4000 ;
	    RECT 106.6000 40.4000 107.8000 40.6000 ;
	    RECT 407.4000 40.4000 408.6000 40.6000 ;
	    RECT 106.6000 1.4000 107.8000 1.6000 ;
	    RECT 407.4000 1.4000 408.6000 1.6000 ;
	    RECT 104.3000 0.6000 110.1000 1.4000 ;
	    RECT 405.1000 0.6000 410.9000 1.4000 ;
	    RECT 106.6000 0.4000 107.8000 0.6000 ;
	    RECT 407.4000 0.4000 408.6000 0.6000 ;
         LAYER metal3 ;
	    RECT 104.2000 320.4000 110.2000 321.6000 ;
	    RECT 405.0000 320.4000 411.0000 321.6000 ;
	    RECT 104.2000 280.4000 110.2000 281.6000 ;
	    RECT 405.0000 280.4000 411.0000 281.6000 ;
	    RECT 104.2000 240.4000 110.2000 241.6000 ;
	    RECT 405.0000 240.4000 411.0000 241.6000 ;
	    RECT 104.2000 200.4000 110.2000 201.6000 ;
	    RECT 405.0000 200.4000 411.0000 201.6000 ;
	    RECT 104.2000 160.4000 110.2000 161.6000 ;
	    RECT 405.0000 160.4000 411.0000 161.6000 ;
	    RECT 104.2000 120.4000 110.2000 121.6000 ;
	    RECT 405.0000 120.4000 411.0000 121.6000 ;
	    RECT 104.2000 80.4000 110.2000 81.6000 ;
	    RECT 405.0000 80.4000 411.0000 81.6000 ;
	    RECT 104.2000 40.4000 110.2000 41.6000 ;
	    RECT 405.0000 40.4000 411.0000 41.6000 ;
	    RECT 104.2000 0.4000 110.2000 1.6000 ;
	    RECT 405.0000 0.4000 411.0000 1.6000 ;
         LAYER metal4 ;
	    RECT 104.0000 -1.0000 110.4000 341.6000 ;
	    RECT 404.8000 -1.0000 411.2000 341.6000 ;
      END
   END vdd
   PIN clock
      PORT
         LAYER metal1 ;
	    RECT 92.4000 333.8000 93.2000 334.4000 ;
	    RECT 91.4000 333.0000 93.2000 333.8000 ;
	    RECT 228.4000 333.8000 229.2000 334.4000 ;
	    RECT 228.4000 333.0000 230.2000 333.8000 ;
	    RECT 22.6000 308.2000 24.4000 309.0000 ;
	    RECT 502.6000 308.2000 504.4000 309.0000 ;
	    RECT 23.6000 307.6000 24.4000 308.2000 ;
	    RECT 503.6000 307.6000 504.4000 308.2000 ;
	    RECT 446.6000 268.2000 448.4000 269.0000 ;
	    RECT 447.6000 267.6000 448.4000 268.2000 ;
	    RECT 49.2000 253.8000 50.0000 254.4000 ;
	    RECT 48.2000 253.0000 50.0000 253.8000 ;
	    RECT 388.4000 174.3000 389.2000 174.4000 ;
	    RECT 390.0000 174.3000 390.8000 174.4000 ;
	    RECT 388.4000 173.8000 390.8000 174.3000 ;
	    RECT 387.4000 173.7000 390.8000 173.8000 ;
	    RECT 387.4000 173.0000 389.2000 173.7000 ;
	    RECT 390.0000 173.6000 390.8000 173.7000 ;
	    RECT 57.2000 68.2000 59.0000 69.0000 ;
	    RECT 443.4000 68.2000 445.2000 69.0000 ;
	    RECT 512.2000 68.2000 514.0000 69.0000 ;
	    RECT 57.2000 67.6000 58.0000 68.2000 ;
	    RECT 444.4000 67.6000 445.2000 68.2000 ;
	    RECT 513.2000 67.6000 514.0000 68.2000 ;
	    RECT 6.0000 53.8000 6.8000 54.4000 ;
	    RECT 6.0000 53.0000 7.8000 53.8000 ;
	    RECT 513.2000 13.8000 514.0000 14.4000 ;
	    RECT 512.2000 13.0000 514.0000 13.8000 ;
         LAYER metal2 ;
	    RECT 268.4000 341.6000 269.2000 342.4000 ;
	    RECT 447.6000 341.6000 448.4000 342.4000 ;
	    RECT 92.4000 339.6000 93.2000 340.4000 ;
	    RECT 228.4000 339.6000 229.2000 340.4000 ;
	    RECT 252.4000 339.6000 253.2000 340.4000 ;
	    RECT 92.5000 334.4000 93.1000 339.6000 ;
	    RECT 228.5000 334.4000 229.1000 339.6000 ;
	    RECT 92.4000 333.6000 93.2000 334.4000 ;
	    RECT 228.4000 333.6000 229.2000 334.4000 ;
	    RECT 92.5000 308.4000 93.1000 333.6000 ;
	    RECT 252.5000 330.4000 253.1000 339.6000 ;
	    RECT 268.5000 330.4000 269.1000 341.6000 ;
	    RECT 252.4000 329.6000 253.2000 330.4000 ;
	    RECT 268.4000 329.6000 269.2000 330.4000 ;
	    RECT 447.7000 314.4000 448.3000 341.6000 ;
	    RECT 447.6000 313.6000 448.4000 314.4000 ;
	    RECT 503.6000 313.6000 504.4000 314.4000 ;
	    RECT 23.6000 307.6000 24.4000 308.4000 ;
	    RECT 50.8000 307.6000 51.6000 308.4000 ;
	    RECT 92.4000 307.6000 93.2000 308.4000 ;
	    RECT 50.9000 256.3000 51.5000 307.6000 ;
	    RECT 447.7000 268.4000 448.3000 313.6000 ;
	    RECT 503.7000 308.4000 504.3000 313.6000 ;
	    RECT 503.6000 307.6000 504.4000 308.4000 ;
	    RECT 447.6000 267.6000 448.4000 268.4000 ;
	    RECT 49.3000 255.7000 51.5000 256.3000 ;
	    RECT 49.3000 254.4000 49.9000 255.7000 ;
	    RECT 49.2000 253.6000 50.0000 254.4000 ;
	    RECT 49.3000 238.4000 49.9000 253.6000 ;
	    RECT 49.2000 237.6000 50.0000 238.4000 ;
	    RECT 390.0000 205.6000 390.8000 206.4000 ;
	    RECT 390.1000 178.4000 390.7000 205.6000 ;
	    RECT 390.0000 177.6000 390.8000 178.4000 ;
	    RECT 390.1000 174.4000 390.7000 177.6000 ;
	    RECT 390.0000 173.6000 390.8000 174.4000 ;
	    RECT 444.4000 77.6000 445.2000 78.4000 ;
	    RECT 513.2000 77.6000 514.0000 78.4000 ;
	    RECT 444.5000 68.4000 445.1000 77.6000 ;
	    RECT 513.3000 68.4000 513.9000 77.6000 ;
	    RECT 6.0000 67.6000 6.8000 68.4000 ;
	    RECT 57.2000 67.6000 58.0000 68.4000 ;
	    RECT 444.4000 67.6000 445.2000 68.4000 ;
	    RECT 513.2000 67.6000 514.0000 68.4000 ;
	    RECT 6.1000 54.4000 6.7000 67.6000 ;
	    RECT 6.0000 53.6000 6.8000 54.4000 ;
	    RECT 513.3000 14.4000 513.9000 67.6000 ;
	    RECT 513.2000 13.6000 514.0000 14.4000 ;
         LAYER metal3 ;
	    RECT 268.4000 342.3000 269.2000 342.4000 ;
	    RECT 385.2000 342.3000 386.0000 342.4000 ;
	    RECT 447.6000 342.3000 448.4000 342.4000 ;
	    RECT 268.4000 341.7000 448.4000 342.3000 ;
	    RECT 268.4000 341.6000 269.2000 341.7000 ;
	    RECT 385.2000 341.6000 386.0000 341.7000 ;
	    RECT 447.6000 341.6000 448.4000 341.7000 ;
	    RECT 92.4000 340.3000 93.2000 340.4000 ;
	    RECT 228.4000 340.3000 229.2000 340.4000 ;
	    RECT 252.4000 340.3000 253.2000 340.4000 ;
	    RECT 92.4000 339.7000 253.2000 340.3000 ;
	    RECT 92.4000 339.6000 93.2000 339.7000 ;
	    RECT 228.4000 339.6000 229.2000 339.7000 ;
	    RECT 252.4000 339.6000 253.2000 339.7000 ;
	    RECT 252.4000 330.3000 253.2000 330.4000 ;
	    RECT 268.4000 330.3000 269.2000 330.4000 ;
	    RECT 252.4000 329.7000 269.2000 330.3000 ;
	    RECT 252.4000 329.6000 253.2000 329.7000 ;
	    RECT 268.4000 329.6000 269.2000 329.7000 ;
	    RECT 447.6000 314.3000 448.4000 314.4000 ;
	    RECT 503.6000 314.3000 504.4000 314.4000 ;
	    RECT 447.6000 313.7000 504.4000 314.3000 ;
	    RECT 447.6000 313.6000 448.4000 313.7000 ;
	    RECT 503.6000 313.6000 504.4000 313.7000 ;
	    RECT 23.6000 308.3000 24.4000 308.4000 ;
	    RECT 50.8000 308.3000 51.6000 308.4000 ;
	    RECT 92.4000 308.3000 93.2000 308.4000 ;
	    RECT 23.6000 307.7000 93.2000 308.3000 ;
	    RECT 23.6000 307.6000 24.4000 307.7000 ;
	    RECT 50.8000 307.6000 51.6000 307.7000 ;
	    RECT 92.4000 307.6000 93.2000 307.7000 ;
	    RECT 49.2000 237.6000 50.0000 238.4000 ;
	    RECT 385.2000 206.3000 386.0000 206.4000 ;
	    RECT 390.0000 206.3000 390.8000 206.4000 ;
	    RECT 385.2000 205.7000 390.8000 206.3000 ;
	    RECT 385.2000 205.6000 386.0000 205.7000 ;
	    RECT 390.0000 205.6000 390.8000 205.7000 ;
	    RECT 390.0000 178.3000 390.8000 178.4000 ;
	    RECT 423.6000 178.3000 424.4000 178.4000 ;
	    RECT 390.0000 177.7000 424.4000 178.3000 ;
	    RECT 390.0000 177.6000 390.8000 177.7000 ;
	    RECT 423.6000 177.6000 424.4000 177.7000 ;
	    RECT 49.2000 170.3000 50.0000 170.4000 ;
	    RECT 55.6000 170.3000 56.4000 170.4000 ;
	    RECT 49.2000 169.7000 56.4000 170.3000 ;
	    RECT 49.2000 169.6000 50.0000 169.7000 ;
	    RECT 55.6000 169.6000 56.4000 169.7000 ;
	    RECT 444.4000 78.3000 445.2000 78.4000 ;
	    RECT 513.2000 78.3000 514.0000 78.4000 ;
	    RECT 444.4000 77.7000 514.0000 78.3000 ;
	    RECT 444.4000 77.6000 445.2000 77.7000 ;
	    RECT 513.2000 77.6000 514.0000 77.7000 ;
	    RECT 6.0000 68.3000 6.8000 68.4000 ;
	    RECT 55.6000 68.3000 56.4000 68.4000 ;
	    RECT 57.2000 68.3000 58.0000 68.4000 ;
	    RECT 6.0000 67.7000 58.0000 68.3000 ;
	    RECT 6.0000 67.6000 6.8000 67.7000 ;
	    RECT 55.6000 67.6000 56.4000 67.7000 ;
	    RECT 57.2000 67.6000 58.0000 67.7000 ;
	    RECT 423.6000 68.3000 424.4000 68.4000 ;
	    RECT 444.4000 68.3000 445.2000 68.4000 ;
	    RECT 423.6000 67.7000 445.2000 68.3000 ;
	    RECT 423.6000 67.6000 424.4000 67.7000 ;
	    RECT 444.4000 67.6000 445.2000 67.7000 ;
	    RECT 513.2000 14.3000 514.0000 14.4000 ;
	    RECT 513.2000 13.7000 518.7000 14.3000 ;
	    RECT 513.2000 13.6000 514.0000 13.7000 ;
         LAYER metal4 ;
	    RECT 49.0000 169.4000 50.2000 238.6000 ;
	    RECT 385.0000 205.4000 386.2000 342.6000 ;
	    RECT 55.4000 67.4000 56.6000 170.6000 ;
	    RECT 423.4000 67.4000 424.6000 178.6000 ;
      END
   END clock
   PIN data_in[15]
      PORT
         LAYER metal1 ;
	    RECT 194.8000 333.6000 195.6000 335.2000 ;
	    RECT 398.0000 329.6000 398.8000 331.2000 ;
	    RECT 417.2000 329.6000 418.0000 332.4000 ;
         LAYER metal2 ;
	    RECT 194.9000 338.4000 195.5000 346.3000 ;
	    RECT 398.0000 339.6000 398.8000 340.4000 ;
	    RECT 194.8000 337.6000 195.6000 338.4000 ;
	    RECT 194.9000 334.4000 195.5000 337.6000 ;
	    RECT 194.8000 333.6000 195.6000 334.4000 ;
	    RECT 398.1000 332.4000 398.7000 339.6000 ;
	    RECT 398.0000 331.6000 398.8000 332.4000 ;
	    RECT 417.2000 331.6000 418.0000 332.4000 ;
	    RECT 398.1000 330.4000 398.7000 331.6000 ;
	    RECT 398.0000 329.6000 398.8000 330.4000 ;
         LAYER metal3 ;
	    RECT 398.0000 340.3000 398.8000 340.4000 ;
	    RECT 262.1000 339.7000 398.8000 340.3000 ;
	    RECT 194.8000 338.3000 195.6000 338.4000 ;
	    RECT 262.1000 338.3000 262.7000 339.7000 ;
	    RECT 398.0000 339.6000 398.8000 339.7000 ;
	    RECT 194.8000 337.7000 262.7000 338.3000 ;
	    RECT 194.8000 337.6000 195.6000 337.7000 ;
	    RECT 398.0000 332.3000 398.8000 332.4000 ;
	    RECT 417.2000 332.3000 418.0000 332.4000 ;
	    RECT 398.0000 331.7000 418.0000 332.3000 ;
	    RECT 398.0000 331.6000 398.8000 331.7000 ;
	    RECT 417.2000 331.6000 418.0000 331.7000 ;
      END
   END data_in[15]
   PIN data_in[14]
      PORT
         LAYER metal1 ;
	    RECT 473.2000 190.8000 474.0000 192.4000 ;
	    RECT 446.0000 186.8000 446.8000 188.4000 ;
	    RECT 479.6000 169.6000 480.4000 172.4000 ;
         LAYER metal2 ;
	    RECT 473.2000 191.6000 474.0000 192.4000 ;
	    RECT 446.0000 187.6000 446.8000 188.4000 ;
	    RECT 446.1000 180.4000 446.7000 187.6000 ;
	    RECT 473.3000 184.4000 473.9000 191.6000 ;
	    RECT 473.2000 183.6000 474.0000 184.4000 ;
	    RECT 479.6000 183.6000 480.4000 184.4000 ;
	    RECT 473.3000 180.4000 473.9000 183.6000 ;
	    RECT 446.0000 179.6000 446.8000 180.4000 ;
	    RECT 473.2000 179.6000 474.0000 180.4000 ;
	    RECT 479.7000 172.4000 480.3000 183.6000 ;
	    RECT 511.6000 179.6000 512.4000 180.4000 ;
	    RECT 511.7000 176.4000 512.3000 179.6000 ;
	    RECT 511.6000 175.6000 512.4000 176.4000 ;
	    RECT 479.6000 171.6000 480.4000 172.4000 ;
         LAYER metal3 ;
	    RECT 473.2000 184.3000 474.0000 184.4000 ;
	    RECT 479.6000 184.3000 480.4000 184.4000 ;
	    RECT 473.2000 183.7000 480.4000 184.3000 ;
	    RECT 473.2000 183.6000 474.0000 183.7000 ;
	    RECT 479.6000 183.6000 480.4000 183.7000 ;
	    RECT 446.0000 180.3000 446.8000 180.4000 ;
	    RECT 473.2000 180.3000 474.0000 180.4000 ;
	    RECT 511.6000 180.3000 512.4000 180.4000 ;
	    RECT 446.0000 179.7000 512.4000 180.3000 ;
	    RECT 446.0000 179.6000 446.8000 179.7000 ;
	    RECT 473.2000 179.6000 474.0000 179.7000 ;
	    RECT 511.6000 179.6000 512.4000 179.7000 ;
	    RECT 511.6000 176.3000 512.4000 176.4000 ;
	    RECT 511.6000 175.7000 518.7000 176.3000 ;
	    RECT 511.6000 175.6000 512.4000 175.7000 ;
      END
   END data_in[14]
   PIN data_in[13]
      PORT
         LAYER metal1 ;
	    RECT 460.4000 190.8000 461.2000 192.4000 ;
	    RECT 454.0000 186.8000 454.8000 188.4000 ;
	    RECT 458.8000 169.6000 459.6000 172.4000 ;
         LAYER metal2 ;
	    RECT 460.4000 191.6000 461.2000 192.4000 ;
	    RECT 454.0000 187.6000 454.8000 188.4000 ;
	    RECT 460.5000 188.3000 461.1000 191.6000 ;
	    RECT 458.9000 187.7000 461.1000 188.3000 ;
	    RECT 454.1000 184.4000 454.7000 187.6000 ;
	    RECT 458.9000 184.4000 459.5000 187.7000 ;
	    RECT 454.0000 183.6000 454.8000 184.4000 ;
	    RECT 458.8000 183.6000 459.6000 184.4000 ;
	    RECT 458.9000 182.4000 459.5000 183.6000 ;
	    RECT 458.8000 181.6000 459.6000 182.4000 ;
	    RECT 458.9000 172.4000 459.5000 181.6000 ;
	    RECT 458.8000 171.6000 459.6000 172.4000 ;
         LAYER metal3 ;
	    RECT 513.2000 188.3000 514.0000 188.4000 ;
	    RECT 518.1000 188.3000 518.7000 190.3000 ;
	    RECT 513.2000 187.7000 518.7000 188.3000 ;
	    RECT 513.2000 187.6000 514.0000 187.7000 ;
	    RECT 454.0000 184.3000 454.8000 184.4000 ;
	    RECT 458.8000 184.3000 459.6000 184.4000 ;
	    RECT 454.0000 183.7000 459.6000 184.3000 ;
	    RECT 454.0000 183.6000 454.8000 183.7000 ;
	    RECT 458.8000 183.6000 459.6000 183.7000 ;
	    RECT 458.8000 182.3000 459.6000 182.4000 ;
	    RECT 513.2000 182.3000 514.0000 182.4000 ;
	    RECT 458.8000 181.7000 514.0000 182.3000 ;
	    RECT 458.8000 181.6000 459.6000 181.7000 ;
	    RECT 513.2000 181.6000 514.0000 181.7000 ;
         LAYER metal4 ;
	    RECT 513.0000 181.4000 514.2000 188.6000 ;
      END
   END data_in[13]
   PIN data_in[12]
      PORT
         LAYER metal1 ;
	    RECT 489.2000 70.8000 490.0000 72.4000 ;
	    RECT 474.8000 53.6000 475.6000 55.2000 ;
	    RECT 474.9000 52.3000 475.5000 53.6000 ;
	    RECT 476.4000 52.3000 477.2000 52.4000 ;
	    RECT 474.9000 51.7000 477.2000 52.3000 ;
	    RECT 476.4000 49.6000 477.2000 51.7000 ;
         LAYER metal2 ;
	    RECT 489.2000 71.6000 490.0000 72.4000 ;
	    RECT 489.3000 70.4000 489.9000 71.6000 ;
	    RECT 476.4000 69.6000 477.2000 70.4000 ;
	    RECT 489.2000 69.6000 490.0000 70.4000 ;
	    RECT 476.5000 52.4000 477.1000 69.6000 ;
	    RECT 476.4000 51.6000 477.2000 52.4000 ;
         LAYER metal3 ;
	    RECT 476.4000 70.3000 477.2000 70.4000 ;
	    RECT 489.2000 70.3000 490.0000 70.4000 ;
	    RECT 476.4000 69.7000 518.7000 70.3000 ;
	    RECT 476.4000 69.6000 477.2000 69.7000 ;
	    RECT 489.2000 69.6000 490.0000 69.7000 ;
      END
   END data_in[12]
   PIN data_in[11]
      PORT
         LAYER metal1 ;
	    RECT 367.6000 333.6000 368.4000 335.2000 ;
	    RECT 410.8000 329.6000 411.6000 331.2000 ;
	    RECT 423.6000 329.6000 424.4000 332.4000 ;
         LAYER metal2 ;
	    RECT 367.7000 336.4000 368.3000 346.3000 ;
	    RECT 367.6000 335.6000 368.4000 336.4000 ;
	    RECT 367.7000 334.4000 368.3000 335.6000 ;
	    RECT 367.6000 333.6000 368.4000 334.4000 ;
	    RECT 410.8000 333.6000 411.6000 334.4000 ;
	    RECT 423.6000 333.6000 424.4000 334.4000 ;
	    RECT 410.9000 330.4000 411.5000 333.6000 ;
	    RECT 423.7000 332.4000 424.3000 333.6000 ;
	    RECT 423.6000 331.6000 424.4000 332.4000 ;
	    RECT 410.8000 329.6000 411.6000 330.4000 ;
         LAYER metal3 ;
	    RECT 367.6000 336.3000 368.4000 336.4000 ;
	    RECT 367.6000 335.7000 411.5000 336.3000 ;
	    RECT 367.6000 335.6000 368.4000 335.7000 ;
	    RECT 410.9000 334.4000 411.5000 335.7000 ;
	    RECT 410.8000 334.3000 411.6000 334.4000 ;
	    RECT 423.6000 334.3000 424.4000 334.4000 ;
	    RECT 410.8000 333.7000 424.4000 334.3000 ;
	    RECT 410.8000 333.6000 411.6000 333.7000 ;
	    RECT 423.6000 333.6000 424.4000 333.7000 ;
      END
   END data_in[11]
   PIN data_in[10]
      PORT
         LAYER metal1 ;
	    RECT 500.4000 110.8000 501.2000 112.4000 ;
	    RECT 484.4000 53.6000 485.2000 55.2000 ;
	    RECT 490.8000 49.6000 491.6000 52.4000 ;
         LAYER metal2 ;
	    RECT 500.4000 115.6000 501.2000 116.4000 ;
	    RECT 500.5000 112.4000 501.1000 115.6000 ;
	    RECT 500.4000 111.6000 501.2000 112.4000 ;
	    RECT 484.4000 53.6000 485.2000 54.4000 ;
	    RECT 490.8000 53.6000 491.6000 54.4000 ;
	    RECT 490.9000 52.4000 491.5000 53.6000 ;
	    RECT 490.8000 51.6000 491.6000 52.4000 ;
         LAYER metal3 ;
	    RECT 500.4000 116.3000 501.2000 116.4000 ;
	    RECT 500.4000 115.7000 518.7000 116.3000 ;
	    RECT 500.4000 115.6000 501.2000 115.7000 ;
	    RECT 494.0000 112.3000 494.8000 112.4000 ;
	    RECT 500.4000 112.3000 501.2000 112.4000 ;
	    RECT 494.0000 111.7000 501.2000 112.3000 ;
	    RECT 494.0000 111.6000 494.8000 111.7000 ;
	    RECT 500.4000 111.6000 501.2000 111.7000 ;
	    RECT 484.4000 54.3000 485.2000 54.4000 ;
	    RECT 490.8000 54.3000 491.6000 54.4000 ;
	    RECT 494.0000 54.3000 494.8000 54.4000 ;
	    RECT 484.4000 53.7000 494.8000 54.3000 ;
	    RECT 484.4000 53.6000 485.2000 53.7000 ;
	    RECT 490.8000 53.6000 491.6000 53.7000 ;
	    RECT 494.0000 53.6000 494.8000 53.7000 ;
         LAYER metal4 ;
	    RECT 493.8000 53.4000 495.0000 112.6000 ;
      END
   END data_in[10]
   PIN data_in[9]
      PORT
         LAYER metal1 ;
	    RECT 503.6000 289.6000 504.4000 291.2000 ;
	    RECT 506.8000 110.8000 507.6000 112.4000 ;
	    RECT 466.8000 106.8000 467.6000 108.4000 ;
         LAYER metal2 ;
	    RECT 503.6000 289.6000 504.4000 290.4000 ;
	    RECT 503.7000 274.4000 504.3000 289.6000 ;
	    RECT 503.6000 273.6000 504.4000 274.4000 ;
	    RECT 466.8000 121.6000 467.6000 122.4000 ;
	    RECT 506.8000 121.6000 507.6000 122.4000 ;
	    RECT 466.9000 108.4000 467.5000 121.6000 ;
	    RECT 506.9000 112.4000 507.5000 121.6000 ;
	    RECT 506.8000 111.6000 507.6000 112.4000 ;
	    RECT 466.8000 107.6000 467.6000 108.4000 ;
         LAYER metal3 ;
	    RECT 497.2000 274.3000 498.0000 274.4000 ;
	    RECT 503.6000 274.3000 504.4000 274.4000 ;
	    RECT 497.2000 273.7000 504.4000 274.3000 ;
	    RECT 497.2000 273.6000 498.0000 273.7000 ;
	    RECT 503.6000 273.6000 504.4000 273.7000 ;
	    RECT 490.8000 248.3000 491.6000 248.4000 ;
	    RECT 497.2000 248.3000 498.0000 248.4000 ;
	    RECT 490.8000 247.7000 498.0000 248.3000 ;
	    RECT 490.8000 247.6000 491.6000 247.7000 ;
	    RECT 497.2000 247.6000 498.0000 247.7000 ;
	    RECT 466.8000 122.3000 467.6000 122.4000 ;
	    RECT 490.8000 122.3000 491.6000 122.4000 ;
	    RECT 506.8000 122.3000 507.6000 122.4000 ;
	    RECT 466.8000 121.7000 518.7000 122.3000 ;
	    RECT 466.8000 121.6000 467.6000 121.7000 ;
	    RECT 490.8000 121.6000 491.6000 121.7000 ;
	    RECT 506.8000 121.6000 507.6000 121.7000 ;
	    RECT 518.1000 119.7000 518.7000 121.7000 ;
         LAYER metal4 ;
	    RECT 490.6000 121.4000 491.8000 248.6000 ;
	    RECT 497.0000 247.4000 498.2000 274.6000 ;
      END
   END data_in[9]
   PIN data_in[8]
      PORT
         LAYER metal1 ;
	    RECT 463.6000 330.3000 464.4000 331.2000 ;
	    RECT 465.2000 330.3000 466.0000 332.4000 ;
	    RECT 463.6000 329.7000 466.0000 330.3000 ;
	    RECT 463.6000 329.6000 464.4000 329.7000 ;
	    RECT 465.2000 329.6000 466.0000 329.7000 ;
	    RECT 457.2000 306.8000 458.0000 308.4000 ;
         LAYER metal2 ;
	    RECT 465.3000 345.7000 467.5000 346.3000 ;
	    RECT 465.3000 332.4000 465.9000 345.7000 ;
	    RECT 465.2000 331.6000 466.0000 332.4000 ;
	    RECT 465.3000 310.4000 465.9000 331.6000 ;
	    RECT 457.2000 309.6000 458.0000 310.4000 ;
	    RECT 465.2000 309.6000 466.0000 310.4000 ;
	    RECT 457.3000 308.4000 457.9000 309.6000 ;
	    RECT 457.2000 307.6000 458.0000 308.4000 ;
         LAYER metal3 ;
	    RECT 457.2000 310.3000 458.0000 310.4000 ;
	    RECT 465.2000 310.3000 466.0000 310.4000 ;
	    RECT 457.2000 309.7000 466.0000 310.3000 ;
	    RECT 457.2000 309.6000 458.0000 309.7000 ;
	    RECT 465.2000 309.6000 466.0000 309.7000 ;
      END
   END data_in[8]
   PIN data_in[7]
      PORT
         LAYER metal1 ;
	    RECT 438.0000 230.8000 438.8000 232.4000 ;
	    RECT 438.0000 213.6000 438.8000 215.2000 ;
	    RECT 442.8000 210.3000 443.6000 210.4000 ;
	    RECT 444.4000 210.3000 445.2000 211.2000 ;
	    RECT 442.8000 209.7000 445.2000 210.3000 ;
	    RECT 442.8000 209.6000 443.6000 209.7000 ;
	    RECT 444.4000 209.6000 445.2000 209.7000 ;
         LAYER metal2 ;
	    RECT 438.0000 231.6000 438.8000 232.4000 ;
	    RECT 438.1000 218.4000 438.7000 231.6000 ;
	    RECT 438.0000 217.6000 438.8000 218.4000 ;
	    RECT 514.8000 217.6000 515.6000 218.4000 ;
	    RECT 438.1000 214.4000 438.7000 217.6000 ;
	    RECT 438.0000 213.6000 438.8000 214.4000 ;
	    RECT 438.1000 210.4000 438.7000 213.6000 ;
	    RECT 514.9000 212.4000 515.5000 217.6000 ;
	    RECT 514.8000 211.6000 515.6000 212.4000 ;
	    RECT 438.0000 209.6000 438.8000 210.4000 ;
	    RECT 442.8000 209.6000 443.6000 210.4000 ;
         LAYER metal3 ;
	    RECT 438.0000 218.3000 438.8000 218.4000 ;
	    RECT 514.8000 218.3000 515.6000 218.4000 ;
	    RECT 438.0000 217.7000 515.6000 218.3000 ;
	    RECT 438.0000 217.6000 438.8000 217.7000 ;
	    RECT 514.8000 217.6000 515.6000 217.7000 ;
	    RECT 514.8000 212.3000 515.6000 212.4000 ;
	    RECT 514.8000 211.7000 518.7000 212.3000 ;
	    RECT 514.8000 211.6000 515.6000 211.7000 ;
	    RECT 438.0000 210.3000 438.8000 210.4000 ;
	    RECT 442.8000 210.3000 443.6000 210.4000 ;
	    RECT 438.0000 209.7000 443.6000 210.3000 ;
	    RECT 438.0000 209.6000 438.8000 209.7000 ;
	    RECT 442.8000 209.6000 443.6000 209.7000 ;
      END
   END data_in[7]
   PIN data_in[6]
      PORT
         LAYER metal1 ;
	    RECT 497.2000 89.6000 498.0000 91.2000 ;
	    RECT 465.2000 53.6000 466.0000 55.2000 ;
	    RECT 471.6000 49.6000 472.4000 52.4000 ;
         LAYER metal2 ;
	    RECT 497.2000 89.6000 498.0000 90.4000 ;
	    RECT 497.3000 66.4000 497.9000 89.6000 ;
	    RECT 471.6000 65.6000 472.4000 66.4000 ;
	    RECT 497.2000 65.6000 498.0000 66.4000 ;
	    RECT 471.7000 54.4000 472.3000 65.6000 ;
	    RECT 465.2000 53.6000 466.0000 54.4000 ;
	    RECT 471.6000 53.6000 472.4000 54.4000 ;
	    RECT 471.7000 52.4000 472.3000 53.6000 ;
	    RECT 471.6000 51.6000 472.4000 52.4000 ;
         LAYER metal3 ;
	    RECT 497.2000 90.3000 498.0000 90.4000 ;
	    RECT 497.2000 89.7000 518.7000 90.3000 ;
	    RECT 497.2000 89.6000 498.0000 89.7000 ;
	    RECT 471.6000 66.3000 472.4000 66.4000 ;
	    RECT 497.2000 66.3000 498.0000 66.4000 ;
	    RECT 471.6000 65.7000 498.0000 66.3000 ;
	    RECT 471.6000 65.6000 472.4000 65.7000 ;
	    RECT 497.2000 65.6000 498.0000 65.7000 ;
	    RECT 465.2000 54.3000 466.0000 54.4000 ;
	    RECT 471.6000 54.3000 472.4000 54.4000 ;
	    RECT 465.2000 53.7000 472.4000 54.3000 ;
	    RECT 465.2000 53.6000 466.0000 53.7000 ;
	    RECT 471.6000 53.6000 472.4000 53.7000 ;
      END
   END data_in[6]
   PIN data_in[5]
      PORT
         LAYER metal1 ;
	    RECT 423.6000 293.6000 424.4000 295.2000 ;
	    RECT 490.8000 290.3000 491.6000 291.2000 ;
	    RECT 492.4000 290.3000 493.2000 290.4000 ;
	    RECT 490.8000 289.7000 493.2000 290.3000 ;
	    RECT 490.8000 289.6000 491.6000 289.7000 ;
	    RECT 492.4000 289.6000 493.2000 289.7000 ;
	    RECT 497.2000 289.6000 498.0000 291.2000 ;
         LAYER metal2 ;
	    RECT 423.6000 293.6000 424.4000 294.4000 ;
	    RECT 423.7000 292.4000 424.3000 293.6000 ;
	    RECT 423.6000 291.6000 424.4000 292.4000 ;
	    RECT 492.4000 289.6000 493.2000 290.4000 ;
	    RECT 497.2000 289.6000 498.0000 290.4000 ;
         LAYER metal3 ;
	    RECT 423.6000 292.3000 424.4000 292.4000 ;
	    RECT 423.6000 291.7000 433.9000 292.3000 ;
	    RECT 423.6000 291.6000 424.4000 291.7000 ;
	    RECT 433.3000 290.3000 433.9000 291.7000 ;
	    RECT 497.3000 291.7000 518.7000 292.3000 ;
	    RECT 497.3000 290.4000 497.9000 291.7000 ;
	    RECT 492.4000 290.3000 493.2000 290.4000 ;
	    RECT 497.2000 290.3000 498.0000 290.4000 ;
	    RECT 433.3000 289.7000 498.0000 290.3000 ;
	    RECT 518.1000 289.7000 518.7000 291.7000 ;
	    RECT 492.4000 289.6000 493.2000 289.7000 ;
	    RECT 497.2000 289.6000 498.0000 289.7000 ;
      END
   END data_in[5]
   PIN data_in[4]
      PORT
         LAYER metal1 ;
	    RECT 426.8000 253.6000 427.6000 255.2000 ;
	    RECT 503.6000 249.6000 504.4000 251.2000 ;
	    RECT 484.4000 230.8000 485.2000 232.4000 ;
         LAYER metal2 ;
	    RECT 426.8000 253.6000 427.6000 254.4000 ;
	    RECT 426.9000 242.4000 427.5000 253.6000 ;
	    RECT 503.6000 249.6000 504.4000 250.4000 ;
	    RECT 503.7000 248.4000 504.3000 249.6000 ;
	    RECT 503.6000 247.6000 504.4000 248.4000 ;
	    RECT 503.7000 242.4000 504.3000 247.6000 ;
	    RECT 426.8000 241.6000 427.6000 242.4000 ;
	    RECT 484.4000 241.6000 485.2000 242.4000 ;
	    RECT 503.6000 241.6000 504.4000 242.4000 ;
	    RECT 484.5000 232.4000 485.1000 241.6000 ;
	    RECT 484.4000 231.6000 485.2000 232.4000 ;
         LAYER metal3 ;
	    RECT 503.6000 248.3000 504.4000 248.4000 ;
	    RECT 518.1000 248.3000 518.7000 250.3000 ;
	    RECT 503.6000 247.7000 518.7000 248.3000 ;
	    RECT 503.6000 247.6000 504.4000 247.7000 ;
	    RECT 426.8000 242.3000 427.6000 242.4000 ;
	    RECT 484.4000 242.3000 485.2000 242.4000 ;
	    RECT 503.6000 242.3000 504.4000 242.4000 ;
	    RECT 426.8000 241.7000 504.4000 242.3000 ;
	    RECT 426.8000 241.6000 427.6000 241.7000 ;
	    RECT 484.4000 241.6000 485.2000 241.7000 ;
	    RECT 503.6000 241.6000 504.4000 241.7000 ;
      END
   END data_in[4]
   PIN data_in[3]
      PORT
         LAYER metal1 ;
	    RECT 466.8000 190.8000 467.6000 192.4000 ;
	    RECT 508.4000 189.6000 509.2000 192.4000 ;
	    RECT 330.8000 173.6000 331.6000 175.2000 ;
         LAYER metal2 ;
	    RECT 466.8000 191.6000 467.6000 192.4000 ;
	    RECT 466.9000 188.4000 467.5000 191.6000 ;
	    RECT 508.4000 189.6000 509.2000 190.4000 ;
	    RECT 330.8000 187.6000 331.6000 188.4000 ;
	    RECT 466.8000 187.6000 467.6000 188.4000 ;
	    RECT 330.9000 174.4000 331.5000 187.6000 ;
	    RECT 508.5000 186.4000 509.1000 189.6000 ;
	    RECT 508.4000 185.6000 509.2000 186.4000 ;
	    RECT 514.8000 185.6000 515.6000 186.4000 ;
	    RECT 330.8000 173.6000 331.6000 174.4000 ;
	    RECT 514.9000 172.4000 515.5000 185.6000 ;
	    RECT 514.8000 171.6000 515.6000 172.4000 ;
         LAYER metal3 ;
	    RECT 330.8000 188.3000 331.6000 188.4000 ;
	    RECT 466.8000 188.3000 467.6000 188.4000 ;
	    RECT 330.8000 187.7000 352.3000 188.3000 ;
	    RECT 330.8000 187.6000 331.6000 187.7000 ;
	    RECT 351.7000 186.3000 352.3000 187.7000 ;
	    RECT 402.9000 187.7000 502.7000 188.3000 ;
	    RECT 402.9000 186.3000 403.5000 187.7000 ;
	    RECT 466.8000 187.6000 467.6000 187.7000 ;
	    RECT 351.7000 185.7000 403.5000 186.3000 ;
	    RECT 502.1000 186.3000 502.7000 187.7000 ;
	    RECT 508.4000 186.3000 509.2000 186.4000 ;
	    RECT 514.8000 186.3000 515.6000 186.4000 ;
	    RECT 502.1000 185.7000 515.6000 186.3000 ;
	    RECT 508.4000 185.6000 509.2000 185.7000 ;
	    RECT 514.8000 185.6000 515.6000 185.7000 ;
	    RECT 514.8000 172.3000 515.6000 172.4000 ;
	    RECT 514.8000 171.7000 518.7000 172.3000 ;
	    RECT 514.8000 171.6000 515.6000 171.7000 ;
      END
   END data_in[3]
   PIN data_in[2]
      PORT
         LAYER metal1 ;
	    RECT 455.6000 270.8000 456.4000 272.4000 ;
	    RECT 444.4000 230.8000 445.2000 232.4000 ;
	    RECT 300.4000 226.8000 301.2000 228.4000 ;
         LAYER metal2 ;
	    RECT 455.7000 340.4000 456.3000 346.3000 ;
	    RECT 449.2000 339.6000 450.0000 340.4000 ;
	    RECT 455.6000 339.6000 456.4000 340.4000 ;
	    RECT 449.3000 272.4000 449.9000 339.6000 ;
	    RECT 444.4000 271.6000 445.2000 272.4000 ;
	    RECT 449.2000 271.6000 450.0000 272.4000 ;
	    RECT 455.6000 271.6000 456.4000 272.4000 ;
	    RECT 444.5000 248.4000 445.1000 271.6000 ;
	    RECT 300.4000 247.6000 301.2000 248.4000 ;
	    RECT 444.4000 247.6000 445.2000 248.4000 ;
	    RECT 300.5000 228.4000 301.1000 247.6000 ;
	    RECT 444.5000 232.4000 445.1000 247.6000 ;
	    RECT 444.4000 231.6000 445.2000 232.4000 ;
	    RECT 300.4000 227.6000 301.2000 228.4000 ;
         LAYER metal3 ;
	    RECT 449.2000 340.3000 450.0000 340.4000 ;
	    RECT 455.6000 340.3000 456.4000 340.4000 ;
	    RECT 449.2000 339.7000 456.4000 340.3000 ;
	    RECT 449.2000 339.6000 450.0000 339.7000 ;
	    RECT 455.6000 339.6000 456.4000 339.7000 ;
	    RECT 444.4000 272.3000 445.2000 272.4000 ;
	    RECT 449.2000 272.3000 450.0000 272.4000 ;
	    RECT 455.6000 272.3000 456.4000 272.4000 ;
	    RECT 444.4000 271.7000 456.4000 272.3000 ;
	    RECT 444.4000 271.6000 445.2000 271.7000 ;
	    RECT 449.2000 271.6000 450.0000 271.7000 ;
	    RECT 455.6000 271.6000 456.4000 271.7000 ;
	    RECT 300.4000 248.3000 301.2000 248.4000 ;
	    RECT 444.4000 248.3000 445.2000 248.4000 ;
	    RECT 300.4000 247.7000 445.2000 248.3000 ;
	    RECT 300.4000 247.6000 301.2000 247.7000 ;
	    RECT 444.4000 247.6000 445.2000 247.7000 ;
      END
   END data_in[2]
   PIN data_in[1]
      PORT
         LAYER metal1 ;
	    RECT 394.8000 310.8000 395.6000 312.4000 ;
	    RECT 382.0000 293.6000 382.8000 295.2000 ;
	    RECT 455.6000 289.6000 456.4000 292.4000 ;
         LAYER metal2 ;
	    RECT 394.9000 312.4000 395.5000 346.3000 ;
	    RECT 394.8000 311.6000 395.6000 312.4000 ;
	    RECT 394.9000 308.4000 395.5000 311.6000 ;
	    RECT 382.0000 307.6000 382.8000 308.4000 ;
	    RECT 394.8000 307.6000 395.6000 308.4000 ;
	    RECT 382.1000 294.4000 382.7000 307.6000 ;
	    RECT 382.0000 293.6000 382.8000 294.4000 ;
	    RECT 455.6000 291.6000 456.4000 292.4000 ;
         LAYER metal3 ;
	    RECT 382.0000 308.3000 382.8000 308.4000 ;
	    RECT 394.8000 308.3000 395.6000 308.4000 ;
	    RECT 446.0000 308.3000 446.8000 308.4000 ;
	    RECT 382.0000 307.7000 446.8000 308.3000 ;
	    RECT 382.0000 307.6000 382.8000 307.7000 ;
	    RECT 394.8000 307.6000 395.6000 307.7000 ;
	    RECT 446.0000 307.6000 446.8000 307.7000 ;
	    RECT 446.0000 292.3000 446.8000 292.4000 ;
	    RECT 455.6000 292.3000 456.4000 292.4000 ;
	    RECT 446.0000 291.7000 456.4000 292.3000 ;
	    RECT 446.0000 291.6000 446.8000 291.7000 ;
	    RECT 455.6000 291.6000 456.4000 291.7000 ;
         LAYER metal4 ;
	    RECT 445.8000 291.4000 447.0000 308.6000 ;
      END
   END data_in[1]
   PIN data_in[0]
      PORT
         LAYER metal1 ;
	    RECT 508.4000 129.6000 509.2000 131.2000 ;
	    RECT 470.0000 106.8000 470.8000 108.4000 ;
	    RECT 508.4000 90.3000 509.2000 91.2000 ;
	    RECT 514.8000 90.3000 515.6000 90.4000 ;
	    RECT 508.4000 89.7000 515.6000 90.3000 ;
	    RECT 508.4000 89.6000 509.2000 89.7000 ;
	    RECT 514.8000 89.6000 515.6000 89.7000 ;
         LAYER metal2 ;
	    RECT 508.4000 129.6000 509.2000 130.4000 ;
	    RECT 508.5000 120.4000 509.1000 129.6000 ;
	    RECT 470.0000 119.6000 470.8000 120.4000 ;
	    RECT 508.4000 119.6000 509.2000 120.4000 ;
	    RECT 514.8000 119.6000 515.6000 120.4000 ;
	    RECT 470.1000 108.4000 470.7000 119.6000 ;
	    RECT 514.9000 112.4000 515.5000 119.6000 ;
	    RECT 514.8000 111.6000 515.6000 112.4000 ;
	    RECT 470.0000 107.6000 470.8000 108.4000 ;
	    RECT 514.9000 90.4000 515.5000 111.6000 ;
	    RECT 514.8000 89.6000 515.6000 90.4000 ;
         LAYER metal3 ;
	    RECT 470.0000 120.3000 470.8000 120.4000 ;
	    RECT 508.4000 120.3000 509.2000 120.4000 ;
	    RECT 514.8000 120.3000 515.6000 120.4000 ;
	    RECT 470.0000 119.7000 515.6000 120.3000 ;
	    RECT 470.0000 119.6000 470.8000 119.7000 ;
	    RECT 508.4000 119.6000 509.2000 119.7000 ;
	    RECT 514.8000 119.6000 515.6000 119.7000 ;
	    RECT 514.8000 112.3000 515.6000 112.4000 ;
	    RECT 514.8000 111.7000 518.7000 112.3000 ;
	    RECT 514.8000 111.6000 515.6000 111.7000 ;
      END
   END data_in[0]
   PIN enable
      PORT
         LAYER metal1 ;
	    RECT 7.6000 174.3000 8.4000 175.2000 ;
	    RECT 9.2000 174.3000 10.0000 174.4000 ;
	    RECT 7.6000 173.7000 10.0000 174.3000 ;
	    RECT 16.0000 173.8000 16.8000 174.0000 ;
	    RECT 7.6000 173.6000 8.4000 173.7000 ;
	    RECT 9.2000 173.6000 10.0000 173.7000 ;
	    RECT 15.8000 173.2000 16.8000 173.8000 ;
	    RECT 15.8000 172.4000 16.4000 173.2000 ;
	    RECT 15.6000 171.6000 16.4000 172.4000 ;
	    RECT 9.2000 168.8000 10.0000 170.4000 ;
         LAYER metal2 ;
	    RECT 9.2000 173.6000 10.0000 174.4000 ;
	    RECT 9.3000 170.4000 9.9000 173.6000 ;
	    RECT 15.6000 171.6000 16.4000 172.4000 ;
	    RECT 15.7000 170.4000 16.3000 171.6000 ;
	    RECT 9.2000 169.6000 10.0000 170.4000 ;
	    RECT 15.6000 169.6000 16.4000 170.4000 ;
         LAYER metal3 ;
	    RECT 9.2000 170.3000 10.0000 170.4000 ;
	    RECT 15.6000 170.3000 16.4000 170.4000 ;
	    RECT -3.5000 169.7000 16.4000 170.3000 ;
	    RECT 9.2000 169.6000 10.0000 169.7000 ;
	    RECT 15.6000 169.6000 16.4000 169.7000 ;
      END
   END enable
   PIN ra_adrs[2]
      PORT
         LAYER metal1 ;
	    RECT 89.2000 188.8000 90.0000 190.4000 ;
	    RECT 82.8000 148.8000 83.6000 150.4000 ;
	    RECT 122.8000 52.3000 123.6000 53.2000 ;
	    RECT 124.4000 52.3000 125.2000 53.2000 ;
	    RECT 122.8000 51.7000 125.2000 52.3000 ;
	    RECT 122.8000 51.6000 123.6000 51.7000 ;
	    RECT 124.4000 51.6000 125.2000 51.7000 ;
         LAYER metal2 ;
	    RECT 89.2000 190.3000 90.0000 190.4000 ;
	    RECT 89.2000 189.7000 91.5000 190.3000 ;
	    RECT 89.2000 189.6000 90.0000 189.7000 ;
	    RECT 90.9000 164.3000 91.5000 189.7000 ;
	    RECT 89.3000 163.7000 91.5000 164.3000 ;
	    RECT 82.8000 149.6000 83.6000 150.4000 ;
	    RECT 82.9000 148.4000 83.5000 149.6000 ;
	    RECT 89.3000 148.4000 89.9000 163.7000 ;
	    RECT 82.8000 147.6000 83.6000 148.4000 ;
	    RECT 89.2000 147.6000 90.0000 148.4000 ;
	    RECT 124.4000 65.6000 125.2000 66.4000 ;
	    RECT 124.5000 52.4000 125.1000 65.6000 ;
	    RECT 122.8000 51.6000 123.6000 52.4000 ;
	    RECT 124.4000 51.6000 125.2000 52.4000 ;
	    RECT 122.9000 -2.3000 123.5000 51.6000 ;
         LAYER metal3 ;
	    RECT 82.8000 148.3000 83.6000 148.4000 ;
	    RECT 89.2000 148.3000 90.0000 148.4000 ;
	    RECT 94.0000 148.3000 94.8000 148.4000 ;
	    RECT 82.8000 147.7000 94.8000 148.3000 ;
	    RECT 82.8000 147.6000 83.6000 147.7000 ;
	    RECT 89.2000 147.6000 90.0000 147.7000 ;
	    RECT 94.0000 147.6000 94.8000 147.7000 ;
	    RECT 94.0000 66.3000 94.8000 66.4000 ;
	    RECT 124.4000 66.3000 125.2000 66.4000 ;
	    RECT 94.0000 65.7000 125.2000 66.3000 ;
	    RECT 94.0000 65.6000 94.8000 65.7000 ;
	    RECT 124.4000 65.6000 125.2000 65.7000 ;
         LAYER metal4 ;
	    RECT 93.8000 65.4000 95.0000 148.6000 ;
      END
   END ra_adrs[2]
   PIN ra_adrs[1]
      PORT
         LAYER metal1 ;
	    RECT 178.8000 251.6000 179.6000 253.2000 ;
	    RECT 311.6000 251.6000 312.4000 253.2000 ;
	    RECT 166.0000 211.6000 166.8000 213.2000 ;
	    RECT 222.0000 188.8000 222.8000 190.4000 ;
	    RECT 188.4000 131.6000 189.2000 133.2000 ;
	    RECT 329.2000 108.8000 330.0000 110.4000 ;
	    RECT 210.8000 68.8000 211.6000 70.4000 ;
	    RECT 268.4000 11.6000 269.2000 13.2000 ;
         LAYER metal2 ;
	    RECT 178.8000 251.6000 179.6000 252.4000 ;
	    RECT 311.6000 251.6000 312.4000 252.4000 ;
	    RECT 311.7000 244.4000 312.3000 251.6000 ;
	    RECT 311.6000 243.6000 312.4000 244.4000 ;
	    RECT 335.6000 243.6000 336.4000 244.4000 ;
	    RECT 166.0000 211.6000 166.8000 212.4000 ;
	    RECT 186.8000 211.6000 187.6000 212.4000 ;
	    RECT 186.9000 196.4000 187.5000 211.6000 ;
	    RECT 190.0000 207.6000 190.8000 208.4000 ;
	    RECT 222.0000 207.6000 222.8000 208.4000 ;
	    RECT 190.1000 196.4000 190.7000 207.6000 ;
	    RECT 186.8000 195.6000 187.6000 196.4000 ;
	    RECT 190.0000 195.6000 190.8000 196.4000 ;
	    RECT 186.9000 140.3000 187.5000 195.6000 ;
	    RECT 222.1000 190.4000 222.7000 207.6000 ;
	    RECT 222.0000 189.6000 222.8000 190.4000 ;
	    RECT 335.7000 184.3000 336.3000 243.6000 ;
	    RECT 335.7000 183.7000 337.9000 184.3000 ;
	    RECT 337.3000 156.4000 337.9000 183.7000 ;
	    RECT 337.2000 155.6000 338.0000 156.4000 ;
	    RECT 186.9000 139.7000 189.1000 140.3000 ;
	    RECT 188.5000 134.4000 189.1000 139.7000 ;
	    RECT 188.4000 133.6000 189.2000 134.4000 ;
	    RECT 191.6000 133.6000 192.4000 134.4000 ;
	    RECT 188.5000 132.4000 189.1000 133.6000 ;
	    RECT 188.4000 131.6000 189.2000 132.4000 ;
	    RECT 191.7000 112.3000 192.3000 133.6000 ;
	    RECT 329.2000 123.6000 330.0000 124.4000 ;
	    RECT 191.7000 111.7000 193.9000 112.3000 ;
	    RECT 193.3000 96.3000 193.9000 111.7000 ;
	    RECT 329.3000 110.4000 329.9000 123.6000 ;
	    RECT 329.2000 109.6000 330.0000 110.4000 ;
	    RECT 191.7000 95.7000 193.9000 96.3000 ;
	    RECT 191.7000 68.4000 192.3000 95.7000 ;
	    RECT 329.3000 76.4000 329.9000 109.6000 ;
	    RECT 329.2000 75.6000 330.0000 76.4000 ;
	    RECT 210.8000 69.6000 211.6000 70.4000 ;
	    RECT 210.9000 68.4000 211.5000 69.6000 ;
	    RECT 191.6000 67.6000 192.4000 68.4000 ;
	    RECT 210.8000 67.6000 211.6000 68.4000 ;
	    RECT 268.4000 11.6000 269.2000 12.4000 ;
	    RECT 268.5000 6.4000 269.1000 11.6000 ;
	    RECT 263.6000 5.6000 264.4000 6.4000 ;
	    RECT 268.4000 5.6000 269.2000 6.4000 ;
	    RECT 263.7000 -2.3000 264.3000 5.6000 ;
         LAYER metal3 ;
	    RECT 178.8000 252.3000 179.6000 252.4000 ;
	    RECT 180.4000 252.3000 181.2000 252.4000 ;
	    RECT 178.8000 251.7000 181.2000 252.3000 ;
	    RECT 178.8000 251.6000 179.6000 251.7000 ;
	    RECT 180.4000 251.6000 181.2000 251.7000 ;
	    RECT 311.6000 244.3000 312.4000 244.4000 ;
	    RECT 335.6000 244.3000 336.4000 244.4000 ;
	    RECT 311.6000 243.7000 336.4000 244.3000 ;
	    RECT 311.6000 243.6000 312.4000 243.7000 ;
	    RECT 335.6000 243.6000 336.4000 243.7000 ;
	    RECT 166.0000 212.3000 166.8000 212.4000 ;
	    RECT 180.4000 212.3000 181.2000 212.4000 ;
	    RECT 186.8000 212.3000 187.6000 212.4000 ;
	    RECT 166.0000 211.7000 187.6000 212.3000 ;
	    RECT 166.0000 211.6000 166.8000 211.7000 ;
	    RECT 180.4000 211.6000 181.2000 211.7000 ;
	    RECT 186.8000 211.6000 187.6000 211.7000 ;
	    RECT 190.0000 208.3000 190.8000 208.4000 ;
	    RECT 222.0000 208.3000 222.8000 208.4000 ;
	    RECT 190.0000 207.7000 222.8000 208.3000 ;
	    RECT 190.0000 207.6000 190.8000 207.7000 ;
	    RECT 222.0000 207.6000 222.8000 207.7000 ;
	    RECT 186.8000 196.3000 187.6000 196.4000 ;
	    RECT 190.0000 196.3000 190.8000 196.4000 ;
	    RECT 186.8000 195.7000 190.8000 196.3000 ;
	    RECT 186.8000 195.6000 187.6000 195.7000 ;
	    RECT 190.0000 195.6000 190.8000 195.7000 ;
	    RECT 337.2000 155.6000 338.0000 156.4000 ;
	    RECT 188.4000 134.3000 189.2000 134.4000 ;
	    RECT 191.6000 134.3000 192.4000 134.4000 ;
	    RECT 188.4000 133.7000 192.4000 134.3000 ;
	    RECT 188.4000 133.6000 189.2000 133.7000 ;
	    RECT 191.6000 133.6000 192.4000 133.7000 ;
	    RECT 329.2000 124.3000 330.0000 124.4000 ;
	    RECT 337.2000 124.3000 338.0000 124.4000 ;
	    RECT 329.2000 123.7000 338.0000 124.3000 ;
	    RECT 329.2000 123.6000 330.0000 123.7000 ;
	    RECT 337.2000 123.6000 338.0000 123.7000 ;
	    RECT 324.4000 76.3000 325.2000 76.4000 ;
	    RECT 329.2000 76.3000 330.0000 76.4000 ;
	    RECT 324.4000 75.7000 330.0000 76.3000 ;
	    RECT 324.4000 75.6000 325.2000 75.7000 ;
	    RECT 329.2000 75.6000 330.0000 75.7000 ;
	    RECT 191.6000 68.3000 192.4000 68.4000 ;
	    RECT 210.8000 68.3000 211.6000 68.4000 ;
	    RECT 215.6000 68.3000 216.4000 68.4000 ;
	    RECT 191.6000 67.7000 216.4000 68.3000 ;
	    RECT 191.6000 67.6000 192.4000 67.7000 ;
	    RECT 210.8000 67.6000 211.6000 67.7000 ;
	    RECT 215.6000 67.6000 216.4000 67.7000 ;
	    RECT 215.6000 6.3000 216.4000 6.4000 ;
	    RECT 263.6000 6.3000 264.4000 6.4000 ;
	    RECT 268.4000 6.3000 269.2000 6.4000 ;
	    RECT 321.2000 6.3000 322.0000 6.4000 ;
	    RECT 215.6000 5.7000 322.0000 6.3000 ;
	    RECT 215.6000 5.6000 216.4000 5.7000 ;
	    RECT 263.6000 5.6000 264.4000 5.7000 ;
	    RECT 268.4000 5.6000 269.2000 5.7000 ;
	    RECT 321.2000 5.6000 322.0000 5.7000 ;
         LAYER metal4 ;
	    RECT 180.2000 211.4000 181.4000 252.6000 ;
	    RECT 337.0000 123.4000 338.2000 156.6000 ;
	    RECT 215.4000 5.4000 216.6000 68.6000 ;
	    RECT 324.2000 52.6000 325.4000 76.6000 ;
	    RECT 321.0000 51.4000 325.4000 52.6000 ;
	    RECT 321.0000 5.4000 322.2000 51.4000 ;
      END
   END ra_adrs[1]
   PIN ra_adrs[0]
      PORT
         LAYER metal1 ;
	    RECT 226.8000 310.3000 227.6000 310.4000 ;
	    RECT 228.4000 310.3000 229.2000 310.4000 ;
	    RECT 226.8000 309.7000 229.2000 310.3000 ;
	    RECT 226.8000 309.6000 227.6000 309.7000 ;
	    RECT 228.4000 308.8000 229.2000 309.7000 ;
	    RECT 180.4000 291.6000 181.2000 293.2000 ;
	    RECT 268.4000 251.6000 269.2000 253.2000 ;
	    RECT 276.4000 211.6000 277.2000 213.2000 ;
	    RECT 183.6000 131.6000 184.4000 133.2000 ;
	    RECT 279.6000 131.6000 280.4000 133.2000 ;
	    RECT 279.6000 91.6000 280.4000 93.2000 ;
	    RECT 287.6000 92.3000 288.4000 92.4000 ;
	    RECT 289.2000 92.3000 290.0000 93.2000 ;
	    RECT 287.6000 91.7000 290.0000 92.3000 ;
	    RECT 287.6000 91.6000 288.4000 91.7000 ;
	    RECT 289.2000 91.6000 290.0000 91.7000 ;
         LAYER metal2 ;
	    RECT 225.3000 336.4000 225.9000 346.3000 ;
	    RECT 225.2000 335.6000 226.0000 336.4000 ;
	    RECT 226.8000 309.6000 227.6000 310.4000 ;
	    RECT 226.9000 292.4000 227.5000 309.6000 ;
	    RECT 180.4000 291.6000 181.2000 292.4000 ;
	    RECT 226.8000 291.6000 227.6000 292.4000 ;
	    RECT 180.5000 290.4000 181.1000 291.6000 ;
	    RECT 180.4000 289.6000 181.2000 290.4000 ;
	    RECT 241.2000 261.6000 242.0000 262.4000 ;
	    RECT 241.3000 242.4000 241.9000 261.6000 ;
	    RECT 268.4000 251.6000 269.2000 252.4000 ;
	    RECT 268.5000 242.4000 269.1000 251.6000 ;
	    RECT 241.2000 241.6000 242.0000 242.4000 ;
	    RECT 268.4000 241.6000 269.2000 242.4000 ;
	    RECT 276.4000 241.6000 277.2000 242.4000 ;
	    RECT 276.5000 212.4000 277.1000 241.6000 ;
	    RECT 276.4000 211.6000 277.2000 212.4000 ;
	    RECT 276.5000 176.4000 277.1000 211.6000 ;
	    RECT 276.4000 175.6000 277.2000 176.4000 ;
	    RECT 279.6000 147.6000 280.4000 148.4000 ;
	    RECT 279.7000 132.4000 280.3000 147.6000 ;
	    RECT 183.6000 131.6000 184.4000 132.4000 ;
	    RECT 279.6000 131.6000 280.4000 132.4000 ;
	    RECT 183.7000 130.4000 184.3000 131.6000 ;
	    RECT 279.7000 130.4000 280.3000 131.6000 ;
	    RECT 183.6000 129.6000 184.4000 130.4000 ;
	    RECT 222.0000 129.6000 222.8000 130.4000 ;
	    RECT 246.0000 129.6000 246.8000 130.4000 ;
	    RECT 279.6000 129.6000 280.4000 130.4000 ;
	    RECT 222.1000 120.4000 222.7000 129.6000 ;
	    RECT 246.1000 120.4000 246.7000 129.6000 ;
	    RECT 222.0000 119.6000 222.8000 120.4000 ;
	    RECT 246.0000 119.6000 246.8000 120.4000 ;
	    RECT 279.7000 92.4000 280.3000 129.6000 ;
	    RECT 279.6000 91.6000 280.4000 92.4000 ;
	    RECT 287.6000 91.6000 288.4000 92.4000 ;
         LAYER metal3 ;
	    RECT 225.2000 335.6000 226.0000 336.4000 ;
	    RECT 225.2000 292.3000 226.0000 292.4000 ;
	    RECT 226.8000 292.3000 227.6000 292.4000 ;
	    RECT 225.2000 291.7000 227.6000 292.3000 ;
	    RECT 225.2000 291.6000 226.0000 291.7000 ;
	    RECT 226.8000 291.6000 227.6000 291.7000 ;
	    RECT 180.4000 290.3000 181.2000 290.4000 ;
	    RECT 225.3000 290.3000 225.9000 291.6000 ;
	    RECT 180.4000 289.7000 225.9000 290.3000 ;
	    RECT 180.4000 289.6000 181.2000 289.7000 ;
	    RECT 225.2000 262.3000 226.0000 262.4000 ;
	    RECT 241.2000 262.3000 242.0000 262.4000 ;
	    RECT 225.2000 261.7000 242.0000 262.3000 ;
	    RECT 225.2000 261.6000 226.0000 261.7000 ;
	    RECT 241.2000 261.6000 242.0000 261.7000 ;
	    RECT 241.2000 242.3000 242.0000 242.4000 ;
	    RECT 268.4000 242.3000 269.2000 242.4000 ;
	    RECT 276.4000 242.3000 277.2000 242.4000 ;
	    RECT 241.2000 241.7000 277.2000 242.3000 ;
	    RECT 241.2000 241.6000 242.0000 241.7000 ;
	    RECT 268.4000 241.6000 269.2000 241.7000 ;
	    RECT 276.4000 241.6000 277.2000 241.7000 ;
	    RECT 276.4000 175.6000 277.2000 176.4000 ;
	    RECT 276.4000 148.3000 277.2000 148.4000 ;
	    RECT 279.6000 148.3000 280.4000 148.4000 ;
	    RECT 276.4000 147.7000 280.4000 148.3000 ;
	    RECT 276.4000 147.6000 277.2000 147.7000 ;
	    RECT 279.6000 147.6000 280.4000 147.7000 ;
	    RECT 183.6000 130.3000 184.4000 130.4000 ;
	    RECT 222.0000 130.3000 222.8000 130.4000 ;
	    RECT 183.6000 129.7000 222.8000 130.3000 ;
	    RECT 183.6000 129.6000 184.4000 129.7000 ;
	    RECT 222.0000 129.6000 222.8000 129.7000 ;
	    RECT 246.0000 130.3000 246.8000 130.4000 ;
	    RECT 279.6000 130.3000 280.4000 130.4000 ;
	    RECT 246.0000 129.7000 280.4000 130.3000 ;
	    RECT 246.0000 129.6000 246.8000 129.7000 ;
	    RECT 279.6000 129.6000 280.4000 129.7000 ;
	    RECT 222.0000 120.3000 222.8000 120.4000 ;
	    RECT 246.0000 120.3000 246.8000 120.4000 ;
	    RECT 222.0000 119.7000 246.8000 120.3000 ;
	    RECT 222.0000 119.6000 222.8000 119.7000 ;
	    RECT 246.0000 119.6000 246.8000 119.7000 ;
	    RECT 279.6000 92.3000 280.4000 92.4000 ;
	    RECT 287.6000 92.3000 288.4000 92.4000 ;
	    RECT 279.6000 91.7000 288.4000 92.3000 ;
	    RECT 279.6000 91.6000 280.4000 91.7000 ;
	    RECT 287.6000 91.6000 288.4000 91.7000 ;
         LAYER metal4 ;
	    RECT 225.0000 261.4000 226.2000 336.6000 ;
	    RECT 276.2000 147.4000 277.4000 176.6000 ;
      END
   END ra_adrs[0]
   PIN ra_out[15]
      PORT
         LAYER metal1 ;
	    RECT 28.4000 332.4000 29.2000 339.8000 ;
	    RECT 28.6000 330.2000 29.2000 332.4000 ;
	    RECT 28.4000 322.2000 29.2000 330.2000 ;
         LAYER metal2 ;
	    RECT 26.9000 345.7000 29.1000 346.3000 ;
	    RECT 28.5000 338.4000 29.1000 345.7000 ;
	    RECT 28.4000 337.6000 29.2000 338.4000 ;
      END
   END ra_out[15]
   PIN ra_out[14]
      PORT
         LAYER metal1 ;
	    RECT 137.2000 12.4000 138.0000 19.8000 ;
	    RECT 137.2000 10.2000 137.8000 12.4000 ;
	    RECT 137.2000 2.2000 138.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 137.2000 3.6000 138.0000 4.4000 ;
	    RECT 137.3000 -1.7000 137.9000 3.6000 ;
	    RECT 137.3000 -2.3000 139.5000 -1.7000 ;
      END
   END ra_out[14]
   PIN ra_out[13]
      PORT
         LAYER metal1 ;
	    RECT 78.0000 12.4000 78.8000 19.8000 ;
	    RECT 78.0000 10.2000 78.6000 12.4000 ;
	    RECT 78.0000 2.2000 78.8000 10.2000 ;
         LAYER metal2 ;
	    RECT 78.0000 3.6000 78.8000 4.4000 ;
	    RECT 78.1000 -1.7000 78.7000 3.6000 ;
	    RECT 78.1000 -2.3000 80.3000 -1.7000 ;
      END
   END ra_out[13]
   PIN ra_out[12]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 12.4000 6.8000 19.8000 ;
	    RECT 6.0000 10.2000 6.6000 12.4000 ;
	    RECT 6.0000 2.2000 6.8000 10.2000 ;
         LAYER metal2 ;
	    RECT 6.0000 13.6000 6.8000 14.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 14.3000 6.8000 14.4000 ;
	    RECT -3.5000 13.7000 6.8000 14.3000 ;
	    RECT 6.0000 13.6000 6.8000 13.7000 ;
      END
   END ra_out[12]
   PIN ra_out[11]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 311.8000 2.0000 319.8000 ;
	    RECT 1.2000 309.6000 1.8000 311.8000 ;
	    RECT 1.2000 302.2000 2.0000 309.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 309.6000 2.0000 310.4000 ;
	    RECT 1.3000 308.4000 1.9000 309.6000 ;
	    RECT 1.2000 307.6000 2.0000 308.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 310.3000 2.0000 310.4000 ;
	    RECT -3.5000 309.7000 2.0000 310.3000 ;
	    RECT 1.2000 309.6000 2.0000 309.7000 ;
      END
   END ra_out[11]
   PIN ra_out[10]
      PORT
         LAYER metal1 ;
	    RECT 102.0000 31.8000 102.8000 39.8000 ;
	    RECT 102.0000 29.6000 102.6000 31.8000 ;
	    RECT 102.0000 22.2000 102.8000 29.6000 ;
         LAYER metal2 ;
	    RECT 102.0000 23.6000 102.8000 24.4000 ;
	    RECT 102.1000 14.3000 102.7000 23.6000 ;
	    RECT 102.1000 13.7000 104.3000 14.3000 ;
	    RECT 103.7000 4.4000 104.3000 13.7000 ;
	    RECT 103.6000 3.6000 104.4000 4.4000 ;
	    RECT 113.2000 3.6000 114.0000 4.4000 ;
	    RECT 113.3000 -2.3000 113.9000 3.6000 ;
         LAYER metal3 ;
	    RECT 103.6000 4.3000 104.4000 4.4000 ;
	    RECT 113.2000 4.3000 114.0000 4.4000 ;
	    RECT 103.6000 3.7000 114.0000 4.3000 ;
	    RECT 103.6000 3.6000 104.4000 3.7000 ;
	    RECT 113.2000 3.6000 114.0000 3.7000 ;
      END
   END ra_out[10]
   PIN ra_out[9]
      PORT
         LAYER metal1 ;
	    RECT 47.6000 12.4000 48.4000 19.8000 ;
	    RECT 47.6000 10.2000 48.2000 12.4000 ;
	    RECT 47.6000 2.2000 48.4000 10.2000 ;
         LAYER metal2 ;
	    RECT 47.6000 3.6000 48.4000 4.4000 ;
	    RECT 47.7000 -1.7000 48.3000 3.6000 ;
	    RECT 47.7000 -2.3000 49.9000 -1.7000 ;
      END
   END ra_out[9]
   PIN ra_out[8]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 252.4000 2.0000 259.8000 ;
	    RECT 1.2000 250.2000 1.8000 252.4000 ;
	    RECT 1.2000 242.2000 2.0000 250.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 249.6000 2.0000 250.4000 ;
	    RECT 1.3000 248.4000 1.9000 249.6000 ;
	    RECT 1.2000 247.6000 2.0000 248.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 250.3000 2.0000 250.4000 ;
	    RECT -3.5000 249.7000 2.0000 250.3000 ;
	    RECT 1.2000 249.6000 2.0000 249.7000 ;
      END
   END ra_out[8]
   PIN ra_out[7]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 71.8000 2.0000 79.8000 ;
	    RECT 1.2000 69.6000 1.8000 71.8000 ;
	    RECT 1.2000 62.2000 2.0000 69.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 73.6000 2.0000 74.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 74.3000 2.0000 74.4000 ;
	    RECT -3.5000 73.7000 2.0000 74.3000 ;
	    RECT 1.2000 73.6000 2.0000 73.7000 ;
      END
   END ra_out[7]
   PIN ra_out[6]
      PORT
         LAYER metal1 ;
	    RECT 105.2000 12.4000 106.0000 19.8000 ;
	    RECT 105.4000 10.2000 106.0000 12.4000 ;
	    RECT 105.2000 4.3000 106.0000 10.2000 ;
	    RECT 111.6000 4.3000 112.4000 4.4000 ;
	    RECT 105.2000 3.7000 112.4000 4.3000 ;
	    RECT 105.2000 2.2000 106.0000 3.7000 ;
	    RECT 111.6000 3.6000 112.4000 3.7000 ;
         LAYER metal2 ;
	    RECT 111.6000 3.6000 112.4000 4.4000 ;
	    RECT 111.7000 2.4000 112.3000 3.6000 ;
	    RECT 111.6000 1.6000 112.4000 2.4000 ;
	    RECT 116.4000 1.6000 117.2000 2.4000 ;
	    RECT 116.5000 -2.3000 117.1000 1.6000 ;
         LAYER metal3 ;
	    RECT 111.6000 2.3000 112.4000 2.4000 ;
	    RECT 116.4000 2.3000 117.2000 2.4000 ;
	    RECT 111.6000 1.7000 117.2000 2.3000 ;
	    RECT 111.6000 1.6000 112.4000 1.7000 ;
	    RECT 116.4000 1.6000 117.2000 1.7000 ;
      END
   END ra_out[6]
   PIN ra_out[5]
      PORT
         LAYER metal1 ;
	    RECT 132.4000 12.4000 133.2000 19.8000 ;
	    RECT 132.4000 10.2000 133.0000 12.4000 ;
	    RECT 132.4000 2.2000 133.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 132.4000 3.6000 133.2000 4.4000 ;
	    RECT 132.5000 -1.7000 133.1000 3.6000 ;
	    RECT 132.5000 -2.3000 134.7000 -1.7000 ;
      END
   END ra_out[5]
   PIN ra_out[4]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 231.8000 6.8000 239.8000 ;
	    RECT 6.0000 229.6000 6.6000 231.8000 ;
	    RECT 6.0000 222.2000 6.8000 229.6000 ;
         LAYER metal2 ;
	    RECT 6.0000 233.6000 6.8000 234.4000 ;
	    RECT 6.1000 230.4000 6.7000 233.6000 ;
	    RECT 6.0000 229.6000 6.8000 230.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 230.3000 6.8000 230.4000 ;
	    RECT -3.5000 229.7000 6.8000 230.3000 ;
	    RECT 6.0000 229.6000 6.8000 229.7000 ;
      END
   END ra_out[4]
   PIN ra_out[3]
      PORT
         LAYER metal1 ;
	    RECT 68.4000 31.8000 69.2000 39.8000 ;
	    RECT 68.6000 29.6000 69.2000 31.8000 ;
	    RECT 68.4000 22.2000 69.2000 29.6000 ;
         LAYER metal2 ;
	    RECT 68.4000 23.6000 69.2000 24.4000 ;
	    RECT 68.5000 -1.7000 69.1000 23.6000 ;
	    RECT 66.9000 -2.3000 69.1000 -1.7000 ;
      END
   END ra_out[3]
   PIN ra_out[2]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 191.8000 2.0000 199.8000 ;
	    RECT 1.2000 189.6000 1.8000 191.8000 ;
	    RECT 1.2000 182.2000 2.0000 189.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 189.6000 2.0000 190.4000 ;
	    RECT 1.3000 188.4000 1.9000 189.6000 ;
	    RECT 1.2000 187.6000 2.0000 188.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 190.3000 2.0000 190.4000 ;
	    RECT -3.5000 189.7000 2.0000 190.3000 ;
	    RECT 1.2000 189.6000 2.0000 189.7000 ;
      END
   END ra_out[2]
   PIN ra_out[1]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 151.8000 2.0000 159.8000 ;
	    RECT 1.2000 149.6000 1.8000 151.8000 ;
	    RECT 1.2000 142.2000 2.0000 149.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 149.6000 2.0000 150.4000 ;
	    RECT 1.3000 148.4000 1.9000 149.6000 ;
	    RECT 1.2000 147.6000 2.0000 148.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 150.3000 2.0000 150.4000 ;
	    RECT -3.5000 149.7000 2.0000 150.3000 ;
	    RECT 1.2000 149.6000 2.0000 149.7000 ;
      END
   END ra_out[1]
   PIN ra_out[0]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 111.8000 2.0000 119.8000 ;
	    RECT 1.2000 109.6000 1.8000 111.8000 ;
	    RECT 1.2000 102.2000 2.0000 109.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 109.6000 2.0000 110.4000 ;
	    RECT 1.3000 108.4000 1.9000 109.6000 ;
	    RECT 1.2000 107.6000 2.0000 108.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 110.3000 2.0000 110.4000 ;
	    RECT -3.5000 109.7000 2.0000 110.3000 ;
	    RECT 1.2000 109.6000 2.0000 109.7000 ;
      END
   END ra_out[0]
   PIN rb_adrs[2]
      PORT
         LAYER metal1 ;
	    RECT 71.6000 310.3000 72.4000 310.4000 ;
	    RECT 73.2000 310.3000 74.0000 310.4000 ;
	    RECT 71.6000 309.7000 74.0000 310.3000 ;
	    RECT 71.6000 308.8000 72.4000 309.7000 ;
	    RECT 73.2000 309.6000 74.0000 309.7000 ;
	    RECT 66.8000 211.6000 67.6000 213.2000 ;
	    RECT 76.4000 70.3000 77.2000 70.4000 ;
	    RECT 78.0000 70.3000 78.8000 70.4000 ;
	    RECT 76.4000 69.7000 78.8000 70.3000 ;
	    RECT 76.4000 69.6000 77.2000 69.7000 ;
	    RECT 78.0000 68.8000 78.8000 69.7000 ;
	    RECT 119.6000 68.8000 120.4000 70.4000 ;
         LAYER metal2 ;
	    RECT 70.1000 328.4000 70.7000 346.3000 ;
	    RECT 70.0000 327.6000 70.8000 328.4000 ;
	    RECT 73.2000 327.6000 74.0000 328.4000 ;
	    RECT 73.3000 310.4000 73.9000 327.6000 ;
	    RECT 73.2000 309.6000 74.0000 310.4000 ;
	    RECT 66.8000 215.6000 67.6000 216.4000 ;
	    RECT 66.9000 212.4000 67.5000 215.6000 ;
	    RECT 66.8000 211.6000 67.6000 212.4000 ;
	    RECT 66.9000 176.4000 67.5000 211.6000 ;
	    RECT 66.8000 175.6000 67.6000 176.4000 ;
	    RECT 76.4000 175.6000 77.2000 176.4000 ;
	    RECT 76.5000 70.4000 77.1000 175.6000 ;
	    RECT 76.4000 69.6000 77.2000 70.4000 ;
	    RECT 119.6000 69.6000 120.4000 70.4000 ;
         LAYER metal3 ;
	    RECT 70.0000 328.3000 70.8000 328.4000 ;
	    RECT 73.2000 328.3000 74.0000 328.4000 ;
	    RECT 70.0000 327.7000 74.0000 328.3000 ;
	    RECT 70.0000 327.6000 70.8000 327.7000 ;
	    RECT 73.2000 327.6000 74.0000 327.7000 ;
	    RECT 73.2000 310.3000 74.0000 310.4000 ;
	    RECT 81.2000 310.3000 82.0000 310.4000 ;
	    RECT 73.2000 309.7000 82.0000 310.3000 ;
	    RECT 73.2000 309.6000 74.0000 309.7000 ;
	    RECT 81.2000 309.6000 82.0000 309.7000 ;
	    RECT 66.8000 216.3000 67.6000 216.4000 ;
	    RECT 81.2000 216.3000 82.0000 216.4000 ;
	    RECT 66.8000 215.7000 82.0000 216.3000 ;
	    RECT 66.8000 215.6000 67.6000 215.7000 ;
	    RECT 81.2000 215.6000 82.0000 215.7000 ;
	    RECT 66.8000 176.3000 67.6000 176.4000 ;
	    RECT 76.4000 176.3000 77.2000 176.4000 ;
	    RECT 66.8000 175.7000 77.2000 176.3000 ;
	    RECT 66.8000 175.6000 67.6000 175.7000 ;
	    RECT 76.4000 175.6000 77.2000 175.7000 ;
	    RECT 76.4000 70.3000 77.2000 70.4000 ;
	    RECT 119.6000 70.3000 120.4000 70.4000 ;
	    RECT 76.4000 69.7000 120.4000 70.3000 ;
	    RECT 76.4000 69.6000 77.2000 69.7000 ;
	    RECT 119.6000 69.6000 120.4000 69.7000 ;
         LAYER metal4 ;
	    RECT 81.0000 215.4000 82.2000 310.6000 ;
      END
   END rb_adrs[2]
   PIN rb_adrs[1]
      PORT
         LAYER metal1 ;
	    RECT 191.6000 251.6000 192.4000 253.2000 ;
	    RECT 303.6000 251.6000 304.4000 253.2000 ;
	    RECT 191.6000 211.6000 192.4000 213.2000 ;
	    RECT 220.4000 148.8000 221.2000 150.4000 ;
	    RECT 282.8000 148.8000 283.6000 150.4000 ;
	    RECT 193.2000 131.6000 194.0000 133.2000 ;
	    RECT 244.4000 51.6000 245.2000 53.2000 ;
	    RECT 209.2000 28.8000 210.0000 30.4000 ;
         LAYER metal2 ;
	    RECT 191.6000 251.6000 192.4000 252.4000 ;
	    RECT 303.6000 251.6000 304.4000 252.4000 ;
	    RECT 191.7000 212.4000 192.3000 251.6000 ;
	    RECT 191.6000 211.6000 192.4000 212.4000 ;
	    RECT 209.2000 211.6000 210.0000 212.4000 ;
	    RECT 209.3000 174.4000 209.9000 211.6000 ;
	    RECT 209.2000 173.6000 210.0000 174.4000 ;
	    RECT 220.4000 173.6000 221.2000 174.4000 ;
	    RECT 231.6000 173.6000 232.4000 174.4000 ;
	    RECT 193.2000 133.6000 194.0000 134.4000 ;
	    RECT 193.3000 132.4000 193.9000 133.6000 ;
	    RECT 209.3000 132.4000 209.9000 173.6000 ;
	    RECT 220.5000 150.4000 221.1000 173.6000 ;
	    RECT 231.7000 170.4000 232.3000 173.6000 ;
	    RECT 231.6000 169.6000 232.4000 170.4000 ;
	    RECT 270.0000 169.6000 270.8000 170.4000 ;
	    RECT 270.1000 162.4000 270.7000 169.6000 ;
	    RECT 270.0000 161.6000 270.8000 162.4000 ;
	    RECT 282.8000 161.6000 283.6000 162.4000 ;
	    RECT 282.9000 150.4000 283.5000 161.6000 ;
	    RECT 220.4000 149.6000 221.2000 150.4000 ;
	    RECT 282.8000 149.6000 283.6000 150.4000 ;
	    RECT 193.2000 131.6000 194.0000 132.4000 ;
	    RECT 209.2000 131.6000 210.0000 132.4000 ;
	    RECT 220.5000 114.4000 221.1000 149.6000 ;
	    RECT 220.4000 113.6000 221.2000 114.4000 ;
	    RECT 209.2000 53.6000 210.0000 54.4000 ;
	    RECT 244.4000 53.6000 245.2000 54.4000 ;
	    RECT 209.3000 30.4000 209.9000 53.6000 ;
	    RECT 244.5000 52.4000 245.1000 53.6000 ;
	    RECT 244.4000 51.6000 245.2000 52.4000 ;
	    RECT 209.2000 30.3000 210.0000 30.4000 ;
	    RECT 209.2000 29.7000 211.5000 30.3000 ;
	    RECT 209.2000 29.6000 210.0000 29.7000 ;
	    RECT 210.9000 -2.3000 211.5000 29.7000 ;
         LAYER metal3 ;
	    RECT 303.6000 252.3000 304.4000 252.4000 ;
	    RECT 305.2000 252.3000 306.0000 252.4000 ;
	    RECT 303.6000 251.7000 306.0000 252.3000 ;
	    RECT 303.6000 251.6000 304.4000 251.7000 ;
	    RECT 305.2000 251.6000 306.0000 251.7000 ;
	    RECT 295.6000 220.3000 296.4000 220.4000 ;
	    RECT 305.2000 220.3000 306.0000 220.4000 ;
	    RECT 295.6000 219.7000 306.0000 220.3000 ;
	    RECT 295.6000 219.6000 296.4000 219.7000 ;
	    RECT 305.2000 219.6000 306.0000 219.7000 ;
	    RECT 191.6000 212.3000 192.4000 212.4000 ;
	    RECT 209.2000 212.3000 210.0000 212.4000 ;
	    RECT 191.6000 211.7000 210.0000 212.3000 ;
	    RECT 191.6000 211.6000 192.4000 211.7000 ;
	    RECT 209.2000 211.6000 210.0000 211.7000 ;
	    RECT 295.6000 188.3000 296.4000 188.4000 ;
	    RECT 298.8000 188.3000 299.6000 188.4000 ;
	    RECT 295.6000 187.7000 299.6000 188.3000 ;
	    RECT 295.6000 187.6000 296.4000 187.7000 ;
	    RECT 298.8000 187.6000 299.6000 187.7000 ;
	    RECT 209.2000 174.3000 210.0000 174.4000 ;
	    RECT 220.4000 174.3000 221.2000 174.4000 ;
	    RECT 231.6000 174.3000 232.4000 174.4000 ;
	    RECT 209.2000 173.7000 232.4000 174.3000 ;
	    RECT 209.2000 173.6000 210.0000 173.7000 ;
	    RECT 220.4000 173.6000 221.2000 173.7000 ;
	    RECT 231.6000 173.6000 232.4000 173.7000 ;
	    RECT 231.6000 170.3000 232.4000 170.4000 ;
	    RECT 270.0000 170.3000 270.8000 170.4000 ;
	    RECT 231.6000 169.7000 270.8000 170.3000 ;
	    RECT 231.6000 169.6000 232.4000 169.7000 ;
	    RECT 270.0000 169.6000 270.8000 169.7000 ;
	    RECT 270.0000 162.3000 270.8000 162.4000 ;
	    RECT 282.8000 162.3000 283.6000 162.4000 ;
	    RECT 298.8000 162.3000 299.6000 162.4000 ;
	    RECT 270.0000 161.7000 299.6000 162.3000 ;
	    RECT 270.0000 161.6000 270.8000 161.7000 ;
	    RECT 282.8000 161.6000 283.6000 161.7000 ;
	    RECT 298.8000 161.6000 299.6000 161.7000 ;
	    RECT 193.2000 134.3000 194.0000 134.4000 ;
	    RECT 193.2000 133.7000 198.7000 134.3000 ;
	    RECT 193.2000 133.6000 194.0000 133.7000 ;
	    RECT 198.1000 132.3000 198.7000 133.7000 ;
	    RECT 209.2000 132.3000 210.0000 132.4000 ;
	    RECT 198.1000 131.7000 210.0000 132.3000 ;
	    RECT 209.2000 131.6000 210.0000 131.7000 ;
	    RECT 220.4000 114.3000 221.2000 114.4000 ;
	    RECT 225.2000 114.3000 226.0000 114.4000 ;
	    RECT 220.4000 113.7000 226.0000 114.3000 ;
	    RECT 220.4000 113.6000 221.2000 113.7000 ;
	    RECT 225.2000 113.6000 226.0000 113.7000 ;
	    RECT 209.2000 54.3000 210.0000 54.4000 ;
	    RECT 225.2000 54.3000 226.0000 54.4000 ;
	    RECT 244.4000 54.3000 245.2000 54.4000 ;
	    RECT 209.2000 53.7000 245.2000 54.3000 ;
	    RECT 209.2000 53.6000 210.0000 53.7000 ;
	    RECT 225.2000 53.6000 226.0000 53.7000 ;
	    RECT 244.4000 53.6000 245.2000 53.7000 ;
         LAYER metal4 ;
	    RECT 295.4000 187.4000 296.6000 220.6000 ;
	    RECT 305.0000 219.4000 306.2000 252.6000 ;
	    RECT 298.6000 161.4000 299.8000 188.6000 ;
	    RECT 225.0000 53.4000 226.2000 114.6000 ;
      END
   END rb_adrs[1]
   PIN rb_adrs[0]
      PORT
         LAYER metal1 ;
	    RECT 153.2000 268.8000 154.0000 270.4000 ;
	    RECT 252.4000 268.8000 253.2000 270.4000 ;
	    RECT 174.0000 251.6000 174.8000 253.2000 ;
	    RECT 327.6000 171.6000 328.4000 173.2000 ;
	    RECT 230.0000 148.8000 230.8000 150.4000 ;
	    RECT 159.6000 131.6000 160.4000 133.2000 ;
	    RECT 327.6000 108.8000 328.4000 110.4000 ;
	    RECT 327.6000 91.6000 328.4000 93.2000 ;
         LAYER metal2 ;
	    RECT 262.1000 345.7000 264.3000 346.3000 ;
	    RECT 262.1000 338.3000 262.7000 345.7000 ;
	    RECT 258.9000 337.7000 262.7000 338.3000 ;
	    RECT 258.9000 328.4000 259.5000 337.7000 ;
	    RECT 258.8000 327.6000 259.6000 328.4000 ;
	    RECT 153.2000 269.6000 154.0000 270.4000 ;
	    RECT 252.4000 269.6000 253.2000 270.4000 ;
	    RECT 153.3000 268.4000 153.9000 269.6000 ;
	    RECT 252.5000 268.4000 253.1000 269.6000 ;
	    RECT 153.2000 267.6000 154.0000 268.4000 ;
	    RECT 174.0000 267.6000 174.8000 268.4000 ;
	    RECT 252.4000 267.6000 253.2000 268.4000 ;
	    RECT 174.1000 252.4000 174.7000 267.6000 ;
	    RECT 174.0000 251.6000 174.8000 252.4000 ;
	    RECT 327.6000 171.6000 328.4000 172.4000 ;
	    RECT 230.0000 149.6000 230.8000 150.4000 ;
	    RECT 159.6000 131.6000 160.4000 132.4000 ;
	    RECT 159.7000 128.4000 160.3000 131.6000 ;
	    RECT 230.1000 128.4000 230.7000 149.6000 ;
	    RECT 159.6000 127.6000 160.4000 128.4000 ;
	    RECT 230.0000 127.6000 230.8000 128.4000 ;
	    RECT 327.6000 109.6000 328.4000 110.4000 ;
	    RECT 327.7000 92.4000 328.3000 109.6000 ;
	    RECT 327.6000 91.6000 328.4000 92.4000 ;
         LAYER metal3 ;
	    RECT 247.6000 328.3000 248.4000 328.4000 ;
	    RECT 258.8000 328.3000 259.6000 328.4000 ;
	    RECT 247.6000 327.7000 259.6000 328.3000 ;
	    RECT 247.6000 327.6000 248.4000 327.7000 ;
	    RECT 258.8000 327.6000 259.6000 327.7000 ;
	    RECT 153.2000 268.3000 154.0000 268.4000 ;
	    RECT 174.0000 268.3000 174.8000 268.4000 ;
	    RECT 247.6000 268.3000 248.4000 268.4000 ;
	    RECT 252.4000 268.3000 253.2000 268.4000 ;
	    RECT 153.2000 267.7000 253.2000 268.3000 ;
	    RECT 153.2000 267.6000 154.0000 267.7000 ;
	    RECT 174.0000 267.6000 174.8000 267.7000 ;
	    RECT 247.6000 267.6000 248.4000 267.7000 ;
	    RECT 252.4000 267.6000 253.2000 267.7000 ;
	    RECT 247.6000 172.3000 248.4000 172.4000 ;
	    RECT 327.6000 172.3000 328.4000 172.4000 ;
	    RECT 247.6000 171.7000 328.4000 172.3000 ;
	    RECT 247.6000 171.6000 248.4000 171.7000 ;
	    RECT 327.6000 171.6000 328.4000 171.7000 ;
	    RECT 230.0000 150.3000 230.8000 150.4000 ;
	    RECT 247.6000 150.3000 248.4000 150.4000 ;
	    RECT 230.0000 149.7000 248.4000 150.3000 ;
	    RECT 230.0000 149.6000 230.8000 149.7000 ;
	    RECT 247.6000 149.6000 248.4000 149.7000 ;
	    RECT 159.6000 128.3000 160.4000 128.4000 ;
	    RECT 230.0000 128.3000 230.8000 128.4000 ;
	    RECT 159.6000 127.7000 230.8000 128.3000 ;
	    RECT 159.6000 127.6000 160.4000 127.7000 ;
	    RECT 230.0000 127.6000 230.8000 127.7000 ;
	    RECT 327.6000 109.6000 328.4000 110.4000 ;
         LAYER metal4 ;
	    RECT 247.4000 149.4000 248.6000 328.6000 ;
	    RECT 327.4000 109.4000 328.6000 172.6000 ;
      END
   END rb_adrs[0]
   PIN rb_out[15]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 311.8000 6.8000 319.8000 ;
	    RECT 6.0000 309.6000 6.6000 311.8000 ;
	    RECT 6.0000 302.2000 6.8000 309.6000 ;
         LAYER metal2 ;
	    RECT 6.0000 313.6000 6.8000 314.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 314.3000 6.8000 314.4000 ;
	    RECT -3.5000 313.7000 6.8000 314.3000 ;
	    RECT 6.0000 313.6000 6.8000 313.7000 ;
      END
   END rb_out[15]
   PIN rb_out[14]
      PORT
         LAYER metal1 ;
	    RECT 188.4000 12.4000 189.2000 19.8000 ;
	    RECT 188.6000 10.2000 189.2000 12.4000 ;
	    RECT 188.4000 2.2000 189.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 188.4000 3.6000 189.2000 4.4000 ;
	    RECT 188.5000 -1.7000 189.1000 3.6000 ;
	    RECT 186.9000 -2.3000 189.1000 -1.7000 ;
      END
   END rb_out[14]
   PIN rb_out[13]
      PORT
         LAYER metal1 ;
	    RECT 36.4000 12.4000 37.2000 19.8000 ;
	    RECT 36.4000 10.2000 37.0000 12.4000 ;
	    RECT 36.4000 2.2000 37.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 36.4000 3.6000 37.2000 4.4000 ;
	    RECT 36.5000 -1.7000 37.1000 3.6000 ;
	    RECT 36.5000 -2.3000 38.7000 -1.7000 ;
      END
   END rb_out[13]
   PIN rb_out[12]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 12.4000 2.0000 19.8000 ;
	    RECT 1.2000 10.2000 1.8000 12.4000 ;
	    RECT 1.2000 2.2000 2.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 9.6000 2.0000 10.4000 ;
	    RECT 1.3000 8.4000 1.9000 9.6000 ;
	    RECT 1.2000 7.6000 2.0000 8.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 10.3000 2.0000 10.4000 ;
	    RECT -3.5000 9.7000 2.0000 10.3000 ;
	    RECT 1.2000 9.6000 2.0000 9.7000 ;
      END
   END rb_out[12]
   PIN rb_out[11]
      PORT
         LAYER metal1 ;
	    RECT 20.4000 332.4000 21.2000 339.8000 ;
	    RECT 20.4000 330.2000 21.0000 332.4000 ;
	    RECT 20.4000 322.2000 21.2000 330.2000 ;
         LAYER metal2 ;
	    RECT 20.5000 345.7000 22.7000 346.3000 ;
	    RECT 20.5000 338.4000 21.1000 345.7000 ;
	    RECT 20.4000 337.6000 21.2000 338.4000 ;
      END
   END rb_out[11]
   PIN rb_out[10]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 92.4000 2.0000 99.8000 ;
	    RECT 1.2000 90.2000 1.8000 92.4000 ;
	    RECT 1.2000 82.2000 2.0000 90.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 89.6000 2.0000 90.4000 ;
	    RECT 1.3000 88.4000 1.9000 89.6000 ;
	    RECT 1.2000 87.6000 2.0000 88.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 90.3000 2.0000 90.4000 ;
	    RECT -3.5000 89.7000 2.0000 90.3000 ;
	    RECT 1.2000 89.6000 2.0000 89.7000 ;
      END
   END rb_out[10]
   PIN rb_out[9]
      PORT
         LAYER metal1 ;
	    RECT 161.2000 12.4000 162.0000 19.8000 ;
	    RECT 161.2000 10.2000 161.8000 12.4000 ;
	    RECT 161.2000 2.2000 162.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 161.2000 3.6000 162.0000 4.4000 ;
	    RECT 161.3000 -1.7000 161.9000 3.6000 ;
	    RECT 161.3000 -2.3000 163.5000 -1.7000 ;
      END
   END rb_out[9]
   PIN rb_out[8]
      PORT
         LAYER metal1 ;
	    RECT 42.8000 332.4000 43.6000 339.8000 ;
	    RECT 42.8000 330.2000 43.4000 332.4000 ;
	    RECT 42.8000 322.2000 43.6000 330.2000 ;
         LAYER metal2 ;
	    RECT 42.9000 345.7000 45.1000 346.3000 ;
	    RECT 42.9000 338.4000 43.5000 345.7000 ;
	    RECT 42.8000 337.6000 43.6000 338.4000 ;
      END
   END rb_out[8]
   PIN rb_out[7]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 132.4000 2.0000 139.8000 ;
	    RECT 1.2000 130.2000 1.8000 132.4000 ;
	    RECT 1.2000 122.2000 2.0000 130.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 133.6000 2.0000 134.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 134.3000 2.0000 134.4000 ;
	    RECT -3.5000 133.7000 2.0000 134.3000 ;
	    RECT 1.2000 133.6000 2.0000 133.7000 ;
      END
   END rb_out[7]
   PIN rb_out[6]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 52.4000 2.0000 59.8000 ;
	    RECT 1.2000 50.2000 1.8000 52.4000 ;
	    RECT 1.2000 42.2000 2.0000 50.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 49.6000 2.0000 50.4000 ;
	    RECT 1.3000 48.4000 1.9000 49.6000 ;
	    RECT 1.2000 47.6000 2.0000 48.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 50.3000 2.0000 50.4000 ;
	    RECT -3.5000 49.7000 2.0000 50.3000 ;
	    RECT 1.2000 49.6000 2.0000 49.7000 ;
      END
   END rb_out[6]
   PIN rb_out[5]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 271.8000 2.0000 279.8000 ;
	    RECT 1.2000 269.6000 1.8000 271.8000 ;
	    RECT 1.2000 262.2000 2.0000 269.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 269.6000 2.0000 270.4000 ;
	    RECT 1.3000 268.4000 1.9000 269.6000 ;
	    RECT 1.2000 267.6000 2.0000 268.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 270.3000 2.0000 270.4000 ;
	    RECT -3.5000 269.7000 2.0000 270.3000 ;
	    RECT 1.2000 269.6000 2.0000 269.7000 ;
      END
   END rb_out[5]
   PIN rb_out[4]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 252.4000 6.8000 259.8000 ;
	    RECT 6.0000 250.2000 6.6000 252.4000 ;
	    RECT 6.0000 242.2000 6.8000 250.2000 ;
         LAYER metal2 ;
	    RECT 6.0000 253.6000 6.8000 254.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 254.3000 6.8000 254.4000 ;
	    RECT -3.5000 253.7000 6.8000 254.3000 ;
	    RECT 6.0000 253.6000 6.8000 253.7000 ;
      END
   END rb_out[4]
   PIN rb_out[3]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 132.4000 6.8000 139.8000 ;
	    RECT 6.0000 130.2000 6.6000 132.4000 ;
	    RECT 6.0000 122.2000 6.8000 130.2000 ;
         LAYER metal2 ;
	    RECT 6.0000 133.6000 6.8000 134.4000 ;
	    RECT 6.1000 130.4000 6.7000 133.6000 ;
	    RECT 6.0000 129.6000 6.8000 130.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 130.3000 6.8000 130.4000 ;
	    RECT -3.5000 129.7000 6.8000 130.3000 ;
	    RECT 6.0000 129.6000 6.8000 129.7000 ;
      END
   END rb_out[3]
   PIN rb_out[2]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 212.4000 2.0000 219.8000 ;
	    RECT 1.2000 210.2000 1.8000 212.4000 ;
	    RECT 1.2000 202.2000 2.0000 210.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 209.6000 2.0000 210.4000 ;
	    RECT 1.3000 208.4000 1.9000 209.6000 ;
	    RECT 1.2000 207.6000 2.0000 208.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 210.3000 2.0000 210.4000 ;
	    RECT -3.5000 209.7000 2.0000 210.3000 ;
	    RECT 1.2000 209.6000 2.0000 209.7000 ;
      END
   END rb_out[2]
   PIN rb_out[1]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 231.8000 2.0000 239.8000 ;
	    RECT 1.2000 229.6000 1.8000 231.8000 ;
	    RECT 1.2000 222.2000 2.0000 229.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 233.6000 2.0000 234.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 234.3000 2.0000 234.4000 ;
	    RECT -3.5000 233.7000 2.0000 234.3000 ;
	    RECT 1.2000 233.6000 2.0000 233.7000 ;
      END
   END rb_out[1]
   PIN rb_out[0]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 92.4000 6.8000 99.8000 ;
	    RECT 6.0000 90.2000 6.6000 92.4000 ;
	    RECT 6.0000 82.2000 6.8000 90.2000 ;
         LAYER metal2 ;
	    RECT 6.0000 93.6000 6.8000 94.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 94.3000 6.8000 94.4000 ;
	    RECT -3.5000 93.7000 6.8000 94.3000 ;
	    RECT 6.0000 93.6000 6.8000 93.7000 ;
      END
   END rb_out[0]
   PIN rd_adrs[2]
      PORT
         LAYER metal1 ;
	    RECT 428.4000 189.6000 429.2000 192.4000 ;
	    RECT 438.0000 186.8000 438.8000 188.4000 ;
	    RECT 442.8000 175.6000 443.6000 177.2000 ;
	    RECT 452.4000 175.6000 453.2000 177.2000 ;
         LAYER metal2 ;
	    RECT 428.4000 189.6000 429.2000 190.4000 ;
	    RECT 428.5000 186.4000 429.1000 189.6000 ;
	    RECT 438.0000 187.6000 438.8000 188.4000 ;
	    RECT 438.1000 186.4000 438.7000 187.6000 ;
	    RECT 428.4000 185.6000 429.2000 186.4000 ;
	    RECT 438.0000 185.6000 438.8000 186.4000 ;
	    RECT 442.8000 185.6000 443.6000 186.4000 ;
	    RECT 442.9000 182.4000 443.5000 185.6000 ;
	    RECT 442.8000 181.6000 443.6000 182.4000 ;
	    RECT 452.4000 181.6000 453.2000 182.4000 ;
	    RECT 442.9000 176.4000 443.5000 181.6000 ;
	    RECT 452.5000 178.4000 453.1000 181.6000 ;
	    RECT 452.4000 177.6000 453.2000 178.4000 ;
	    RECT 452.5000 176.4000 453.1000 177.6000 ;
	    RECT 442.8000 175.6000 443.6000 176.4000 ;
	    RECT 452.4000 175.6000 453.2000 176.4000 ;
         LAYER metal3 ;
	    RECT 428.4000 186.3000 429.2000 186.4000 ;
	    RECT 438.0000 186.3000 438.8000 186.4000 ;
	    RECT 442.8000 186.3000 443.6000 186.4000 ;
	    RECT 428.4000 185.7000 443.6000 186.3000 ;
	    RECT 428.4000 185.6000 429.2000 185.7000 ;
	    RECT 438.0000 185.6000 438.8000 185.7000 ;
	    RECT 442.8000 185.6000 443.6000 185.7000 ;
	    RECT 442.8000 182.3000 443.6000 182.4000 ;
	    RECT 452.4000 182.3000 453.2000 182.4000 ;
	    RECT 442.8000 181.7000 453.2000 182.3000 ;
	    RECT 518.1000 182.3000 518.7000 184.3000 ;
	    RECT 518.1000 181.7000 520.3000 182.3000 ;
	    RECT 442.8000 181.6000 443.6000 181.7000 ;
	    RECT 452.4000 181.6000 453.2000 181.7000 ;
	    RECT 452.4000 178.3000 453.2000 178.4000 ;
	    RECT 519.7000 178.3000 520.3000 181.7000 ;
	    RECT 452.4000 177.7000 520.3000 178.3000 ;
	    RECT 452.4000 177.6000 453.2000 177.7000 ;
      END
   END rd_adrs[2]
   PIN rd_adrs[1]
      PORT
         LAYER metal1 ;
	    RECT 434.8000 191.6000 435.6000 193.2000 ;
	    RECT 430.0000 189.6000 431.6000 190.4000 ;
	    RECT 433.2000 175.6000 434.0000 177.2000 ;
	    RECT 447.6000 176.3000 448.4000 177.2000 ;
	    RECT 449.2000 176.3000 450.0000 176.4000 ;
	    RECT 447.6000 175.7000 450.0000 176.3000 ;
	    RECT 447.6000 175.6000 448.4000 175.7000 ;
	    RECT 449.2000 175.6000 450.0000 175.7000 ;
         LAYER metal2 ;
	    RECT 434.8000 192.3000 435.6000 192.4000 ;
	    RECT 433.3000 191.7000 435.6000 192.3000 ;
	    RECT 430.0000 189.6000 430.8000 190.4000 ;
	    RECT 430.1000 178.4000 430.7000 189.6000 ;
	    RECT 433.3000 178.4000 433.9000 191.7000 ;
	    RECT 434.8000 191.6000 435.6000 191.7000 ;
	    RECT 449.2000 185.6000 450.0000 186.4000 ;
	    RECT 449.3000 178.4000 449.9000 185.6000 ;
	    RECT 513.2000 183.6000 514.0000 184.4000 ;
	    RECT 513.3000 180.4000 513.9000 183.6000 ;
	    RECT 513.2000 179.6000 514.0000 180.4000 ;
	    RECT 430.0000 177.6000 430.8000 178.4000 ;
	    RECT 433.2000 177.6000 434.0000 178.4000 ;
	    RECT 449.2000 177.6000 450.0000 178.4000 ;
	    RECT 433.3000 176.4000 433.9000 177.6000 ;
	    RECT 449.3000 176.4000 449.9000 177.6000 ;
	    RECT 433.2000 175.6000 434.0000 176.4000 ;
	    RECT 449.2000 175.6000 450.0000 176.4000 ;
         LAYER metal3 ;
	    RECT 449.2000 186.3000 450.0000 186.4000 ;
	    RECT 449.2000 185.7000 501.1000 186.3000 ;
	    RECT 449.2000 185.6000 450.0000 185.7000 ;
	    RECT 500.5000 184.3000 501.1000 185.7000 ;
	    RECT 513.2000 184.3000 514.0000 184.4000 ;
	    RECT 500.5000 183.7000 514.0000 184.3000 ;
	    RECT 513.2000 183.6000 514.0000 183.7000 ;
	    RECT 513.2000 180.3000 514.0000 180.4000 ;
	    RECT 513.2000 179.7000 518.7000 180.3000 ;
	    RECT 513.2000 179.6000 514.0000 179.7000 ;
	    RECT 430.0000 178.3000 430.8000 178.4000 ;
	    RECT 433.2000 178.3000 434.0000 178.4000 ;
	    RECT 449.2000 178.3000 450.0000 178.4000 ;
	    RECT 430.0000 177.7000 450.0000 178.3000 ;
	    RECT 430.0000 177.6000 430.8000 177.7000 ;
	    RECT 433.2000 177.6000 434.0000 177.7000 ;
	    RECT 449.2000 177.6000 450.0000 177.7000 ;
      END
   END rd_adrs[1]
   PIN rd_adrs[0]
      PORT
         LAYER metal1 ;
	    RECT 23.6000 175.6000 24.4000 177.2000 ;
	    RECT 23.7000 174.4000 24.3000 175.6000 ;
	    RECT 23.6000 174.3000 24.4000 174.4000 ;
	    RECT 25.2000 174.3000 26.0000 175.2000 ;
	    RECT 23.6000 173.7000 26.0000 174.3000 ;
	    RECT 23.6000 173.6000 24.4000 173.7000 ;
	    RECT 25.2000 173.6000 26.0000 173.7000 ;
         LAYER metal2 ;
	    RECT 23.6000 173.6000 24.4000 174.4000 ;
         LAYER metal3 ;
	    RECT 23.6000 174.3000 24.4000 174.4000 ;
	    RECT -3.5000 173.7000 24.4000 174.3000 ;
	    RECT 23.6000 173.6000 24.4000 173.7000 ;
      END
   END rd_adrs[0]
   PIN wr_en
      PORT
         LAYER metal1 ;
	    RECT 6.0000 211.6000 6.8000 213.2000 ;
	    RECT 10.8000 188.8000 11.6000 190.4000 ;
	    RECT 10.8000 148.8000 11.6000 150.4000 ;
	    RECT 6.0000 68.8000 6.8000 70.4000 ;
	    RECT 10.8000 68.8000 11.6000 70.4000 ;
         LAYER metal2 ;
	    RECT 6.0000 211.6000 6.8000 212.4000 ;
	    RECT 6.1000 210.4000 6.7000 211.6000 ;
	    RECT 6.0000 209.6000 6.8000 210.4000 ;
	    RECT 10.8000 209.6000 11.6000 210.4000 ;
	    RECT 10.9000 190.4000 11.5000 209.6000 ;
	    RECT 10.8000 189.6000 11.6000 190.4000 ;
	    RECT 10.9000 150.4000 11.5000 189.6000 ;
	    RECT 10.8000 149.6000 11.6000 150.4000 ;
	    RECT 10.9000 140.4000 11.5000 149.6000 ;
	    RECT 10.8000 139.6000 11.6000 140.4000 ;
	    RECT 6.0000 69.6000 6.8000 70.4000 ;
	    RECT 10.8000 69.6000 11.6000 70.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 210.3000 6.8000 210.4000 ;
	    RECT 10.8000 210.3000 11.6000 210.4000 ;
	    RECT 6.0000 209.7000 11.6000 210.3000 ;
	    RECT 6.0000 209.6000 6.8000 209.7000 ;
	    RECT 10.8000 209.6000 11.6000 209.7000 ;
	    RECT 1.2000 140.3000 2.0000 140.4000 ;
	    RECT 10.8000 140.3000 11.6000 140.4000 ;
	    RECT 1.2000 139.7000 11.6000 140.3000 ;
	    RECT 1.2000 139.6000 2.0000 139.7000 ;
	    RECT 10.8000 139.6000 11.6000 139.7000 ;
	    RECT 1.2000 70.3000 2.0000 70.4000 ;
	    RECT 6.0000 70.3000 6.8000 70.4000 ;
	    RECT 10.8000 70.3000 11.6000 70.4000 ;
	    RECT -3.5000 69.7000 11.6000 70.3000 ;
	    RECT 1.2000 69.6000 2.0000 69.7000 ;
	    RECT 6.0000 69.6000 6.8000 69.7000 ;
	    RECT 10.8000 69.6000 11.6000 69.7000 ;
         LAYER metal4 ;
	    RECT 1.0000 69.4000 2.2000 140.6000 ;
      END
   END wr_en
   OBS
         LAYER metal1 ;
	    RECT 1.2000 335.4000 2.0000 339.8000 ;
	    RECT 5.4000 338.4000 6.6000 339.8000 ;
	    RECT 5.4000 337.8000 6.8000 338.4000 ;
	    RECT 10.0000 337.8000 10.8000 339.8000 ;
	    RECT 14.4000 338.4000 15.2000 339.8000 ;
	    RECT 14.4000 337.8000 16.4000 338.4000 ;
	    RECT 6.0000 337.0000 6.8000 337.8000 ;
	    RECT 10.2000 337.2000 10.8000 337.8000 ;
	    RECT 10.2000 336.6000 13.0000 337.2000 ;
	    RECT 12.2000 336.4000 13.0000 336.6000 ;
	    RECT 14.0000 336.4000 14.8000 337.2000 ;
	    RECT 15.6000 337.0000 16.4000 337.8000 ;
	    RECT 4.2000 335.4000 5.0000 335.6000 ;
	    RECT 1.2000 334.8000 5.0000 335.4000 ;
	    RECT 1.2000 331.4000 2.0000 334.8000 ;
	    RECT 8.2000 334.2000 9.0000 334.4000 ;
	    RECT 12.4000 334.2000 13.2000 334.4000 ;
	    RECT 14.0000 334.2000 14.6000 336.4000 ;
	    RECT 18.8000 335.0000 19.6000 339.8000 ;
	    RECT 23.6000 335.2000 24.4000 339.8000 ;
	    RECT 22.2000 334.6000 24.4000 335.2000 ;
	    RECT 25.2000 335.2000 26.0000 339.8000 ;
	    RECT 30.0000 335.8000 30.8000 339.8000 ;
	    RECT 31.6000 336.0000 32.4000 339.8000 ;
	    RECT 34.8000 336.0000 35.6000 339.8000 ;
	    RECT 31.6000 335.8000 35.6000 336.0000 ;
	    RECT 25.2000 334.6000 27.4000 335.2000 ;
	    RECT 17.2000 334.2000 18.8000 334.4000 ;
	    RECT 7.8000 333.6000 18.8000 334.2000 ;
	    RECT 6.0000 332.8000 6.8000 333.0000 ;
	    RECT 3.0000 332.2000 6.8000 332.8000 ;
	    RECT 3.0000 332.0000 3.8000 332.2000 ;
	    RECT 4.6000 331.4000 5.4000 331.6000 ;
	    RECT 1.2000 330.8000 5.4000 331.4000 ;
	    RECT 1.2000 322.2000 2.0000 330.8000 ;
	    RECT 7.8000 330.4000 8.4000 333.6000 ;
	    RECT 15.0000 333.4000 15.8000 333.6000 ;
	    RECT 14.0000 332.4000 14.8000 332.6000 ;
	    RECT 16.6000 332.4000 17.4000 332.6000 ;
	    RECT 12.4000 331.8000 17.4000 332.4000 ;
	    RECT 12.4000 331.6000 13.2000 331.8000 ;
	    RECT 22.2000 331.6000 22.8000 334.6000 ;
	    RECT 23.6000 331.6000 24.4000 333.2000 ;
	    RECT 25.2000 331.6000 26.0000 333.2000 ;
	    RECT 26.8000 331.6000 27.4000 334.6000 ;
	    RECT 30.2000 334.4000 30.8000 335.8000 ;
	    RECT 31.8000 335.4000 35.4000 335.8000 ;
	    RECT 36.4000 335.6000 37.2000 339.8000 ;
	    RECT 38.0000 336.0000 38.8000 339.8000 ;
	    RECT 41.2000 336.0000 42.0000 339.8000 ;
	    RECT 38.0000 335.8000 42.0000 336.0000 ;
	    RECT 34.0000 334.4000 34.8000 334.8000 ;
	    RECT 36.6000 334.4000 37.2000 335.6000 ;
	    RECT 38.2000 335.4000 41.8000 335.8000 ;
	    RECT 46.0000 335.2000 46.8000 339.8000 ;
	    RECT 47.6000 336.0000 48.4000 339.8000 ;
	    RECT 50.8000 336.0000 51.6000 339.8000 ;
	    RECT 47.6000 335.8000 51.6000 336.0000 ;
	    RECT 52.4000 335.8000 53.2000 339.8000 ;
	    RECT 47.8000 335.4000 51.4000 335.8000 ;
	    RECT 40.4000 334.4000 41.2000 334.8000 ;
	    RECT 44.6000 334.6000 46.8000 335.2000 ;
	    RECT 30.0000 333.6000 32.6000 334.4000 ;
	    RECT 34.0000 333.8000 35.6000 334.4000 ;
	    RECT 34.8000 333.6000 35.6000 333.8000 ;
	    RECT 36.4000 333.6000 39.0000 334.4000 ;
	    RECT 40.4000 333.8000 42.0000 334.4000 ;
	    RECT 41.2000 333.6000 42.0000 333.8000 ;
	    RECT 14.0000 331.0000 19.6000 331.2000 ;
	    RECT 13.8000 330.8000 19.6000 331.0000 ;
	    RECT 21.6000 330.8000 22.8000 331.6000 ;
	    RECT 6.0000 329.8000 8.4000 330.4000 ;
	    RECT 9.8000 330.6000 19.6000 330.8000 ;
	    RECT 9.8000 330.2000 14.6000 330.6000 ;
	    RECT 6.0000 328.8000 6.6000 329.8000 ;
	    RECT 5.2000 328.0000 6.6000 328.8000 ;
	    RECT 8.2000 329.0000 9.0000 329.2000 ;
	    RECT 9.8000 329.0000 10.4000 330.2000 ;
	    RECT 8.2000 328.4000 10.4000 329.0000 ;
	    RECT 11.0000 329.0000 16.4000 329.6000 ;
	    RECT 11.0000 328.8000 11.8000 329.0000 ;
	    RECT 15.6000 328.8000 16.4000 329.0000 ;
	    RECT 9.4000 327.4000 10.2000 327.6000 ;
	    RECT 12.2000 327.4000 13.0000 327.6000 ;
	    RECT 6.0000 326.2000 6.8000 327.0000 ;
	    RECT 9.4000 326.8000 13.0000 327.4000 ;
	    RECT 10.2000 326.2000 10.8000 326.8000 ;
	    RECT 15.6000 326.2000 16.4000 327.0000 ;
	    RECT 5.4000 322.2000 6.6000 326.2000 ;
	    RECT 10.0000 322.2000 10.8000 326.2000 ;
	    RECT 14.4000 325.6000 16.4000 326.2000 ;
	    RECT 14.4000 322.2000 15.2000 325.6000 ;
	    RECT 18.8000 322.2000 19.6000 330.6000 ;
	    RECT 22.2000 330.2000 22.8000 330.8000 ;
	    RECT 26.8000 330.8000 28.0000 331.6000 ;
	    RECT 26.8000 330.2000 27.4000 330.8000 ;
	    RECT 32.0000 330.4000 32.6000 333.6000 ;
	    RECT 33.2000 332.3000 34.0000 333.2000 ;
	    RECT 34.8000 332.3000 35.6000 332.4000 ;
	    RECT 33.2000 331.7000 35.6000 332.3000 ;
	    RECT 33.2000 331.6000 34.0000 331.7000 ;
	    RECT 34.8000 331.6000 35.6000 331.7000 ;
	    RECT 22.2000 329.6000 24.4000 330.2000 ;
	    RECT 23.6000 322.2000 24.4000 329.6000 ;
	    RECT 25.2000 329.6000 27.4000 330.2000 ;
	    RECT 30.0000 330.2000 30.8000 330.4000 ;
	    RECT 30.0000 329.6000 31.4000 330.2000 ;
	    RECT 32.0000 329.6000 34.0000 330.4000 ;
	    RECT 36.4000 330.2000 37.2000 330.4000 ;
	    RECT 38.4000 330.2000 39.0000 333.6000 ;
	    RECT 39.6000 331.6000 40.4000 333.2000 ;
	    RECT 44.6000 331.6000 45.2000 334.6000 ;
	    RECT 48.4000 334.4000 49.2000 334.8000 ;
	    RECT 52.4000 334.4000 53.0000 335.8000 ;
	    RECT 54.0000 335.4000 54.8000 339.8000 ;
	    RECT 58.2000 338.4000 59.4000 339.8000 ;
	    RECT 58.2000 337.8000 59.6000 338.4000 ;
	    RECT 62.8000 337.8000 63.6000 339.8000 ;
	    RECT 67.2000 338.4000 68.0000 339.8000 ;
	    RECT 67.2000 337.8000 69.2000 338.4000 ;
	    RECT 58.8000 337.0000 59.6000 337.8000 ;
	    RECT 63.0000 337.2000 63.6000 337.8000 ;
	    RECT 63.0000 336.6000 65.8000 337.2000 ;
	    RECT 65.0000 336.4000 65.8000 336.6000 ;
	    RECT 66.8000 336.4000 67.6000 337.2000 ;
	    RECT 68.4000 337.0000 69.2000 337.8000 ;
	    RECT 57.0000 335.4000 57.8000 335.6000 ;
	    RECT 54.0000 334.8000 57.8000 335.4000 ;
	    RECT 47.6000 333.8000 49.2000 334.4000 ;
	    RECT 47.6000 333.6000 48.4000 333.8000 ;
	    RECT 50.6000 333.6000 53.2000 334.4000 ;
	    RECT 46.0000 331.6000 46.8000 333.2000 ;
	    RECT 49.2000 331.6000 50.0000 333.2000 ;
	    RECT 50.6000 332.3000 51.2000 333.6000 ;
	    RECT 52.4000 332.3000 53.2000 332.4000 ;
	    RECT 50.6000 331.7000 53.2000 332.3000 ;
	    RECT 44.0000 330.8000 45.2000 331.6000 ;
	    RECT 44.6000 330.2000 45.2000 330.8000 ;
	    RECT 50.6000 330.2000 51.2000 331.7000 ;
	    RECT 52.4000 331.6000 53.2000 331.7000 ;
	    RECT 54.0000 331.4000 54.8000 334.8000 ;
	    RECT 61.0000 334.2000 61.8000 334.4000 ;
	    RECT 66.8000 334.2000 67.4000 336.4000 ;
	    RECT 71.6000 335.0000 72.4000 339.8000 ;
	    RECT 73.2000 335.8000 74.0000 339.8000 ;
	    RECT 74.8000 336.0000 75.6000 339.8000 ;
	    RECT 78.0000 336.0000 78.8000 339.8000 ;
	    RECT 74.8000 335.8000 78.8000 336.0000 ;
	    RECT 73.4000 334.4000 74.0000 335.8000 ;
	    RECT 75.0000 335.4000 78.6000 335.8000 ;
	    RECT 81.2000 335.2000 82.0000 339.8000 ;
	    RECT 84.4000 335.2000 85.2000 339.8000 ;
	    RECT 87.6000 335.2000 88.4000 339.8000 ;
	    RECT 90.8000 335.2000 91.6000 339.8000 ;
	    RECT 77.2000 334.4000 78.0000 334.8000 ;
	    RECT 79.6000 334.4000 82.0000 335.2000 ;
	    RECT 83.0000 334.4000 85.2000 335.2000 ;
	    RECT 86.2000 334.4000 88.4000 335.2000 ;
	    RECT 89.8000 334.4000 91.6000 335.2000 ;
	    RECT 94.0000 335.4000 94.8000 339.8000 ;
	    RECT 98.2000 338.4000 99.4000 339.8000 ;
	    RECT 98.2000 337.8000 99.6000 338.4000 ;
	    RECT 102.8000 337.8000 103.6000 339.8000 ;
	    RECT 107.2000 338.4000 108.0000 339.8000 ;
	    RECT 107.2000 337.8000 109.2000 338.4000 ;
	    RECT 98.8000 337.0000 99.6000 337.8000 ;
	    RECT 103.0000 337.2000 103.6000 337.8000 ;
	    RECT 103.0000 336.6000 105.8000 337.2000 ;
	    RECT 105.0000 336.4000 105.8000 336.6000 ;
	    RECT 106.8000 336.4000 107.6000 337.2000 ;
	    RECT 108.4000 337.0000 109.2000 337.8000 ;
	    RECT 97.0000 335.4000 97.8000 335.6000 ;
	    RECT 94.0000 334.8000 97.8000 335.4000 ;
	    RECT 70.0000 334.2000 71.6000 334.4000 ;
	    RECT 60.6000 333.6000 71.6000 334.2000 ;
	    RECT 73.2000 333.6000 75.8000 334.4000 ;
	    RECT 77.2000 333.8000 78.8000 334.4000 ;
	    RECT 78.0000 333.6000 78.8000 333.8000 ;
	    RECT 58.8000 332.8000 59.6000 333.0000 ;
	    RECT 55.8000 332.2000 59.6000 332.8000 ;
	    RECT 60.6000 332.4000 61.2000 333.6000 ;
	    RECT 67.8000 333.4000 68.6000 333.6000 ;
	    RECT 66.8000 332.4000 67.6000 332.6000 ;
	    RECT 69.4000 332.4000 70.2000 332.6000 ;
	    RECT 55.8000 332.0000 56.6000 332.2000 ;
	    RECT 60.4000 331.6000 61.2000 332.4000 ;
	    RECT 65.2000 331.8000 70.2000 332.4000 ;
	    RECT 65.2000 331.6000 66.0000 331.8000 ;
	    RECT 57.4000 331.4000 58.2000 331.6000 ;
	    RECT 54.0000 330.8000 58.2000 331.4000 ;
	    RECT 52.4000 330.2000 53.2000 330.4000 ;
	    RECT 36.4000 329.6000 37.8000 330.2000 ;
	    RECT 38.4000 329.6000 39.4000 330.2000 ;
	    RECT 44.6000 329.6000 46.8000 330.2000 ;
	    RECT 25.2000 322.2000 26.0000 329.6000 ;
	    RECT 30.8000 328.4000 31.4000 329.6000 ;
	    RECT 30.8000 327.6000 31.6000 328.4000 ;
	    RECT 32.2000 322.2000 33.0000 329.6000 ;
	    RECT 37.2000 328.4000 37.8000 329.6000 ;
	    RECT 37.2000 327.6000 38.0000 328.4000 ;
	    RECT 38.6000 322.2000 39.4000 329.6000 ;
	    RECT 46.0000 322.2000 46.8000 329.6000 ;
	    RECT 50.2000 329.6000 51.2000 330.2000 ;
	    RECT 51.8000 329.6000 53.2000 330.2000 ;
	    RECT 50.2000 322.2000 51.0000 329.6000 ;
	    RECT 51.8000 328.4000 52.4000 329.6000 ;
	    RECT 51.6000 328.3000 52.4000 328.4000 ;
	    RECT 54.0000 328.3000 54.8000 330.8000 ;
	    RECT 60.6000 330.4000 61.2000 331.6000 ;
	    RECT 66.8000 331.0000 72.4000 331.2000 ;
	    RECT 66.6000 330.8000 72.4000 331.0000 ;
	    RECT 58.8000 329.8000 61.2000 330.4000 ;
	    RECT 62.6000 330.6000 72.4000 330.8000 ;
	    RECT 62.6000 330.2000 67.4000 330.6000 ;
	    RECT 58.8000 328.8000 59.4000 329.8000 ;
	    RECT 51.6000 327.7000 54.8000 328.3000 ;
	    RECT 58.0000 328.0000 59.4000 328.8000 ;
	    RECT 61.0000 329.0000 61.8000 329.2000 ;
	    RECT 62.6000 329.0000 63.2000 330.2000 ;
	    RECT 61.0000 328.4000 63.2000 329.0000 ;
	    RECT 63.8000 329.0000 69.2000 329.6000 ;
	    RECT 63.8000 328.8000 64.6000 329.0000 ;
	    RECT 68.4000 328.8000 69.2000 329.0000 ;
	    RECT 51.6000 327.6000 52.4000 327.7000 ;
	    RECT 54.0000 322.2000 54.8000 327.7000 ;
	    RECT 62.2000 327.4000 63.0000 327.6000 ;
	    RECT 65.0000 327.4000 65.8000 327.6000 ;
	    RECT 58.8000 326.2000 59.6000 327.0000 ;
	    RECT 62.2000 326.8000 65.8000 327.4000 ;
	    RECT 63.0000 326.2000 63.6000 326.8000 ;
	    RECT 68.4000 326.2000 69.2000 327.0000 ;
	    RECT 58.2000 322.2000 59.4000 326.2000 ;
	    RECT 62.8000 322.2000 63.6000 326.2000 ;
	    RECT 67.2000 325.6000 69.2000 326.2000 ;
	    RECT 67.2000 322.2000 68.0000 325.6000 ;
	    RECT 71.6000 322.2000 72.4000 330.6000 ;
	    RECT 73.2000 330.2000 74.0000 330.4000 ;
	    RECT 75.2000 330.2000 75.8000 333.6000 ;
	    RECT 76.4000 331.6000 77.2000 333.2000 ;
	    RECT 79.6000 331.6000 80.4000 334.4000 ;
	    RECT 83.0000 333.8000 83.8000 334.4000 ;
	    RECT 86.2000 333.8000 87.0000 334.4000 ;
	    RECT 89.8000 333.8000 90.6000 334.4000 ;
	    RECT 81.2000 333.0000 83.8000 333.8000 ;
	    RECT 84.6000 333.0000 87.0000 333.8000 ;
	    RECT 88.0000 333.0000 90.6000 333.8000 ;
	    RECT 83.0000 331.6000 83.8000 333.0000 ;
	    RECT 86.2000 331.6000 87.0000 333.0000 ;
	    RECT 89.8000 331.6000 90.6000 333.0000 ;
	    RECT 79.6000 330.8000 82.0000 331.6000 ;
	    RECT 83.0000 330.8000 85.2000 331.6000 ;
	    RECT 86.2000 330.8000 88.4000 331.6000 ;
	    RECT 89.8000 330.8000 91.6000 331.6000 ;
	    RECT 73.2000 329.6000 74.6000 330.2000 ;
	    RECT 75.2000 329.6000 76.2000 330.2000 ;
	    RECT 74.0000 328.4000 74.6000 329.6000 ;
	    RECT 74.0000 327.6000 74.8000 328.4000 ;
	    RECT 75.4000 322.2000 76.2000 329.6000 ;
	    RECT 81.2000 322.2000 82.0000 330.8000 ;
	    RECT 84.4000 322.2000 85.2000 330.8000 ;
	    RECT 87.6000 322.2000 88.4000 330.8000 ;
	    RECT 90.8000 322.2000 91.6000 330.8000 ;
	    RECT 94.0000 331.4000 94.8000 334.8000 ;
	    RECT 101.0000 334.2000 101.8000 334.4000 ;
	    RECT 106.8000 334.2000 107.4000 336.4000 ;
	    RECT 111.6000 335.0000 112.4000 339.8000 ;
	    RECT 122.2000 336.4000 123.0000 339.8000 ;
	    RECT 121.2000 335.8000 123.0000 336.4000 ;
	    RECT 124.4000 335.8000 125.2000 339.8000 ;
	    RECT 126.0000 336.0000 126.8000 339.8000 ;
	    RECT 129.2000 336.0000 130.0000 339.8000 ;
	    RECT 126.0000 335.8000 130.0000 336.0000 ;
	    RECT 110.0000 334.2000 111.6000 334.4000 ;
	    RECT 100.6000 333.6000 111.6000 334.2000 ;
	    RECT 116.4000 334.3000 117.2000 334.4000 ;
	    RECT 119.6000 334.3000 120.4000 335.2000 ;
	    RECT 116.4000 333.7000 120.4000 334.3000 ;
	    RECT 116.4000 333.6000 117.2000 333.7000 ;
	    RECT 119.6000 333.6000 120.4000 333.7000 ;
	    RECT 98.8000 332.8000 99.6000 333.0000 ;
	    RECT 95.8000 332.2000 99.6000 332.8000 ;
	    RECT 100.6000 332.4000 101.2000 333.6000 ;
	    RECT 107.8000 333.4000 108.6000 333.6000 ;
	    RECT 106.8000 332.4000 107.6000 332.6000 ;
	    RECT 109.4000 332.4000 110.2000 332.6000 ;
	    RECT 95.8000 332.0000 96.6000 332.2000 ;
	    RECT 100.4000 331.6000 101.2000 332.4000 ;
	    RECT 105.2000 331.8000 110.2000 332.4000 ;
	    RECT 121.2000 332.3000 122.0000 335.8000 ;
	    RECT 124.6000 334.4000 125.2000 335.8000 ;
	    RECT 126.2000 335.4000 129.8000 335.8000 ;
	    RECT 130.8000 335.4000 131.6000 339.8000 ;
	    RECT 135.0000 338.4000 136.2000 339.8000 ;
	    RECT 135.0000 337.8000 136.4000 338.4000 ;
	    RECT 139.6000 337.8000 140.4000 339.8000 ;
	    RECT 144.0000 338.4000 144.8000 339.8000 ;
	    RECT 144.0000 337.8000 146.0000 338.4000 ;
	    RECT 135.6000 337.0000 136.4000 337.8000 ;
	    RECT 139.8000 337.2000 140.4000 337.8000 ;
	    RECT 139.8000 336.6000 142.6000 337.2000 ;
	    RECT 141.8000 336.4000 142.6000 336.6000 ;
	    RECT 143.6000 336.4000 144.4000 337.2000 ;
	    RECT 145.2000 337.0000 146.0000 337.8000 ;
	    RECT 133.8000 335.4000 134.6000 335.6000 ;
	    RECT 130.8000 334.8000 134.6000 335.4000 ;
	    RECT 128.4000 334.4000 129.2000 334.8000 ;
	    RECT 122.8000 334.3000 123.6000 334.4000 ;
	    RECT 124.4000 334.3000 127.0000 334.4000 ;
	    RECT 122.8000 333.7000 127.0000 334.3000 ;
	    RECT 128.4000 333.8000 130.0000 334.4000 ;
	    RECT 122.8000 333.6000 123.6000 333.7000 ;
	    RECT 124.4000 333.6000 127.0000 333.7000 ;
	    RECT 129.2000 333.6000 130.0000 333.8000 ;
	    RECT 105.2000 331.6000 106.0000 331.8000 ;
	    RECT 121.2000 331.7000 125.1000 332.3000 ;
	    RECT 97.4000 331.4000 98.2000 331.6000 ;
	    RECT 94.0000 330.8000 98.2000 331.4000 ;
	    RECT 94.0000 322.2000 94.8000 330.8000 ;
	    RECT 100.6000 330.4000 101.2000 331.6000 ;
	    RECT 106.8000 331.0000 112.4000 331.2000 ;
	    RECT 106.6000 330.8000 112.4000 331.0000 ;
	    RECT 98.8000 329.8000 101.2000 330.4000 ;
	    RECT 102.6000 330.6000 112.4000 330.8000 ;
	    RECT 102.6000 330.2000 107.4000 330.6000 ;
	    RECT 98.8000 328.8000 99.4000 329.8000 ;
	    RECT 98.0000 328.0000 99.4000 328.8000 ;
	    RECT 101.0000 329.0000 101.8000 329.2000 ;
	    RECT 102.6000 329.0000 103.2000 330.2000 ;
	    RECT 101.0000 328.4000 103.2000 329.0000 ;
	    RECT 103.8000 329.0000 109.2000 329.6000 ;
	    RECT 103.8000 328.8000 104.6000 329.0000 ;
	    RECT 108.4000 328.8000 109.2000 329.0000 ;
	    RECT 102.2000 327.4000 103.0000 327.6000 ;
	    RECT 105.0000 327.4000 105.8000 327.6000 ;
	    RECT 98.8000 326.2000 99.6000 327.0000 ;
	    RECT 102.2000 326.8000 105.8000 327.4000 ;
	    RECT 103.0000 326.2000 103.6000 326.8000 ;
	    RECT 108.4000 326.2000 109.2000 327.0000 ;
	    RECT 98.2000 322.2000 99.4000 326.2000 ;
	    RECT 102.8000 322.2000 103.6000 326.2000 ;
	    RECT 107.2000 325.6000 109.2000 326.2000 ;
	    RECT 107.2000 322.2000 108.0000 325.6000 ;
	    RECT 111.6000 322.2000 112.4000 330.6000 ;
	    RECT 121.2000 322.2000 122.0000 331.7000 ;
	    RECT 124.5000 330.4000 125.1000 331.7000 ;
	    RECT 122.8000 328.8000 123.6000 330.4000 ;
	    RECT 124.4000 330.2000 125.2000 330.4000 ;
	    RECT 126.4000 330.2000 127.0000 333.6000 ;
	    RECT 127.6000 331.6000 128.4000 333.2000 ;
	    RECT 130.8000 331.4000 131.6000 334.8000 ;
	    RECT 137.8000 334.2000 138.6000 334.4000 ;
	    RECT 143.6000 334.2000 144.2000 336.4000 ;
	    RECT 148.4000 335.0000 149.2000 339.8000 ;
	    RECT 152.6000 336.4000 153.4000 339.8000 ;
	    RECT 151.6000 335.8000 153.4000 336.4000 ;
	    RECT 154.8000 335.8000 155.6000 339.8000 ;
	    RECT 156.4000 336.0000 157.2000 339.8000 ;
	    RECT 159.6000 336.0000 160.4000 339.8000 ;
	    RECT 156.4000 335.8000 160.4000 336.0000 ;
	    RECT 146.8000 334.2000 148.4000 334.4000 ;
	    RECT 137.4000 333.6000 148.4000 334.2000 ;
	    RECT 150.0000 333.6000 150.8000 335.2000 ;
	    RECT 135.6000 332.8000 136.4000 333.0000 ;
	    RECT 132.6000 332.2000 136.4000 332.8000 ;
	    RECT 137.4000 332.4000 138.0000 333.6000 ;
	    RECT 144.6000 333.4000 145.4000 333.6000 ;
	    RECT 143.6000 332.4000 144.4000 332.6000 ;
	    RECT 146.2000 332.4000 147.0000 332.6000 ;
	    RECT 132.6000 332.0000 133.4000 332.2000 ;
	    RECT 137.2000 331.6000 138.0000 332.4000 ;
	    RECT 142.0000 331.8000 147.0000 332.4000 ;
	    RECT 151.6000 332.3000 152.4000 335.8000 ;
	    RECT 155.0000 334.4000 155.6000 335.8000 ;
	    RECT 156.6000 335.4000 160.2000 335.8000 ;
	    RECT 161.2000 335.4000 162.0000 339.8000 ;
	    RECT 165.4000 338.4000 166.6000 339.8000 ;
	    RECT 165.4000 337.8000 166.8000 338.4000 ;
	    RECT 170.0000 337.8000 170.8000 339.8000 ;
	    RECT 174.4000 338.4000 175.2000 339.8000 ;
	    RECT 174.4000 337.8000 176.4000 338.4000 ;
	    RECT 166.0000 337.0000 166.8000 337.8000 ;
	    RECT 170.2000 337.2000 170.8000 337.8000 ;
	    RECT 170.2000 336.6000 173.0000 337.2000 ;
	    RECT 172.2000 336.4000 173.0000 336.6000 ;
	    RECT 174.0000 336.4000 174.8000 337.2000 ;
	    RECT 175.6000 337.0000 176.4000 337.8000 ;
	    RECT 164.2000 335.4000 165.0000 335.6000 ;
	    RECT 161.2000 334.8000 165.0000 335.4000 ;
	    RECT 158.8000 334.4000 159.6000 334.8000 ;
	    RECT 153.2000 334.3000 154.0000 334.4000 ;
	    RECT 154.8000 334.3000 157.4000 334.4000 ;
	    RECT 153.2000 333.7000 157.4000 334.3000 ;
	    RECT 158.8000 333.8000 160.4000 334.4000 ;
	    RECT 153.2000 333.6000 154.0000 333.7000 ;
	    RECT 154.8000 333.6000 157.4000 333.7000 ;
	    RECT 159.6000 333.6000 160.4000 333.8000 ;
	    RECT 142.0000 331.6000 142.8000 331.8000 ;
	    RECT 151.6000 331.7000 155.5000 332.3000 ;
	    RECT 134.2000 331.4000 135.0000 331.6000 ;
	    RECT 130.8000 330.8000 135.0000 331.4000 ;
	    RECT 124.4000 329.6000 125.8000 330.2000 ;
	    RECT 126.4000 329.6000 127.4000 330.2000 ;
	    RECT 125.2000 328.4000 125.8000 329.6000 ;
	    RECT 125.2000 327.6000 126.0000 328.4000 ;
	    RECT 126.6000 322.2000 127.4000 329.6000 ;
	    RECT 130.8000 322.2000 131.6000 330.8000 ;
	    RECT 134.0000 329.6000 134.8000 330.8000 ;
	    RECT 137.4000 330.4000 138.0000 331.6000 ;
	    RECT 143.6000 331.0000 149.2000 331.2000 ;
	    RECT 143.4000 330.8000 149.2000 331.0000 ;
	    RECT 135.6000 329.8000 138.0000 330.4000 ;
	    RECT 139.4000 330.6000 149.2000 330.8000 ;
	    RECT 139.4000 330.2000 144.2000 330.6000 ;
	    RECT 135.6000 328.8000 136.2000 329.8000 ;
	    RECT 134.8000 328.0000 136.2000 328.8000 ;
	    RECT 137.8000 329.0000 138.6000 329.2000 ;
	    RECT 139.4000 329.0000 140.0000 330.2000 ;
	    RECT 137.8000 328.4000 140.0000 329.0000 ;
	    RECT 140.6000 329.0000 146.0000 329.6000 ;
	    RECT 140.6000 328.8000 141.4000 329.0000 ;
	    RECT 145.2000 328.8000 146.0000 329.0000 ;
	    RECT 139.0000 327.4000 139.8000 327.6000 ;
	    RECT 141.8000 327.4000 142.6000 327.6000 ;
	    RECT 135.6000 326.2000 136.4000 327.0000 ;
	    RECT 139.0000 326.8000 142.6000 327.4000 ;
	    RECT 139.8000 326.2000 140.4000 326.8000 ;
	    RECT 145.2000 326.2000 146.0000 327.0000 ;
	    RECT 135.0000 322.2000 136.2000 326.2000 ;
	    RECT 139.6000 322.2000 140.4000 326.2000 ;
	    RECT 144.0000 325.6000 146.0000 326.2000 ;
	    RECT 144.0000 322.2000 144.8000 325.6000 ;
	    RECT 148.4000 322.2000 149.2000 330.6000 ;
	    RECT 151.6000 322.2000 152.4000 331.7000 ;
	    RECT 154.9000 330.4000 155.5000 331.7000 ;
	    RECT 153.2000 328.8000 154.0000 330.4000 ;
	    RECT 154.8000 330.2000 155.6000 330.4000 ;
	    RECT 156.8000 330.2000 157.4000 333.6000 ;
	    RECT 158.0000 331.6000 158.8000 333.2000 ;
	    RECT 161.2000 331.4000 162.0000 334.8000 ;
	    RECT 168.2000 334.2000 169.0000 334.4000 ;
	    RECT 170.8000 334.2000 171.6000 334.4000 ;
	    RECT 174.0000 334.2000 174.6000 336.4000 ;
	    RECT 178.8000 335.0000 179.6000 339.8000 ;
	    RECT 180.4000 335.8000 181.2000 339.8000 ;
	    RECT 182.0000 336.0000 182.8000 339.8000 ;
	    RECT 185.2000 336.0000 186.0000 339.8000 ;
	    RECT 182.0000 335.8000 186.0000 336.0000 ;
	    RECT 186.8000 335.8000 187.6000 339.8000 ;
	    RECT 188.4000 336.0000 189.2000 339.8000 ;
	    RECT 191.6000 336.0000 192.4000 339.8000 ;
	    RECT 188.4000 335.8000 192.4000 336.0000 ;
	    RECT 180.6000 334.4000 181.2000 335.8000 ;
	    RECT 182.2000 335.4000 185.8000 335.8000 ;
	    RECT 184.4000 334.4000 185.2000 334.8000 ;
	    RECT 187.0000 334.4000 187.6000 335.8000 ;
	    RECT 188.6000 335.4000 192.2000 335.8000 ;
	    RECT 190.8000 334.4000 191.6000 334.8000 ;
	    RECT 177.2000 334.2000 178.8000 334.4000 ;
	    RECT 167.8000 333.6000 178.8000 334.2000 ;
	    RECT 180.4000 333.6000 183.0000 334.4000 ;
	    RECT 184.4000 333.8000 186.0000 334.4000 ;
	    RECT 185.2000 333.6000 186.0000 333.8000 ;
	    RECT 186.8000 333.6000 189.4000 334.4000 ;
	    RECT 190.8000 334.3000 192.4000 334.4000 ;
	    RECT 193.2000 334.3000 194.0000 339.8000 ;
	    RECT 196.4000 335.0000 197.2000 339.8000 ;
	    RECT 200.8000 338.4000 201.6000 339.8000 ;
	    RECT 199.6000 337.8000 201.6000 338.4000 ;
	    RECT 205.2000 337.8000 206.0000 339.8000 ;
	    RECT 209.4000 338.4000 210.6000 339.8000 ;
	    RECT 209.2000 337.8000 210.6000 338.4000 ;
	    RECT 199.6000 337.0000 200.4000 337.8000 ;
	    RECT 205.2000 337.2000 205.8000 337.8000 ;
	    RECT 201.2000 336.4000 202.0000 337.2000 ;
	    RECT 203.0000 336.6000 205.8000 337.2000 ;
	    RECT 209.2000 337.0000 210.0000 337.8000 ;
	    RECT 203.0000 336.4000 203.8000 336.6000 ;
	    RECT 190.8000 333.8000 194.0000 334.3000 ;
	    RECT 191.6000 333.7000 194.0000 333.8000 ;
	    RECT 191.6000 333.6000 192.4000 333.7000 ;
	    RECT 166.0000 332.8000 166.8000 333.0000 ;
	    RECT 163.0000 332.2000 166.8000 332.8000 ;
	    RECT 163.0000 332.0000 163.8000 332.2000 ;
	    RECT 164.6000 331.4000 165.4000 331.6000 ;
	    RECT 161.2000 330.8000 165.4000 331.4000 ;
	    RECT 154.8000 329.6000 156.2000 330.2000 ;
	    RECT 156.8000 329.6000 157.8000 330.2000 ;
	    RECT 155.6000 328.4000 156.2000 329.6000 ;
	    RECT 155.6000 327.6000 156.4000 328.4000 ;
	    RECT 157.0000 322.2000 157.8000 329.6000 ;
	    RECT 161.2000 322.2000 162.0000 330.8000 ;
	    RECT 167.8000 330.4000 168.4000 333.6000 ;
	    RECT 175.0000 333.4000 175.8000 333.6000 ;
	    RECT 174.0000 332.4000 174.8000 332.6000 ;
	    RECT 176.6000 332.4000 177.4000 332.6000 ;
	    RECT 172.4000 331.8000 177.4000 332.4000 ;
	    RECT 172.4000 331.6000 173.2000 331.8000 ;
	    RECT 174.0000 331.0000 179.6000 331.2000 ;
	    RECT 173.8000 330.8000 179.6000 331.0000 ;
	    RECT 166.0000 329.8000 168.4000 330.4000 ;
	    RECT 169.8000 330.6000 179.6000 330.8000 ;
	    RECT 169.8000 330.2000 174.6000 330.6000 ;
	    RECT 166.0000 328.8000 166.6000 329.8000 ;
	    RECT 165.2000 328.0000 166.6000 328.8000 ;
	    RECT 168.2000 329.0000 169.0000 329.2000 ;
	    RECT 169.8000 329.0000 170.4000 330.2000 ;
	    RECT 168.2000 328.4000 170.4000 329.0000 ;
	    RECT 171.0000 329.0000 176.4000 329.6000 ;
	    RECT 171.0000 328.8000 171.8000 329.0000 ;
	    RECT 175.6000 328.8000 176.4000 329.0000 ;
	    RECT 169.4000 327.4000 170.2000 327.6000 ;
	    RECT 172.2000 327.4000 173.0000 327.6000 ;
	    RECT 166.0000 326.2000 166.8000 327.0000 ;
	    RECT 169.4000 326.8000 173.0000 327.4000 ;
	    RECT 170.2000 326.2000 170.8000 326.8000 ;
	    RECT 175.6000 326.2000 176.4000 327.0000 ;
	    RECT 165.4000 322.2000 166.6000 326.2000 ;
	    RECT 170.0000 322.2000 170.8000 326.2000 ;
	    RECT 174.4000 325.6000 176.4000 326.2000 ;
	    RECT 174.4000 322.2000 175.2000 325.6000 ;
	    RECT 178.8000 322.2000 179.6000 330.6000 ;
	    RECT 182.4000 330.4000 183.0000 333.6000 ;
	    RECT 183.6000 331.6000 184.4000 333.2000 ;
	    RECT 180.4000 330.2000 181.2000 330.4000 ;
	    RECT 180.4000 329.6000 181.8000 330.2000 ;
	    RECT 182.4000 329.6000 184.4000 330.4000 ;
	    RECT 186.8000 330.2000 187.6000 330.4000 ;
	    RECT 188.8000 330.2000 189.4000 333.6000 ;
	    RECT 190.0000 331.6000 190.8000 333.2000 ;
	    RECT 186.8000 329.6000 188.2000 330.2000 ;
	    RECT 188.8000 329.6000 189.8000 330.2000 ;
	    RECT 181.2000 328.4000 181.8000 329.6000 ;
	    RECT 180.4000 327.6000 182.0000 328.4000 ;
	    RECT 182.6000 322.2000 183.4000 329.6000 ;
	    RECT 187.6000 328.4000 188.2000 329.6000 ;
	    RECT 187.6000 327.6000 188.4000 328.4000 ;
	    RECT 189.0000 322.2000 189.8000 329.6000 ;
	    RECT 193.2000 322.2000 194.0000 333.7000 ;
	    RECT 197.2000 334.2000 198.8000 334.4000 ;
	    RECT 201.4000 334.2000 202.0000 336.4000 ;
	    RECT 211.0000 335.4000 211.8000 335.6000 ;
	    RECT 214.0000 335.4000 214.8000 339.8000 ;
	    RECT 215.6000 336.0000 216.4000 339.8000 ;
	    RECT 218.8000 336.0000 219.6000 339.8000 ;
	    RECT 215.6000 335.8000 219.6000 336.0000 ;
	    RECT 220.4000 335.8000 221.2000 339.8000 ;
	    RECT 222.0000 335.8000 222.8000 339.8000 ;
	    RECT 223.6000 336.0000 224.4000 339.8000 ;
	    RECT 226.8000 336.0000 227.6000 339.8000 ;
	    RECT 223.6000 335.8000 227.6000 336.0000 ;
	    RECT 215.8000 335.4000 219.4000 335.8000 ;
	    RECT 211.0000 334.8000 214.8000 335.4000 ;
	    RECT 207.0000 334.2000 207.8000 334.4000 ;
	    RECT 197.2000 333.6000 208.2000 334.2000 ;
	    RECT 200.2000 333.4000 201.0000 333.6000 ;
	    RECT 198.6000 332.4000 199.4000 332.6000 ;
	    RECT 207.6000 332.4000 208.2000 333.6000 ;
	    RECT 209.2000 332.8000 210.0000 333.0000 ;
	    RECT 198.6000 331.8000 203.6000 332.4000 ;
	    RECT 202.8000 331.6000 203.6000 331.8000 ;
	    RECT 207.6000 331.6000 208.4000 332.4000 ;
	    RECT 209.2000 332.2000 213.0000 332.8000 ;
	    RECT 212.2000 332.0000 213.0000 332.2000 ;
	    RECT 196.4000 331.0000 202.0000 331.2000 ;
	    RECT 196.4000 330.8000 202.2000 331.0000 ;
	    RECT 196.4000 330.6000 206.2000 330.8000 ;
	    RECT 196.4000 322.2000 197.2000 330.6000 ;
	    RECT 201.4000 330.2000 206.2000 330.6000 ;
	    RECT 199.6000 329.0000 205.0000 329.6000 ;
	    RECT 199.6000 328.8000 200.4000 329.0000 ;
	    RECT 204.2000 328.8000 205.0000 329.0000 ;
	    RECT 205.6000 329.0000 206.2000 330.2000 ;
	    RECT 207.6000 330.4000 208.2000 331.6000 ;
	    RECT 210.6000 331.4000 211.4000 331.6000 ;
	    RECT 214.0000 331.4000 214.8000 334.8000 ;
	    RECT 216.4000 334.4000 217.2000 334.8000 ;
	    RECT 220.4000 334.4000 221.0000 335.8000 ;
	    RECT 222.2000 334.4000 222.8000 335.8000 ;
	    RECT 223.8000 335.4000 227.4000 335.8000 ;
	    RECT 230.0000 335.2000 230.8000 339.8000 ;
	    RECT 233.2000 335.2000 234.0000 339.8000 ;
	    RECT 236.4000 335.2000 237.2000 339.8000 ;
	    RECT 239.6000 335.2000 240.4000 339.8000 ;
	    RECT 242.8000 335.4000 243.6000 339.8000 ;
	    RECT 247.0000 338.4000 248.2000 339.8000 ;
	    RECT 247.0000 337.8000 248.4000 338.4000 ;
	    RECT 251.6000 337.8000 252.4000 339.8000 ;
	    RECT 256.0000 338.4000 256.8000 339.8000 ;
	    RECT 256.0000 337.8000 258.0000 338.4000 ;
	    RECT 247.6000 337.0000 248.4000 337.8000 ;
	    RECT 251.8000 337.2000 252.4000 337.8000 ;
	    RECT 251.8000 336.6000 254.6000 337.2000 ;
	    RECT 253.8000 336.4000 254.6000 336.6000 ;
	    RECT 255.6000 336.4000 256.4000 337.2000 ;
	    RECT 257.2000 337.0000 258.0000 337.8000 ;
	    RECT 245.8000 335.4000 246.6000 335.6000 ;
	    RECT 226.0000 334.4000 226.8000 334.8000 ;
	    RECT 230.0000 334.4000 231.8000 335.2000 ;
	    RECT 233.2000 334.4000 235.4000 335.2000 ;
	    RECT 236.4000 334.4000 238.6000 335.2000 ;
	    RECT 239.6000 334.4000 242.0000 335.2000 ;
	    RECT 215.6000 333.8000 217.2000 334.4000 ;
	    RECT 215.6000 333.6000 216.4000 333.8000 ;
	    RECT 218.6000 333.6000 221.2000 334.4000 ;
	    RECT 222.0000 333.6000 224.6000 334.4000 ;
	    RECT 226.0000 333.8000 227.6000 334.4000 ;
	    RECT 226.8000 333.6000 227.6000 333.8000 ;
	    RECT 231.0000 333.8000 231.8000 334.4000 ;
	    RECT 234.6000 333.8000 235.4000 334.4000 ;
	    RECT 237.8000 333.8000 238.6000 334.4000 ;
	    RECT 217.2000 331.6000 218.0000 333.2000 ;
	    RECT 218.6000 332.3000 219.2000 333.6000 ;
	    RECT 218.6000 331.7000 222.7000 332.3000 ;
	    RECT 210.6000 330.8000 214.8000 331.4000 ;
	    RECT 207.6000 329.8000 210.0000 330.4000 ;
	    RECT 207.0000 329.0000 207.8000 329.2000 ;
	    RECT 205.6000 328.4000 207.8000 329.0000 ;
	    RECT 209.4000 328.8000 210.0000 329.8000 ;
	    RECT 209.4000 328.0000 210.8000 328.8000 ;
	    RECT 203.0000 327.4000 203.8000 327.6000 ;
	    RECT 205.8000 327.4000 206.6000 327.6000 ;
	    RECT 199.6000 326.2000 200.4000 327.0000 ;
	    RECT 203.0000 326.8000 206.6000 327.4000 ;
	    RECT 205.2000 326.2000 205.8000 326.8000 ;
	    RECT 209.2000 326.2000 210.0000 327.0000 ;
	    RECT 199.6000 325.6000 201.6000 326.2000 ;
	    RECT 200.8000 322.2000 201.6000 325.6000 ;
	    RECT 205.2000 322.2000 206.0000 326.2000 ;
	    RECT 209.4000 322.2000 210.6000 326.2000 ;
	    RECT 214.0000 322.2000 214.8000 330.8000 ;
	    RECT 218.6000 330.2000 219.2000 331.7000 ;
	    RECT 222.1000 330.4000 222.7000 331.7000 ;
	    RECT 220.4000 330.2000 221.2000 330.4000 ;
	    RECT 218.2000 329.6000 219.2000 330.2000 ;
	    RECT 219.8000 329.6000 221.2000 330.2000 ;
	    RECT 222.0000 330.2000 222.8000 330.4000 ;
	    RECT 224.0000 330.2000 224.6000 333.6000 ;
	    RECT 225.2000 331.6000 226.0000 333.2000 ;
	    RECT 231.0000 333.0000 233.6000 333.8000 ;
	    RECT 234.6000 333.0000 237.0000 333.8000 ;
	    RECT 237.8000 333.0000 240.4000 333.8000 ;
	    RECT 231.0000 331.6000 231.8000 333.0000 ;
	    RECT 234.6000 331.6000 235.4000 333.0000 ;
	    RECT 237.8000 331.6000 238.6000 333.0000 ;
	    RECT 241.2000 331.6000 242.0000 334.4000 ;
	    RECT 230.0000 330.8000 231.8000 331.6000 ;
	    RECT 233.2000 330.8000 235.4000 331.6000 ;
	    RECT 236.4000 330.8000 238.6000 331.6000 ;
	    RECT 239.6000 330.8000 242.0000 331.6000 ;
	    RECT 242.8000 334.8000 246.6000 335.4000 ;
	    RECT 242.8000 331.4000 243.6000 334.8000 ;
	    RECT 249.8000 334.2000 250.6000 334.4000 ;
	    RECT 255.6000 334.2000 256.2000 336.4000 ;
	    RECT 260.4000 335.0000 261.2000 339.8000 ;
	    RECT 262.0000 336.3000 262.8000 336.4000 ;
	    RECT 268.4000 336.3000 269.2000 337.2000 ;
	    RECT 262.0000 335.7000 269.2000 336.3000 ;
	    RECT 262.0000 335.6000 262.8000 335.7000 ;
	    RECT 268.4000 335.6000 269.2000 335.7000 ;
	    RECT 258.8000 334.2000 260.4000 334.4000 ;
	    RECT 249.4000 333.6000 260.4000 334.2000 ;
	    RECT 270.0000 334.3000 270.8000 339.8000 ;
	    RECT 271.6000 336.0000 272.4000 339.8000 ;
	    RECT 274.8000 336.0000 275.6000 339.8000 ;
	    RECT 271.6000 335.8000 275.6000 336.0000 ;
	    RECT 276.4000 335.8000 277.2000 339.8000 ;
	    RECT 281.8000 336.0000 282.6000 339.0000 ;
	    RECT 286.0000 337.0000 286.8000 339.0000 ;
	    RECT 271.8000 335.4000 275.4000 335.8000 ;
	    RECT 272.4000 334.4000 273.2000 334.8000 ;
	    RECT 276.4000 334.4000 277.0000 335.8000 ;
	    RECT 281.0000 335.4000 282.6000 336.0000 ;
	    RECT 281.0000 335.0000 281.8000 335.4000 ;
	    RECT 281.0000 334.4000 281.6000 335.0000 ;
	    RECT 286.2000 334.8000 286.8000 337.0000 ;
	    RECT 291.4000 336.0000 292.2000 339.0000 ;
	    RECT 295.6000 337.0000 296.4000 339.0000 ;
	    RECT 271.6000 334.3000 273.2000 334.4000 ;
	    RECT 270.0000 333.8000 273.2000 334.3000 ;
	    RECT 270.0000 333.7000 272.4000 333.8000 ;
	    RECT 247.6000 332.8000 248.4000 333.0000 ;
	    RECT 244.6000 332.2000 248.4000 332.8000 ;
	    RECT 249.4000 332.4000 250.0000 333.6000 ;
	    RECT 256.6000 333.4000 257.4000 333.6000 ;
	    RECT 255.6000 332.4000 256.4000 332.6000 ;
	    RECT 258.2000 332.4000 259.0000 332.6000 ;
	    RECT 244.6000 332.0000 245.4000 332.2000 ;
	    RECT 249.2000 331.6000 250.0000 332.4000 ;
	    RECT 254.0000 331.8000 259.0000 332.4000 ;
	    RECT 254.0000 331.6000 254.8000 331.8000 ;
	    RECT 246.2000 331.4000 247.0000 331.6000 ;
	    RECT 242.8000 330.8000 247.0000 331.4000 ;
	    RECT 222.0000 329.6000 223.4000 330.2000 ;
	    RECT 224.0000 329.6000 225.0000 330.2000 ;
	    RECT 218.2000 322.2000 219.0000 329.6000 ;
	    RECT 219.8000 328.4000 220.4000 329.6000 ;
	    RECT 222.8000 328.4000 223.4000 329.6000 ;
	    RECT 219.6000 327.6000 221.2000 328.4000 ;
	    RECT 222.8000 327.6000 223.6000 328.4000 ;
	    RECT 224.2000 322.2000 225.0000 329.6000 ;
	    RECT 230.0000 322.2000 230.8000 330.8000 ;
	    RECT 233.2000 322.2000 234.0000 330.8000 ;
	    RECT 236.4000 322.2000 237.2000 330.8000 ;
	    RECT 239.6000 322.2000 240.4000 330.8000 ;
	    RECT 242.8000 322.2000 243.6000 330.8000 ;
	    RECT 249.4000 330.4000 250.0000 331.6000 ;
	    RECT 255.6000 331.0000 261.2000 331.2000 ;
	    RECT 255.4000 330.8000 261.2000 331.0000 ;
	    RECT 247.6000 329.8000 250.0000 330.4000 ;
	    RECT 251.4000 330.6000 261.2000 330.8000 ;
	    RECT 251.4000 330.2000 256.2000 330.6000 ;
	    RECT 247.6000 328.8000 248.2000 329.8000 ;
	    RECT 246.8000 328.0000 248.2000 328.8000 ;
	    RECT 249.8000 329.0000 250.6000 329.2000 ;
	    RECT 251.4000 329.0000 252.0000 330.2000 ;
	    RECT 249.8000 328.4000 252.0000 329.0000 ;
	    RECT 252.6000 329.0000 258.0000 329.6000 ;
	    RECT 252.6000 328.8000 253.4000 329.0000 ;
	    RECT 257.2000 328.8000 258.0000 329.0000 ;
	    RECT 251.0000 327.4000 251.8000 327.6000 ;
	    RECT 253.8000 327.4000 254.6000 327.6000 ;
	    RECT 247.6000 326.2000 248.4000 327.0000 ;
	    RECT 251.0000 326.8000 254.6000 327.4000 ;
	    RECT 251.8000 326.2000 252.4000 326.8000 ;
	    RECT 257.2000 326.2000 258.0000 327.0000 ;
	    RECT 247.0000 322.2000 248.2000 326.2000 ;
	    RECT 251.6000 322.2000 252.4000 326.2000 ;
	    RECT 256.0000 325.6000 258.0000 326.2000 ;
	    RECT 256.0000 322.2000 256.8000 325.6000 ;
	    RECT 260.4000 322.2000 261.2000 330.6000 ;
	    RECT 270.0000 322.2000 270.8000 333.7000 ;
	    RECT 271.6000 333.6000 272.4000 333.7000 ;
	    RECT 274.6000 333.6000 277.2000 334.4000 ;
	    RECT 279.6000 333.6000 281.6000 334.4000 ;
	    RECT 282.6000 334.2000 286.8000 334.8000 ;
	    RECT 290.6000 335.4000 292.2000 336.0000 ;
	    RECT 290.6000 335.0000 291.4000 335.4000 ;
	    RECT 290.6000 334.4000 291.2000 335.0000 ;
	    RECT 295.8000 334.8000 296.4000 337.0000 ;
	    RECT 282.6000 333.8000 283.6000 334.2000 ;
	    RECT 273.2000 331.6000 274.0000 333.2000 ;
	    RECT 274.6000 330.2000 275.2000 333.6000 ;
	    RECT 278.0000 332.3000 278.8000 332.4000 ;
	    RECT 279.6000 332.3000 280.4000 332.4000 ;
	    RECT 278.0000 331.7000 280.4000 332.3000 ;
	    RECT 278.0000 331.6000 278.8000 331.7000 ;
	    RECT 279.6000 330.8000 280.4000 331.7000 ;
	    RECT 276.4000 330.2000 277.2000 330.4000 ;
	    RECT 274.2000 329.6000 275.2000 330.2000 ;
	    RECT 275.8000 329.6000 277.2000 330.2000 ;
	    RECT 281.0000 329.8000 281.6000 333.6000 ;
	    RECT 282.2000 333.0000 283.6000 333.8000 ;
	    RECT 289.2000 333.6000 291.2000 334.4000 ;
	    RECT 292.2000 334.2000 296.4000 334.8000 ;
	    RECT 297.2000 337.0000 298.0000 339.0000 ;
	    RECT 297.2000 334.8000 297.8000 337.0000 ;
	    RECT 301.4000 336.0000 302.2000 339.0000 ;
	    RECT 306.8000 337.0000 307.6000 339.0000 ;
	    RECT 301.4000 335.4000 303.0000 336.0000 ;
	    RECT 302.2000 335.0000 303.0000 335.4000 ;
	    RECT 297.2000 334.2000 301.4000 334.8000 ;
	    RECT 292.2000 333.8000 293.2000 334.2000 ;
	    RECT 283.0000 331.0000 283.6000 333.0000 ;
	    RECT 284.4000 331.6000 285.2000 333.2000 ;
	    RECT 286.0000 331.6000 286.8000 333.2000 ;
	    RECT 283.0000 330.4000 286.8000 331.0000 ;
	    RECT 289.2000 330.8000 290.0000 332.4000 ;
	    RECT 274.2000 322.2000 275.0000 329.6000 ;
	    RECT 275.8000 328.4000 276.4000 329.6000 ;
	    RECT 281.0000 329.2000 282.6000 329.8000 ;
	    RECT 275.6000 327.6000 276.4000 328.4000 ;
	    RECT 281.8000 322.2000 282.6000 329.2000 ;
	    RECT 286.2000 327.0000 286.8000 330.4000 ;
	    RECT 290.6000 329.8000 291.2000 333.6000 ;
	    RECT 291.8000 333.0000 293.2000 333.8000 ;
	    RECT 300.4000 333.8000 301.4000 334.2000 ;
	    RECT 302.4000 334.4000 303.0000 335.0000 ;
	    RECT 306.8000 334.8000 307.4000 337.0000 ;
	    RECT 311.0000 336.0000 311.8000 339.0000 ;
	    RECT 311.0000 335.4000 312.6000 336.0000 ;
	    RECT 311.8000 335.0000 312.6000 335.4000 ;
	    RECT 292.6000 331.0000 293.2000 333.0000 ;
	    RECT 294.0000 331.6000 294.8000 333.2000 ;
	    RECT 295.6000 331.6000 296.4000 333.2000 ;
	    RECT 297.2000 331.6000 298.0000 333.2000 ;
	    RECT 298.8000 331.6000 299.6000 333.2000 ;
	    RECT 300.4000 333.0000 301.8000 333.8000 ;
	    RECT 302.4000 333.6000 304.4000 334.4000 ;
	    RECT 306.8000 334.2000 311.0000 334.8000 ;
	    RECT 310.0000 333.8000 311.0000 334.2000 ;
	    RECT 312.0000 334.4000 312.6000 335.0000 ;
	    RECT 316.4000 335.4000 317.2000 339.8000 ;
	    RECT 320.6000 338.4000 321.8000 339.8000 ;
	    RECT 320.6000 337.8000 322.0000 338.4000 ;
	    RECT 325.2000 337.8000 326.0000 339.8000 ;
	    RECT 329.6000 338.4000 330.4000 339.8000 ;
	    RECT 329.6000 337.8000 331.6000 338.4000 ;
	    RECT 321.2000 337.0000 322.0000 337.8000 ;
	    RECT 325.4000 337.2000 326.0000 337.8000 ;
	    RECT 325.4000 336.6000 328.2000 337.2000 ;
	    RECT 327.4000 336.4000 328.2000 336.6000 ;
	    RECT 329.2000 336.4000 330.0000 337.2000 ;
	    RECT 330.8000 337.0000 331.6000 337.8000 ;
	    RECT 319.4000 335.4000 320.2000 335.6000 ;
	    RECT 316.4000 334.8000 320.2000 335.4000 ;
	    RECT 300.4000 331.0000 301.0000 333.0000 ;
	    RECT 292.6000 330.4000 296.4000 331.0000 ;
	    RECT 290.6000 329.2000 292.2000 329.8000 ;
	    RECT 286.0000 323.0000 286.8000 327.0000 ;
	    RECT 291.4000 324.4000 292.2000 329.2000 ;
	    RECT 295.8000 327.0000 296.4000 330.4000 ;
	    RECT 290.8000 323.6000 292.2000 324.4000 ;
	    RECT 291.4000 322.2000 292.2000 323.6000 ;
	    RECT 295.6000 323.0000 296.4000 327.0000 ;
	    RECT 297.2000 330.4000 301.0000 331.0000 ;
	    RECT 297.2000 327.0000 297.8000 330.4000 ;
	    RECT 302.4000 329.8000 303.0000 333.6000 ;
	    RECT 303.6000 330.8000 304.4000 332.4000 ;
	    RECT 305.2000 332.3000 306.0000 332.4000 ;
	    RECT 306.8000 332.3000 307.6000 333.2000 ;
	    RECT 305.2000 331.7000 307.6000 332.3000 ;
	    RECT 305.2000 331.6000 306.0000 331.7000 ;
	    RECT 306.8000 331.6000 307.6000 331.7000 ;
	    RECT 308.4000 331.6000 309.2000 333.2000 ;
	    RECT 310.0000 333.0000 311.4000 333.8000 ;
	    RECT 312.0000 333.6000 314.0000 334.4000 ;
	    RECT 310.0000 331.0000 310.6000 333.0000 ;
	    RECT 301.4000 329.2000 303.0000 329.8000 ;
	    RECT 306.8000 330.4000 310.6000 331.0000 ;
	    RECT 297.2000 323.0000 298.0000 327.0000 ;
	    RECT 301.4000 324.4000 302.2000 329.2000 ;
	    RECT 300.4000 323.6000 302.2000 324.4000 ;
	    RECT 301.4000 322.2000 302.2000 323.6000 ;
	    RECT 306.8000 327.0000 307.4000 330.4000 ;
	    RECT 312.0000 329.8000 312.6000 333.6000 ;
	    RECT 313.2000 330.8000 314.0000 332.4000 ;
	    RECT 316.4000 331.4000 317.2000 334.8000 ;
	    RECT 323.4000 334.2000 324.2000 334.4000 ;
	    RECT 329.2000 334.2000 329.8000 336.4000 ;
	    RECT 334.0000 335.0000 334.8000 339.8000 ;
	    RECT 338.2000 336.4000 339.0000 339.8000 ;
	    RECT 337.2000 335.8000 339.0000 336.4000 ;
	    RECT 340.4000 335.8000 341.2000 339.8000 ;
	    RECT 342.0000 336.0000 342.8000 339.8000 ;
	    RECT 345.2000 336.0000 346.0000 339.8000 ;
	    RECT 342.0000 335.8000 346.0000 336.0000 ;
	    RECT 332.4000 334.2000 334.0000 334.4000 ;
	    RECT 323.0000 333.6000 334.0000 334.2000 ;
	    RECT 335.6000 333.6000 336.4000 335.2000 ;
	    RECT 321.2000 332.8000 322.0000 333.0000 ;
	    RECT 318.2000 332.2000 322.0000 332.8000 ;
	    RECT 318.2000 332.0000 319.0000 332.2000 ;
	    RECT 319.8000 331.4000 320.6000 331.6000 ;
	    RECT 316.4000 330.8000 320.6000 331.4000 ;
	    RECT 311.0000 329.2000 312.6000 329.8000 ;
	    RECT 306.8000 323.0000 307.6000 327.0000 ;
	    RECT 311.0000 324.4000 311.8000 329.2000 ;
	    RECT 311.0000 323.6000 312.4000 324.4000 ;
	    RECT 311.0000 322.2000 311.8000 323.6000 ;
	    RECT 316.4000 322.2000 317.2000 330.8000 ;
	    RECT 323.0000 330.4000 323.6000 333.6000 ;
	    RECT 330.2000 333.4000 331.0000 333.6000 ;
	    RECT 329.2000 332.4000 330.0000 332.6000 ;
	    RECT 331.8000 332.4000 332.6000 332.6000 ;
	    RECT 327.6000 331.8000 332.6000 332.4000 ;
	    RECT 337.2000 332.3000 338.0000 335.8000 ;
	    RECT 340.6000 334.4000 341.2000 335.8000 ;
	    RECT 342.2000 335.4000 345.8000 335.8000 ;
	    RECT 346.8000 335.4000 347.6000 339.8000 ;
	    RECT 351.0000 338.4000 352.2000 339.8000 ;
	    RECT 351.0000 337.8000 352.4000 338.4000 ;
	    RECT 355.6000 337.8000 356.4000 339.8000 ;
	    RECT 360.0000 338.4000 360.8000 339.8000 ;
	    RECT 360.0000 337.8000 362.0000 338.4000 ;
	    RECT 351.6000 337.0000 352.4000 337.8000 ;
	    RECT 355.8000 337.2000 356.4000 337.8000 ;
	    RECT 355.8000 336.6000 358.6000 337.2000 ;
	    RECT 357.8000 336.4000 358.6000 336.6000 ;
	    RECT 359.6000 336.4000 360.4000 337.2000 ;
	    RECT 361.2000 337.0000 362.0000 337.8000 ;
	    RECT 349.8000 335.4000 350.6000 335.6000 ;
	    RECT 346.8000 334.8000 350.6000 335.4000 ;
	    RECT 344.4000 334.4000 345.2000 334.8000 ;
	    RECT 340.4000 333.6000 343.0000 334.4000 ;
	    RECT 344.4000 333.8000 346.0000 334.4000 ;
	    RECT 345.2000 333.6000 346.0000 333.8000 ;
	    RECT 327.6000 331.6000 328.4000 331.8000 ;
	    RECT 337.2000 331.7000 341.1000 332.3000 ;
	    RECT 329.2000 331.0000 334.8000 331.2000 ;
	    RECT 329.0000 330.8000 334.8000 331.0000 ;
	    RECT 321.2000 329.8000 323.6000 330.4000 ;
	    RECT 325.0000 330.6000 334.8000 330.8000 ;
	    RECT 325.0000 330.2000 329.8000 330.6000 ;
	    RECT 321.2000 328.8000 321.8000 329.8000 ;
	    RECT 320.4000 328.0000 321.8000 328.8000 ;
	    RECT 323.4000 329.0000 324.2000 329.2000 ;
	    RECT 325.0000 329.0000 325.6000 330.2000 ;
	    RECT 323.4000 328.4000 325.6000 329.0000 ;
	    RECT 326.2000 329.0000 331.6000 329.6000 ;
	    RECT 326.2000 328.8000 327.0000 329.0000 ;
	    RECT 330.8000 328.8000 331.6000 329.0000 ;
	    RECT 324.6000 327.4000 325.4000 327.6000 ;
	    RECT 327.4000 327.4000 328.2000 327.6000 ;
	    RECT 321.2000 326.2000 322.0000 327.0000 ;
	    RECT 324.6000 326.8000 328.2000 327.4000 ;
	    RECT 325.4000 326.2000 326.0000 326.8000 ;
	    RECT 330.8000 326.2000 331.6000 327.0000 ;
	    RECT 320.6000 322.2000 321.8000 326.2000 ;
	    RECT 325.2000 322.2000 326.0000 326.2000 ;
	    RECT 329.6000 325.6000 331.6000 326.2000 ;
	    RECT 329.6000 322.2000 330.4000 325.6000 ;
	    RECT 334.0000 322.2000 334.8000 330.6000 ;
	    RECT 337.2000 322.2000 338.0000 331.7000 ;
	    RECT 340.5000 330.4000 341.1000 331.7000 ;
	    RECT 338.8000 328.8000 339.6000 330.4000 ;
	    RECT 340.4000 330.2000 341.2000 330.4000 ;
	    RECT 342.4000 330.2000 343.0000 333.6000 ;
	    RECT 343.6000 331.6000 344.4000 333.2000 ;
	    RECT 346.8000 331.4000 347.6000 334.8000 ;
	    RECT 353.8000 334.2000 354.6000 334.4000 ;
	    RECT 359.6000 334.2000 360.2000 336.4000 ;
	    RECT 364.4000 335.0000 365.2000 339.8000 ;
	    RECT 362.8000 334.2000 364.4000 334.4000 ;
	    RECT 353.4000 333.6000 364.4000 334.2000 ;
	    RECT 351.6000 332.8000 352.4000 333.0000 ;
	    RECT 348.6000 332.2000 352.4000 332.8000 ;
	    RECT 353.4000 332.4000 354.0000 333.6000 ;
	    RECT 360.6000 333.4000 361.4000 333.6000 ;
	    RECT 362.2000 332.4000 363.0000 332.6000 ;
	    RECT 348.6000 332.0000 349.4000 332.2000 ;
	    RECT 353.2000 331.6000 354.0000 332.4000 ;
	    RECT 358.0000 331.8000 363.0000 332.4000 ;
	    RECT 358.0000 331.6000 358.8000 331.8000 ;
	    RECT 350.2000 331.4000 351.0000 331.6000 ;
	    RECT 346.8000 330.8000 351.0000 331.4000 ;
	    RECT 340.4000 329.6000 341.8000 330.2000 ;
	    RECT 342.4000 329.6000 343.4000 330.2000 ;
	    RECT 341.2000 328.4000 341.8000 329.6000 ;
	    RECT 342.6000 328.4000 343.4000 329.6000 ;
	    RECT 341.2000 327.6000 342.0000 328.4000 ;
	    RECT 342.6000 327.6000 344.4000 328.4000 ;
	    RECT 342.6000 322.2000 343.4000 327.6000 ;
	    RECT 346.8000 322.2000 347.6000 330.8000 ;
	    RECT 353.4000 330.4000 354.0000 331.6000 ;
	    RECT 359.6000 331.0000 365.2000 331.2000 ;
	    RECT 359.4000 330.8000 365.2000 331.0000 ;
	    RECT 351.6000 329.8000 354.0000 330.4000 ;
	    RECT 355.4000 330.6000 365.2000 330.8000 ;
	    RECT 355.4000 330.2000 360.2000 330.6000 ;
	    RECT 351.6000 328.8000 352.2000 329.8000 ;
	    RECT 350.8000 328.0000 352.2000 328.8000 ;
	    RECT 353.8000 329.0000 354.6000 329.2000 ;
	    RECT 355.4000 329.0000 356.0000 330.2000 ;
	    RECT 353.8000 328.4000 356.0000 329.0000 ;
	    RECT 356.6000 329.0000 362.0000 329.6000 ;
	    RECT 356.6000 328.8000 357.4000 329.0000 ;
	    RECT 361.2000 328.8000 362.0000 329.0000 ;
	    RECT 355.0000 327.4000 355.8000 327.6000 ;
	    RECT 357.8000 327.4000 358.6000 327.6000 ;
	    RECT 351.6000 326.2000 352.4000 327.0000 ;
	    RECT 355.0000 326.8000 358.6000 327.4000 ;
	    RECT 355.8000 326.2000 356.4000 326.8000 ;
	    RECT 361.2000 326.2000 362.0000 327.0000 ;
	    RECT 351.0000 322.2000 352.2000 326.2000 ;
	    RECT 355.6000 322.2000 356.4000 326.2000 ;
	    RECT 360.0000 325.6000 362.0000 326.2000 ;
	    RECT 360.0000 322.2000 360.8000 325.6000 ;
	    RECT 364.4000 322.2000 365.2000 330.6000 ;
	    RECT 366.0000 322.2000 366.8000 339.8000 ;
	    RECT 369.2000 335.4000 370.0000 339.8000 ;
	    RECT 373.4000 338.4000 374.6000 339.8000 ;
	    RECT 373.4000 337.8000 374.8000 338.4000 ;
	    RECT 378.0000 337.8000 378.8000 339.8000 ;
	    RECT 382.4000 338.4000 383.2000 339.8000 ;
	    RECT 382.4000 337.8000 384.4000 338.4000 ;
	    RECT 374.0000 337.0000 374.8000 337.8000 ;
	    RECT 378.2000 337.2000 378.8000 337.8000 ;
	    RECT 378.2000 336.6000 381.0000 337.2000 ;
	    RECT 380.2000 336.4000 381.0000 336.6000 ;
	    RECT 382.0000 336.4000 382.8000 337.2000 ;
	    RECT 383.6000 337.0000 384.4000 337.8000 ;
	    RECT 372.2000 335.4000 373.0000 335.6000 ;
	    RECT 369.2000 334.8000 373.0000 335.4000 ;
	    RECT 369.2000 331.4000 370.0000 334.8000 ;
	    RECT 376.2000 334.2000 377.0000 334.4000 ;
	    RECT 378.8000 334.2000 379.6000 334.4000 ;
	    RECT 382.0000 334.2000 382.6000 336.4000 ;
	    RECT 386.8000 335.0000 387.6000 339.8000 ;
	    RECT 388.4000 335.6000 389.2000 337.2000 ;
	    RECT 385.2000 334.2000 386.8000 334.4000 ;
	    RECT 375.8000 333.6000 386.8000 334.2000 ;
	    RECT 390.0000 334.3000 390.8000 339.8000 ;
	    RECT 391.6000 336.0000 392.4000 339.8000 ;
	    RECT 394.8000 336.0000 395.6000 339.8000 ;
	    RECT 391.6000 335.8000 395.6000 336.0000 ;
	    RECT 396.4000 335.8000 397.2000 339.8000 ;
	    RECT 391.8000 335.4000 395.4000 335.8000 ;
	    RECT 392.4000 334.4000 393.2000 334.8000 ;
	    RECT 396.4000 334.4000 397.0000 335.8000 ;
	    RECT 391.6000 334.3000 393.2000 334.4000 ;
	    RECT 390.0000 333.8000 393.2000 334.3000 ;
	    RECT 390.0000 333.7000 392.4000 333.8000 ;
	    RECT 374.0000 332.8000 374.8000 333.0000 ;
	    RECT 371.0000 332.2000 374.8000 332.8000 ;
	    RECT 371.0000 332.0000 371.8000 332.2000 ;
	    RECT 372.6000 331.4000 373.4000 331.6000 ;
	    RECT 369.2000 330.8000 373.4000 331.4000 ;
	    RECT 369.2000 322.2000 370.0000 330.8000 ;
	    RECT 375.8000 330.4000 376.4000 333.6000 ;
	    RECT 383.0000 333.4000 383.8000 333.6000 ;
	    RECT 382.0000 332.4000 382.8000 332.6000 ;
	    RECT 384.6000 332.4000 385.4000 332.6000 ;
	    RECT 380.4000 331.8000 385.4000 332.4000 ;
	    RECT 380.4000 331.6000 381.2000 331.8000 ;
	    RECT 382.0000 331.0000 387.6000 331.2000 ;
	    RECT 381.8000 330.8000 387.6000 331.0000 ;
	    RECT 374.0000 329.8000 376.4000 330.4000 ;
	    RECT 377.8000 330.6000 387.6000 330.8000 ;
	    RECT 377.8000 330.2000 382.6000 330.6000 ;
	    RECT 374.0000 328.8000 374.6000 329.8000 ;
	    RECT 373.2000 328.0000 374.6000 328.8000 ;
	    RECT 376.2000 329.0000 377.0000 329.2000 ;
	    RECT 377.8000 329.0000 378.4000 330.2000 ;
	    RECT 376.2000 328.4000 378.4000 329.0000 ;
	    RECT 379.0000 329.0000 384.4000 329.6000 ;
	    RECT 379.0000 328.8000 379.8000 329.0000 ;
	    RECT 383.6000 328.8000 384.4000 329.0000 ;
	    RECT 377.4000 327.4000 378.2000 327.6000 ;
	    RECT 380.2000 327.4000 381.0000 327.6000 ;
	    RECT 374.0000 326.2000 374.8000 327.0000 ;
	    RECT 377.4000 326.8000 381.0000 327.4000 ;
	    RECT 378.2000 326.2000 378.8000 326.8000 ;
	    RECT 383.6000 326.2000 384.4000 327.0000 ;
	    RECT 373.4000 322.2000 374.6000 326.2000 ;
	    RECT 378.0000 322.2000 378.8000 326.2000 ;
	    RECT 382.4000 325.6000 384.4000 326.2000 ;
	    RECT 382.4000 322.2000 383.2000 325.6000 ;
	    RECT 386.8000 322.2000 387.6000 330.6000 ;
	    RECT 390.0000 322.2000 390.8000 333.7000 ;
	    RECT 391.6000 333.6000 392.4000 333.7000 ;
	    RECT 394.6000 333.6000 397.2000 334.4000 ;
	    RECT 401.6000 334.2000 402.4000 339.8000 ;
	    RECT 414.4000 334.2000 415.2000 339.8000 ;
	    RECT 420.8000 334.2000 421.6000 339.8000 ;
	    RECT 427.2000 334.2000 428.0000 339.8000 ;
	    RECT 430.0000 335.6000 430.8000 337.2000 ;
	    RECT 431.6000 334.3000 432.4000 339.8000 ;
	    RECT 433.2000 336.0000 434.0000 339.8000 ;
	    RECT 436.4000 336.0000 437.2000 339.8000 ;
	    RECT 433.2000 335.8000 437.2000 336.0000 ;
	    RECT 438.0000 335.8000 438.8000 339.8000 ;
	    RECT 433.4000 335.4000 437.0000 335.8000 ;
	    RECT 434.0000 334.4000 434.8000 334.8000 ;
	    RECT 438.0000 334.4000 438.6000 335.8000 ;
	    RECT 439.6000 335.4000 440.4000 339.8000 ;
	    RECT 443.8000 338.4000 445.0000 339.8000 ;
	    RECT 443.8000 337.8000 445.2000 338.4000 ;
	    RECT 448.4000 337.8000 449.2000 339.8000 ;
	    RECT 452.8000 338.4000 453.6000 339.8000 ;
	    RECT 452.8000 337.8000 454.8000 338.4000 ;
	    RECT 444.4000 337.0000 445.2000 337.8000 ;
	    RECT 448.6000 337.2000 449.2000 337.8000 ;
	    RECT 448.6000 336.6000 451.4000 337.2000 ;
	    RECT 450.6000 336.4000 451.4000 336.6000 ;
	    RECT 452.4000 336.4000 453.2000 337.2000 ;
	    RECT 454.0000 337.0000 454.8000 337.8000 ;
	    RECT 442.6000 335.4000 443.4000 335.6000 ;
	    RECT 439.6000 334.8000 443.4000 335.4000 ;
	    RECT 433.2000 334.3000 434.8000 334.4000 ;
	    RECT 401.6000 333.8000 403.4000 334.2000 ;
	    RECT 414.4000 333.8000 416.2000 334.2000 ;
	    RECT 420.8000 333.8000 422.6000 334.2000 ;
	    RECT 427.2000 333.8000 429.0000 334.2000 ;
	    RECT 401.8000 333.6000 403.4000 333.8000 ;
	    RECT 414.6000 333.6000 416.2000 333.8000 ;
	    RECT 421.0000 333.6000 422.6000 333.8000 ;
	    RECT 427.4000 333.6000 429.0000 333.8000 ;
	    RECT 393.2000 331.6000 394.0000 333.2000 ;
	    RECT 394.6000 330.4000 395.2000 333.6000 ;
	    RECT 399.6000 331.6000 401.2000 332.4000 ;
	    RECT 402.8000 330.4000 403.4000 333.6000 ;
	    RECT 412.4000 331.6000 414.0000 332.4000 ;
	    RECT 415.6000 330.4000 416.2000 333.6000 ;
	    RECT 418.8000 331.6000 420.4000 332.4000 ;
	    RECT 422.0000 330.4000 422.6000 333.6000 ;
	    RECT 425.2000 331.6000 426.8000 332.4000 ;
	    RECT 428.4000 330.4000 429.0000 333.6000 ;
	    RECT 431.6000 333.8000 434.8000 334.3000 ;
	    RECT 431.6000 333.7000 434.0000 333.8000 ;
	    RECT 393.2000 329.6000 395.2000 330.4000 ;
	    RECT 396.4000 330.2000 397.2000 330.4000 ;
	    RECT 395.8000 329.6000 397.2000 330.2000 ;
	    RECT 402.8000 329.6000 403.6000 330.4000 ;
	    RECT 415.6000 329.6000 416.4000 330.4000 ;
	    RECT 422.0000 329.6000 422.8000 330.4000 ;
	    RECT 428.4000 330.3000 429.2000 330.4000 ;
	    RECT 430.0000 330.3000 430.8000 330.4000 ;
	    RECT 428.4000 329.7000 430.8000 330.3000 ;
	    RECT 428.4000 329.6000 429.2000 329.7000 ;
	    RECT 430.0000 329.6000 430.8000 329.7000 ;
	    RECT 394.2000 322.2000 395.0000 329.6000 ;
	    RECT 395.8000 328.4000 396.4000 329.6000 ;
	    RECT 395.6000 327.6000 396.4000 328.4000 ;
	    RECT 401.2000 327.6000 402.0000 329.2000 ;
	    RECT 402.8000 327.0000 403.4000 329.6000 ;
	    RECT 414.0000 327.6000 414.8000 329.2000 ;
	    RECT 415.6000 327.0000 416.2000 329.6000 ;
	    RECT 417.2000 328.3000 418.0000 328.4000 ;
	    RECT 420.4000 328.3000 421.2000 329.2000 ;
	    RECT 417.2000 327.7000 421.2000 328.3000 ;
	    RECT 417.2000 327.6000 418.0000 327.7000 ;
	    RECT 420.4000 327.6000 421.2000 327.7000 ;
	    RECT 422.0000 328.3000 422.6000 329.6000 ;
	    RECT 425.2000 328.3000 426.0000 328.4000 ;
	    RECT 422.0000 327.7000 426.0000 328.3000 ;
	    RECT 422.0000 327.0000 422.6000 327.7000 ;
	    RECT 425.2000 327.6000 426.0000 327.7000 ;
	    RECT 426.8000 327.6000 427.6000 329.2000 ;
	    RECT 428.4000 327.0000 429.0000 329.6000 ;
	    RECT 399.8000 326.4000 403.4000 327.0000 ;
	    RECT 399.8000 326.2000 400.4000 326.4000 ;
	    RECT 399.6000 322.2000 400.4000 326.2000 ;
	    RECT 402.8000 326.2000 403.4000 326.4000 ;
	    RECT 412.6000 326.4000 416.2000 327.0000 ;
	    RECT 412.6000 326.2000 413.2000 326.4000 ;
	    RECT 402.8000 322.2000 403.6000 326.2000 ;
	    RECT 412.4000 322.2000 413.2000 326.2000 ;
	    RECT 415.6000 326.2000 416.2000 326.4000 ;
	    RECT 419.0000 326.4000 422.6000 327.0000 ;
	    RECT 419.0000 326.2000 419.6000 326.4000 ;
	    RECT 415.6000 322.2000 416.4000 326.2000 ;
	    RECT 418.8000 322.2000 419.6000 326.2000 ;
	    RECT 422.0000 326.2000 422.6000 326.4000 ;
	    RECT 425.4000 326.4000 429.0000 327.0000 ;
	    RECT 425.4000 326.2000 426.0000 326.4000 ;
	    RECT 422.0000 322.2000 422.8000 326.2000 ;
	    RECT 425.2000 322.2000 426.0000 326.2000 ;
	    RECT 428.4000 326.2000 429.0000 326.4000 ;
	    RECT 428.4000 322.2000 429.2000 326.2000 ;
	    RECT 431.6000 322.2000 432.4000 333.7000 ;
	    RECT 433.2000 333.6000 434.0000 333.7000 ;
	    RECT 436.2000 333.6000 438.8000 334.4000 ;
	    RECT 434.8000 331.6000 435.6000 333.2000 ;
	    RECT 436.2000 330.2000 436.8000 333.6000 ;
	    RECT 439.6000 331.4000 440.4000 334.8000 ;
	    RECT 452.4000 334.4000 453.0000 336.4000 ;
	    RECT 457.2000 335.0000 458.0000 339.8000 ;
	    RECT 446.6000 334.2000 447.4000 334.4000 ;
	    RECT 452.4000 334.2000 453.2000 334.4000 ;
	    RECT 455.6000 334.2000 457.2000 334.4000 ;
	    RECT 460.0000 334.2000 460.8000 339.8000 ;
	    RECT 446.2000 333.6000 457.2000 334.2000 ;
	    RECT 459.0000 333.8000 460.8000 334.2000 ;
	    RECT 468.8000 334.2000 469.6000 339.8000 ;
	    RECT 471.6000 335.8000 472.4000 339.8000 ;
	    RECT 473.2000 336.0000 474.0000 339.8000 ;
	    RECT 476.4000 336.0000 477.2000 339.8000 ;
	    RECT 473.2000 335.8000 477.2000 336.0000 ;
	    RECT 471.8000 334.4000 472.4000 335.8000 ;
	    RECT 473.4000 335.4000 477.0000 335.8000 ;
	    RECT 475.6000 334.4000 476.4000 334.8000 ;
	    RECT 468.8000 333.8000 470.6000 334.2000 ;
	    RECT 459.0000 333.6000 460.6000 333.8000 ;
	    RECT 469.0000 333.6000 470.6000 333.8000 ;
	    RECT 471.6000 333.6000 474.2000 334.4000 ;
	    RECT 475.6000 334.3000 477.2000 334.4000 ;
	    RECT 478.0000 334.3000 478.8000 339.8000 ;
	    RECT 479.6000 335.6000 480.4000 337.2000 ;
	    RECT 475.6000 333.8000 478.8000 334.3000 ;
	    RECT 476.4000 333.7000 478.8000 333.8000 ;
	    RECT 476.4000 333.6000 477.2000 333.7000 ;
	    RECT 444.4000 332.8000 445.2000 333.0000 ;
	    RECT 441.4000 332.2000 445.2000 332.8000 ;
	    RECT 441.4000 332.0000 442.2000 332.2000 ;
	    RECT 443.0000 331.4000 443.8000 331.6000 ;
	    RECT 439.6000 330.8000 443.8000 331.4000 ;
	    RECT 438.0000 330.2000 438.8000 330.4000 ;
	    RECT 435.8000 329.6000 436.8000 330.2000 ;
	    RECT 437.4000 329.6000 438.8000 330.2000 ;
	    RECT 435.8000 322.2000 436.6000 329.6000 ;
	    RECT 437.4000 328.4000 438.0000 329.6000 ;
	    RECT 437.2000 327.6000 438.0000 328.4000 ;
	    RECT 439.6000 322.2000 440.4000 330.8000 ;
	    RECT 446.2000 330.4000 446.8000 333.6000 ;
	    RECT 453.4000 333.4000 454.2000 333.6000 ;
	    RECT 455.0000 332.4000 455.8000 332.6000 ;
	    RECT 450.8000 331.8000 455.8000 332.4000 ;
	    RECT 450.8000 331.6000 451.6000 331.8000 ;
	    RECT 452.4000 331.0000 458.0000 331.2000 ;
	    RECT 452.2000 330.8000 458.0000 331.0000 ;
	    RECT 444.4000 329.8000 446.8000 330.4000 ;
	    RECT 448.2000 330.6000 458.0000 330.8000 ;
	    RECT 448.2000 330.2000 453.0000 330.6000 ;
	    RECT 444.4000 328.8000 445.0000 329.8000 ;
	    RECT 443.6000 328.0000 445.0000 328.8000 ;
	    RECT 446.6000 329.0000 447.4000 329.2000 ;
	    RECT 448.2000 329.0000 448.8000 330.2000 ;
	    RECT 446.6000 328.4000 448.8000 329.0000 ;
	    RECT 449.4000 329.0000 454.8000 329.6000 ;
	    RECT 449.4000 328.8000 450.2000 329.0000 ;
	    RECT 454.0000 328.8000 454.8000 329.0000 ;
	    RECT 447.8000 327.4000 448.6000 327.6000 ;
	    RECT 450.6000 327.4000 451.4000 327.6000 ;
	    RECT 444.4000 326.2000 445.2000 327.0000 ;
	    RECT 447.8000 326.8000 451.4000 327.4000 ;
	    RECT 448.6000 326.2000 449.2000 326.8000 ;
	    RECT 454.0000 326.2000 454.8000 327.0000 ;
	    RECT 443.8000 322.2000 445.0000 326.2000 ;
	    RECT 448.4000 322.2000 449.2000 326.2000 ;
	    RECT 452.8000 325.6000 454.8000 326.2000 ;
	    RECT 452.8000 322.2000 453.6000 325.6000 ;
	    RECT 457.2000 322.2000 458.0000 330.6000 ;
	    RECT 459.0000 330.4000 459.6000 333.6000 ;
	    RECT 461.2000 331.6000 462.8000 332.4000 ;
	    RECT 466.8000 331.6000 468.4000 332.4000 ;
	    RECT 458.8000 329.6000 459.6000 330.4000 ;
	    RECT 459.0000 327.0000 459.6000 329.6000 ;
	    RECT 470.0000 330.4000 470.6000 333.6000 ;
	    RECT 473.6000 332.4000 474.2000 333.6000 ;
	    RECT 473.2000 331.6000 474.2000 332.4000 ;
	    RECT 474.8000 331.6000 475.6000 333.2000 ;
	    RECT 470.0000 329.6000 470.8000 330.4000 ;
	    RECT 471.6000 330.2000 472.4000 330.4000 ;
	    RECT 473.6000 330.2000 474.2000 331.6000 ;
	    RECT 471.6000 329.6000 473.0000 330.2000 ;
	    RECT 473.6000 329.6000 474.6000 330.2000 ;
	    RECT 460.4000 328.3000 461.2000 329.2000 ;
	    RECT 468.4000 328.3000 469.2000 329.2000 ;
	    RECT 460.4000 327.7000 469.2000 328.3000 ;
	    RECT 460.4000 327.6000 461.2000 327.7000 ;
	    RECT 468.4000 327.6000 469.2000 327.7000 ;
	    RECT 470.0000 327.0000 470.6000 329.6000 ;
	    RECT 472.4000 328.4000 473.0000 329.6000 ;
	    RECT 472.4000 327.6000 473.2000 328.4000 ;
	    RECT 459.0000 326.4000 462.6000 327.0000 ;
	    RECT 459.0000 326.2000 459.6000 326.4000 ;
	    RECT 458.8000 322.2000 459.6000 326.2000 ;
	    RECT 462.0000 326.2000 462.6000 326.4000 ;
	    RECT 467.0000 326.4000 470.6000 327.0000 ;
	    RECT 467.0000 326.2000 467.6000 326.4000 ;
	    RECT 462.0000 322.2000 462.8000 326.2000 ;
	    RECT 466.8000 322.2000 467.6000 326.2000 ;
	    RECT 470.0000 326.2000 470.6000 326.4000 ;
	    RECT 470.0000 322.2000 470.8000 326.2000 ;
	    RECT 473.8000 322.2000 474.6000 329.6000 ;
	    RECT 478.0000 322.2000 478.8000 333.7000 ;
	    RECT 481.2000 335.4000 482.0000 339.8000 ;
	    RECT 485.4000 338.4000 486.6000 339.8000 ;
	    RECT 485.4000 337.8000 486.8000 338.4000 ;
	    RECT 490.0000 337.8000 490.8000 339.8000 ;
	    RECT 494.4000 338.4000 495.2000 339.8000 ;
	    RECT 494.4000 337.8000 496.4000 338.4000 ;
	    RECT 486.0000 337.0000 486.8000 337.8000 ;
	    RECT 490.2000 337.2000 490.8000 337.8000 ;
	    RECT 490.2000 336.6000 493.0000 337.2000 ;
	    RECT 492.2000 336.4000 493.0000 336.6000 ;
	    RECT 494.0000 336.4000 494.8000 337.2000 ;
	    RECT 495.6000 337.0000 496.4000 337.8000 ;
	    RECT 484.2000 335.4000 485.0000 335.6000 ;
	    RECT 481.2000 334.8000 485.0000 335.4000 ;
	    RECT 481.2000 331.4000 482.0000 334.8000 ;
	    RECT 488.2000 334.2000 489.0000 334.4000 ;
	    RECT 492.4000 334.2000 493.2000 334.4000 ;
	    RECT 494.0000 334.2000 494.6000 336.4000 ;
	    RECT 498.8000 335.0000 499.6000 339.8000 ;
	    RECT 500.4000 335.6000 501.2000 337.2000 ;
	    RECT 497.2000 334.2000 498.8000 334.4000 ;
	    RECT 487.8000 333.6000 498.8000 334.2000 ;
	    RECT 486.0000 332.8000 486.8000 333.0000 ;
	    RECT 483.0000 332.2000 486.8000 332.8000 ;
	    RECT 483.0000 332.0000 483.8000 332.2000 ;
	    RECT 484.6000 331.4000 485.4000 331.6000 ;
	    RECT 481.2000 330.8000 485.4000 331.4000 ;
	    RECT 479.6000 328.3000 480.4000 328.4000 ;
	    RECT 481.2000 328.3000 482.0000 330.8000 ;
	    RECT 487.8000 330.4000 488.4000 333.6000 ;
	    RECT 495.0000 333.4000 495.8000 333.6000 ;
	    RECT 496.6000 332.4000 497.4000 332.6000 ;
	    RECT 490.8000 332.3000 491.6000 332.4000 ;
	    RECT 492.4000 332.3000 497.4000 332.4000 ;
	    RECT 490.8000 331.8000 497.4000 332.3000 ;
	    RECT 490.8000 331.7000 493.2000 331.8000 ;
	    RECT 490.8000 331.6000 491.6000 331.7000 ;
	    RECT 492.4000 331.6000 493.2000 331.7000 ;
	    RECT 494.0000 331.0000 499.6000 331.2000 ;
	    RECT 493.8000 330.8000 499.6000 331.0000 ;
	    RECT 486.0000 329.8000 488.4000 330.4000 ;
	    RECT 489.8000 330.6000 499.6000 330.8000 ;
	    RECT 489.8000 330.2000 494.6000 330.6000 ;
	    RECT 486.0000 328.8000 486.6000 329.8000 ;
	    RECT 479.6000 327.7000 482.0000 328.3000 ;
	    RECT 485.2000 328.0000 486.6000 328.8000 ;
	    RECT 488.2000 329.0000 489.0000 329.2000 ;
	    RECT 489.8000 329.0000 490.4000 330.2000 ;
	    RECT 488.2000 328.4000 490.4000 329.0000 ;
	    RECT 491.0000 329.0000 496.4000 329.6000 ;
	    RECT 491.0000 328.8000 491.8000 329.0000 ;
	    RECT 495.6000 328.8000 496.4000 329.0000 ;
	    RECT 479.6000 327.6000 480.4000 327.7000 ;
	    RECT 481.2000 322.2000 482.0000 327.7000 ;
	    RECT 489.4000 327.4000 490.2000 327.6000 ;
	    RECT 492.2000 327.4000 493.0000 327.6000 ;
	    RECT 486.0000 326.2000 486.8000 327.0000 ;
	    RECT 489.4000 326.8000 493.0000 327.4000 ;
	    RECT 490.2000 326.2000 490.8000 326.8000 ;
	    RECT 495.6000 326.2000 496.4000 327.0000 ;
	    RECT 485.4000 322.2000 486.6000 326.2000 ;
	    RECT 490.0000 322.2000 490.8000 326.2000 ;
	    RECT 494.4000 325.6000 496.4000 326.2000 ;
	    RECT 494.4000 322.2000 495.2000 325.6000 ;
	    RECT 498.8000 322.2000 499.6000 330.6000 ;
	    RECT 502.0000 322.2000 502.8000 339.8000 ;
	    RECT 503.6000 332.4000 504.4000 339.8000 ;
	    RECT 506.8000 335.2000 507.6000 339.8000 ;
	    RECT 508.4000 335.8000 509.2000 339.8000 ;
	    RECT 512.6000 336.8000 513.4000 339.8000 ;
	    RECT 512.6000 335.8000 514.0000 336.8000 ;
	    RECT 505.4000 334.6000 507.6000 335.2000 ;
	    RECT 508.6000 335.6000 509.2000 335.8000 ;
	    RECT 508.6000 335.2000 510.4000 335.6000 ;
	    RECT 508.6000 335.0000 512.8000 335.2000 ;
	    RECT 509.8000 334.6000 512.8000 335.0000 ;
	    RECT 503.6000 330.2000 504.2000 332.4000 ;
	    RECT 505.4000 331.6000 506.0000 334.6000 ;
	    RECT 512.0000 334.4000 512.8000 334.6000 ;
	    RECT 506.8000 331.6000 507.6000 333.2000 ;
	    RECT 508.4000 332.8000 509.2000 334.4000 ;
	    RECT 510.4000 333.8000 511.2000 334.0000 ;
	    RECT 510.2000 333.2000 511.2000 333.8000 ;
	    RECT 510.2000 332.4000 510.8000 333.2000 ;
	    RECT 510.0000 331.6000 510.8000 332.4000 ;
	    RECT 504.8000 330.8000 506.0000 331.6000 ;
	    RECT 512.0000 331.0000 512.6000 334.4000 ;
	    RECT 513.4000 332.4000 514.0000 335.8000 ;
	    RECT 513.2000 331.6000 514.0000 332.4000 ;
	    RECT 505.4000 330.2000 506.0000 330.8000 ;
	    RECT 510.2000 330.4000 512.6000 331.0000 ;
	    RECT 503.6000 322.2000 504.4000 330.2000 ;
	    RECT 505.4000 329.6000 507.6000 330.2000 ;
	    RECT 506.8000 322.2000 507.6000 329.6000 ;
	    RECT 510.2000 326.2000 510.8000 330.4000 ;
	    RECT 513.4000 330.2000 514.0000 331.6000 ;
	    RECT 510.0000 322.2000 510.8000 326.2000 ;
	    RECT 513.2000 322.2000 514.0000 330.2000 ;
	    RECT 4.4000 312.4000 5.2000 319.8000 ;
	    RECT 9.2000 312.4000 10.0000 319.8000 ;
	    RECT 3.0000 311.8000 5.2000 312.4000 ;
	    RECT 7.8000 311.8000 10.0000 312.4000 ;
	    RECT 3.0000 311.2000 3.6000 311.8000 ;
	    RECT 7.8000 311.2000 8.4000 311.8000 ;
	    RECT 12.4000 311.2000 13.2000 319.8000 ;
	    RECT 15.6000 311.2000 16.4000 319.8000 ;
	    RECT 18.8000 311.2000 19.6000 319.8000 ;
	    RECT 22.0000 311.2000 22.8000 319.8000 ;
	    RECT 2.4000 310.4000 3.6000 311.2000 ;
	    RECT 7.2000 310.4000 8.4000 311.2000 ;
	    RECT 10.8000 310.4000 13.2000 311.2000 ;
	    RECT 14.2000 310.4000 16.4000 311.2000 ;
	    RECT 17.4000 310.4000 19.6000 311.2000 ;
	    RECT 21.0000 310.4000 22.8000 311.2000 ;
	    RECT 25.2000 311.2000 26.0000 319.8000 ;
	    RECT 29.4000 315.8000 30.6000 319.8000 ;
	    RECT 34.0000 315.8000 34.8000 319.8000 ;
	    RECT 38.4000 316.4000 39.2000 319.8000 ;
	    RECT 38.4000 315.8000 40.4000 316.4000 ;
	    RECT 30.0000 315.0000 30.8000 315.8000 ;
	    RECT 34.2000 315.2000 34.8000 315.8000 ;
	    RECT 33.4000 314.6000 37.0000 315.2000 ;
	    RECT 39.6000 315.0000 40.4000 315.8000 ;
	    RECT 33.4000 314.4000 34.2000 314.6000 ;
	    RECT 36.2000 314.4000 37.0000 314.6000 ;
	    RECT 29.2000 313.2000 30.6000 314.0000 ;
	    RECT 30.0000 312.2000 30.6000 313.2000 ;
	    RECT 32.2000 313.0000 34.4000 313.6000 ;
	    RECT 32.2000 312.8000 33.0000 313.0000 ;
	    RECT 30.0000 311.6000 32.4000 312.2000 ;
	    RECT 25.2000 310.6000 29.4000 311.2000 ;
	    RECT 3.0000 307.4000 3.6000 310.4000 ;
	    RECT 4.4000 308.8000 5.2000 310.4000 ;
	    RECT 7.8000 307.4000 8.4000 310.4000 ;
	    RECT 9.2000 308.8000 10.0000 310.4000 ;
	    RECT 10.8000 307.6000 11.6000 310.4000 ;
	    RECT 14.2000 309.0000 15.0000 310.4000 ;
	    RECT 17.4000 309.0000 18.2000 310.4000 ;
	    RECT 21.0000 309.0000 21.8000 310.4000 ;
	    RECT 12.4000 308.2000 15.0000 309.0000 ;
	    RECT 15.8000 308.2000 18.2000 309.0000 ;
	    RECT 19.2000 308.2000 21.8000 309.0000 ;
	    RECT 14.2000 307.6000 15.0000 308.2000 ;
	    RECT 17.4000 307.6000 18.2000 308.2000 ;
	    RECT 21.0000 307.6000 21.8000 308.2000 ;
	    RECT 3.0000 306.8000 5.2000 307.4000 ;
	    RECT 7.8000 306.8000 10.0000 307.4000 ;
	    RECT 10.8000 306.8000 13.2000 307.6000 ;
	    RECT 14.2000 306.8000 16.4000 307.6000 ;
	    RECT 17.4000 306.8000 19.6000 307.6000 ;
	    RECT 21.0000 306.8000 22.8000 307.6000 ;
	    RECT 4.4000 302.2000 5.2000 306.8000 ;
	    RECT 9.2000 302.2000 10.0000 306.8000 ;
	    RECT 12.4000 302.2000 13.2000 306.8000 ;
	    RECT 15.6000 302.2000 16.4000 306.8000 ;
	    RECT 18.8000 302.2000 19.6000 306.8000 ;
	    RECT 22.0000 302.2000 22.8000 306.8000 ;
	    RECT 25.2000 307.2000 26.0000 310.6000 ;
	    RECT 28.6000 310.4000 29.4000 310.6000 ;
	    RECT 27.0000 309.8000 27.8000 310.0000 ;
	    RECT 27.0000 309.2000 30.8000 309.8000 ;
	    RECT 30.0000 309.0000 30.8000 309.2000 ;
	    RECT 31.8000 308.4000 32.4000 311.6000 ;
	    RECT 33.8000 311.8000 34.4000 313.0000 ;
	    RECT 35.0000 313.0000 35.8000 313.2000 ;
	    RECT 39.6000 313.0000 40.4000 313.2000 ;
	    RECT 35.0000 312.4000 40.4000 313.0000 ;
	    RECT 33.8000 311.4000 38.6000 311.8000 ;
	    RECT 42.8000 311.4000 43.6000 319.8000 ;
	    RECT 44.4000 313.6000 46.0000 314.4000 ;
	    RECT 45.2000 312.4000 45.8000 313.6000 ;
	    RECT 46.6000 312.4000 47.4000 319.8000 ;
	    RECT 53.0000 316.4000 53.8000 319.8000 ;
	    RECT 59.8000 318.4000 60.6000 319.8000 ;
	    RECT 58.8000 317.6000 60.6000 318.4000 ;
	    RECT 53.0000 315.6000 54.8000 316.4000 ;
	    RECT 51.6000 313.6000 52.4000 314.4000 ;
	    RECT 51.6000 312.4000 52.2000 313.6000 ;
	    RECT 53.0000 312.4000 53.8000 315.6000 ;
	    RECT 59.8000 312.6000 60.6000 317.6000 ;
	    RECT 64.2000 318.4000 65.0000 319.8000 ;
	    RECT 64.2000 317.6000 66.0000 318.4000 ;
	    RECT 44.4000 311.8000 45.8000 312.4000 ;
	    RECT 44.4000 311.6000 45.2000 311.8000 ;
	    RECT 46.4000 311.6000 48.4000 312.4000 ;
	    RECT 50.8000 311.8000 52.2000 312.4000 ;
	    RECT 52.8000 311.8000 53.8000 312.4000 ;
	    RECT 58.8000 311.8000 60.6000 312.6000 ;
	    RECT 62.8000 313.6000 63.6000 314.4000 ;
	    RECT 62.8000 312.4000 63.4000 313.6000 ;
	    RECT 64.2000 312.4000 65.0000 317.6000 ;
	    RECT 62.0000 311.8000 63.4000 312.4000 ;
	    RECT 64.0000 311.8000 65.0000 312.4000 ;
	    RECT 68.4000 311.8000 69.2000 319.8000 ;
	    RECT 71.6000 312.4000 72.4000 319.8000 ;
	    RECT 75.8000 318.4000 76.6000 319.8000 ;
	    RECT 74.8000 317.6000 76.6000 318.4000 ;
	    RECT 70.2000 311.8000 72.4000 312.4000 ;
	    RECT 75.8000 312.4000 76.6000 317.6000 ;
	    RECT 82.2000 314.4000 83.0000 319.8000 ;
	    RECT 77.2000 313.6000 78.0000 314.4000 ;
	    RECT 81.2000 313.6000 83.0000 314.4000 ;
	    RECT 77.4000 312.4000 78.0000 313.6000 ;
	    RECT 82.2000 312.6000 83.0000 313.6000 ;
	    RECT 75.8000 311.8000 76.8000 312.4000 ;
	    RECT 77.4000 311.8000 78.8000 312.4000 ;
	    RECT 81.2000 311.8000 83.0000 312.6000 ;
	    RECT 50.8000 311.6000 51.6000 311.8000 ;
	    RECT 33.8000 311.2000 43.6000 311.4000 ;
	    RECT 37.8000 311.0000 43.6000 311.2000 ;
	    RECT 38.0000 310.8000 43.6000 311.0000 ;
	    RECT 36.4000 310.2000 37.2000 310.4000 ;
	    RECT 36.4000 309.6000 41.4000 310.2000 ;
	    RECT 38.0000 309.4000 38.8000 309.6000 ;
	    RECT 40.6000 309.4000 41.4000 309.6000 ;
	    RECT 39.0000 308.4000 39.8000 308.6000 ;
	    RECT 46.4000 308.4000 47.0000 311.6000 ;
	    RECT 47.6000 308.8000 48.4000 310.4000 ;
	    RECT 52.8000 308.4000 53.4000 311.8000 ;
	    RECT 54.0000 308.8000 54.8000 310.4000 ;
	    RECT 59.0000 308.4000 59.6000 311.8000 ;
	    RECT 62.0000 311.6000 62.8000 311.8000 ;
	    RECT 60.4000 309.6000 61.2000 311.2000 ;
	    RECT 64.0000 308.4000 64.6000 311.8000 ;
	    RECT 65.2000 310.3000 66.0000 310.4000 ;
	    RECT 66.8000 310.3000 67.6000 310.4000 ;
	    RECT 65.2000 309.7000 67.6000 310.3000 ;
	    RECT 65.2000 308.8000 66.0000 309.7000 ;
	    RECT 66.8000 309.6000 67.6000 309.7000 ;
	    RECT 68.4000 309.6000 69.0000 311.8000 ;
	    RECT 70.2000 311.2000 70.8000 311.8000 ;
	    RECT 69.6000 310.4000 70.8000 311.2000 ;
	    RECT 31.8000 307.8000 42.8000 308.4000 ;
	    RECT 32.2000 307.6000 33.0000 307.8000 ;
	    RECT 36.4000 307.6000 37.2000 307.8000 ;
	    RECT 25.2000 306.6000 29.0000 307.2000 ;
	    RECT 25.2000 302.2000 26.0000 306.6000 ;
	    RECT 28.2000 306.4000 29.0000 306.6000 ;
	    RECT 38.0000 305.6000 38.6000 307.8000 ;
	    RECT 41.2000 307.6000 42.8000 307.8000 ;
	    RECT 44.4000 307.6000 47.0000 308.4000 ;
	    RECT 49.2000 308.2000 50.0000 308.4000 ;
	    RECT 48.4000 307.6000 50.0000 308.2000 ;
	    RECT 50.8000 307.6000 53.4000 308.4000 ;
	    RECT 55.6000 308.2000 56.4000 308.4000 ;
	    RECT 54.8000 307.6000 56.4000 308.2000 ;
	    RECT 58.8000 307.6000 59.6000 308.4000 ;
	    RECT 62.0000 307.6000 64.6000 308.4000 ;
	    RECT 66.8000 308.3000 67.6000 308.4000 ;
	    RECT 68.4000 308.3000 69.2000 309.6000 ;
	    RECT 66.8000 308.2000 69.2000 308.3000 ;
	    RECT 66.0000 307.7000 69.2000 308.2000 ;
	    RECT 66.0000 307.6000 67.6000 307.7000 ;
	    RECT 36.2000 305.4000 37.0000 305.6000 ;
	    RECT 30.0000 304.2000 30.8000 305.0000 ;
	    RECT 34.2000 304.8000 37.0000 305.4000 ;
	    RECT 38.0000 304.8000 38.8000 305.6000 ;
	    RECT 34.2000 304.2000 34.8000 304.8000 ;
	    RECT 39.6000 304.2000 40.4000 305.0000 ;
	    RECT 29.4000 303.6000 30.8000 304.2000 ;
	    RECT 29.4000 302.2000 30.6000 303.6000 ;
	    RECT 34.0000 302.2000 34.8000 304.2000 ;
	    RECT 38.4000 303.6000 40.4000 304.2000 ;
	    RECT 38.4000 302.2000 39.2000 303.6000 ;
	    RECT 42.8000 302.2000 43.6000 307.0000 ;
	    RECT 44.6000 306.2000 45.2000 307.6000 ;
	    RECT 48.4000 307.2000 49.2000 307.6000 ;
	    RECT 46.2000 306.2000 49.8000 306.6000 ;
	    RECT 51.0000 306.2000 51.6000 307.6000 ;
	    RECT 54.8000 307.2000 55.6000 307.6000 ;
	    RECT 52.6000 306.2000 56.2000 306.6000 ;
	    RECT 44.4000 302.2000 45.2000 306.2000 ;
	    RECT 46.0000 306.0000 50.0000 306.2000 ;
	    RECT 46.0000 302.2000 46.8000 306.0000 ;
	    RECT 49.2000 302.2000 50.0000 306.0000 ;
	    RECT 50.8000 302.2000 51.6000 306.2000 ;
	    RECT 52.4000 306.0000 56.4000 306.2000 ;
	    RECT 52.4000 302.2000 53.2000 306.0000 ;
	    RECT 55.6000 302.2000 56.4000 306.0000 ;
	    RECT 57.2000 304.8000 58.0000 306.4000 ;
	    RECT 59.0000 304.2000 59.6000 307.6000 ;
	    RECT 62.2000 306.2000 62.8000 307.6000 ;
	    RECT 66.0000 307.2000 66.8000 307.6000 ;
	    RECT 63.8000 306.2000 67.4000 306.6000 ;
	    RECT 58.8000 302.2000 59.6000 304.2000 ;
	    RECT 62.0000 302.2000 62.8000 306.2000 ;
	    RECT 63.6000 306.0000 67.6000 306.2000 ;
	    RECT 63.6000 302.2000 64.4000 306.0000 ;
	    RECT 66.8000 302.2000 67.6000 306.0000 ;
	    RECT 68.4000 302.2000 69.2000 307.7000 ;
	    RECT 70.2000 307.4000 70.8000 310.4000 ;
	    RECT 74.8000 308.8000 75.6000 310.4000 ;
	    RECT 76.2000 308.4000 76.8000 311.8000 ;
	    RECT 78.0000 311.6000 78.8000 311.8000 ;
	    RECT 81.4000 308.4000 82.0000 311.8000 ;
	    RECT 84.4000 311.4000 85.2000 319.8000 ;
	    RECT 88.8000 316.4000 89.6000 319.8000 ;
	    RECT 87.6000 315.8000 89.6000 316.4000 ;
	    RECT 93.2000 315.8000 94.0000 319.8000 ;
	    RECT 97.4000 315.8000 98.6000 319.8000 ;
	    RECT 87.6000 315.0000 88.4000 315.8000 ;
	    RECT 93.2000 315.2000 93.8000 315.8000 ;
	    RECT 91.0000 314.6000 94.6000 315.2000 ;
	    RECT 97.2000 315.0000 98.0000 315.8000 ;
	    RECT 91.0000 314.4000 91.8000 314.6000 ;
	    RECT 93.8000 314.4000 94.6000 314.6000 ;
	    RECT 87.6000 313.0000 88.4000 313.2000 ;
	    RECT 92.2000 313.0000 93.0000 313.2000 ;
	    RECT 87.6000 312.4000 93.0000 313.0000 ;
	    RECT 93.6000 313.0000 95.8000 313.6000 ;
	    RECT 93.6000 311.8000 94.2000 313.0000 ;
	    RECT 95.0000 312.8000 95.8000 313.0000 ;
	    RECT 97.4000 313.2000 98.8000 314.0000 ;
	    RECT 97.4000 312.2000 98.0000 313.2000 ;
	    RECT 89.4000 311.4000 94.2000 311.8000 ;
	    RECT 84.4000 311.2000 94.2000 311.4000 ;
	    RECT 95.6000 311.6000 98.0000 312.2000 ;
	    RECT 82.8000 309.6000 83.6000 311.2000 ;
	    RECT 84.4000 311.0000 90.2000 311.2000 ;
	    RECT 84.4000 310.8000 90.0000 311.0000 ;
	    RECT 90.8000 310.2000 91.6000 310.4000 ;
	    RECT 86.6000 309.6000 91.6000 310.2000 ;
	    RECT 86.6000 309.4000 87.4000 309.6000 ;
	    RECT 88.2000 308.4000 89.0000 308.6000 ;
	    RECT 95.6000 308.4000 96.2000 311.6000 ;
	    RECT 102.0000 311.2000 102.8000 319.8000 ;
	    RECT 98.6000 310.6000 102.8000 311.2000 ;
	    RECT 98.6000 310.4000 99.4000 310.6000 ;
	    RECT 100.2000 309.8000 101.0000 310.0000 ;
	    RECT 97.2000 309.2000 101.0000 309.8000 ;
	    RECT 97.2000 309.0000 98.0000 309.2000 ;
	    RECT 73.2000 308.2000 74.0000 308.4000 ;
	    RECT 73.2000 307.6000 74.8000 308.2000 ;
	    RECT 76.2000 307.6000 78.8000 308.4000 ;
	    RECT 81.2000 307.6000 82.0000 308.4000 ;
	    RECT 85.2000 307.8000 96.2000 308.4000 ;
	    RECT 85.2000 307.6000 86.8000 307.8000 ;
	    RECT 70.2000 306.8000 72.4000 307.4000 ;
	    RECT 74.0000 307.2000 74.8000 307.6000 ;
	    RECT 71.6000 302.2000 72.4000 306.8000 ;
	    RECT 73.4000 306.2000 77.0000 306.6000 ;
	    RECT 78.0000 306.2000 78.6000 307.6000 ;
	    RECT 73.2000 306.0000 77.2000 306.2000 ;
	    RECT 73.2000 302.2000 74.0000 306.0000 ;
	    RECT 76.4000 302.2000 77.2000 306.0000 ;
	    RECT 78.0000 302.2000 78.8000 306.2000 ;
	    RECT 79.6000 304.8000 80.4000 306.4000 ;
	    RECT 81.4000 304.2000 82.0000 307.6000 ;
	    RECT 81.2000 302.2000 82.0000 304.2000 ;
	    RECT 84.4000 302.2000 85.2000 307.0000 ;
	    RECT 89.4000 306.4000 90.0000 307.8000 ;
	    RECT 95.0000 307.6000 95.8000 307.8000 ;
	    RECT 102.0000 307.2000 102.8000 310.6000 ;
	    RECT 111.6000 310.3000 112.4000 319.8000 ;
	    RECT 115.6000 313.6000 116.4000 314.4000 ;
	    RECT 113.2000 311.6000 114.0000 313.2000 ;
	    RECT 115.6000 312.4000 116.2000 313.6000 ;
	    RECT 117.0000 312.4000 117.8000 319.8000 ;
	    RECT 123.8000 318.4000 125.8000 319.8000 ;
	    RECT 122.8000 317.6000 125.8000 318.4000 ;
	    RECT 114.8000 311.8000 116.2000 312.4000 ;
	    RECT 116.8000 311.8000 117.8000 312.4000 ;
	    RECT 123.8000 311.8000 125.8000 317.6000 ;
	    RECT 130.0000 313.6000 130.8000 314.4000 ;
	    RECT 130.0000 312.4000 130.6000 313.6000 ;
	    RECT 131.4000 312.4000 132.2000 319.8000 ;
	    RECT 129.2000 311.8000 130.6000 312.4000 ;
	    RECT 131.2000 311.8000 132.2000 312.4000 ;
	    RECT 135.6000 315.0000 136.4000 319.0000 ;
	    RECT 114.8000 311.6000 115.6000 311.8000 ;
	    RECT 114.9000 310.3000 115.5000 311.6000 ;
	    RECT 111.6000 309.7000 115.5000 310.3000 ;
	    RECT 103.6000 308.3000 104.4000 308.4000 ;
	    RECT 110.0000 308.3000 110.8000 308.4000 ;
	    RECT 103.6000 307.7000 110.8000 308.3000 ;
	    RECT 103.6000 307.6000 104.4000 307.7000 ;
	    RECT 99.0000 306.6000 102.8000 307.2000 ;
	    RECT 110.0000 306.8000 110.8000 307.7000 ;
	    RECT 99.0000 306.4000 99.8000 306.6000 ;
	    RECT 87.6000 304.2000 88.4000 305.0000 ;
	    RECT 89.2000 304.8000 90.0000 306.4000 ;
	    RECT 91.0000 305.4000 91.8000 305.6000 ;
	    RECT 91.0000 304.8000 93.8000 305.4000 ;
	    RECT 93.2000 304.2000 93.8000 304.8000 ;
	    RECT 97.2000 304.2000 98.0000 305.0000 ;
	    RECT 102.0000 304.3000 102.8000 306.6000 ;
	    RECT 111.6000 306.2000 112.4000 309.7000 ;
	    RECT 116.8000 308.4000 117.4000 311.8000 ;
	    RECT 118.0000 308.8000 118.8000 310.4000 ;
	    RECT 114.8000 307.6000 117.4000 308.4000 ;
	    RECT 119.6000 308.2000 120.4000 308.4000 ;
	    RECT 118.8000 307.6000 120.4000 308.2000 ;
	    RECT 121.2000 307.6000 122.0000 309.2000 ;
	    RECT 122.8000 308.8000 123.6000 310.4000 ;
	    RECT 124.6000 308.4000 125.2000 311.8000 ;
	    RECT 129.2000 311.6000 130.0000 311.8000 ;
	    RECT 126.0000 308.8000 126.8000 310.4000 ;
	    RECT 131.2000 308.4000 131.8000 311.8000 ;
	    RECT 135.6000 311.6000 136.2000 315.0000 ;
	    RECT 139.8000 312.8000 140.6000 319.8000 ;
	    RECT 139.8000 312.2000 141.4000 312.8000 ;
	    RECT 135.6000 311.0000 139.4000 311.6000 ;
	    RECT 132.4000 310.3000 133.2000 310.4000 ;
	    RECT 135.6000 310.3000 136.4000 310.4000 ;
	    RECT 132.4000 309.7000 136.4000 310.3000 ;
	    RECT 132.4000 308.8000 133.2000 309.7000 ;
	    RECT 135.6000 308.8000 136.4000 309.7000 ;
	    RECT 137.2000 308.8000 138.0000 310.4000 ;
	    RECT 138.8000 309.0000 139.4000 311.0000 ;
	    RECT 124.4000 308.2000 125.2000 308.4000 ;
	    RECT 127.6000 308.3000 128.4000 308.4000 ;
	    RECT 129.2000 308.3000 131.8000 308.4000 ;
	    RECT 127.6000 308.2000 131.8000 308.3000 ;
	    RECT 134.0000 308.2000 134.8000 308.4000 ;
	    RECT 122.8000 307.6000 125.2000 308.2000 ;
	    RECT 126.8000 307.7000 131.8000 308.2000 ;
	    RECT 126.8000 307.6000 128.4000 307.7000 ;
	    RECT 129.2000 307.6000 131.8000 307.7000 ;
	    RECT 133.2000 307.6000 134.8000 308.2000 ;
	    RECT 138.8000 308.2000 140.2000 309.0000 ;
	    RECT 140.8000 308.4000 141.4000 312.2000 ;
	    RECT 145.8000 312.6000 146.6000 319.8000 ;
	    RECT 145.8000 311.8000 147.6000 312.6000 ;
	    RECT 142.0000 309.6000 142.8000 311.2000 ;
	    RECT 143.6000 310.3000 144.4000 310.4000 ;
	    RECT 145.2000 310.3000 146.0000 311.2000 ;
	    RECT 143.6000 309.7000 146.0000 310.3000 ;
	    RECT 143.6000 309.6000 144.4000 309.7000 ;
	    RECT 145.2000 309.6000 146.0000 309.7000 ;
	    RECT 146.8000 310.4000 147.4000 311.8000 ;
	    RECT 150.0000 311.2000 150.8000 319.8000 ;
	    RECT 154.2000 315.8000 155.4000 319.8000 ;
	    RECT 158.8000 315.8000 159.6000 319.8000 ;
	    RECT 163.2000 316.4000 164.0000 319.8000 ;
	    RECT 163.2000 315.8000 165.2000 316.4000 ;
	    RECT 154.8000 315.0000 155.6000 315.8000 ;
	    RECT 159.0000 315.2000 159.6000 315.8000 ;
	    RECT 158.2000 314.6000 161.8000 315.2000 ;
	    RECT 164.4000 315.0000 165.2000 315.8000 ;
	    RECT 158.2000 314.4000 159.0000 314.6000 ;
	    RECT 161.0000 314.4000 161.8000 314.6000 ;
	    RECT 154.0000 313.2000 155.4000 314.0000 ;
	    RECT 154.8000 312.2000 155.4000 313.2000 ;
	    RECT 157.0000 313.0000 159.2000 313.6000 ;
	    RECT 157.0000 312.8000 157.8000 313.0000 ;
	    RECT 154.8000 311.6000 157.2000 312.2000 ;
	    RECT 150.0000 310.6000 154.2000 311.2000 ;
	    RECT 146.8000 309.6000 147.6000 310.4000 ;
	    RECT 146.8000 308.4000 147.4000 309.6000 ;
	    RECT 138.8000 307.8000 139.8000 308.2000 ;
	    RECT 115.0000 306.2000 115.6000 307.6000 ;
	    RECT 118.8000 307.2000 119.6000 307.6000 ;
	    RECT 116.6000 306.2000 120.2000 306.6000 ;
	    RECT 122.8000 306.2000 123.4000 307.6000 ;
	    RECT 126.8000 307.2000 127.6000 307.6000 ;
	    RECT 124.6000 306.2000 128.2000 306.6000 ;
	    RECT 129.4000 306.2000 130.0000 307.6000 ;
	    RECT 133.2000 307.2000 134.0000 307.6000 ;
	    RECT 135.6000 307.2000 139.8000 307.8000 ;
	    RECT 140.8000 307.6000 142.8000 308.4000 ;
	    RECT 146.8000 307.6000 147.6000 308.4000 ;
	    RECT 131.0000 306.2000 134.6000 306.6000 ;
	    RECT 111.6000 305.6000 113.4000 306.2000 ;
	    RECT 103.6000 304.3000 104.4000 304.4000 ;
	    RECT 87.6000 303.6000 89.6000 304.2000 ;
	    RECT 88.8000 302.2000 89.6000 303.6000 ;
	    RECT 93.2000 302.2000 94.0000 304.2000 ;
	    RECT 97.2000 303.6000 98.6000 304.2000 ;
	    RECT 97.4000 302.2000 98.6000 303.6000 ;
	    RECT 102.0000 303.7000 104.4000 304.3000 ;
	    RECT 102.0000 302.2000 102.8000 303.7000 ;
	    RECT 103.6000 303.6000 104.4000 303.7000 ;
	    RECT 112.6000 302.2000 113.4000 305.6000 ;
	    RECT 114.8000 302.2000 115.6000 306.2000 ;
	    RECT 116.4000 306.0000 120.4000 306.2000 ;
	    RECT 116.4000 302.2000 117.2000 306.0000 ;
	    RECT 119.6000 302.2000 120.4000 306.0000 ;
	    RECT 121.2000 302.8000 122.0000 306.2000 ;
	    RECT 122.8000 303.4000 123.6000 306.2000 ;
	    RECT 124.4000 306.0000 128.4000 306.2000 ;
	    RECT 124.4000 302.8000 125.2000 306.0000 ;
	    RECT 121.2000 302.2000 125.2000 302.8000 ;
	    RECT 127.6000 302.2000 128.4000 306.0000 ;
	    RECT 129.2000 302.2000 130.0000 306.2000 ;
	    RECT 130.8000 306.0000 134.8000 306.2000 ;
	    RECT 130.8000 302.2000 131.6000 306.0000 ;
	    RECT 134.0000 302.2000 134.8000 306.0000 ;
	    RECT 135.6000 305.0000 136.2000 307.2000 ;
	    RECT 140.8000 307.0000 141.4000 307.6000 ;
	    RECT 140.6000 306.6000 141.4000 307.0000 ;
	    RECT 139.8000 306.0000 141.4000 306.6000 ;
	    RECT 135.6000 303.0000 136.4000 305.0000 ;
	    RECT 139.8000 304.4000 140.6000 306.0000 ;
	    RECT 138.8000 303.6000 140.6000 304.4000 ;
	    RECT 139.8000 303.0000 140.6000 303.6000 ;
	    RECT 146.8000 304.2000 147.4000 307.6000 ;
	    RECT 150.0000 307.2000 150.8000 310.6000 ;
	    RECT 153.4000 310.4000 154.2000 310.6000 ;
	    RECT 156.6000 310.4000 157.2000 311.6000 ;
	    RECT 158.6000 311.8000 159.2000 313.0000 ;
	    RECT 159.8000 313.0000 160.6000 313.2000 ;
	    RECT 164.4000 313.0000 165.2000 313.2000 ;
	    RECT 159.8000 312.4000 165.2000 313.0000 ;
	    RECT 158.6000 311.4000 163.4000 311.8000 ;
	    RECT 167.6000 311.4000 168.4000 319.8000 ;
	    RECT 158.6000 311.2000 168.4000 311.4000 ;
	    RECT 162.6000 311.0000 168.4000 311.2000 ;
	    RECT 162.8000 310.8000 168.4000 311.0000 ;
	    RECT 169.2000 311.2000 170.0000 319.8000 ;
	    RECT 173.4000 315.8000 174.6000 319.8000 ;
	    RECT 178.0000 315.8000 178.8000 319.8000 ;
	    RECT 182.4000 316.4000 183.2000 319.8000 ;
	    RECT 182.4000 315.8000 184.4000 316.4000 ;
	    RECT 174.0000 315.0000 174.8000 315.8000 ;
	    RECT 178.2000 315.2000 178.8000 315.8000 ;
	    RECT 177.4000 314.6000 181.0000 315.2000 ;
	    RECT 183.6000 315.0000 184.4000 315.8000 ;
	    RECT 177.4000 314.4000 178.2000 314.6000 ;
	    RECT 180.2000 314.4000 181.0000 314.6000 ;
	    RECT 173.2000 313.2000 174.6000 314.0000 ;
	    RECT 174.0000 312.2000 174.6000 313.2000 ;
	    RECT 176.2000 313.0000 178.4000 313.6000 ;
	    RECT 176.2000 312.8000 177.0000 313.0000 ;
	    RECT 174.0000 311.6000 176.4000 312.2000 ;
	    RECT 169.2000 310.6000 173.4000 311.2000 ;
	    RECT 151.8000 309.8000 152.6000 310.0000 ;
	    RECT 151.8000 309.2000 155.6000 309.8000 ;
	    RECT 156.4000 309.6000 157.2000 310.4000 ;
	    RECT 161.2000 310.2000 162.0000 310.4000 ;
	    RECT 161.2000 309.6000 166.2000 310.2000 ;
	    RECT 154.8000 309.0000 155.6000 309.2000 ;
	    RECT 156.6000 308.4000 157.2000 309.6000 ;
	    RECT 162.8000 309.4000 163.6000 309.6000 ;
	    RECT 165.4000 309.4000 166.2000 309.6000 ;
	    RECT 163.8000 308.4000 164.6000 308.6000 ;
	    RECT 156.6000 307.8000 167.6000 308.4000 ;
	    RECT 157.0000 307.6000 157.8000 307.8000 ;
	    RECT 150.0000 306.6000 153.8000 307.2000 ;
	    RECT 148.4000 304.8000 149.2000 306.4000 ;
	    RECT 146.8000 302.2000 147.6000 304.2000 ;
	    RECT 150.0000 302.2000 150.8000 306.6000 ;
	    RECT 153.0000 306.4000 153.8000 306.6000 ;
	    RECT 162.8000 305.6000 163.4000 307.8000 ;
	    RECT 166.0000 307.6000 167.6000 307.8000 ;
	    RECT 169.2000 307.2000 170.0000 310.6000 ;
	    RECT 172.6000 310.4000 173.4000 310.6000 ;
	    RECT 175.8000 310.4000 176.4000 311.6000 ;
	    RECT 177.8000 311.8000 178.4000 313.0000 ;
	    RECT 179.0000 313.0000 179.8000 313.2000 ;
	    RECT 183.6000 313.0000 184.4000 313.2000 ;
	    RECT 179.0000 312.4000 184.4000 313.0000 ;
	    RECT 177.8000 311.4000 182.6000 311.8000 ;
	    RECT 186.8000 311.4000 187.6000 319.8000 ;
	    RECT 177.8000 311.2000 187.6000 311.4000 ;
	    RECT 181.8000 311.0000 187.6000 311.2000 ;
	    RECT 182.0000 310.8000 187.6000 311.0000 ;
	    RECT 171.0000 309.8000 171.8000 310.0000 ;
	    RECT 171.0000 309.2000 174.8000 309.8000 ;
	    RECT 175.6000 309.6000 176.4000 310.4000 ;
	    RECT 180.4000 310.2000 181.2000 310.4000 ;
	    RECT 180.4000 309.6000 185.4000 310.2000 ;
	    RECT 174.0000 309.0000 174.8000 309.2000 ;
	    RECT 175.8000 308.4000 176.4000 309.6000 ;
	    RECT 182.0000 309.4000 182.8000 309.6000 ;
	    RECT 184.6000 309.4000 185.4000 309.6000 ;
	    RECT 183.0000 308.4000 183.8000 308.6000 ;
	    RECT 175.8000 307.8000 186.8000 308.4000 ;
	    RECT 176.2000 307.6000 177.0000 307.8000 ;
	    RECT 161.0000 305.4000 161.8000 305.6000 ;
	    RECT 154.8000 304.2000 155.6000 305.0000 ;
	    RECT 159.0000 304.8000 161.8000 305.4000 ;
	    RECT 162.8000 304.8000 163.6000 305.6000 ;
	    RECT 159.0000 304.2000 159.6000 304.8000 ;
	    RECT 164.4000 304.2000 165.2000 305.0000 ;
	    RECT 154.2000 303.6000 155.6000 304.2000 ;
	    RECT 154.2000 302.2000 155.4000 303.6000 ;
	    RECT 158.8000 302.2000 159.6000 304.2000 ;
	    RECT 163.2000 303.6000 165.2000 304.2000 ;
	    RECT 163.2000 302.2000 164.0000 303.6000 ;
	    RECT 167.6000 302.2000 168.4000 307.0000 ;
	    RECT 169.2000 306.6000 173.0000 307.2000 ;
	    RECT 169.2000 302.2000 170.0000 306.6000 ;
	    RECT 172.2000 306.4000 173.0000 306.6000 ;
	    RECT 182.0000 305.6000 182.6000 307.8000 ;
	    RECT 185.2000 307.6000 186.8000 307.8000 ;
	    RECT 180.2000 305.4000 181.0000 305.6000 ;
	    RECT 174.0000 304.2000 174.8000 305.0000 ;
	    RECT 178.2000 304.8000 181.0000 305.4000 ;
	    RECT 182.0000 304.8000 182.8000 305.6000 ;
	    RECT 178.2000 304.2000 178.8000 304.8000 ;
	    RECT 183.6000 304.2000 184.4000 305.0000 ;
	    RECT 173.4000 303.6000 174.8000 304.2000 ;
	    RECT 173.4000 302.2000 174.6000 303.6000 ;
	    RECT 178.0000 302.2000 178.8000 304.2000 ;
	    RECT 182.4000 303.6000 184.4000 304.2000 ;
	    RECT 182.4000 302.2000 183.2000 303.6000 ;
	    RECT 186.8000 302.2000 187.6000 307.0000 ;
	    RECT 188.4000 304.8000 189.2000 306.4000 ;
	    RECT 190.0000 302.2000 190.8000 319.8000 ;
	    RECT 193.2000 310.3000 194.0000 319.8000 ;
	    RECT 197.2000 313.6000 198.0000 314.4000 ;
	    RECT 194.8000 311.6000 195.6000 313.2000 ;
	    RECT 197.2000 312.4000 197.8000 313.6000 ;
	    RECT 198.6000 312.4000 199.4000 319.8000 ;
	    RECT 196.4000 311.8000 197.8000 312.4000 ;
	    RECT 196.4000 311.6000 197.2000 311.8000 ;
	    RECT 198.4000 311.6000 200.4000 312.4000 ;
	    RECT 196.5000 310.3000 197.1000 311.6000 ;
	    RECT 193.2000 309.7000 197.1000 310.3000 ;
	    RECT 191.6000 306.8000 192.4000 308.4000 ;
	    RECT 193.2000 306.2000 194.0000 309.7000 ;
	    RECT 198.4000 308.4000 199.0000 311.6000 ;
	    RECT 202.8000 311.4000 203.6000 319.8000 ;
	    RECT 207.2000 316.4000 208.0000 319.8000 ;
	    RECT 206.0000 315.8000 208.0000 316.4000 ;
	    RECT 211.6000 315.8000 212.4000 319.8000 ;
	    RECT 215.8000 315.8000 217.0000 319.8000 ;
	    RECT 206.0000 315.0000 206.8000 315.8000 ;
	    RECT 211.6000 315.2000 212.2000 315.8000 ;
	    RECT 209.4000 314.6000 213.0000 315.2000 ;
	    RECT 215.6000 315.0000 216.4000 315.8000 ;
	    RECT 209.4000 314.4000 210.2000 314.6000 ;
	    RECT 212.2000 314.4000 213.0000 314.6000 ;
	    RECT 206.0000 313.0000 206.8000 313.2000 ;
	    RECT 210.6000 313.0000 211.4000 313.2000 ;
	    RECT 206.0000 312.4000 211.4000 313.0000 ;
	    RECT 212.0000 313.0000 214.2000 313.6000 ;
	    RECT 212.0000 311.8000 212.6000 313.0000 ;
	    RECT 213.4000 312.8000 214.2000 313.0000 ;
	    RECT 215.8000 313.2000 217.2000 314.0000 ;
	    RECT 215.8000 312.2000 216.4000 313.2000 ;
	    RECT 207.8000 311.4000 212.6000 311.8000 ;
	    RECT 202.8000 311.2000 212.6000 311.4000 ;
	    RECT 214.0000 311.6000 216.4000 312.2000 ;
	    RECT 202.8000 311.0000 208.6000 311.2000 ;
	    RECT 202.8000 310.8000 208.4000 311.0000 ;
	    RECT 214.0000 310.4000 214.6000 311.6000 ;
	    RECT 220.4000 311.2000 221.2000 319.8000 ;
	    RECT 224.6000 314.4000 225.4000 319.8000 ;
	    RECT 223.6000 313.6000 225.4000 314.4000 ;
	    RECT 226.0000 313.6000 226.8000 314.4000 ;
	    RECT 224.6000 312.4000 225.4000 313.6000 ;
	    RECT 226.2000 312.4000 226.8000 313.6000 ;
	    RECT 228.4000 312.4000 229.2000 319.8000 ;
	    RECT 224.6000 311.8000 225.6000 312.4000 ;
	    RECT 226.2000 311.8000 227.6000 312.4000 ;
	    RECT 228.4000 311.8000 230.6000 312.4000 ;
	    RECT 231.6000 311.8000 232.4000 319.8000 ;
	    RECT 235.8000 314.4000 236.6000 319.8000 ;
	    RECT 235.8000 313.6000 237.2000 314.4000 ;
	    RECT 235.8000 312.6000 236.6000 313.6000 ;
	    RECT 234.8000 311.8000 236.6000 312.6000 ;
	    RECT 240.6000 311.8000 242.6000 319.8000 ;
	    RECT 248.6000 311.8000 250.6000 319.8000 ;
	    RECT 261.0000 312.6000 261.8000 319.8000 ;
	    RECT 267.4000 318.4000 268.2000 319.8000 ;
	    RECT 267.4000 317.6000 269.2000 318.4000 ;
	    RECT 266.0000 313.6000 266.8000 314.4000 ;
	    RECT 261.0000 311.8000 262.8000 312.6000 ;
	    RECT 266.0000 312.4000 266.6000 313.6000 ;
	    RECT 267.4000 312.4000 268.2000 317.6000 ;
	    RECT 275.4000 312.8000 276.2000 319.8000 ;
	    RECT 279.6000 315.0000 280.4000 319.0000 ;
	    RECT 265.2000 311.8000 266.6000 312.4000 ;
	    RECT 267.2000 311.8000 268.2000 312.4000 ;
	    RECT 274.6000 312.2000 276.2000 312.8000 ;
	    RECT 217.0000 310.6000 221.2000 311.2000 ;
	    RECT 217.0000 310.4000 217.8000 310.6000 ;
	    RECT 199.6000 308.8000 200.4000 310.4000 ;
	    RECT 209.2000 310.2000 210.0000 310.4000 ;
	    RECT 205.0000 309.6000 210.0000 310.2000 ;
	    RECT 214.0000 309.6000 214.8000 310.4000 ;
	    RECT 218.6000 309.8000 219.4000 310.0000 ;
	    RECT 205.0000 309.4000 205.8000 309.6000 ;
	    RECT 207.6000 309.4000 208.4000 309.6000 ;
	    RECT 206.6000 308.4000 207.4000 308.6000 ;
	    RECT 214.0000 308.4000 214.6000 309.6000 ;
	    RECT 215.6000 309.2000 219.4000 309.8000 ;
	    RECT 215.6000 309.0000 216.4000 309.2000 ;
	    RECT 196.4000 307.6000 199.0000 308.4000 ;
	    RECT 201.2000 308.2000 202.0000 308.4000 ;
	    RECT 200.4000 307.6000 202.0000 308.2000 ;
	    RECT 203.6000 307.8000 214.6000 308.4000 ;
	    RECT 203.6000 307.6000 205.2000 307.8000 ;
	    RECT 196.6000 306.2000 197.2000 307.6000 ;
	    RECT 200.4000 307.2000 201.2000 307.6000 ;
	    RECT 198.2000 306.2000 201.8000 306.6000 ;
	    RECT 193.2000 305.6000 195.0000 306.2000 ;
	    RECT 194.2000 302.2000 195.0000 305.6000 ;
	    RECT 196.4000 302.2000 197.2000 306.2000 ;
	    RECT 198.0000 306.0000 202.0000 306.2000 ;
	    RECT 198.0000 302.2000 198.8000 306.0000 ;
	    RECT 201.2000 302.2000 202.0000 306.0000 ;
	    RECT 202.8000 302.2000 203.6000 307.0000 ;
	    RECT 207.8000 305.6000 208.4000 307.8000 ;
	    RECT 213.4000 307.6000 214.2000 307.8000 ;
	    RECT 220.4000 307.2000 221.2000 310.6000 ;
	    RECT 223.6000 308.8000 224.4000 310.4000 ;
	    RECT 225.0000 308.4000 225.6000 311.8000 ;
	    RECT 226.8000 311.6000 227.6000 311.8000 ;
	    RECT 230.0000 311.2000 230.6000 311.8000 ;
	    RECT 230.0000 310.4000 231.2000 311.2000 ;
	    RECT 222.0000 308.2000 222.8000 308.4000 ;
	    RECT 222.0000 307.6000 223.6000 308.2000 ;
	    RECT 225.0000 307.6000 227.6000 308.4000 ;
	    RECT 222.8000 307.2000 223.6000 307.6000 ;
	    RECT 217.4000 306.6000 221.2000 307.2000 ;
	    RECT 217.4000 306.4000 218.2000 306.6000 ;
	    RECT 206.0000 304.2000 206.8000 305.0000 ;
	    RECT 207.6000 304.8000 208.4000 305.6000 ;
	    RECT 209.4000 305.4000 210.2000 305.6000 ;
	    RECT 209.4000 304.8000 212.2000 305.4000 ;
	    RECT 211.6000 304.2000 212.2000 304.8000 ;
	    RECT 215.6000 304.2000 216.4000 305.0000 ;
	    RECT 206.0000 303.6000 208.0000 304.2000 ;
	    RECT 207.2000 302.2000 208.0000 303.6000 ;
	    RECT 211.6000 302.2000 212.4000 304.2000 ;
	    RECT 215.6000 303.6000 217.0000 304.2000 ;
	    RECT 215.8000 302.2000 217.0000 303.6000 ;
	    RECT 220.4000 302.2000 221.2000 306.6000 ;
	    RECT 222.2000 306.2000 225.8000 306.6000 ;
	    RECT 226.8000 306.2000 227.4000 307.6000 ;
	    RECT 230.0000 307.4000 230.6000 310.4000 ;
	    RECT 231.8000 309.6000 232.4000 311.8000 ;
	    RECT 228.4000 306.8000 230.6000 307.4000 ;
	    RECT 222.0000 306.0000 226.0000 306.2000 ;
	    RECT 222.0000 302.2000 222.8000 306.0000 ;
	    RECT 225.2000 302.2000 226.0000 306.0000 ;
	    RECT 226.8000 302.2000 227.6000 306.2000 ;
	    RECT 228.4000 302.2000 229.2000 306.8000 ;
	    RECT 231.6000 302.2000 232.4000 309.6000 ;
	    RECT 235.0000 308.4000 235.6000 311.8000 ;
	    RECT 236.4000 309.6000 237.2000 311.2000 ;
	    RECT 238.0000 310.3000 238.8000 310.4000 ;
	    RECT 239.6000 310.3000 240.4000 310.4000 ;
	    RECT 238.0000 309.7000 240.4000 310.3000 ;
	    RECT 238.0000 309.6000 238.8000 309.7000 ;
	    RECT 239.6000 308.8000 240.4000 309.7000 ;
	    RECT 241.2000 308.4000 241.8000 311.8000 ;
	    RECT 242.8000 308.8000 243.6000 310.4000 ;
	    RECT 234.8000 307.6000 235.6000 308.4000 ;
	    RECT 238.0000 308.2000 238.8000 308.4000 ;
	    RECT 241.2000 308.2000 242.0000 308.4000 ;
	    RECT 244.4000 308.3000 245.2000 309.2000 ;
	    RECT 246.0000 308.3000 246.8000 309.2000 ;
	    RECT 247.6000 308.8000 248.4000 310.4000 ;
	    RECT 249.4000 308.4000 250.0000 311.8000 ;
	    RECT 250.8000 310.3000 251.6000 310.4000 ;
	    RECT 250.8000 309.7000 254.7000 310.3000 ;
	    RECT 250.8000 308.8000 251.6000 309.7000 ;
	    RECT 238.0000 307.6000 239.6000 308.2000 ;
	    RECT 241.2000 307.6000 243.6000 308.2000 ;
	    RECT 244.4000 307.7000 246.8000 308.3000 ;
	    RECT 249.2000 308.2000 250.0000 308.4000 ;
	    RECT 252.4000 308.2000 253.2000 308.4000 ;
	    RECT 244.4000 307.6000 245.2000 307.7000 ;
	    RECT 246.0000 307.6000 246.8000 307.7000 ;
	    RECT 247.6000 307.6000 250.0000 308.2000 ;
	    RECT 251.6000 307.6000 253.2000 308.2000 ;
	    RECT 254.1000 308.3000 254.7000 309.7000 ;
	    RECT 260.4000 309.6000 261.2000 311.2000 ;
	    RECT 262.0000 308.4000 262.6000 311.8000 ;
	    RECT 265.2000 311.6000 266.0000 311.8000 ;
	    RECT 267.2000 308.4000 267.8000 311.8000 ;
	    RECT 268.4000 308.8000 269.2000 310.4000 ;
	    RECT 271.6000 310.3000 272.4000 310.4000 ;
	    RECT 273.2000 310.3000 274.0000 311.2000 ;
	    RECT 271.6000 309.7000 274.0000 310.3000 ;
	    RECT 271.6000 309.6000 272.4000 309.7000 ;
	    RECT 273.2000 309.6000 274.0000 309.7000 ;
	    RECT 274.6000 308.4000 275.2000 312.2000 ;
	    RECT 279.8000 311.6000 280.4000 315.0000 ;
	    RECT 276.6000 311.0000 280.4000 311.6000 ;
	    RECT 281.2000 315.0000 282.0000 319.0000 ;
	    RECT 281.2000 311.6000 281.8000 315.0000 ;
	    RECT 285.4000 312.8000 286.2000 319.8000 ;
	    RECT 285.4000 312.2000 287.0000 312.8000 ;
	    RECT 293.4000 312.4000 295.4000 319.8000 ;
	    RECT 281.2000 311.0000 285.0000 311.6000 ;
	    RECT 276.6000 309.0000 277.2000 311.0000 ;
	    RECT 262.0000 308.3000 262.8000 308.4000 ;
	    RECT 254.1000 307.7000 262.8000 308.3000 ;
	    RECT 262.0000 307.6000 262.8000 307.7000 ;
	    RECT 265.2000 307.6000 267.8000 308.4000 ;
	    RECT 270.0000 308.2000 270.8000 308.4000 ;
	    RECT 269.2000 307.6000 270.8000 308.2000 ;
	    RECT 273.2000 307.6000 275.2000 308.4000 ;
	    RECT 275.8000 308.2000 277.2000 309.0000 ;
	    RECT 278.0000 308.8000 278.8000 310.4000 ;
	    RECT 279.6000 308.8000 280.4000 310.4000 ;
	    RECT 281.2000 308.8000 282.0000 310.4000 ;
	    RECT 282.8000 308.8000 283.6000 310.4000 ;
	    RECT 284.4000 309.0000 285.0000 311.0000 ;
	    RECT 233.2000 304.8000 234.0000 306.4000 ;
	    RECT 235.0000 304.2000 235.6000 307.6000 ;
	    RECT 238.8000 307.2000 239.6000 307.6000 ;
	    RECT 238.2000 306.2000 241.8000 306.6000 ;
	    RECT 243.0000 306.2000 243.6000 307.6000 ;
	    RECT 247.6000 306.2000 248.2000 307.6000 ;
	    RECT 251.6000 307.2000 252.4000 307.6000 ;
	    RECT 249.4000 306.2000 253.0000 306.6000 ;
	    RECT 234.8000 302.2000 235.6000 304.2000 ;
	    RECT 238.0000 306.0000 242.0000 306.2000 ;
	    RECT 238.0000 302.2000 238.8000 306.0000 ;
	    RECT 241.2000 302.8000 242.0000 306.0000 ;
	    RECT 242.8000 303.4000 243.6000 306.2000 ;
	    RECT 244.4000 302.8000 245.2000 306.2000 ;
	    RECT 241.2000 302.2000 245.2000 302.8000 ;
	    RECT 246.0000 302.8000 246.8000 306.2000 ;
	    RECT 247.6000 303.4000 248.4000 306.2000 ;
	    RECT 249.2000 306.0000 253.2000 306.2000 ;
	    RECT 249.2000 302.8000 250.0000 306.0000 ;
	    RECT 246.0000 302.2000 250.0000 302.8000 ;
	    RECT 252.4000 302.2000 253.2000 306.0000 ;
	    RECT 262.0000 304.2000 262.6000 307.6000 ;
	    RECT 263.6000 304.8000 264.4000 306.4000 ;
	    RECT 265.4000 306.2000 266.0000 307.6000 ;
	    RECT 269.2000 307.2000 270.0000 307.6000 ;
	    RECT 274.6000 307.0000 275.2000 307.6000 ;
	    RECT 276.2000 307.8000 277.2000 308.2000 ;
	    RECT 284.4000 308.2000 285.8000 309.0000 ;
	    RECT 286.4000 308.4000 287.0000 312.2000 ;
	    RECT 292.4000 311.8000 295.4000 312.4000 ;
	    RECT 299.4000 312.6000 300.2000 319.8000 ;
	    RECT 299.4000 311.8000 301.2000 312.6000 ;
	    RECT 292.4000 311.6000 294.6000 311.8000 ;
	    RECT 287.6000 310.3000 288.4000 311.2000 ;
	    RECT 289.2000 310.3000 290.0000 310.4000 ;
	    RECT 287.6000 309.7000 290.0000 310.3000 ;
	    RECT 287.6000 309.6000 288.4000 309.7000 ;
	    RECT 289.2000 309.6000 290.0000 309.7000 ;
	    RECT 292.4000 308.8000 293.2000 310.4000 ;
	    RECT 294.0000 308.4000 294.6000 311.6000 ;
	    RECT 295.6000 308.8000 296.4000 310.4000 ;
	    RECT 298.8000 309.6000 299.6000 311.2000 ;
	    RECT 284.4000 307.8000 285.4000 308.2000 ;
	    RECT 276.2000 307.2000 280.4000 307.8000 ;
	    RECT 274.6000 306.6000 275.4000 307.0000 ;
	    RECT 267.0000 306.2000 270.6000 306.6000 ;
	    RECT 262.0000 302.2000 262.8000 304.2000 ;
	    RECT 265.2000 302.2000 266.0000 306.2000 ;
	    RECT 266.8000 306.0000 270.8000 306.2000 ;
	    RECT 274.6000 306.0000 276.2000 306.6000 ;
	    RECT 266.8000 302.2000 267.6000 306.0000 ;
	    RECT 270.0000 302.2000 270.8000 306.0000 ;
	    RECT 275.4000 303.0000 276.2000 306.0000 ;
	    RECT 279.8000 305.0000 280.4000 307.2000 ;
	    RECT 279.6000 303.0000 280.4000 305.0000 ;
	    RECT 281.2000 307.2000 285.4000 307.8000 ;
	    RECT 286.4000 307.6000 288.4000 308.4000 ;
	    RECT 290.8000 308.2000 291.6000 308.4000 ;
	    RECT 294.0000 308.2000 294.8000 308.4000 ;
	    RECT 290.8000 307.6000 292.4000 308.2000 ;
	    RECT 294.0000 307.6000 296.4000 308.2000 ;
	    RECT 297.2000 307.6000 298.0000 309.2000 ;
	    RECT 300.4000 308.4000 301.0000 311.8000 ;
	    RECT 303.6000 311.2000 304.4000 319.8000 ;
	    RECT 307.8000 315.8000 309.0000 319.8000 ;
	    RECT 312.4000 315.8000 313.2000 319.8000 ;
	    RECT 316.8000 316.4000 317.6000 319.8000 ;
	    RECT 316.8000 315.8000 318.8000 316.4000 ;
	    RECT 308.4000 315.0000 309.2000 315.8000 ;
	    RECT 312.6000 315.2000 313.2000 315.8000 ;
	    RECT 311.8000 314.6000 315.4000 315.2000 ;
	    RECT 318.0000 315.0000 318.8000 315.8000 ;
	    RECT 311.8000 314.4000 312.6000 314.6000 ;
	    RECT 314.6000 314.4000 315.4000 314.6000 ;
	    RECT 307.6000 313.2000 309.0000 314.0000 ;
	    RECT 308.4000 312.2000 309.0000 313.2000 ;
	    RECT 310.6000 313.0000 312.8000 313.6000 ;
	    RECT 310.6000 312.8000 311.4000 313.0000 ;
	    RECT 308.4000 311.6000 310.8000 312.2000 ;
	    RECT 303.6000 310.6000 307.8000 311.2000 ;
	    RECT 298.8000 308.3000 299.6000 308.4000 ;
	    RECT 300.4000 308.3000 301.2000 308.4000 ;
	    RECT 298.8000 307.7000 301.2000 308.3000 ;
	    RECT 298.8000 307.6000 299.6000 307.7000 ;
	    RECT 300.4000 307.6000 301.2000 307.7000 ;
	    RECT 281.2000 305.0000 281.8000 307.2000 ;
	    RECT 286.4000 307.0000 287.0000 307.6000 ;
	    RECT 291.6000 307.2000 292.4000 307.6000 ;
	    RECT 286.2000 306.6000 287.0000 307.0000 ;
	    RECT 285.4000 306.0000 287.0000 306.6000 ;
	    RECT 291.0000 306.2000 294.6000 306.6000 ;
	    RECT 295.8000 306.2000 296.4000 307.6000 ;
	    RECT 290.8000 306.0000 294.8000 306.2000 ;
	    RECT 281.2000 303.0000 282.0000 305.0000 ;
	    RECT 285.4000 303.0000 286.2000 306.0000 ;
	    RECT 290.8000 302.2000 291.6000 306.0000 ;
	    RECT 294.0000 302.8000 294.8000 306.0000 ;
	    RECT 295.6000 303.4000 296.4000 306.2000 ;
	    RECT 297.2000 302.8000 298.0000 306.2000 ;
	    RECT 294.0000 302.2000 298.0000 302.8000 ;
	    RECT 300.4000 304.2000 301.0000 307.6000 ;
	    RECT 303.6000 307.2000 304.4000 310.6000 ;
	    RECT 307.0000 310.4000 307.8000 310.6000 ;
	    RECT 305.4000 309.8000 306.2000 310.0000 ;
	    RECT 305.4000 309.2000 309.2000 309.8000 ;
	    RECT 308.4000 309.0000 309.2000 309.2000 ;
	    RECT 310.2000 308.4000 310.8000 311.6000 ;
	    RECT 312.2000 311.8000 312.8000 313.0000 ;
	    RECT 313.4000 313.0000 314.2000 313.2000 ;
	    RECT 318.0000 313.0000 318.8000 313.2000 ;
	    RECT 313.4000 312.4000 318.8000 313.0000 ;
	    RECT 312.2000 311.4000 317.0000 311.8000 ;
	    RECT 321.2000 311.4000 322.0000 319.8000 ;
	    RECT 312.2000 311.2000 322.0000 311.4000 ;
	    RECT 316.2000 311.0000 322.0000 311.2000 ;
	    RECT 316.4000 310.8000 322.0000 311.0000 ;
	    RECT 314.8000 310.2000 315.6000 310.4000 ;
	    RECT 324.4000 310.3000 325.2000 319.8000 ;
	    RECT 328.4000 313.6000 329.2000 314.4000 ;
	    RECT 326.0000 311.6000 326.8000 313.2000 ;
	    RECT 328.4000 312.4000 329.0000 313.6000 ;
	    RECT 329.8000 312.4000 330.6000 319.8000 ;
	    RECT 327.6000 311.8000 329.0000 312.4000 ;
	    RECT 329.6000 311.8000 330.6000 312.4000 ;
	    RECT 327.6000 311.6000 328.4000 311.8000 ;
	    RECT 327.7000 310.3000 328.3000 311.6000 ;
	    RECT 314.8000 309.6000 319.8000 310.2000 ;
	    RECT 316.4000 309.4000 317.2000 309.6000 ;
	    RECT 319.0000 309.4000 319.8000 309.6000 ;
	    RECT 324.4000 309.7000 328.3000 310.3000 ;
	    RECT 317.4000 308.4000 318.2000 308.6000 ;
	    RECT 310.2000 307.8000 321.2000 308.4000 ;
	    RECT 310.6000 307.6000 311.4000 307.8000 ;
	    RECT 303.6000 306.6000 307.4000 307.2000 ;
	    RECT 302.0000 304.8000 302.8000 306.4000 ;
	    RECT 300.4000 302.2000 301.2000 304.2000 ;
	    RECT 303.6000 302.2000 304.4000 306.6000 ;
	    RECT 306.6000 306.4000 307.4000 306.6000 ;
	    RECT 316.4000 306.4000 317.0000 307.8000 ;
	    RECT 319.6000 307.6000 321.2000 307.8000 ;
	    RECT 314.6000 305.4000 315.4000 305.6000 ;
	    RECT 308.4000 304.2000 309.2000 305.0000 ;
	    RECT 312.6000 304.8000 315.4000 305.4000 ;
	    RECT 316.4000 304.8000 317.2000 306.4000 ;
	    RECT 312.6000 304.2000 313.2000 304.8000 ;
	    RECT 318.0000 304.2000 318.8000 305.0000 ;
	    RECT 307.8000 303.6000 309.2000 304.2000 ;
	    RECT 307.8000 302.2000 309.0000 303.6000 ;
	    RECT 312.4000 302.2000 313.2000 304.2000 ;
	    RECT 316.8000 303.6000 318.8000 304.2000 ;
	    RECT 316.8000 302.2000 317.6000 303.6000 ;
	    RECT 321.2000 302.2000 322.0000 307.0000 ;
	    RECT 322.8000 306.8000 323.6000 308.4000 ;
	    RECT 324.4000 306.2000 325.2000 309.7000 ;
	    RECT 329.6000 308.4000 330.2000 311.8000 ;
	    RECT 330.8000 308.8000 331.6000 310.4000 ;
	    RECT 335.6000 310.3000 336.4000 319.8000 ;
	    RECT 339.6000 313.6000 340.4000 314.4000 ;
	    RECT 337.2000 311.6000 338.0000 313.2000 ;
	    RECT 339.6000 312.4000 340.2000 313.6000 ;
	    RECT 341.0000 312.4000 341.8000 319.8000 ;
	    RECT 338.8000 311.8000 340.2000 312.4000 ;
	    RECT 340.8000 311.8000 341.8000 312.4000 ;
	    RECT 338.8000 311.6000 339.6000 311.8000 ;
	    RECT 338.9000 310.3000 339.5000 311.6000 ;
	    RECT 340.8000 310.4000 341.4000 311.8000 ;
	    RECT 345.2000 311.2000 346.0000 319.8000 ;
	    RECT 349.4000 315.8000 350.6000 319.8000 ;
	    RECT 354.0000 315.8000 354.8000 319.8000 ;
	    RECT 358.4000 316.4000 359.2000 319.8000 ;
	    RECT 358.4000 315.8000 360.4000 316.4000 ;
	    RECT 350.0000 315.0000 350.8000 315.8000 ;
	    RECT 354.2000 315.2000 354.8000 315.8000 ;
	    RECT 353.4000 314.6000 357.0000 315.2000 ;
	    RECT 359.6000 315.0000 360.4000 315.8000 ;
	    RECT 353.4000 314.4000 354.2000 314.6000 ;
	    RECT 356.2000 314.4000 357.0000 314.6000 ;
	    RECT 349.2000 313.2000 350.6000 314.0000 ;
	    RECT 350.0000 312.2000 350.6000 313.2000 ;
	    RECT 352.2000 313.0000 354.4000 313.6000 ;
	    RECT 352.2000 312.8000 353.0000 313.0000 ;
	    RECT 350.0000 311.6000 352.4000 312.2000 ;
	    RECT 345.2000 310.6000 349.4000 311.2000 ;
	    RECT 335.6000 309.7000 339.5000 310.3000 ;
	    RECT 327.6000 307.6000 330.2000 308.4000 ;
	    RECT 332.4000 308.2000 333.2000 308.4000 ;
	    RECT 331.6000 307.6000 333.2000 308.2000 ;
	    RECT 327.8000 306.2000 328.4000 307.6000 ;
	    RECT 331.6000 307.2000 332.4000 307.6000 ;
	    RECT 334.0000 306.8000 334.8000 308.4000 ;
	    RECT 329.4000 306.2000 333.0000 306.6000 ;
	    RECT 335.6000 306.2000 336.4000 309.7000 ;
	    RECT 340.4000 309.6000 341.4000 310.4000 ;
	    RECT 340.8000 308.4000 341.4000 309.6000 ;
	    RECT 342.0000 308.8000 342.8000 310.4000 ;
	    RECT 338.8000 307.6000 341.4000 308.4000 ;
	    RECT 343.6000 308.2000 344.4000 308.4000 ;
	    RECT 342.8000 307.6000 344.4000 308.2000 ;
	    RECT 339.0000 306.2000 339.6000 307.6000 ;
	    RECT 342.8000 307.2000 343.6000 307.6000 ;
	    RECT 345.2000 307.2000 346.0000 310.6000 ;
	    RECT 348.6000 310.4000 349.4000 310.6000 ;
	    RECT 351.8000 310.3000 352.4000 311.6000 ;
	    RECT 353.8000 311.8000 354.4000 313.0000 ;
	    RECT 355.0000 313.0000 355.8000 313.2000 ;
	    RECT 359.6000 313.0000 360.4000 313.2000 ;
	    RECT 355.0000 312.4000 360.4000 313.0000 ;
	    RECT 353.8000 311.4000 358.6000 311.8000 ;
	    RECT 362.8000 311.4000 363.6000 319.8000 ;
	    RECT 353.8000 311.2000 363.6000 311.4000 ;
	    RECT 357.8000 311.0000 363.6000 311.2000 ;
	    RECT 358.0000 310.8000 363.6000 311.0000 ;
	    RECT 353.2000 310.3000 354.0000 310.4000 ;
	    RECT 347.0000 309.8000 347.8000 310.0000 ;
	    RECT 347.0000 309.2000 350.8000 309.8000 ;
	    RECT 351.7000 309.7000 354.0000 310.3000 ;
	    RECT 350.0000 309.0000 350.8000 309.2000 ;
	    RECT 351.8000 308.4000 352.4000 309.7000 ;
	    RECT 353.2000 309.6000 354.0000 309.7000 ;
	    RECT 356.4000 310.2000 357.2000 310.4000 ;
	    RECT 366.0000 310.3000 366.8000 319.8000 ;
	    RECT 370.0000 313.6000 370.8000 314.4000 ;
	    RECT 367.6000 311.6000 368.4000 313.2000 ;
	    RECT 370.0000 312.4000 370.6000 313.6000 ;
	    RECT 371.4000 312.4000 372.2000 319.8000 ;
	    RECT 369.2000 311.8000 370.6000 312.4000 ;
	    RECT 371.2000 311.8000 372.2000 312.4000 ;
	    RECT 369.2000 311.6000 370.0000 311.8000 ;
	    RECT 369.3000 310.3000 369.9000 311.6000 ;
	    RECT 356.4000 309.6000 361.4000 310.2000 ;
	    RECT 358.0000 309.4000 358.8000 309.6000 ;
	    RECT 360.6000 309.4000 361.4000 309.6000 ;
	    RECT 366.0000 309.7000 369.9000 310.3000 ;
	    RECT 359.0000 308.4000 359.8000 308.6000 ;
	    RECT 351.8000 307.8000 362.8000 308.4000 ;
	    RECT 352.2000 307.6000 353.0000 307.8000 ;
	    RECT 345.2000 306.6000 349.0000 307.2000 ;
	    RECT 340.6000 306.2000 344.2000 306.6000 ;
	    RECT 324.4000 305.6000 326.2000 306.2000 ;
	    RECT 325.4000 302.2000 326.2000 305.6000 ;
	    RECT 327.6000 302.2000 328.4000 306.2000 ;
	    RECT 329.2000 306.0000 333.2000 306.2000 ;
	    RECT 329.2000 302.2000 330.0000 306.0000 ;
	    RECT 332.4000 302.2000 333.2000 306.0000 ;
	    RECT 335.6000 305.6000 337.4000 306.2000 ;
	    RECT 336.6000 302.2000 337.4000 305.6000 ;
	    RECT 338.8000 302.2000 339.6000 306.2000 ;
	    RECT 340.4000 306.0000 344.4000 306.2000 ;
	    RECT 340.4000 302.2000 341.2000 306.0000 ;
	    RECT 343.6000 302.2000 344.4000 306.0000 ;
	    RECT 345.2000 302.2000 346.0000 306.6000 ;
	    RECT 348.2000 306.4000 349.0000 306.6000 ;
	    RECT 358.0000 305.6000 358.6000 307.8000 ;
	    RECT 361.2000 307.6000 362.8000 307.8000 ;
	    RECT 356.2000 305.4000 357.0000 305.6000 ;
	    RECT 350.0000 304.2000 350.8000 305.0000 ;
	    RECT 354.2000 304.8000 357.0000 305.4000 ;
	    RECT 358.0000 304.8000 358.8000 305.6000 ;
	    RECT 354.2000 304.2000 354.8000 304.8000 ;
	    RECT 359.6000 304.2000 360.4000 305.0000 ;
	    RECT 349.4000 303.6000 350.8000 304.2000 ;
	    RECT 349.4000 302.2000 350.6000 303.6000 ;
	    RECT 354.0000 302.2000 354.8000 304.2000 ;
	    RECT 358.4000 303.6000 360.4000 304.2000 ;
	    RECT 358.4000 302.2000 359.2000 303.6000 ;
	    RECT 362.8000 302.2000 363.6000 307.0000 ;
	    RECT 364.4000 306.8000 365.2000 308.4000 ;
	    RECT 366.0000 306.2000 366.8000 309.7000 ;
	    RECT 371.2000 308.4000 371.8000 311.8000 ;
	    RECT 375.6000 311.2000 376.4000 319.8000 ;
	    RECT 379.8000 315.8000 381.0000 319.8000 ;
	    RECT 384.4000 315.8000 385.2000 319.8000 ;
	    RECT 388.8000 316.4000 389.6000 319.8000 ;
	    RECT 388.8000 315.8000 390.8000 316.4000 ;
	    RECT 380.4000 315.0000 381.2000 315.8000 ;
	    RECT 384.6000 315.2000 385.2000 315.8000 ;
	    RECT 383.8000 314.6000 387.4000 315.2000 ;
	    RECT 390.0000 315.0000 390.8000 315.8000 ;
	    RECT 383.8000 314.4000 384.6000 314.6000 ;
	    RECT 386.6000 314.4000 387.4000 314.6000 ;
	    RECT 378.8000 314.0000 380.2000 314.4000 ;
	    RECT 378.8000 313.6000 381.0000 314.0000 ;
	    RECT 379.6000 313.2000 381.0000 313.6000 ;
	    RECT 380.4000 312.2000 381.0000 313.2000 ;
	    RECT 382.6000 313.0000 384.8000 313.6000 ;
	    RECT 382.6000 312.8000 383.4000 313.0000 ;
	    RECT 380.4000 311.6000 382.8000 312.2000 ;
	    RECT 375.6000 310.6000 379.8000 311.2000 ;
	    RECT 372.4000 308.8000 373.2000 310.4000 ;
	    RECT 367.6000 308.3000 368.4000 308.4000 ;
	    RECT 369.2000 308.3000 371.8000 308.4000 ;
	    RECT 367.6000 307.7000 371.8000 308.3000 ;
	    RECT 374.0000 308.2000 374.8000 308.4000 ;
	    RECT 367.6000 307.6000 368.4000 307.7000 ;
	    RECT 369.2000 307.6000 371.8000 307.7000 ;
	    RECT 373.2000 307.6000 374.8000 308.2000 ;
	    RECT 369.4000 306.2000 370.0000 307.6000 ;
	    RECT 373.2000 307.2000 374.0000 307.6000 ;
	    RECT 375.6000 307.2000 376.4000 310.6000 ;
	    RECT 379.0000 310.4000 379.8000 310.6000 ;
	    RECT 377.4000 309.8000 378.2000 310.0000 ;
	    RECT 377.4000 309.2000 381.2000 309.8000 ;
	    RECT 380.4000 309.0000 381.2000 309.2000 ;
	    RECT 382.2000 308.4000 382.8000 311.6000 ;
	    RECT 384.2000 311.8000 384.8000 313.0000 ;
	    RECT 385.4000 313.0000 386.2000 313.2000 ;
	    RECT 390.0000 313.0000 390.8000 313.2000 ;
	    RECT 385.4000 312.4000 390.8000 313.0000 ;
	    RECT 384.2000 311.4000 389.0000 311.8000 ;
	    RECT 393.2000 311.4000 394.0000 319.8000 ;
	    RECT 396.4000 315.8000 397.2000 319.8000 ;
	    RECT 396.6000 315.6000 397.2000 315.8000 ;
	    RECT 399.6000 315.8000 400.4000 319.8000 ;
	    RECT 399.6000 315.6000 400.2000 315.8000 ;
	    RECT 396.6000 315.0000 400.2000 315.6000 ;
	    RECT 398.0000 312.8000 398.8000 314.4000 ;
	    RECT 384.2000 311.2000 394.0000 311.4000 ;
	    RECT 388.2000 311.0000 394.0000 311.2000 ;
	    RECT 388.4000 310.8000 394.0000 311.0000 ;
	    RECT 399.6000 312.4000 400.2000 315.0000 ;
	    RECT 399.6000 311.6000 400.4000 312.4000 ;
	    RECT 386.8000 310.2000 387.6000 310.4000 ;
	    RECT 386.8000 309.6000 391.8000 310.2000 ;
	    RECT 396.4000 309.6000 398.0000 310.4000 ;
	    RECT 388.4000 309.4000 389.2000 309.6000 ;
	    RECT 391.0000 309.4000 391.8000 309.6000 ;
	    RECT 389.4000 308.4000 390.2000 308.6000 ;
	    RECT 399.6000 308.4000 400.2000 311.6000 ;
	    RECT 382.2000 307.8000 393.2000 308.4000 ;
	    RECT 398.6000 308.2000 400.2000 308.4000 ;
	    RECT 382.6000 307.6000 383.4000 307.8000 ;
	    RECT 375.6000 306.6000 379.4000 307.2000 ;
	    RECT 371.0000 306.2000 374.6000 306.6000 ;
	    RECT 366.0000 305.6000 367.8000 306.2000 ;
	    RECT 367.0000 302.2000 367.8000 305.6000 ;
	    RECT 369.2000 302.2000 370.0000 306.2000 ;
	    RECT 370.8000 306.0000 374.8000 306.2000 ;
	    RECT 370.8000 302.2000 371.6000 306.0000 ;
	    RECT 374.0000 302.2000 374.8000 306.0000 ;
	    RECT 375.6000 302.2000 376.4000 306.6000 ;
	    RECT 378.6000 306.4000 379.4000 306.6000 ;
	    RECT 388.4000 305.6000 389.0000 307.8000 ;
	    RECT 391.6000 307.6000 393.2000 307.8000 ;
	    RECT 398.4000 307.8000 400.2000 308.2000 ;
	    RECT 407.6000 311.2000 408.4000 319.8000 ;
	    RECT 411.8000 315.8000 413.0000 319.8000 ;
	    RECT 416.4000 315.8000 417.2000 319.8000 ;
	    RECT 420.8000 316.4000 421.6000 319.8000 ;
	    RECT 420.8000 315.8000 422.8000 316.4000 ;
	    RECT 412.4000 315.0000 413.2000 315.8000 ;
	    RECT 416.6000 315.2000 417.2000 315.8000 ;
	    RECT 415.8000 314.6000 419.4000 315.2000 ;
	    RECT 422.0000 315.0000 422.8000 315.8000 ;
	    RECT 415.8000 314.4000 416.6000 314.6000 ;
	    RECT 418.6000 314.4000 419.4000 314.6000 ;
	    RECT 411.6000 313.2000 413.0000 314.0000 ;
	    RECT 412.4000 312.2000 413.0000 313.2000 ;
	    RECT 414.6000 313.0000 416.8000 313.6000 ;
	    RECT 414.6000 312.8000 415.4000 313.0000 ;
	    RECT 412.4000 311.6000 414.8000 312.2000 ;
	    RECT 407.6000 310.6000 411.8000 311.2000 ;
	    RECT 386.6000 305.4000 387.4000 305.6000 ;
	    RECT 380.4000 304.2000 381.2000 305.0000 ;
	    RECT 384.6000 304.8000 387.4000 305.4000 ;
	    RECT 388.4000 304.8000 389.2000 305.6000 ;
	    RECT 384.6000 304.2000 385.2000 304.8000 ;
	    RECT 390.0000 304.2000 390.8000 305.0000 ;
	    RECT 379.8000 303.6000 381.2000 304.2000 ;
	    RECT 379.8000 302.2000 381.0000 303.6000 ;
	    RECT 384.4000 302.2000 385.2000 304.2000 ;
	    RECT 388.8000 303.6000 390.8000 304.2000 ;
	    RECT 388.8000 302.2000 389.6000 303.6000 ;
	    RECT 393.2000 302.2000 394.0000 307.0000 ;
	    RECT 398.4000 302.2000 399.2000 307.8000 ;
	    RECT 407.6000 307.2000 408.4000 310.6000 ;
	    RECT 411.0000 310.4000 411.8000 310.6000 ;
	    RECT 409.4000 309.8000 410.2000 310.0000 ;
	    RECT 409.4000 309.2000 413.2000 309.8000 ;
	    RECT 412.4000 309.0000 413.2000 309.2000 ;
	    RECT 414.2000 308.4000 414.8000 311.6000 ;
	    RECT 416.2000 311.8000 416.8000 313.0000 ;
	    RECT 417.4000 313.0000 418.2000 313.2000 ;
	    RECT 422.0000 313.0000 422.8000 313.2000 ;
	    RECT 417.4000 312.4000 422.8000 313.0000 ;
	    RECT 416.2000 311.4000 421.0000 311.8000 ;
	    RECT 425.2000 311.4000 426.0000 319.8000 ;
	    RECT 427.6000 313.6000 428.4000 314.4000 ;
	    RECT 427.6000 312.4000 428.2000 313.6000 ;
	    RECT 429.0000 312.4000 429.8000 319.8000 ;
	    RECT 426.8000 311.8000 428.2000 312.4000 ;
	    RECT 426.8000 311.6000 427.6000 311.8000 ;
	    RECT 428.8000 311.6000 430.8000 312.4000 ;
	    RECT 416.2000 311.2000 426.0000 311.4000 ;
	    RECT 420.2000 311.0000 426.0000 311.2000 ;
	    RECT 420.4000 310.8000 426.0000 311.0000 ;
	    RECT 418.8000 310.2000 419.6000 310.4000 ;
	    RECT 418.8000 309.6000 423.8000 310.2000 ;
	    RECT 420.4000 309.4000 421.2000 309.6000 ;
	    RECT 423.0000 309.4000 423.8000 309.6000 ;
	    RECT 421.4000 308.4000 422.2000 308.6000 ;
	    RECT 428.8000 308.4000 429.4000 311.6000 ;
	    RECT 430.0000 310.3000 430.8000 310.4000 ;
	    RECT 431.6000 310.3000 432.4000 310.4000 ;
	    RECT 430.0000 309.7000 432.4000 310.3000 ;
	    RECT 430.0000 308.8000 430.8000 309.7000 ;
	    RECT 431.6000 309.6000 432.4000 309.7000 ;
	    RECT 414.2000 307.8000 425.2000 308.4000 ;
	    RECT 414.6000 307.6000 415.4000 307.8000 ;
	    RECT 418.8000 307.6000 419.6000 307.8000 ;
	    RECT 407.6000 306.6000 411.4000 307.2000 ;
	    RECT 407.6000 302.2000 408.4000 306.6000 ;
	    RECT 410.6000 306.4000 411.4000 306.6000 ;
	    RECT 420.4000 305.6000 421.0000 307.8000 ;
	    RECT 423.6000 307.6000 425.2000 307.8000 ;
	    RECT 426.8000 307.6000 429.4000 308.4000 ;
	    RECT 431.6000 308.3000 432.4000 308.4000 ;
	    RECT 433.2000 308.3000 434.0000 319.8000 ;
	    RECT 434.8000 314.3000 435.6000 314.4000 ;
	    RECT 436.4000 314.3000 437.2000 319.8000 ;
	    RECT 440.6000 315.8000 441.8000 319.8000 ;
	    RECT 445.2000 315.8000 446.0000 319.8000 ;
	    RECT 449.6000 316.4000 450.4000 319.8000 ;
	    RECT 449.6000 315.8000 451.6000 316.4000 ;
	    RECT 441.2000 315.0000 442.0000 315.8000 ;
	    RECT 445.4000 315.2000 446.0000 315.8000 ;
	    RECT 444.6000 314.6000 448.2000 315.2000 ;
	    RECT 450.8000 315.0000 451.6000 315.8000 ;
	    RECT 444.6000 314.4000 445.4000 314.6000 ;
	    RECT 447.4000 314.4000 448.2000 314.6000 ;
	    RECT 434.8000 313.7000 437.2000 314.3000 ;
	    RECT 434.8000 313.6000 435.6000 313.7000 ;
	    RECT 431.6000 308.2000 434.0000 308.3000 ;
	    RECT 430.8000 307.7000 434.0000 308.2000 ;
	    RECT 430.8000 307.6000 432.4000 307.7000 ;
	    RECT 418.6000 305.4000 419.4000 305.6000 ;
	    RECT 412.4000 304.2000 413.2000 305.0000 ;
	    RECT 416.6000 304.8000 419.4000 305.4000 ;
	    RECT 420.4000 304.8000 421.2000 305.6000 ;
	    RECT 416.6000 304.2000 417.2000 304.8000 ;
	    RECT 422.0000 304.2000 422.8000 305.0000 ;
	    RECT 411.8000 303.6000 413.2000 304.2000 ;
	    RECT 411.8000 302.2000 413.0000 303.6000 ;
	    RECT 416.4000 302.2000 417.2000 304.2000 ;
	    RECT 420.8000 303.6000 422.8000 304.2000 ;
	    RECT 420.8000 302.2000 421.6000 303.6000 ;
	    RECT 425.2000 302.2000 426.0000 307.0000 ;
	    RECT 427.0000 306.2000 427.6000 307.6000 ;
	    RECT 430.8000 307.2000 431.6000 307.6000 ;
	    RECT 428.6000 306.2000 432.2000 306.6000 ;
	    RECT 426.8000 302.2000 427.6000 306.2000 ;
	    RECT 428.4000 306.0000 432.4000 306.2000 ;
	    RECT 428.4000 302.2000 429.2000 306.0000 ;
	    RECT 431.6000 302.2000 432.4000 306.0000 ;
	    RECT 433.2000 302.2000 434.0000 307.7000 ;
	    RECT 436.4000 311.2000 437.2000 313.7000 ;
	    RECT 440.4000 313.2000 441.8000 314.0000 ;
	    RECT 441.2000 312.2000 441.8000 313.2000 ;
	    RECT 443.4000 313.0000 445.6000 313.6000 ;
	    RECT 443.4000 312.8000 444.2000 313.0000 ;
	    RECT 441.2000 311.6000 443.6000 312.2000 ;
	    RECT 436.4000 310.6000 440.6000 311.2000 ;
	    RECT 436.4000 307.2000 437.2000 310.6000 ;
	    RECT 439.8000 310.4000 440.6000 310.6000 ;
	    RECT 438.2000 309.8000 439.0000 310.0000 ;
	    RECT 438.2000 309.2000 442.0000 309.8000 ;
	    RECT 441.2000 309.0000 442.0000 309.2000 ;
	    RECT 443.0000 308.4000 443.6000 311.6000 ;
	    RECT 445.0000 311.8000 445.6000 313.0000 ;
	    RECT 446.2000 313.0000 447.0000 313.2000 ;
	    RECT 450.8000 313.0000 451.6000 313.2000 ;
	    RECT 446.2000 312.4000 451.6000 313.0000 ;
	    RECT 445.0000 311.4000 449.8000 311.8000 ;
	    RECT 454.0000 311.4000 454.8000 319.8000 ;
	    RECT 445.0000 311.2000 454.8000 311.4000 ;
	    RECT 449.0000 311.0000 454.8000 311.2000 ;
	    RECT 449.2000 310.8000 454.8000 311.0000 ;
	    RECT 446.0000 310.3000 446.8000 310.4000 ;
	    RECT 447.6000 310.3000 448.4000 310.4000 ;
	    RECT 446.0000 310.2000 448.4000 310.3000 ;
	    RECT 446.0000 309.7000 452.6000 310.2000 ;
	    RECT 446.0000 309.6000 446.8000 309.7000 ;
	    RECT 447.6000 309.6000 452.6000 309.7000 ;
	    RECT 451.8000 309.4000 452.6000 309.6000 ;
	    RECT 450.2000 308.4000 451.0000 308.6000 ;
	    RECT 443.0000 307.8000 454.0000 308.4000 ;
	    RECT 443.4000 307.6000 444.2000 307.8000 ;
	    RECT 436.4000 306.6000 440.2000 307.2000 ;
	    RECT 434.8000 304.8000 435.6000 306.4000 ;
	    RECT 436.4000 302.2000 437.2000 306.6000 ;
	    RECT 439.4000 306.4000 440.2000 306.6000 ;
	    RECT 449.2000 305.6000 449.8000 307.8000 ;
	    RECT 452.4000 307.6000 454.0000 307.8000 ;
	    RECT 447.4000 305.4000 448.2000 305.6000 ;
	    RECT 441.2000 304.2000 442.0000 305.0000 ;
	    RECT 445.4000 304.8000 448.2000 305.4000 ;
	    RECT 449.2000 304.8000 450.0000 305.6000 ;
	    RECT 445.4000 304.2000 446.0000 304.8000 ;
	    RECT 450.8000 304.2000 451.6000 305.0000 ;
	    RECT 440.6000 303.6000 442.0000 304.2000 ;
	    RECT 440.6000 302.2000 441.8000 303.6000 ;
	    RECT 445.2000 302.2000 446.0000 304.2000 ;
	    RECT 449.6000 303.6000 451.6000 304.2000 ;
	    RECT 449.6000 302.2000 450.4000 303.6000 ;
	    RECT 454.0000 302.2000 454.8000 307.0000 ;
	    RECT 455.6000 302.2000 456.4000 319.8000 ;
	    RECT 458.8000 311.2000 459.6000 319.8000 ;
	    RECT 463.0000 315.8000 464.2000 319.8000 ;
	    RECT 467.6000 315.8000 468.4000 319.8000 ;
	    RECT 472.0000 316.4000 472.8000 319.8000 ;
	    RECT 472.0000 315.8000 474.0000 316.4000 ;
	    RECT 463.6000 315.0000 464.4000 315.8000 ;
	    RECT 467.8000 315.2000 468.4000 315.8000 ;
	    RECT 467.0000 314.6000 470.6000 315.2000 ;
	    RECT 473.2000 315.0000 474.0000 315.8000 ;
	    RECT 467.0000 314.4000 467.8000 314.6000 ;
	    RECT 469.8000 314.4000 470.6000 314.6000 ;
	    RECT 462.8000 313.2000 464.2000 314.0000 ;
	    RECT 463.6000 312.2000 464.2000 313.2000 ;
	    RECT 465.8000 313.0000 468.0000 313.6000 ;
	    RECT 465.8000 312.8000 466.6000 313.0000 ;
	    RECT 463.6000 311.6000 466.0000 312.2000 ;
	    RECT 458.8000 310.6000 463.0000 311.2000 ;
	    RECT 458.8000 307.2000 459.6000 310.6000 ;
	    RECT 462.2000 310.4000 463.0000 310.6000 ;
	    RECT 460.6000 309.8000 461.4000 310.0000 ;
	    RECT 460.6000 309.2000 464.4000 309.8000 ;
	    RECT 463.6000 309.0000 464.4000 309.2000 ;
	    RECT 465.4000 308.4000 466.0000 311.6000 ;
	    RECT 467.4000 311.8000 468.0000 313.0000 ;
	    RECT 468.6000 313.0000 469.4000 313.2000 ;
	    RECT 473.2000 313.0000 474.0000 313.2000 ;
	    RECT 468.6000 312.4000 474.0000 313.0000 ;
	    RECT 467.4000 311.4000 472.2000 311.8000 ;
	    RECT 476.4000 311.4000 477.2000 319.8000 ;
	    RECT 478.8000 313.6000 479.6000 314.4000 ;
	    RECT 478.8000 312.4000 479.4000 313.6000 ;
	    RECT 480.2000 312.4000 481.0000 319.8000 ;
	    RECT 478.0000 311.8000 479.4000 312.4000 ;
	    RECT 480.0000 311.8000 481.0000 312.4000 ;
	    RECT 478.0000 311.6000 478.8000 311.8000 ;
	    RECT 467.4000 311.2000 477.2000 311.4000 ;
	    RECT 471.4000 311.0000 477.2000 311.2000 ;
	    RECT 471.6000 310.8000 477.2000 311.0000 ;
	    RECT 470.0000 310.2000 470.8000 310.4000 ;
	    RECT 478.0000 310.3000 478.8000 310.4000 ;
	    RECT 480.0000 310.3000 480.6000 311.8000 ;
	    RECT 470.0000 309.6000 475.0000 310.2000 ;
	    RECT 478.0000 309.7000 480.6000 310.3000 ;
	    RECT 478.0000 309.6000 478.8000 309.7000 ;
	    RECT 471.6000 309.4000 472.4000 309.6000 ;
	    RECT 474.2000 309.4000 475.0000 309.6000 ;
	    RECT 472.6000 308.4000 473.4000 308.6000 ;
	    RECT 480.0000 308.4000 480.6000 309.7000 ;
	    RECT 481.2000 310.3000 482.0000 310.4000 ;
	    RECT 482.8000 310.3000 483.6000 310.4000 ;
	    RECT 481.2000 309.7000 483.6000 310.3000 ;
	    RECT 481.2000 308.8000 482.0000 309.7000 ;
	    RECT 482.8000 309.6000 483.6000 309.7000 ;
	    RECT 465.2000 307.8000 476.4000 308.4000 ;
	    RECT 465.2000 307.6000 466.6000 307.8000 ;
	    RECT 458.8000 306.6000 462.6000 307.2000 ;
	    RECT 458.8000 302.2000 459.6000 306.6000 ;
	    RECT 461.8000 306.4000 462.6000 306.6000 ;
	    RECT 471.6000 305.6000 472.2000 307.8000 ;
	    RECT 474.8000 307.6000 476.4000 307.8000 ;
	    RECT 478.0000 307.6000 480.6000 308.4000 ;
	    RECT 482.8000 308.3000 483.6000 308.4000 ;
	    RECT 484.4000 308.3000 485.2000 319.8000 ;
	    RECT 482.8000 308.2000 485.2000 308.3000 ;
	    RECT 482.0000 307.7000 485.2000 308.2000 ;
	    RECT 482.0000 307.6000 483.6000 307.7000 ;
	    RECT 469.8000 305.4000 470.6000 305.6000 ;
	    RECT 463.6000 304.2000 464.4000 305.0000 ;
	    RECT 467.8000 304.8000 470.6000 305.4000 ;
	    RECT 471.6000 304.8000 472.4000 305.6000 ;
	    RECT 467.8000 304.2000 468.4000 304.8000 ;
	    RECT 473.2000 304.2000 474.0000 305.0000 ;
	    RECT 463.0000 303.6000 464.4000 304.2000 ;
	    RECT 463.0000 302.2000 464.2000 303.6000 ;
	    RECT 467.6000 302.2000 468.4000 304.2000 ;
	    RECT 472.0000 303.6000 474.0000 304.2000 ;
	    RECT 472.0000 302.2000 472.8000 303.6000 ;
	    RECT 476.4000 302.2000 477.2000 307.0000 ;
	    RECT 478.2000 306.2000 478.8000 307.6000 ;
	    RECT 482.0000 307.2000 482.8000 307.6000 ;
	    RECT 479.8000 306.2000 483.4000 306.6000 ;
	    RECT 478.0000 302.2000 478.8000 306.2000 ;
	    RECT 479.6000 306.0000 483.6000 306.2000 ;
	    RECT 479.6000 302.2000 480.4000 306.0000 ;
	    RECT 482.8000 302.2000 483.6000 306.0000 ;
	    RECT 484.4000 302.2000 485.2000 307.7000 ;
	    RECT 486.0000 304.8000 486.8000 306.4000 ;
	    RECT 487.6000 304.8000 488.4000 306.4000 ;
	    RECT 489.2000 302.2000 490.0000 319.8000 ;
	    RECT 492.4000 311.2000 493.2000 319.8000 ;
	    RECT 495.6000 311.2000 496.4000 319.8000 ;
	    RECT 498.8000 311.2000 499.6000 319.8000 ;
	    RECT 502.0000 311.2000 502.8000 319.8000 ;
	    RECT 505.2000 312.4000 506.0000 319.8000 ;
	    RECT 505.2000 311.8000 507.4000 312.4000 ;
	    RECT 508.4000 311.8000 509.2000 319.8000 ;
	    RECT 490.8000 310.4000 493.2000 311.2000 ;
	    RECT 494.2000 310.4000 496.4000 311.2000 ;
	    RECT 497.4000 310.4000 499.6000 311.2000 ;
	    RECT 501.0000 310.4000 502.8000 311.2000 ;
	    RECT 506.8000 311.2000 507.4000 311.8000 ;
	    RECT 506.8000 310.4000 508.0000 311.2000 ;
	    RECT 490.8000 307.6000 491.6000 310.4000 ;
	    RECT 494.2000 309.0000 495.0000 310.4000 ;
	    RECT 497.4000 309.0000 498.2000 310.4000 ;
	    RECT 501.0000 309.0000 501.8000 310.4000 ;
	    RECT 492.4000 308.2000 495.0000 309.0000 ;
	    RECT 495.8000 308.2000 498.2000 309.0000 ;
	    RECT 499.2000 308.2000 501.8000 309.0000 ;
	    RECT 505.2000 308.8000 506.0000 310.4000 ;
	    RECT 494.2000 307.6000 495.0000 308.2000 ;
	    RECT 497.4000 307.6000 498.2000 308.2000 ;
	    RECT 501.0000 307.6000 501.8000 308.2000 ;
	    RECT 490.8000 306.8000 493.2000 307.6000 ;
	    RECT 494.2000 306.8000 496.4000 307.6000 ;
	    RECT 497.4000 306.8000 499.6000 307.6000 ;
	    RECT 501.0000 306.8000 502.8000 307.6000 ;
	    RECT 506.8000 307.4000 507.4000 310.4000 ;
	    RECT 508.6000 309.6000 509.2000 311.8000 ;
	    RECT 492.4000 302.2000 493.2000 306.8000 ;
	    RECT 495.6000 302.2000 496.4000 306.8000 ;
	    RECT 498.8000 302.2000 499.6000 306.8000 ;
	    RECT 502.0000 302.2000 502.8000 306.8000 ;
	    RECT 505.2000 306.8000 507.4000 307.4000 ;
	    RECT 505.2000 302.2000 506.0000 306.8000 ;
	    RECT 508.4000 302.2000 509.2000 309.6000 ;
	    RECT 1.2000 295.4000 2.0000 299.8000 ;
	    RECT 5.4000 298.4000 6.6000 299.8000 ;
	    RECT 5.4000 297.8000 6.8000 298.4000 ;
	    RECT 10.0000 297.8000 10.8000 299.8000 ;
	    RECT 14.4000 298.4000 15.2000 299.8000 ;
	    RECT 14.4000 297.8000 16.4000 298.4000 ;
	    RECT 6.0000 297.0000 6.8000 297.8000 ;
	    RECT 10.2000 297.2000 10.8000 297.8000 ;
	    RECT 10.2000 296.6000 13.0000 297.2000 ;
	    RECT 12.2000 296.4000 13.0000 296.6000 ;
	    RECT 14.0000 296.4000 14.8000 297.2000 ;
	    RECT 15.6000 297.0000 16.4000 297.8000 ;
	    RECT 4.2000 295.4000 5.0000 295.6000 ;
	    RECT 1.2000 294.8000 5.0000 295.4000 ;
	    RECT 1.2000 291.4000 2.0000 294.8000 ;
	    RECT 8.2000 294.2000 9.0000 294.4000 ;
	    RECT 12.4000 294.2000 13.2000 294.4000 ;
	    RECT 14.0000 294.2000 14.6000 296.4000 ;
	    RECT 18.8000 295.0000 19.6000 299.8000 ;
	    RECT 20.4000 295.4000 21.2000 299.8000 ;
	    RECT 24.6000 298.4000 25.8000 299.8000 ;
	    RECT 24.6000 297.8000 26.0000 298.4000 ;
	    RECT 29.2000 297.8000 30.0000 299.8000 ;
	    RECT 33.6000 298.4000 34.4000 299.8000 ;
	    RECT 33.6000 297.8000 35.6000 298.4000 ;
	    RECT 25.2000 297.0000 26.0000 297.8000 ;
	    RECT 29.4000 297.2000 30.0000 297.8000 ;
	    RECT 29.4000 296.6000 32.2000 297.2000 ;
	    RECT 31.4000 296.4000 32.2000 296.6000 ;
	    RECT 33.2000 296.4000 34.0000 297.2000 ;
	    RECT 34.8000 297.0000 35.6000 297.8000 ;
	    RECT 23.4000 295.4000 24.2000 295.6000 ;
	    RECT 20.4000 294.8000 24.2000 295.4000 ;
	    RECT 17.2000 294.2000 18.8000 294.4000 ;
	    RECT 7.8000 293.6000 18.8000 294.2000 ;
	    RECT 6.0000 292.8000 6.8000 293.0000 ;
	    RECT 3.0000 292.2000 6.8000 292.8000 ;
	    RECT 3.0000 292.0000 3.8000 292.2000 ;
	    RECT 4.6000 291.4000 5.4000 291.6000 ;
	    RECT 1.2000 290.8000 5.4000 291.4000 ;
	    RECT 1.2000 282.2000 2.0000 290.8000 ;
	    RECT 7.8000 290.4000 8.4000 293.6000 ;
	    RECT 15.0000 293.4000 15.8000 293.6000 ;
	    RECT 14.0000 292.4000 14.8000 292.6000 ;
	    RECT 16.6000 292.4000 17.4000 292.6000 ;
	    RECT 12.4000 291.8000 17.4000 292.4000 ;
	    RECT 12.4000 291.6000 13.2000 291.8000 ;
	    RECT 20.4000 291.4000 21.2000 294.8000 ;
	    RECT 27.4000 294.2000 28.2000 294.4000 ;
	    RECT 33.2000 294.2000 33.8000 296.4000 ;
	    RECT 38.0000 295.0000 38.8000 299.8000 ;
	    RECT 39.6000 295.4000 40.4000 299.8000 ;
	    RECT 43.8000 298.4000 45.0000 299.8000 ;
	    RECT 43.8000 297.8000 45.2000 298.4000 ;
	    RECT 48.4000 297.8000 49.2000 299.8000 ;
	    RECT 52.8000 298.4000 53.6000 299.8000 ;
	    RECT 52.8000 297.8000 54.8000 298.4000 ;
	    RECT 44.4000 297.0000 45.2000 297.8000 ;
	    RECT 48.6000 297.2000 49.2000 297.8000 ;
	    RECT 48.6000 296.6000 51.4000 297.2000 ;
	    RECT 50.6000 296.4000 51.4000 296.6000 ;
	    RECT 52.4000 296.4000 53.2000 297.2000 ;
	    RECT 54.0000 297.0000 54.8000 297.8000 ;
	    RECT 42.6000 295.4000 43.4000 295.6000 ;
	    RECT 39.6000 294.8000 43.4000 295.4000 ;
	    RECT 36.4000 294.2000 38.0000 294.4000 ;
	    RECT 27.0000 293.6000 38.0000 294.2000 ;
	    RECT 25.2000 292.8000 26.0000 293.0000 ;
	    RECT 22.2000 292.2000 26.0000 292.8000 ;
	    RECT 27.0000 292.4000 27.6000 293.6000 ;
	    RECT 34.2000 293.4000 35.0000 293.6000 ;
	    RECT 33.2000 292.4000 34.0000 292.6000 ;
	    RECT 35.8000 292.4000 36.6000 292.6000 ;
	    RECT 22.2000 292.0000 23.0000 292.2000 ;
	    RECT 26.8000 291.6000 27.6000 292.4000 ;
	    RECT 31.6000 291.8000 36.6000 292.4000 ;
	    RECT 31.6000 291.6000 32.4000 291.8000 ;
	    RECT 23.8000 291.4000 24.6000 291.6000 ;
	    RECT 14.0000 291.0000 19.6000 291.2000 ;
	    RECT 13.8000 290.8000 19.6000 291.0000 ;
	    RECT 6.0000 289.8000 8.4000 290.4000 ;
	    RECT 9.8000 290.6000 19.6000 290.8000 ;
	    RECT 9.8000 290.2000 14.6000 290.6000 ;
	    RECT 6.0000 288.8000 6.6000 289.8000 ;
	    RECT 5.2000 288.0000 6.6000 288.8000 ;
	    RECT 8.2000 289.0000 9.0000 289.2000 ;
	    RECT 9.8000 289.0000 10.4000 290.2000 ;
	    RECT 8.2000 288.4000 10.4000 289.0000 ;
	    RECT 11.0000 289.0000 16.4000 289.6000 ;
	    RECT 11.0000 288.8000 11.8000 289.0000 ;
	    RECT 15.6000 288.8000 16.4000 289.0000 ;
	    RECT 9.4000 287.4000 10.2000 287.6000 ;
	    RECT 12.2000 287.4000 13.0000 287.6000 ;
	    RECT 6.0000 286.2000 6.8000 287.0000 ;
	    RECT 9.4000 286.8000 13.0000 287.4000 ;
	    RECT 10.2000 286.2000 10.8000 286.8000 ;
	    RECT 15.6000 286.2000 16.4000 287.0000 ;
	    RECT 5.4000 282.2000 6.6000 286.2000 ;
	    RECT 10.0000 282.2000 10.8000 286.2000 ;
	    RECT 14.4000 285.6000 16.4000 286.2000 ;
	    RECT 14.4000 282.2000 15.2000 285.6000 ;
	    RECT 18.8000 282.2000 19.6000 290.6000 ;
	    RECT 20.4000 290.8000 24.6000 291.4000 ;
	    RECT 20.4000 282.2000 21.2000 290.8000 ;
	    RECT 27.0000 290.4000 27.6000 291.6000 ;
	    RECT 39.6000 291.4000 40.4000 294.8000 ;
	    RECT 46.6000 294.2000 47.4000 294.4000 ;
	    RECT 52.4000 294.2000 53.0000 296.4000 ;
	    RECT 57.2000 295.0000 58.0000 299.8000 ;
	    RECT 55.6000 294.2000 57.2000 294.4000 ;
	    RECT 46.2000 293.6000 57.2000 294.2000 ;
	    RECT 58.8000 294.3000 59.6000 294.4000 ;
	    RECT 60.4000 294.3000 61.2000 299.8000 ;
	    RECT 63.6000 295.8000 64.4000 299.8000 ;
	    RECT 65.2000 296.0000 66.0000 299.8000 ;
	    RECT 68.4000 296.0000 69.2000 299.8000 ;
	    RECT 71.6000 297.6000 72.4000 299.8000 ;
	    RECT 65.2000 295.8000 69.2000 296.0000 ;
	    RECT 58.8000 293.7000 61.2000 294.3000 ;
	    RECT 58.8000 293.6000 59.6000 293.7000 ;
	    RECT 44.4000 292.8000 45.2000 293.0000 ;
	    RECT 41.4000 292.2000 45.2000 292.8000 ;
	    RECT 46.2000 292.4000 46.8000 293.6000 ;
	    RECT 53.4000 293.4000 54.2000 293.6000 ;
	    RECT 52.4000 292.4000 53.2000 292.6000 ;
	    RECT 55.0000 292.4000 55.8000 292.6000 ;
	    RECT 41.4000 292.0000 42.2000 292.2000 ;
	    RECT 46.0000 291.6000 46.8000 292.4000 ;
	    RECT 50.8000 291.8000 55.8000 292.4000 ;
	    RECT 50.8000 291.6000 51.6000 291.8000 ;
	    RECT 43.0000 291.4000 43.8000 291.6000 ;
	    RECT 33.2000 291.0000 38.8000 291.2000 ;
	    RECT 33.0000 290.8000 38.8000 291.0000 ;
	    RECT 25.2000 289.8000 27.6000 290.4000 ;
	    RECT 29.0000 290.6000 38.8000 290.8000 ;
	    RECT 29.0000 290.2000 33.8000 290.6000 ;
	    RECT 25.2000 288.8000 25.8000 289.8000 ;
	    RECT 24.4000 288.0000 25.8000 288.8000 ;
	    RECT 27.4000 289.0000 28.2000 289.2000 ;
	    RECT 29.0000 289.0000 29.6000 290.2000 ;
	    RECT 27.4000 288.4000 29.6000 289.0000 ;
	    RECT 30.2000 289.0000 35.6000 289.6000 ;
	    RECT 30.2000 288.8000 31.0000 289.0000 ;
	    RECT 34.8000 288.8000 35.6000 289.0000 ;
	    RECT 28.6000 287.4000 29.4000 287.6000 ;
	    RECT 31.4000 287.4000 32.2000 287.6000 ;
	    RECT 25.2000 286.2000 26.0000 287.0000 ;
	    RECT 28.6000 286.8000 32.2000 287.4000 ;
	    RECT 29.4000 286.2000 30.0000 286.8000 ;
	    RECT 34.8000 286.2000 35.6000 287.0000 ;
	    RECT 24.6000 282.2000 25.8000 286.2000 ;
	    RECT 29.2000 282.2000 30.0000 286.2000 ;
	    RECT 33.6000 285.6000 35.6000 286.2000 ;
	    RECT 33.6000 282.2000 34.4000 285.6000 ;
	    RECT 38.0000 282.2000 38.8000 290.6000 ;
	    RECT 39.6000 290.8000 43.8000 291.4000 ;
	    RECT 39.6000 282.2000 40.4000 290.8000 ;
	    RECT 42.8000 289.6000 43.6000 290.8000 ;
	    RECT 46.2000 290.4000 46.8000 291.6000 ;
	    RECT 52.4000 291.0000 58.0000 291.2000 ;
	    RECT 52.2000 290.8000 58.0000 291.0000 ;
	    RECT 44.4000 289.8000 46.8000 290.4000 ;
	    RECT 48.2000 290.6000 58.0000 290.8000 ;
	    RECT 48.2000 290.2000 53.0000 290.6000 ;
	    RECT 44.4000 288.8000 45.0000 289.8000 ;
	    RECT 43.6000 288.0000 45.0000 288.8000 ;
	    RECT 46.6000 289.0000 47.4000 289.2000 ;
	    RECT 48.2000 289.0000 48.8000 290.2000 ;
	    RECT 46.6000 288.4000 48.8000 289.0000 ;
	    RECT 49.4000 289.0000 54.8000 289.6000 ;
	    RECT 49.4000 288.8000 50.2000 289.0000 ;
	    RECT 54.0000 288.8000 54.8000 289.0000 ;
	    RECT 47.8000 287.4000 48.6000 287.6000 ;
	    RECT 50.6000 287.4000 51.4000 287.6000 ;
	    RECT 44.4000 286.2000 45.2000 287.0000 ;
	    RECT 47.8000 286.8000 51.4000 287.4000 ;
	    RECT 48.6000 286.2000 49.2000 286.8000 ;
	    RECT 54.0000 286.2000 54.8000 287.0000 ;
	    RECT 43.8000 282.2000 45.0000 286.2000 ;
	    RECT 48.4000 282.2000 49.2000 286.2000 ;
	    RECT 52.8000 285.6000 54.8000 286.2000 ;
	    RECT 52.8000 282.2000 53.6000 285.6000 ;
	    RECT 57.2000 282.2000 58.0000 290.6000 ;
	    RECT 60.4000 282.2000 61.2000 293.7000 ;
	    RECT 62.0000 293.6000 62.8000 295.2000 ;
	    RECT 63.8000 294.4000 64.4000 295.8000 ;
	    RECT 65.4000 295.4000 69.0000 295.8000 ;
	    RECT 70.0000 295.6000 70.8000 297.2000 ;
	    RECT 67.6000 294.4000 68.4000 294.8000 ;
	    RECT 71.8000 294.4000 72.4000 297.6000 ;
	    RECT 77.4000 296.4000 78.2000 299.8000 ;
	    RECT 76.4000 295.8000 78.2000 296.4000 ;
	    RECT 79.6000 295.8000 80.4000 299.8000 ;
	    RECT 81.2000 296.0000 82.0000 299.8000 ;
	    RECT 84.4000 296.0000 85.2000 299.8000 ;
	    RECT 81.2000 295.8000 85.2000 296.0000 ;
	    RECT 86.0000 296.0000 86.8000 299.8000 ;
	    RECT 89.2000 296.0000 90.0000 299.8000 ;
	    RECT 86.0000 295.8000 90.0000 296.0000 ;
	    RECT 90.8000 295.8000 91.6000 299.8000 ;
	    RECT 92.4000 296.0000 93.2000 299.8000 ;
	    RECT 95.6000 299.2000 99.6000 299.8000 ;
	    RECT 95.6000 296.0000 96.4000 299.2000 ;
	    RECT 92.4000 295.8000 96.4000 296.0000 ;
	    RECT 97.2000 295.8000 98.0000 298.6000 ;
	    RECT 98.8000 295.8000 99.6000 299.2000 ;
	    RECT 100.4000 297.0000 101.2000 299.0000 ;
	    RECT 63.6000 293.6000 66.2000 294.4000 ;
	    RECT 67.6000 293.8000 69.2000 294.4000 ;
	    RECT 68.4000 293.6000 69.2000 293.8000 ;
	    RECT 71.6000 293.6000 72.4000 294.4000 ;
	    RECT 74.8000 293.6000 75.6000 295.2000 ;
	    RECT 63.6000 290.2000 64.4000 290.4000 ;
	    RECT 65.6000 290.2000 66.2000 293.6000 ;
	    RECT 66.8000 292.3000 67.6000 293.2000 ;
	    RECT 70.0000 292.3000 70.8000 292.4000 ;
	    RECT 66.8000 291.7000 70.8000 292.3000 ;
	    RECT 66.8000 291.6000 67.6000 291.7000 ;
	    RECT 70.0000 291.6000 70.8000 291.7000 ;
	    RECT 71.8000 290.2000 72.4000 293.6000 ;
	    RECT 73.2000 290.8000 74.0000 292.4000 ;
	    RECT 76.4000 292.3000 77.2000 295.8000 ;
	    RECT 79.8000 294.4000 80.4000 295.8000 ;
	    RECT 81.4000 295.4000 85.0000 295.8000 ;
	    RECT 86.2000 295.4000 89.8000 295.8000 ;
	    RECT 83.6000 294.4000 84.4000 294.8000 ;
	    RECT 86.8000 294.4000 87.6000 294.8000 ;
	    RECT 90.8000 294.4000 91.4000 295.8000 ;
	    RECT 92.6000 295.4000 96.2000 295.8000 ;
	    RECT 93.2000 294.4000 94.0000 294.8000 ;
	    RECT 97.4000 294.4000 98.0000 295.8000 ;
	    RECT 100.4000 294.8000 101.0000 297.0000 ;
	    RECT 104.6000 296.4000 105.4000 299.0000 ;
	    RECT 103.6000 296.0000 105.4000 296.4000 ;
	    RECT 120.2000 296.0000 121.0000 299.0000 ;
	    RECT 124.4000 297.0000 125.2000 299.0000 ;
	    RECT 103.6000 295.6000 106.2000 296.0000 ;
	    RECT 104.6000 295.4000 106.2000 295.6000 ;
	    RECT 105.4000 295.0000 106.2000 295.4000 ;
	    RECT 79.6000 293.6000 82.2000 294.4000 ;
	    RECT 83.6000 293.8000 85.2000 294.4000 ;
	    RECT 84.4000 293.6000 85.2000 293.8000 ;
	    RECT 86.0000 293.8000 87.6000 294.4000 ;
	    RECT 89.0000 294.3000 91.6000 294.4000 ;
	    RECT 92.4000 294.3000 94.0000 294.4000 ;
	    RECT 89.0000 293.8000 94.0000 294.3000 ;
	    RECT 95.6000 293.8000 98.0000 294.4000 ;
	    RECT 86.0000 293.6000 86.8000 293.8000 ;
	    RECT 89.0000 293.7000 93.2000 293.8000 ;
	    RECT 89.0000 293.6000 91.6000 293.7000 ;
	    RECT 92.4000 293.6000 93.2000 293.7000 ;
	    RECT 95.6000 293.6000 96.4000 293.8000 ;
	    RECT 81.6000 292.4000 82.2000 293.6000 ;
	    RECT 76.4000 291.7000 80.3000 292.3000 ;
	    RECT 63.6000 289.6000 65.0000 290.2000 ;
	    RECT 65.6000 289.6000 66.6000 290.2000 ;
	    RECT 64.4000 288.4000 65.0000 289.6000 ;
	    RECT 64.4000 287.6000 65.2000 288.4000 ;
	    RECT 65.8000 282.2000 66.6000 289.6000 ;
	    RECT 71.6000 289.4000 73.4000 290.2000 ;
	    RECT 72.6000 282.2000 73.4000 289.4000 ;
	    RECT 76.4000 282.2000 77.2000 291.7000 ;
	    RECT 79.7000 290.4000 80.3000 291.7000 ;
	    RECT 81.2000 291.6000 82.2000 292.4000 ;
	    RECT 82.8000 291.6000 83.6000 293.2000 ;
	    RECT 86.0000 292.3000 86.8000 292.4000 ;
	    RECT 87.6000 292.3000 88.4000 293.2000 ;
	    RECT 86.0000 291.7000 88.4000 292.3000 ;
	    RECT 86.0000 291.6000 86.8000 291.7000 ;
	    RECT 87.6000 291.6000 88.4000 291.7000 ;
	    RECT 78.0000 288.8000 78.8000 290.4000 ;
	    RECT 79.6000 290.2000 80.4000 290.4000 ;
	    RECT 81.6000 290.2000 82.2000 291.6000 ;
	    RECT 89.0000 290.2000 89.6000 293.6000 ;
	    RECT 94.0000 291.6000 94.8000 293.2000 ;
	    RECT 90.8000 290.2000 91.6000 290.4000 ;
	    RECT 95.6000 290.2000 96.2000 293.6000 ;
	    RECT 97.2000 291.6000 98.0000 293.2000 ;
	    RECT 98.8000 292.8000 99.6000 294.4000 ;
	    RECT 100.4000 294.2000 104.6000 294.8000 ;
	    RECT 103.6000 293.8000 104.6000 294.2000 ;
	    RECT 105.6000 294.4000 106.2000 295.0000 ;
	    RECT 119.4000 295.4000 121.0000 296.0000 ;
	    RECT 119.4000 295.0000 120.2000 295.4000 ;
	    RECT 119.4000 294.4000 120.0000 295.0000 ;
	    RECT 124.6000 294.8000 125.2000 297.0000 ;
	    RECT 100.4000 291.6000 101.2000 293.2000 ;
	    RECT 102.0000 291.6000 102.8000 293.2000 ;
	    RECT 103.6000 293.0000 105.0000 293.8000 ;
	    RECT 105.6000 293.6000 107.6000 294.4000 ;
	    RECT 118.0000 293.6000 120.0000 294.4000 ;
	    RECT 121.0000 294.2000 125.2000 294.8000 ;
	    RECT 127.6000 297.8000 128.4000 299.8000 ;
	    RECT 132.4000 297.8000 133.2000 299.8000 ;
	    RECT 145.2000 299.2000 149.2000 299.8000 ;
	    RECT 127.6000 294.4000 128.2000 297.8000 ;
	    RECT 129.2000 296.3000 130.0000 297.2000 ;
	    RECT 130.8000 296.3000 131.6000 297.2000 ;
	    RECT 129.2000 295.7000 131.6000 296.3000 ;
	    RECT 129.2000 295.6000 130.0000 295.7000 ;
	    RECT 130.8000 295.6000 131.6000 295.7000 ;
	    RECT 132.6000 294.4000 133.2000 297.8000 ;
	    RECT 126.0000 294.3000 126.8000 294.4000 ;
	    RECT 127.6000 294.3000 128.4000 294.4000 ;
	    RECT 121.0000 293.8000 122.0000 294.2000 ;
	    RECT 103.6000 291.0000 104.2000 293.0000 ;
	    RECT 100.4000 290.4000 104.2000 291.0000 ;
	    RECT 79.6000 289.6000 81.0000 290.2000 ;
	    RECT 81.6000 289.6000 82.6000 290.2000 ;
	    RECT 80.4000 288.4000 81.0000 289.6000 ;
	    RECT 80.4000 287.6000 81.2000 288.4000 ;
	    RECT 81.8000 282.2000 82.6000 289.6000 ;
	    RECT 88.6000 289.6000 89.6000 290.2000 ;
	    RECT 90.2000 289.6000 91.6000 290.2000 ;
	    RECT 88.6000 282.2000 89.4000 289.6000 ;
	    RECT 90.2000 288.4000 90.8000 289.6000 ;
	    RECT 90.0000 287.6000 90.8000 288.4000 ;
	    RECT 95.0000 282.2000 97.0000 290.2000 ;
	    RECT 100.4000 287.0000 101.0000 290.4000 ;
	    RECT 105.6000 289.8000 106.2000 293.6000 ;
	    RECT 106.8000 292.3000 107.6000 292.4000 ;
	    RECT 118.0000 292.3000 118.8000 292.4000 ;
	    RECT 106.8000 291.7000 118.8000 292.3000 ;
	    RECT 106.8000 290.8000 107.6000 291.7000 ;
	    RECT 118.0000 290.8000 118.8000 291.7000 ;
	    RECT 104.6000 289.2000 106.2000 289.8000 ;
	    RECT 119.4000 289.8000 120.0000 293.6000 ;
	    RECT 120.6000 293.0000 122.0000 293.8000 ;
	    RECT 126.0000 293.7000 128.4000 294.3000 ;
	    RECT 126.0000 293.6000 126.8000 293.7000 ;
	    RECT 127.6000 293.6000 128.4000 293.7000 ;
	    RECT 132.4000 293.6000 133.2000 294.4000 ;
	    RECT 135.6000 297.0000 136.4000 299.0000 ;
	    RECT 139.8000 298.4000 140.6000 299.0000 ;
	    RECT 139.8000 297.6000 141.2000 298.4000 ;
	    RECT 135.6000 294.8000 136.2000 297.0000 ;
	    RECT 139.8000 296.0000 140.6000 297.6000 ;
	    RECT 139.8000 295.4000 141.4000 296.0000 ;
	    RECT 145.2000 295.8000 146.0000 299.2000 ;
	    RECT 146.8000 295.8000 147.6000 298.6000 ;
	    RECT 148.4000 296.0000 149.2000 299.2000 ;
	    RECT 151.6000 296.0000 152.4000 299.8000 ;
	    RECT 148.4000 295.8000 152.4000 296.0000 ;
	    RECT 153.2000 296.0000 154.0000 299.8000 ;
	    RECT 156.4000 296.0000 157.2000 299.8000 ;
	    RECT 153.2000 295.8000 157.2000 296.0000 ;
	    RECT 158.0000 295.8000 158.8000 299.8000 ;
	    RECT 161.2000 297.8000 162.0000 299.8000 ;
	    RECT 140.6000 295.0000 141.4000 295.4000 ;
	    RECT 135.6000 294.2000 139.8000 294.8000 ;
	    RECT 121.4000 291.0000 122.0000 293.0000 ;
	    RECT 122.8000 291.6000 123.6000 293.2000 ;
	    RECT 124.4000 291.6000 125.2000 293.2000 ;
	    RECT 121.4000 290.4000 125.2000 291.0000 ;
	    RECT 126.0000 290.8000 126.8000 292.4000 ;
	    RECT 119.4000 289.2000 121.0000 289.8000 ;
	    RECT 100.4000 283.0000 101.2000 287.0000 ;
	    RECT 104.6000 282.2000 105.4000 289.2000 ;
	    RECT 120.2000 284.4000 121.0000 289.2000 ;
	    RECT 124.6000 287.0000 125.2000 290.4000 ;
	    RECT 127.6000 290.2000 128.2000 293.6000 ;
	    RECT 132.6000 290.2000 133.2000 293.6000 ;
	    RECT 138.8000 293.8000 139.8000 294.2000 ;
	    RECT 140.8000 294.4000 141.4000 295.0000 ;
	    RECT 146.8000 294.4000 147.4000 295.8000 ;
	    RECT 148.6000 295.4000 152.2000 295.8000 ;
	    RECT 153.4000 295.4000 157.0000 295.8000 ;
	    RECT 150.8000 294.4000 151.6000 294.8000 ;
	    RECT 154.0000 294.4000 154.8000 294.8000 ;
	    RECT 158.0000 294.4000 158.6000 295.8000 ;
	    RECT 159.6000 295.6000 160.4000 297.2000 ;
	    RECT 161.4000 294.4000 162.0000 297.8000 ;
	    RECT 164.4000 296.0000 165.2000 299.8000 ;
	    RECT 167.6000 296.0000 168.4000 299.8000 ;
	    RECT 164.4000 295.8000 168.4000 296.0000 ;
	    RECT 169.2000 295.8000 170.0000 299.8000 ;
	    RECT 170.8000 295.8000 171.6000 299.8000 ;
	    RECT 172.4000 296.0000 173.2000 299.8000 ;
	    RECT 175.6000 296.0000 176.4000 299.8000 ;
	    RECT 172.4000 295.8000 176.4000 296.0000 ;
	    RECT 164.6000 295.4000 168.2000 295.8000 ;
	    RECT 165.2000 294.4000 166.0000 294.8000 ;
	    RECT 169.2000 294.4000 169.8000 295.8000 ;
	    RECT 171.0000 294.4000 171.6000 295.8000 ;
	    RECT 172.6000 295.4000 176.2000 295.8000 ;
	    RECT 174.8000 294.4000 175.6000 294.8000 ;
	    RECT 134.0000 290.8000 134.8000 292.4000 ;
	    RECT 135.6000 291.6000 136.4000 293.2000 ;
	    RECT 137.2000 291.6000 138.0000 293.2000 ;
	    RECT 138.8000 293.0000 140.2000 293.8000 ;
	    RECT 140.8000 293.6000 142.8000 294.4000 ;
	    RECT 138.8000 291.0000 139.4000 293.0000 ;
	    RECT 135.6000 290.4000 139.4000 291.0000 ;
	    RECT 119.6000 283.6000 121.0000 284.4000 ;
	    RECT 120.2000 282.2000 121.0000 283.6000 ;
	    RECT 124.4000 283.0000 125.2000 287.0000 ;
	    RECT 126.6000 289.4000 128.4000 290.2000 ;
	    RECT 132.4000 289.4000 134.2000 290.2000 ;
	    RECT 126.6000 282.2000 127.4000 289.4000 ;
	    RECT 133.4000 284.4000 134.2000 289.4000 ;
	    RECT 135.6000 287.0000 136.2000 290.4000 ;
	    RECT 140.8000 289.8000 141.4000 293.6000 ;
	    RECT 145.2000 292.8000 146.0000 294.4000 ;
	    RECT 146.8000 293.8000 149.2000 294.4000 ;
	    RECT 150.8000 293.8000 152.4000 294.4000 ;
	    RECT 148.4000 293.6000 149.2000 293.8000 ;
	    RECT 151.6000 293.6000 152.4000 293.8000 ;
	    RECT 153.2000 293.8000 154.8000 294.4000 ;
	    RECT 153.2000 293.6000 154.0000 293.8000 ;
	    RECT 156.2000 293.6000 158.8000 294.4000 ;
	    RECT 161.2000 293.6000 162.0000 294.4000 ;
	    RECT 164.4000 293.8000 166.0000 294.4000 ;
	    RECT 164.4000 293.6000 165.2000 293.8000 ;
	    RECT 167.4000 293.6000 170.0000 294.4000 ;
	    RECT 170.8000 293.6000 173.4000 294.4000 ;
	    RECT 174.8000 293.8000 176.4000 294.4000 ;
	    RECT 175.6000 293.6000 176.4000 293.8000 ;
	    RECT 142.0000 290.8000 142.8000 292.4000 ;
	    RECT 146.8000 291.6000 147.6000 293.2000 ;
	    RECT 148.6000 290.2000 149.2000 293.6000 ;
	    RECT 150.0000 291.6000 150.8000 293.2000 ;
	    RECT 154.8000 291.6000 155.6000 293.2000 ;
	    RECT 156.2000 290.2000 156.8000 293.6000 ;
	    RECT 161.4000 290.4000 162.0000 293.6000 ;
	    RECT 162.8000 290.8000 163.6000 292.4000 ;
	    RECT 164.4000 292.3000 165.2000 292.4000 ;
	    RECT 166.0000 292.3000 166.8000 293.2000 ;
	    RECT 164.4000 291.7000 166.8000 292.3000 ;
	    RECT 164.4000 291.6000 165.2000 291.7000 ;
	    RECT 166.0000 291.6000 166.8000 291.7000 ;
	    RECT 158.0000 290.2000 158.8000 290.4000 ;
	    RECT 139.8000 289.2000 141.4000 289.8000 ;
	    RECT 133.4000 283.6000 134.8000 284.4000 ;
	    RECT 133.4000 282.2000 134.2000 283.6000 ;
	    RECT 135.6000 283.0000 136.4000 287.0000 ;
	    RECT 139.8000 282.2000 140.6000 289.2000 ;
	    RECT 147.8000 284.4000 149.8000 290.2000 ;
	    RECT 146.8000 283.6000 149.8000 284.4000 ;
	    RECT 147.8000 282.2000 149.8000 283.6000 ;
	    RECT 155.8000 289.6000 156.8000 290.2000 ;
	    RECT 157.4000 289.6000 158.8000 290.2000 ;
	    RECT 161.2000 290.2000 162.0000 290.4000 ;
	    RECT 167.4000 290.2000 168.0000 293.6000 ;
	    RECT 172.8000 292.3000 173.4000 293.6000 ;
	    RECT 169.3000 291.7000 173.4000 292.3000 ;
	    RECT 169.3000 290.4000 169.9000 291.7000 ;
	    RECT 169.2000 290.2000 170.0000 290.4000 ;
	    RECT 155.8000 282.2000 156.6000 289.6000 ;
	    RECT 157.4000 288.4000 158.0000 289.6000 ;
	    RECT 161.2000 289.4000 163.0000 290.2000 ;
	    RECT 157.2000 287.6000 158.0000 288.4000 ;
	    RECT 162.2000 282.2000 163.0000 289.4000 ;
	    RECT 167.0000 289.6000 168.0000 290.2000 ;
	    RECT 168.6000 289.6000 170.0000 290.2000 ;
	    RECT 170.8000 290.2000 171.6000 290.4000 ;
	    RECT 172.8000 290.2000 173.4000 291.7000 ;
	    RECT 174.0000 291.6000 174.8000 293.2000 ;
	    RECT 177.2000 292.4000 178.0000 299.8000 ;
	    RECT 180.4000 295.2000 181.2000 299.8000 ;
	    RECT 179.0000 294.6000 181.2000 295.2000 ;
	    RECT 182.0000 295.4000 182.8000 299.8000 ;
	    RECT 186.2000 298.4000 187.4000 299.8000 ;
	    RECT 186.2000 297.8000 187.6000 298.4000 ;
	    RECT 190.8000 297.8000 191.6000 299.8000 ;
	    RECT 195.2000 298.4000 196.0000 299.8000 ;
	    RECT 195.2000 297.8000 197.2000 298.4000 ;
	    RECT 186.8000 297.0000 187.6000 297.8000 ;
	    RECT 191.0000 297.2000 191.6000 297.8000 ;
	    RECT 191.0000 296.6000 193.8000 297.2000 ;
	    RECT 193.0000 296.4000 193.8000 296.6000 ;
	    RECT 194.8000 296.4000 195.6000 297.2000 ;
	    RECT 196.4000 297.0000 197.2000 297.8000 ;
	    RECT 185.0000 295.4000 185.8000 295.6000 ;
	    RECT 182.0000 294.8000 185.8000 295.4000 ;
	    RECT 177.2000 290.2000 177.8000 292.4000 ;
	    RECT 179.0000 291.6000 179.6000 294.6000 ;
	    RECT 178.4000 290.8000 179.6000 291.6000 ;
	    RECT 179.0000 290.2000 179.6000 290.8000 ;
	    RECT 182.0000 291.4000 182.8000 294.8000 ;
	    RECT 189.0000 294.2000 189.8000 294.4000 ;
	    RECT 194.8000 294.2000 195.4000 296.4000 ;
	    RECT 199.6000 295.0000 200.4000 299.8000 ;
	    RECT 201.2000 296.0000 202.0000 299.8000 ;
	    RECT 204.4000 296.0000 205.2000 299.8000 ;
	    RECT 201.2000 295.8000 205.2000 296.0000 ;
	    RECT 206.0000 295.8000 206.8000 299.8000 ;
	    RECT 208.2000 296.4000 209.0000 299.8000 ;
	    RECT 208.2000 295.8000 210.0000 296.4000 ;
	    RECT 212.4000 296.0000 213.2000 299.8000 ;
	    RECT 215.6000 296.0000 216.4000 299.8000 ;
	    RECT 212.4000 295.8000 216.4000 296.0000 ;
	    RECT 217.2000 295.8000 218.0000 299.8000 ;
	    RECT 218.8000 295.8000 219.6000 299.8000 ;
	    RECT 220.4000 296.0000 221.2000 299.8000 ;
	    RECT 223.6000 296.0000 224.4000 299.8000 ;
	    RECT 220.4000 295.8000 224.4000 296.0000 ;
	    RECT 201.4000 295.4000 205.0000 295.8000 ;
	    RECT 202.0000 294.4000 202.8000 294.8000 ;
	    RECT 206.0000 294.4000 206.6000 295.8000 ;
	    RECT 198.0000 294.2000 199.6000 294.4000 ;
	    RECT 188.6000 293.6000 199.6000 294.2000 ;
	    RECT 201.2000 293.8000 202.8000 294.4000 ;
	    RECT 201.2000 293.6000 202.0000 293.8000 ;
	    RECT 204.2000 293.6000 206.8000 294.4000 ;
	    RECT 186.8000 292.8000 187.6000 293.0000 ;
	    RECT 183.8000 292.2000 187.6000 292.8000 ;
	    RECT 183.8000 292.0000 184.6000 292.2000 ;
	    RECT 185.4000 291.4000 186.2000 291.6000 ;
	    RECT 182.0000 290.8000 186.2000 291.4000 ;
	    RECT 170.8000 289.6000 172.2000 290.2000 ;
	    RECT 172.8000 289.6000 173.8000 290.2000 ;
	    RECT 167.0000 282.2000 167.8000 289.6000 ;
	    RECT 168.6000 288.4000 169.2000 289.6000 ;
	    RECT 168.4000 287.6000 169.2000 288.4000 ;
	    RECT 171.6000 288.4000 172.2000 289.6000 ;
	    RECT 171.6000 287.6000 172.4000 288.4000 ;
	    RECT 173.0000 282.2000 173.8000 289.6000 ;
	    RECT 177.2000 282.2000 178.0000 290.2000 ;
	    RECT 179.0000 289.6000 181.2000 290.2000 ;
	    RECT 180.4000 282.2000 181.2000 289.6000 ;
	    RECT 182.0000 282.2000 182.8000 290.8000 ;
	    RECT 188.6000 290.4000 189.2000 293.6000 ;
	    RECT 195.8000 293.4000 196.6000 293.6000 ;
	    RECT 194.8000 292.4000 195.6000 292.6000 ;
	    RECT 197.4000 292.4000 198.2000 292.6000 ;
	    RECT 193.2000 291.8000 198.2000 292.4000 ;
	    RECT 193.2000 291.6000 194.0000 291.8000 ;
	    RECT 202.8000 291.6000 203.6000 293.2000 ;
	    RECT 194.8000 291.0000 200.4000 291.2000 ;
	    RECT 194.6000 290.8000 200.4000 291.0000 ;
	    RECT 186.8000 289.8000 189.2000 290.4000 ;
	    RECT 190.6000 290.6000 200.4000 290.8000 ;
	    RECT 190.6000 290.2000 195.4000 290.6000 ;
	    RECT 186.8000 288.8000 187.4000 289.8000 ;
	    RECT 186.0000 288.0000 187.4000 288.8000 ;
	    RECT 189.0000 289.0000 189.8000 289.2000 ;
	    RECT 190.6000 289.0000 191.2000 290.2000 ;
	    RECT 189.0000 288.4000 191.2000 289.0000 ;
	    RECT 191.8000 289.0000 197.2000 289.6000 ;
	    RECT 191.8000 288.8000 192.6000 289.0000 ;
	    RECT 196.4000 288.8000 197.2000 289.0000 ;
	    RECT 190.2000 287.4000 191.0000 287.6000 ;
	    RECT 193.0000 287.4000 193.8000 287.6000 ;
	    RECT 186.8000 286.2000 187.6000 287.0000 ;
	    RECT 190.2000 286.8000 193.8000 287.4000 ;
	    RECT 191.0000 286.2000 191.6000 286.8000 ;
	    RECT 196.4000 286.2000 197.2000 287.0000 ;
	    RECT 186.2000 282.2000 187.4000 286.2000 ;
	    RECT 190.8000 282.2000 191.6000 286.2000 ;
	    RECT 195.2000 285.6000 197.2000 286.2000 ;
	    RECT 195.2000 282.2000 196.0000 285.6000 ;
	    RECT 199.6000 282.2000 200.4000 290.6000 ;
	    RECT 204.2000 290.2000 204.8000 293.6000 ;
	    RECT 209.2000 292.3000 210.0000 295.8000 ;
	    RECT 212.6000 295.4000 216.2000 295.8000 ;
	    RECT 210.8000 293.6000 211.6000 295.2000 ;
	    RECT 213.2000 294.4000 214.0000 294.8000 ;
	    RECT 217.2000 294.4000 217.8000 295.8000 ;
	    RECT 219.0000 294.4000 219.6000 295.8000 ;
	    RECT 220.6000 295.4000 224.2000 295.8000 ;
	    RECT 225.2000 295.4000 226.0000 299.8000 ;
	    RECT 229.4000 298.4000 230.6000 299.8000 ;
	    RECT 229.4000 297.8000 230.8000 298.4000 ;
	    RECT 234.0000 297.8000 234.8000 299.8000 ;
	    RECT 238.4000 298.4000 239.2000 299.8000 ;
	    RECT 238.4000 297.8000 240.4000 298.4000 ;
	    RECT 230.0000 297.0000 230.8000 297.8000 ;
	    RECT 234.2000 297.2000 234.8000 297.8000 ;
	    RECT 234.2000 296.6000 237.0000 297.2000 ;
	    RECT 236.2000 296.4000 237.0000 296.6000 ;
	    RECT 238.0000 296.4000 238.8000 297.2000 ;
	    RECT 239.6000 297.0000 240.4000 297.8000 ;
	    RECT 228.2000 295.4000 229.0000 295.6000 ;
	    RECT 225.2000 294.8000 229.0000 295.4000 ;
	    RECT 222.8000 294.4000 223.6000 294.8000 ;
	    RECT 212.4000 293.8000 214.0000 294.4000 ;
	    RECT 212.4000 293.6000 213.2000 293.8000 ;
	    RECT 215.4000 293.6000 218.0000 294.4000 ;
	    RECT 218.8000 293.6000 221.4000 294.4000 ;
	    RECT 222.8000 293.8000 224.4000 294.4000 ;
	    RECT 223.6000 293.6000 224.4000 293.8000 ;
	    RECT 206.1000 291.7000 210.0000 292.3000 ;
	    RECT 206.1000 290.4000 206.7000 291.7000 ;
	    RECT 206.0000 290.2000 206.8000 290.4000 ;
	    RECT 203.8000 289.6000 204.8000 290.2000 ;
	    RECT 205.4000 289.6000 206.8000 290.2000 ;
	    RECT 203.8000 282.2000 204.6000 289.6000 ;
	    RECT 205.4000 288.4000 206.0000 289.6000 ;
	    RECT 207.6000 288.8000 208.4000 290.4000 ;
	    RECT 205.2000 287.6000 206.0000 288.4000 ;
	    RECT 209.2000 282.2000 210.0000 291.7000 ;
	    RECT 214.0000 291.6000 214.8000 293.2000 ;
	    RECT 215.4000 292.3000 216.0000 293.6000 ;
	    RECT 220.8000 292.4000 221.4000 293.6000 ;
	    RECT 215.4000 291.7000 219.5000 292.3000 ;
	    RECT 215.4000 290.2000 216.0000 291.7000 ;
	    RECT 218.9000 290.4000 219.5000 291.7000 ;
	    RECT 220.4000 291.6000 221.4000 292.4000 ;
	    RECT 222.0000 291.6000 222.8000 293.2000 ;
	    RECT 217.2000 290.2000 218.0000 290.4000 ;
	    RECT 215.0000 289.6000 216.0000 290.2000 ;
	    RECT 216.6000 289.6000 218.0000 290.2000 ;
	    RECT 218.8000 290.2000 219.6000 290.4000 ;
	    RECT 220.8000 290.2000 221.4000 291.6000 ;
	    RECT 225.2000 291.4000 226.0000 294.8000 ;
	    RECT 232.2000 294.2000 233.0000 294.4000 ;
	    RECT 234.8000 294.2000 235.6000 294.4000 ;
	    RECT 238.0000 294.2000 238.6000 296.4000 ;
	    RECT 242.8000 295.0000 243.6000 299.8000 ;
	    RECT 244.4000 297.0000 245.2000 299.0000 ;
	    RECT 244.4000 294.8000 245.0000 297.0000 ;
	    RECT 248.6000 296.0000 249.4000 299.0000 ;
	    RECT 248.6000 295.4000 250.2000 296.0000 ;
	    RECT 260.4000 295.8000 261.2000 299.8000 ;
	    RECT 262.0000 296.0000 262.8000 299.8000 ;
	    RECT 265.2000 296.0000 266.0000 299.8000 ;
	    RECT 268.4000 297.8000 269.2000 299.8000 ;
	    RECT 262.0000 295.8000 266.0000 296.0000 ;
	    RECT 249.4000 295.0000 250.2000 295.4000 ;
	    RECT 241.2000 294.2000 242.8000 294.4000 ;
	    RECT 244.4000 294.2000 248.6000 294.8000 ;
	    RECT 231.8000 293.6000 242.8000 294.2000 ;
	    RECT 247.6000 293.8000 248.6000 294.2000 ;
	    RECT 249.6000 294.4000 250.2000 295.0000 ;
	    RECT 260.6000 294.4000 261.2000 295.8000 ;
	    RECT 262.2000 295.4000 265.8000 295.8000 ;
	    RECT 266.8000 295.6000 267.6000 297.2000 ;
	    RECT 264.4000 294.4000 265.2000 294.8000 ;
	    RECT 268.6000 294.4000 269.2000 297.8000 ;
	    RECT 271.6000 296.0000 272.4000 299.8000 ;
	    RECT 274.8000 299.2000 278.8000 299.8000 ;
	    RECT 274.8000 296.0000 275.6000 299.2000 ;
	    RECT 271.6000 295.8000 275.6000 296.0000 ;
	    RECT 276.4000 295.8000 277.2000 298.6000 ;
	    RECT 278.0000 295.8000 278.8000 299.2000 ;
	    RECT 279.6000 296.0000 280.4000 299.8000 ;
	    RECT 282.8000 296.0000 283.6000 299.8000 ;
	    RECT 279.6000 295.8000 283.6000 296.0000 ;
	    RECT 284.4000 295.8000 285.2000 299.8000 ;
	    RECT 286.0000 299.2000 290.0000 299.8000 ;
	    RECT 286.0000 295.8000 286.8000 299.2000 ;
	    RECT 287.6000 295.8000 288.4000 298.6000 ;
	    RECT 289.2000 296.0000 290.0000 299.2000 ;
	    RECT 292.4000 296.0000 293.2000 299.8000 ;
	    RECT 295.6000 297.8000 296.4000 299.8000 ;
	    RECT 289.2000 295.8000 293.2000 296.0000 ;
	    RECT 271.8000 295.4000 275.4000 295.8000 ;
	    RECT 272.4000 294.4000 273.2000 294.8000 ;
	    RECT 276.6000 294.4000 277.2000 295.8000 ;
	    RECT 279.8000 295.4000 283.4000 295.8000 ;
	    RECT 280.4000 294.4000 281.2000 294.8000 ;
	    RECT 284.4000 294.4000 285.0000 295.8000 ;
	    RECT 287.6000 294.4000 288.2000 295.8000 ;
	    RECT 289.4000 295.4000 293.0000 295.8000 ;
	    RECT 294.0000 295.6000 294.8000 297.2000 ;
	    RECT 291.6000 294.4000 292.4000 294.8000 ;
	    RECT 295.8000 294.4000 296.4000 297.8000 ;
	    RECT 298.8000 295.8000 299.6000 299.8000 ;
	    RECT 300.4000 296.0000 301.2000 299.8000 ;
	    RECT 303.6000 296.0000 304.4000 299.8000 ;
	    RECT 300.4000 295.8000 304.4000 296.0000 ;
	    RECT 306.8000 297.6000 307.6000 299.8000 ;
	    RECT 310.0000 299.2000 314.0000 299.8000 ;
	    RECT 299.0000 294.4000 299.6000 295.8000 ;
	    RECT 300.6000 295.4000 304.2000 295.8000 ;
	    RECT 302.8000 294.4000 303.6000 294.8000 ;
	    RECT 306.8000 294.4000 307.4000 297.6000 ;
	    RECT 308.4000 295.6000 309.2000 297.2000 ;
	    RECT 310.0000 295.8000 310.8000 299.2000 ;
	    RECT 311.6000 295.8000 312.4000 298.6000 ;
	    RECT 313.2000 296.0000 314.0000 299.2000 ;
	    RECT 316.4000 296.0000 317.2000 299.8000 ;
	    RECT 313.2000 295.8000 317.2000 296.0000 ;
	    RECT 318.0000 295.8000 318.8000 299.8000 ;
	    RECT 319.6000 296.0000 320.4000 299.8000 ;
	    RECT 322.8000 296.0000 323.6000 299.8000 ;
	    RECT 319.6000 295.8000 323.6000 296.0000 ;
	    RECT 324.4000 295.8000 325.2000 299.8000 ;
	    RECT 326.0000 296.0000 326.8000 299.8000 ;
	    RECT 329.2000 296.0000 330.0000 299.8000 ;
	    RECT 326.0000 295.8000 330.0000 296.0000 ;
	    RECT 330.8000 297.0000 331.6000 299.0000 ;
	    RECT 311.6000 294.4000 312.2000 295.8000 ;
	    RECT 313.4000 295.4000 317.0000 295.8000 ;
	    RECT 315.6000 294.4000 316.4000 294.8000 ;
	    RECT 318.2000 294.4000 318.8000 295.8000 ;
	    RECT 319.8000 295.4000 323.4000 295.8000 ;
	    RECT 322.0000 294.4000 322.8000 294.8000 ;
	    RECT 324.6000 294.4000 325.2000 295.8000 ;
	    RECT 326.2000 295.4000 329.8000 295.8000 ;
	    RECT 330.8000 294.8000 331.4000 297.0000 ;
	    RECT 335.0000 296.0000 335.8000 299.0000 ;
	    RECT 340.4000 297.0000 341.2000 299.0000 ;
	    RECT 335.0000 295.4000 336.6000 296.0000 ;
	    RECT 335.8000 295.0000 336.6000 295.4000 ;
	    RECT 328.4000 294.4000 329.2000 294.8000 ;
	    RECT 230.0000 292.8000 230.8000 293.0000 ;
	    RECT 227.0000 292.2000 230.8000 292.8000 ;
	    RECT 227.0000 292.0000 227.8000 292.2000 ;
	    RECT 228.6000 291.4000 229.4000 291.6000 ;
	    RECT 225.2000 290.8000 229.4000 291.4000 ;
	    RECT 218.8000 289.6000 220.2000 290.2000 ;
	    RECT 220.8000 289.6000 221.8000 290.2000 ;
	    RECT 215.0000 282.2000 215.8000 289.6000 ;
	    RECT 216.6000 288.4000 217.2000 289.6000 ;
	    RECT 216.4000 287.6000 217.2000 288.4000 ;
	    RECT 219.6000 288.4000 220.2000 289.6000 ;
	    RECT 219.6000 287.6000 220.4000 288.4000 ;
	    RECT 221.0000 282.2000 221.8000 289.6000 ;
	    RECT 225.2000 282.2000 226.0000 290.8000 ;
	    RECT 231.8000 290.4000 232.4000 293.6000 ;
	    RECT 239.0000 293.4000 239.8000 293.6000 ;
	    RECT 240.6000 292.4000 241.4000 292.6000 ;
	    RECT 233.2000 292.3000 234.0000 292.4000 ;
	    RECT 236.4000 292.3000 241.4000 292.4000 ;
	    RECT 233.2000 291.8000 241.4000 292.3000 ;
	    RECT 233.2000 291.7000 237.2000 291.8000 ;
	    RECT 233.2000 291.6000 234.0000 291.7000 ;
	    RECT 236.4000 291.6000 237.2000 291.7000 ;
	    RECT 244.4000 291.6000 245.2000 293.2000 ;
	    RECT 246.0000 291.6000 246.8000 293.2000 ;
	    RECT 247.6000 293.0000 249.0000 293.8000 ;
	    RECT 249.6000 293.6000 251.6000 294.4000 ;
	    RECT 252.4000 294.3000 253.2000 294.4000 ;
	    RECT 260.4000 294.3000 263.0000 294.4000 ;
	    RECT 252.4000 293.7000 263.0000 294.3000 ;
	    RECT 264.4000 294.3000 266.0000 294.4000 ;
	    RECT 266.8000 294.3000 267.6000 294.4000 ;
	    RECT 264.4000 293.8000 267.6000 294.3000 ;
	    RECT 252.4000 293.6000 253.2000 293.7000 ;
	    RECT 260.4000 293.6000 263.0000 293.7000 ;
	    RECT 265.2000 293.7000 267.6000 293.8000 ;
	    RECT 265.2000 293.6000 266.0000 293.7000 ;
	    RECT 266.8000 293.6000 267.6000 293.7000 ;
	    RECT 268.4000 293.6000 269.2000 294.4000 ;
	    RECT 271.6000 293.8000 273.2000 294.4000 ;
	    RECT 274.8000 293.8000 277.2000 294.4000 ;
	    RECT 271.6000 293.6000 272.4000 293.8000 ;
	    RECT 274.8000 293.6000 275.6000 293.8000 ;
	    RECT 238.0000 291.0000 243.6000 291.2000 ;
	    RECT 247.6000 291.0000 248.2000 293.0000 ;
	    RECT 237.8000 290.8000 243.6000 291.0000 ;
	    RECT 230.0000 289.8000 232.4000 290.4000 ;
	    RECT 233.8000 290.6000 243.6000 290.8000 ;
	    RECT 233.8000 290.2000 238.6000 290.6000 ;
	    RECT 230.0000 288.8000 230.6000 289.8000 ;
	    RECT 229.2000 288.0000 230.6000 288.8000 ;
	    RECT 232.2000 289.0000 233.0000 289.2000 ;
	    RECT 233.8000 289.0000 234.4000 290.2000 ;
	    RECT 232.2000 288.4000 234.4000 289.0000 ;
	    RECT 235.0000 289.0000 240.4000 289.6000 ;
	    RECT 235.0000 288.8000 235.8000 289.0000 ;
	    RECT 239.6000 288.8000 240.4000 289.0000 ;
	    RECT 233.4000 287.4000 234.2000 287.6000 ;
	    RECT 236.2000 287.4000 237.0000 287.6000 ;
	    RECT 230.0000 286.2000 230.8000 287.0000 ;
	    RECT 233.4000 286.8000 237.0000 287.4000 ;
	    RECT 234.2000 286.2000 234.8000 286.8000 ;
	    RECT 239.6000 286.2000 240.4000 287.0000 ;
	    RECT 229.4000 282.2000 230.6000 286.2000 ;
	    RECT 234.0000 282.2000 234.8000 286.2000 ;
	    RECT 238.4000 285.6000 240.4000 286.2000 ;
	    RECT 238.4000 282.2000 239.2000 285.6000 ;
	    RECT 242.8000 282.2000 243.6000 290.6000 ;
	    RECT 244.4000 290.4000 248.2000 291.0000 ;
	    RECT 244.4000 287.0000 245.0000 290.4000 ;
	    RECT 249.6000 289.8000 250.2000 293.6000 ;
	    RECT 250.8000 290.8000 251.6000 292.4000 ;
	    RECT 248.6000 289.2000 250.2000 289.8000 ;
	    RECT 260.4000 290.2000 261.2000 290.4000 ;
	    RECT 262.4000 290.2000 263.0000 293.6000 ;
	    RECT 263.6000 291.6000 264.4000 293.2000 ;
	    RECT 268.6000 290.2000 269.2000 293.6000 ;
	    RECT 270.0000 290.8000 270.8000 292.4000 ;
	    RECT 271.6000 292.3000 272.4000 292.4000 ;
	    RECT 273.2000 292.3000 274.0000 293.2000 ;
	    RECT 271.6000 291.7000 274.0000 292.3000 ;
	    RECT 271.6000 291.6000 272.4000 291.7000 ;
	    RECT 273.2000 291.6000 274.0000 291.7000 ;
	    RECT 274.8000 290.2000 275.4000 293.6000 ;
	    RECT 276.4000 291.6000 277.2000 293.2000 ;
	    RECT 278.0000 292.8000 278.8000 294.4000 ;
	    RECT 279.6000 293.8000 281.2000 294.4000 ;
	    RECT 279.6000 293.6000 280.4000 293.8000 ;
	    RECT 282.6000 293.6000 285.2000 294.4000 ;
	    RECT 281.2000 291.6000 282.0000 293.2000 ;
	    RECT 282.6000 290.2000 283.2000 293.6000 ;
	    RECT 286.0000 292.8000 286.8000 294.4000 ;
	    RECT 287.6000 293.8000 290.0000 294.4000 ;
	    RECT 291.6000 294.3000 293.2000 294.4000 ;
	    RECT 294.0000 294.3000 294.8000 294.4000 ;
	    RECT 291.6000 293.8000 294.8000 294.3000 ;
	    RECT 289.2000 293.6000 290.0000 293.8000 ;
	    RECT 292.4000 293.7000 294.8000 293.8000 ;
	    RECT 292.4000 293.6000 293.2000 293.7000 ;
	    RECT 294.0000 293.6000 294.8000 293.7000 ;
	    RECT 295.6000 293.6000 296.4000 294.4000 ;
	    RECT 298.8000 293.6000 301.4000 294.4000 ;
	    RECT 302.8000 293.8000 304.4000 294.4000 ;
	    RECT 303.6000 293.6000 304.4000 293.8000 ;
	    RECT 306.8000 293.6000 307.6000 294.4000 ;
	    RECT 308.4000 294.3000 309.2000 294.4000 ;
	    RECT 310.0000 294.3000 310.8000 294.4000 ;
	    RECT 308.4000 293.7000 310.8000 294.3000 ;
	    RECT 311.6000 293.8000 314.0000 294.4000 ;
	    RECT 315.6000 294.3000 317.2000 294.4000 ;
	    RECT 318.0000 294.3000 320.6000 294.4000 ;
	    RECT 315.6000 293.8000 320.6000 294.3000 ;
	    RECT 322.0000 293.8000 323.6000 294.4000 ;
	    RECT 308.4000 293.6000 309.2000 293.7000 ;
	    RECT 287.6000 291.6000 288.4000 293.2000 ;
	    RECT 284.4000 290.2000 285.2000 290.4000 ;
	    RECT 289.4000 290.2000 290.0000 293.6000 ;
	    RECT 290.8000 292.3000 291.6000 293.2000 ;
	    RECT 295.8000 292.3000 296.4000 293.6000 ;
	    RECT 300.8000 292.4000 301.4000 293.6000 ;
	    RECT 290.8000 291.7000 296.4000 292.3000 ;
	    RECT 290.8000 291.6000 291.6000 291.7000 ;
	    RECT 295.8000 290.2000 296.4000 291.7000 ;
	    RECT 297.2000 290.8000 298.0000 292.4000 ;
	    RECT 300.4000 291.6000 301.4000 292.4000 ;
	    RECT 302.0000 291.6000 302.8000 293.2000 ;
	    RECT 298.8000 290.2000 299.6000 290.4000 ;
	    RECT 300.8000 290.2000 301.4000 291.6000 ;
	    RECT 305.2000 290.8000 306.0000 292.4000 ;
	    RECT 306.8000 290.2000 307.4000 293.6000 ;
	    RECT 310.0000 292.8000 310.8000 293.7000 ;
	    RECT 313.2000 293.6000 314.0000 293.8000 ;
	    RECT 316.4000 293.7000 320.6000 293.8000 ;
	    RECT 316.4000 293.6000 317.2000 293.7000 ;
	    RECT 318.0000 293.6000 320.6000 293.7000 ;
	    RECT 322.8000 293.6000 323.6000 293.8000 ;
	    RECT 324.4000 293.6000 327.0000 294.4000 ;
	    RECT 328.4000 293.8000 330.0000 294.4000 ;
	    RECT 330.8000 294.2000 335.0000 294.8000 ;
	    RECT 329.2000 293.6000 330.0000 293.8000 ;
	    RECT 334.0000 293.8000 335.0000 294.2000 ;
	    RECT 336.0000 294.4000 336.6000 295.0000 ;
	    RECT 340.4000 294.8000 341.0000 297.0000 ;
	    RECT 344.6000 296.0000 345.4000 299.0000 ;
	    RECT 344.6000 295.4000 346.2000 296.0000 ;
	    RECT 345.4000 295.0000 346.2000 295.4000 ;
	    RECT 311.6000 291.6000 312.4000 293.2000 ;
	    RECT 313.4000 290.2000 314.0000 293.6000 ;
	    RECT 314.8000 291.6000 315.6000 293.2000 ;
	    RECT 318.0000 290.2000 318.8000 290.4000 ;
	    RECT 320.0000 290.2000 320.6000 293.6000 ;
	    RECT 321.2000 291.6000 322.0000 293.2000 ;
	    RECT 324.4000 290.2000 325.2000 290.4000 ;
	    RECT 326.4000 290.2000 327.0000 293.6000 ;
	    RECT 327.6000 292.3000 328.4000 293.2000 ;
	    RECT 329.2000 292.3000 330.0000 292.4000 ;
	    RECT 330.8000 292.3000 331.6000 293.2000 ;
	    RECT 327.6000 291.7000 331.6000 292.3000 ;
	    RECT 327.6000 291.6000 328.4000 291.7000 ;
	    RECT 329.2000 291.6000 330.0000 291.7000 ;
	    RECT 330.8000 291.6000 331.6000 291.7000 ;
	    RECT 332.4000 291.6000 333.2000 293.2000 ;
	    RECT 334.0000 293.0000 335.4000 293.8000 ;
	    RECT 336.0000 293.6000 338.0000 294.4000 ;
	    RECT 340.4000 294.2000 344.6000 294.8000 ;
	    RECT 343.6000 293.8000 344.6000 294.2000 ;
	    RECT 345.6000 294.4000 346.2000 295.0000 ;
	    RECT 350.0000 295.4000 350.8000 299.8000 ;
	    RECT 354.2000 298.4000 355.4000 299.8000 ;
	    RECT 354.2000 297.8000 355.6000 298.4000 ;
	    RECT 358.8000 297.8000 359.6000 299.8000 ;
	    RECT 363.2000 298.4000 364.0000 299.8000 ;
	    RECT 363.2000 297.8000 365.2000 298.4000 ;
	    RECT 354.8000 297.0000 355.6000 297.8000 ;
	    RECT 359.0000 297.2000 359.6000 297.8000 ;
	    RECT 359.0000 296.6000 361.8000 297.2000 ;
	    RECT 361.0000 296.4000 361.8000 296.6000 ;
	    RECT 362.8000 296.4000 363.6000 297.2000 ;
	    RECT 364.4000 297.0000 365.2000 297.8000 ;
	    RECT 353.0000 295.4000 353.8000 295.6000 ;
	    RECT 350.0000 294.8000 353.8000 295.4000 ;
	    RECT 334.0000 291.0000 334.6000 293.0000 ;
	    RECT 330.8000 290.4000 334.6000 291.0000 ;
	    RECT 336.0000 290.4000 336.6000 293.6000 ;
	    RECT 337.2000 290.8000 338.0000 292.4000 ;
	    RECT 340.4000 291.6000 341.2000 293.2000 ;
	    RECT 342.0000 291.6000 342.8000 293.2000 ;
	    RECT 343.6000 293.0000 345.0000 293.8000 ;
	    RECT 345.6000 293.6000 347.6000 294.4000 ;
	    RECT 343.6000 291.0000 344.2000 293.0000 ;
	    RECT 260.4000 289.6000 261.8000 290.2000 ;
	    RECT 262.4000 289.6000 263.4000 290.2000 ;
	    RECT 244.4000 283.0000 245.2000 287.0000 ;
	    RECT 248.6000 284.4000 249.4000 289.2000 ;
	    RECT 261.2000 288.4000 261.8000 289.6000 ;
	    RECT 261.2000 287.6000 262.0000 288.4000 ;
	    RECT 247.6000 283.6000 249.4000 284.4000 ;
	    RECT 248.6000 282.2000 249.4000 283.6000 ;
	    RECT 262.6000 282.2000 263.4000 289.6000 ;
	    RECT 268.4000 289.4000 270.2000 290.2000 ;
	    RECT 269.4000 288.4000 270.2000 289.4000 ;
	    RECT 269.4000 287.6000 270.8000 288.4000 ;
	    RECT 269.4000 282.2000 270.2000 287.6000 ;
	    RECT 274.2000 284.4000 276.2000 290.2000 ;
	    RECT 273.2000 283.6000 276.2000 284.4000 ;
	    RECT 274.2000 282.2000 276.2000 283.6000 ;
	    RECT 282.2000 289.6000 283.2000 290.2000 ;
	    RECT 283.8000 289.6000 285.2000 290.2000 ;
	    RECT 282.2000 282.2000 283.0000 289.6000 ;
	    RECT 283.8000 288.4000 284.4000 289.6000 ;
	    RECT 288.6000 288.4000 290.6000 290.2000 ;
	    RECT 295.6000 289.4000 297.4000 290.2000 ;
	    RECT 298.8000 289.6000 300.2000 290.2000 ;
	    RECT 300.8000 289.6000 301.8000 290.2000 ;
	    RECT 283.6000 287.6000 284.4000 288.4000 ;
	    RECT 287.6000 287.6000 290.6000 288.4000 ;
	    RECT 288.6000 282.2000 290.6000 287.6000 ;
	    RECT 296.6000 282.2000 297.4000 289.4000 ;
	    RECT 299.6000 288.4000 300.2000 289.6000 ;
	    RECT 299.6000 287.6000 300.4000 288.4000 ;
	    RECT 301.0000 282.2000 301.8000 289.6000 ;
	    RECT 305.8000 289.4000 307.6000 290.2000 ;
	    RECT 305.8000 282.2000 306.6000 289.4000 ;
	    RECT 312.6000 282.2000 314.6000 290.2000 ;
	    RECT 318.0000 289.6000 319.4000 290.2000 ;
	    RECT 320.0000 289.6000 321.0000 290.2000 ;
	    RECT 324.4000 289.6000 325.8000 290.2000 ;
	    RECT 326.4000 289.6000 327.4000 290.2000 ;
	    RECT 318.8000 288.4000 319.4000 289.6000 ;
	    RECT 318.8000 287.6000 319.6000 288.4000 ;
	    RECT 320.2000 282.2000 321.0000 289.6000 ;
	    RECT 325.2000 288.4000 325.8000 289.6000 ;
	    RECT 325.2000 287.6000 326.0000 288.4000 ;
	    RECT 326.6000 286.4000 327.4000 289.6000 ;
	    RECT 330.8000 287.0000 331.4000 290.4000 ;
	    RECT 335.6000 289.8000 336.6000 290.4000 ;
	    RECT 335.0000 289.2000 336.6000 289.8000 ;
	    RECT 340.4000 290.4000 344.2000 291.0000 ;
	    RECT 326.6000 285.6000 328.4000 286.4000 ;
	    RECT 326.6000 282.2000 327.4000 285.6000 ;
	    RECT 330.8000 283.0000 331.6000 287.0000 ;
	    RECT 335.0000 282.2000 335.8000 289.2000 ;
	    RECT 340.4000 287.0000 341.0000 290.4000 ;
	    RECT 345.6000 289.8000 346.2000 293.6000 ;
	    RECT 346.8000 290.8000 347.6000 292.4000 ;
	    RECT 350.0000 291.4000 350.8000 294.8000 ;
	    RECT 357.0000 294.2000 357.8000 294.4000 ;
	    RECT 361.2000 294.2000 362.0000 294.4000 ;
	    RECT 362.8000 294.2000 363.4000 296.4000 ;
	    RECT 367.6000 295.0000 368.4000 299.8000 ;
	    RECT 371.8000 296.4000 372.6000 299.8000 ;
	    RECT 370.8000 295.8000 372.6000 296.4000 ;
	    RECT 374.0000 295.8000 374.8000 299.8000 ;
	    RECT 375.6000 296.0000 376.4000 299.8000 ;
	    RECT 378.8000 296.0000 379.6000 299.8000 ;
	    RECT 375.6000 295.8000 379.6000 296.0000 ;
	    RECT 366.0000 294.2000 367.6000 294.4000 ;
	    RECT 356.6000 293.6000 367.6000 294.2000 ;
	    RECT 369.2000 293.6000 370.0000 295.2000 ;
	    RECT 354.8000 292.8000 355.6000 293.0000 ;
	    RECT 351.8000 292.2000 355.6000 292.8000 ;
	    RECT 351.8000 292.0000 352.6000 292.2000 ;
	    RECT 353.4000 291.4000 354.2000 291.6000 ;
	    RECT 350.0000 290.8000 354.2000 291.4000 ;
	    RECT 344.6000 289.2000 346.2000 289.8000 ;
	    RECT 340.4000 283.0000 341.2000 287.0000 ;
	    RECT 344.6000 284.4000 345.4000 289.2000 ;
	    RECT 343.6000 283.6000 345.4000 284.4000 ;
	    RECT 344.6000 282.2000 345.4000 283.6000 ;
	    RECT 350.0000 282.2000 350.8000 290.8000 ;
	    RECT 356.6000 290.4000 357.2000 293.6000 ;
	    RECT 363.8000 293.4000 364.6000 293.6000 ;
	    RECT 365.4000 292.4000 366.2000 292.6000 ;
	    RECT 361.2000 291.8000 366.2000 292.4000 ;
	    RECT 370.8000 292.3000 371.6000 295.8000 ;
	    RECT 374.2000 294.4000 374.8000 295.8000 ;
	    RECT 375.8000 295.4000 379.4000 295.8000 ;
	    RECT 378.0000 294.4000 378.8000 294.8000 ;
	    RECT 374.0000 293.6000 376.6000 294.4000 ;
	    RECT 378.0000 293.8000 379.6000 294.4000 ;
	    RECT 378.8000 293.6000 379.6000 293.8000 ;
	    RECT 376.0000 292.4000 376.6000 293.6000 ;
	    RECT 361.2000 291.6000 362.0000 291.8000 ;
	    RECT 370.8000 291.7000 374.7000 292.3000 ;
	    RECT 362.8000 291.0000 368.4000 291.2000 ;
	    RECT 362.6000 290.8000 368.4000 291.0000 ;
	    RECT 354.8000 289.8000 357.2000 290.4000 ;
	    RECT 358.6000 290.6000 368.4000 290.8000 ;
	    RECT 358.6000 290.2000 363.4000 290.6000 ;
	    RECT 354.8000 288.8000 355.4000 289.8000 ;
	    RECT 354.0000 288.0000 355.4000 288.8000 ;
	    RECT 357.0000 289.0000 357.8000 289.2000 ;
	    RECT 358.6000 289.0000 359.2000 290.2000 ;
	    RECT 357.0000 288.4000 359.2000 289.0000 ;
	    RECT 359.8000 289.0000 365.2000 289.6000 ;
	    RECT 359.8000 288.8000 360.6000 289.0000 ;
	    RECT 364.4000 288.8000 365.2000 289.0000 ;
	    RECT 358.2000 287.4000 359.0000 287.6000 ;
	    RECT 361.0000 287.4000 361.8000 287.6000 ;
	    RECT 354.8000 286.2000 355.6000 287.0000 ;
	    RECT 358.2000 286.8000 361.8000 287.4000 ;
	    RECT 359.0000 286.2000 359.6000 286.8000 ;
	    RECT 364.4000 286.2000 365.2000 287.0000 ;
	    RECT 354.2000 282.2000 355.4000 286.2000 ;
	    RECT 358.8000 282.2000 359.6000 286.2000 ;
	    RECT 363.2000 285.6000 365.2000 286.2000 ;
	    RECT 363.2000 282.2000 364.0000 285.6000 ;
	    RECT 367.6000 282.2000 368.4000 290.6000 ;
	    RECT 370.8000 282.2000 371.6000 291.7000 ;
	    RECT 374.1000 290.4000 374.7000 291.7000 ;
	    RECT 375.6000 291.6000 376.6000 292.4000 ;
	    RECT 377.2000 292.3000 378.0000 293.2000 ;
	    RECT 378.8000 292.3000 379.6000 292.4000 ;
	    RECT 377.2000 291.7000 379.6000 292.3000 ;
	    RECT 377.2000 291.6000 378.0000 291.7000 ;
	    RECT 378.8000 291.6000 379.6000 291.7000 ;
	    RECT 372.4000 288.8000 373.2000 290.4000 ;
	    RECT 374.0000 290.2000 374.8000 290.4000 ;
	    RECT 376.0000 290.2000 376.6000 291.6000 ;
	    RECT 374.0000 289.6000 375.4000 290.2000 ;
	    RECT 376.0000 289.6000 377.0000 290.2000 ;
	    RECT 374.8000 288.4000 375.4000 289.6000 ;
	    RECT 374.8000 287.6000 375.6000 288.4000 ;
	    RECT 376.2000 282.2000 377.0000 289.6000 ;
	    RECT 380.4000 282.2000 381.2000 299.8000 ;
	    RECT 383.6000 295.4000 384.4000 299.8000 ;
	    RECT 387.8000 298.4000 389.0000 299.8000 ;
	    RECT 387.8000 297.8000 389.2000 298.4000 ;
	    RECT 392.4000 297.8000 393.2000 299.8000 ;
	    RECT 396.8000 298.4000 397.6000 299.8000 ;
	    RECT 396.8000 297.8000 398.8000 298.4000 ;
	    RECT 388.4000 297.0000 389.2000 297.8000 ;
	    RECT 392.6000 297.2000 393.2000 297.8000 ;
	    RECT 392.6000 296.6000 395.4000 297.2000 ;
	    RECT 394.6000 296.4000 395.4000 296.6000 ;
	    RECT 396.4000 296.4000 397.2000 297.2000 ;
	    RECT 398.0000 297.0000 398.8000 297.8000 ;
	    RECT 386.6000 295.4000 387.4000 295.6000 ;
	    RECT 383.6000 294.8000 387.4000 295.4000 ;
	    RECT 383.6000 291.4000 384.4000 294.8000 ;
	    RECT 390.6000 294.2000 392.4000 294.4000 ;
	    RECT 394.8000 294.2000 395.6000 294.4000 ;
	    RECT 396.4000 294.2000 397.0000 296.4000 ;
	    RECT 401.2000 295.0000 402.0000 299.8000 ;
	    RECT 402.8000 295.8000 403.6000 299.8000 ;
	    RECT 404.4000 296.0000 405.2000 299.8000 ;
	    RECT 407.6000 296.0000 408.4000 299.8000 ;
	    RECT 404.4000 295.8000 408.4000 296.0000 ;
	    RECT 415.6000 296.0000 416.4000 299.8000 ;
	    RECT 418.8000 296.0000 419.6000 299.8000 ;
	    RECT 415.6000 295.8000 419.6000 296.0000 ;
	    RECT 420.4000 295.8000 421.2000 299.8000 ;
	    RECT 403.0000 294.4000 403.6000 295.8000 ;
	    RECT 404.6000 295.4000 408.2000 295.8000 ;
	    RECT 415.8000 295.4000 419.4000 295.8000 ;
	    RECT 406.8000 294.4000 407.6000 294.8000 ;
	    RECT 416.4000 294.4000 417.2000 294.8000 ;
	    RECT 420.4000 294.4000 421.0000 295.8000 ;
	    RECT 399.6000 294.2000 401.2000 294.4000 ;
	    RECT 390.2000 293.6000 401.2000 294.2000 ;
	    RECT 402.8000 293.6000 405.4000 294.4000 ;
	    RECT 406.8000 293.8000 408.4000 294.4000 ;
	    RECT 407.6000 293.6000 408.4000 293.8000 ;
	    RECT 415.6000 293.8000 417.2000 294.4000 ;
	    RECT 415.6000 293.6000 416.4000 293.8000 ;
	    RECT 418.6000 293.6000 421.2000 294.4000 ;
	    RECT 388.4000 292.8000 389.2000 293.0000 ;
	    RECT 385.4000 292.2000 389.2000 292.8000 ;
	    RECT 385.4000 292.0000 386.2000 292.2000 ;
	    RECT 387.0000 291.4000 387.8000 291.6000 ;
	    RECT 383.6000 290.8000 387.8000 291.4000 ;
	    RECT 383.6000 282.2000 384.4000 290.8000 ;
	    RECT 390.2000 290.4000 390.8000 293.6000 ;
	    RECT 397.4000 293.4000 398.2000 293.6000 ;
	    RECT 396.4000 292.4000 397.2000 292.6000 ;
	    RECT 399.0000 292.4000 399.8000 292.6000 ;
	    RECT 394.8000 291.8000 399.8000 292.4000 ;
	    RECT 394.8000 291.6000 395.6000 291.8000 ;
	    RECT 396.4000 291.0000 402.0000 291.2000 ;
	    RECT 396.2000 290.8000 402.0000 291.0000 ;
	    RECT 388.4000 289.8000 390.8000 290.4000 ;
	    RECT 392.2000 290.6000 402.0000 290.8000 ;
	    RECT 392.2000 290.2000 397.0000 290.6000 ;
	    RECT 388.4000 288.8000 389.0000 289.8000 ;
	    RECT 387.6000 288.0000 389.0000 288.8000 ;
	    RECT 390.6000 289.0000 391.4000 289.2000 ;
	    RECT 392.2000 289.0000 392.8000 290.2000 ;
	    RECT 390.6000 288.4000 392.8000 289.0000 ;
	    RECT 393.4000 289.0000 398.8000 289.6000 ;
	    RECT 393.4000 288.8000 394.2000 289.0000 ;
	    RECT 398.0000 288.8000 398.8000 289.0000 ;
	    RECT 391.8000 287.4000 392.6000 287.6000 ;
	    RECT 394.6000 287.4000 395.4000 287.6000 ;
	    RECT 388.4000 286.2000 389.2000 287.0000 ;
	    RECT 391.8000 286.8000 395.4000 287.4000 ;
	    RECT 392.6000 286.2000 393.2000 286.8000 ;
	    RECT 398.0000 286.2000 398.8000 287.0000 ;
	    RECT 387.8000 282.2000 389.0000 286.2000 ;
	    RECT 392.4000 282.2000 393.2000 286.2000 ;
	    RECT 396.8000 285.6000 398.8000 286.2000 ;
	    RECT 396.8000 282.2000 397.6000 285.6000 ;
	    RECT 401.2000 282.2000 402.0000 290.6000 ;
	    RECT 402.8000 290.2000 403.6000 290.4000 ;
	    RECT 404.8000 290.2000 405.4000 293.6000 ;
	    RECT 406.0000 292.3000 406.8000 293.2000 ;
	    RECT 417.2000 292.3000 418.0000 293.2000 ;
	    RECT 406.0000 291.7000 418.0000 292.3000 ;
	    RECT 406.0000 291.6000 406.8000 291.7000 ;
	    RECT 417.2000 291.6000 418.0000 291.7000 ;
	    RECT 418.6000 290.2000 419.2000 293.6000 ;
	    RECT 420.4000 290.2000 421.2000 290.4000 ;
	    RECT 402.8000 289.6000 404.2000 290.2000 ;
	    RECT 404.8000 289.6000 405.8000 290.2000 ;
	    RECT 403.6000 288.4000 404.2000 289.6000 ;
	    RECT 403.6000 287.6000 404.4000 288.4000 ;
	    RECT 405.0000 282.2000 405.8000 289.6000 ;
	    RECT 418.2000 289.6000 419.2000 290.2000 ;
	    RECT 419.8000 289.6000 421.2000 290.2000 ;
	    RECT 418.2000 282.2000 419.0000 289.6000 ;
	    RECT 419.8000 288.4000 420.4000 289.6000 ;
	    RECT 419.6000 287.6000 420.4000 288.4000 ;
	    RECT 422.0000 282.2000 422.8000 299.8000 ;
	    RECT 425.2000 296.0000 426.0000 299.8000 ;
	    RECT 428.4000 296.0000 429.2000 299.8000 ;
	    RECT 425.2000 295.8000 429.2000 296.0000 ;
	    RECT 430.0000 295.8000 430.8000 299.8000 ;
	    RECT 432.2000 296.4000 433.0000 299.8000 ;
	    RECT 432.2000 295.8000 434.0000 296.4000 ;
	    RECT 425.4000 295.4000 429.0000 295.8000 ;
	    RECT 426.0000 294.4000 426.8000 294.8000 ;
	    RECT 430.0000 294.4000 430.6000 295.8000 ;
	    RECT 425.2000 293.8000 426.8000 294.4000 ;
	    RECT 428.2000 294.3000 430.8000 294.4000 ;
	    RECT 431.6000 294.3000 432.4000 294.4000 ;
	    RECT 425.2000 293.6000 426.0000 293.8000 ;
	    RECT 428.2000 293.7000 432.4000 294.3000 ;
	    RECT 428.2000 293.6000 430.8000 293.7000 ;
	    RECT 431.6000 293.6000 432.4000 293.7000 ;
	    RECT 426.8000 291.6000 427.6000 293.2000 ;
	    RECT 428.2000 290.2000 428.8000 293.6000 ;
	    RECT 433.2000 292.3000 434.0000 295.8000 ;
	    RECT 436.4000 295.4000 437.2000 299.8000 ;
	    RECT 440.6000 298.4000 441.8000 299.8000 ;
	    RECT 440.6000 297.8000 442.0000 298.4000 ;
	    RECT 445.2000 297.8000 446.0000 299.8000 ;
	    RECT 449.6000 298.4000 450.4000 299.8000 ;
	    RECT 449.6000 297.8000 451.6000 298.4000 ;
	    RECT 441.2000 297.0000 442.0000 297.8000 ;
	    RECT 445.4000 297.2000 446.0000 297.8000 ;
	    RECT 445.4000 296.6000 448.2000 297.2000 ;
	    RECT 447.4000 296.4000 448.2000 296.6000 ;
	    RECT 449.2000 296.4000 450.0000 297.2000 ;
	    RECT 450.8000 297.0000 451.6000 297.8000 ;
	    RECT 439.4000 295.4000 440.2000 295.6000 ;
	    RECT 434.8000 293.6000 435.6000 295.2000 ;
	    RECT 436.4000 294.8000 440.2000 295.4000 ;
	    RECT 430.1000 291.7000 434.0000 292.3000 ;
	    RECT 430.1000 290.4000 430.7000 291.7000 ;
	    RECT 430.0000 290.2000 430.8000 290.4000 ;
	    RECT 427.8000 289.6000 428.8000 290.2000 ;
	    RECT 429.4000 289.6000 430.8000 290.2000 ;
	    RECT 427.8000 282.2000 428.6000 289.6000 ;
	    RECT 429.4000 288.4000 430.0000 289.6000 ;
	    RECT 431.6000 288.8000 432.4000 290.4000 ;
	    RECT 429.2000 287.6000 430.0000 288.4000 ;
	    RECT 433.2000 282.2000 434.0000 291.7000 ;
	    RECT 436.4000 291.4000 437.2000 294.8000 ;
	    RECT 443.4000 294.2000 444.2000 294.4000 ;
	    RECT 449.2000 294.2000 449.8000 296.4000 ;
	    RECT 454.0000 295.0000 454.8000 299.8000 ;
	    RECT 452.4000 294.2000 454.0000 294.4000 ;
	    RECT 443.0000 293.6000 454.0000 294.2000 ;
	    RECT 459.2000 294.2000 460.0000 299.8000 ;
	    RECT 462.0000 295.6000 462.8000 297.2000 ;
	    RECT 463.6000 294.3000 464.4000 299.8000 ;
	    RECT 465.2000 296.0000 466.0000 299.8000 ;
	    RECT 468.4000 296.0000 469.2000 299.8000 ;
	    RECT 465.2000 295.8000 469.2000 296.0000 ;
	    RECT 470.0000 295.8000 470.8000 299.8000 ;
	    RECT 465.4000 295.4000 469.0000 295.8000 ;
	    RECT 466.0000 294.4000 466.8000 294.8000 ;
	    RECT 470.0000 294.4000 470.6000 295.8000 ;
	    RECT 471.6000 295.4000 472.4000 299.8000 ;
	    RECT 475.8000 298.4000 477.0000 299.8000 ;
	    RECT 475.8000 297.8000 477.2000 298.4000 ;
	    RECT 480.4000 297.8000 481.2000 299.8000 ;
	    RECT 484.8000 298.4000 485.6000 299.8000 ;
	    RECT 484.8000 297.8000 486.8000 298.4000 ;
	    RECT 476.4000 297.0000 477.2000 297.8000 ;
	    RECT 480.6000 297.2000 481.2000 297.8000 ;
	    RECT 480.6000 296.6000 483.4000 297.2000 ;
	    RECT 482.6000 296.4000 483.4000 296.6000 ;
	    RECT 484.4000 296.4000 485.2000 297.2000 ;
	    RECT 486.0000 297.0000 486.8000 297.8000 ;
	    RECT 474.6000 295.4000 475.4000 295.6000 ;
	    RECT 471.6000 294.8000 475.4000 295.4000 ;
	    RECT 465.2000 294.3000 466.8000 294.4000 ;
	    RECT 459.2000 293.8000 461.0000 294.2000 ;
	    RECT 459.4000 293.6000 461.0000 293.8000 ;
	    RECT 441.2000 292.8000 442.0000 293.0000 ;
	    RECT 438.2000 292.2000 442.0000 292.8000 ;
	    RECT 438.2000 292.0000 439.0000 292.2000 ;
	    RECT 439.8000 291.4000 440.6000 291.6000 ;
	    RECT 436.4000 290.8000 440.6000 291.4000 ;
	    RECT 436.4000 282.2000 437.2000 290.8000 ;
	    RECT 443.0000 290.4000 443.6000 293.6000 ;
	    RECT 450.2000 293.4000 451.0000 293.6000 ;
	    RECT 451.8000 292.4000 452.6000 292.6000 ;
	    RECT 444.4000 292.3000 445.2000 292.4000 ;
	    RECT 447.6000 292.3000 452.6000 292.4000 ;
	    RECT 444.4000 291.8000 452.6000 292.3000 ;
	    RECT 444.4000 291.7000 448.4000 291.8000 ;
	    RECT 444.4000 291.6000 445.2000 291.7000 ;
	    RECT 447.6000 291.6000 448.4000 291.7000 ;
	    RECT 457.2000 291.6000 458.8000 292.4000 ;
	    RECT 449.2000 291.0000 454.8000 291.2000 ;
	    RECT 449.0000 290.8000 454.8000 291.0000 ;
	    RECT 441.2000 289.8000 443.6000 290.4000 ;
	    RECT 445.0000 290.6000 454.8000 290.8000 ;
	    RECT 445.0000 290.2000 449.8000 290.6000 ;
	    RECT 441.2000 288.8000 441.8000 289.8000 ;
	    RECT 440.4000 288.0000 441.8000 288.8000 ;
	    RECT 443.4000 289.0000 444.2000 289.2000 ;
	    RECT 445.0000 289.0000 445.6000 290.2000 ;
	    RECT 443.4000 288.4000 445.6000 289.0000 ;
	    RECT 446.2000 289.0000 451.6000 289.6000 ;
	    RECT 446.2000 288.8000 447.0000 289.0000 ;
	    RECT 450.8000 288.8000 451.6000 289.0000 ;
	    RECT 444.6000 287.4000 445.4000 287.6000 ;
	    RECT 447.4000 287.4000 448.2000 287.6000 ;
	    RECT 441.2000 286.2000 442.0000 287.0000 ;
	    RECT 444.6000 286.8000 448.2000 287.4000 ;
	    RECT 445.4000 286.2000 446.0000 286.8000 ;
	    RECT 450.8000 286.2000 451.6000 287.0000 ;
	    RECT 440.6000 282.2000 441.8000 286.2000 ;
	    RECT 445.2000 282.2000 446.0000 286.2000 ;
	    RECT 449.6000 285.6000 451.6000 286.2000 ;
	    RECT 449.6000 282.2000 450.4000 285.6000 ;
	    RECT 454.0000 282.2000 454.8000 290.6000 ;
	    RECT 460.4000 290.4000 461.0000 293.6000 ;
	    RECT 463.6000 293.8000 466.8000 294.3000 ;
	    RECT 463.6000 293.7000 466.0000 293.8000 ;
	    RECT 460.4000 289.6000 461.2000 290.4000 ;
	    RECT 458.8000 287.6000 459.6000 289.2000 ;
	    RECT 460.4000 288.3000 461.0000 289.6000 ;
	    RECT 462.0000 288.3000 462.8000 288.4000 ;
	    RECT 460.4000 287.7000 462.8000 288.3000 ;
	    RECT 460.4000 287.0000 461.0000 287.7000 ;
	    RECT 462.0000 287.6000 462.8000 287.7000 ;
	    RECT 457.4000 286.4000 461.0000 287.0000 ;
	    RECT 457.4000 286.2000 458.0000 286.4000 ;
	    RECT 457.2000 282.2000 458.0000 286.2000 ;
	    RECT 460.4000 286.2000 461.0000 286.4000 ;
	    RECT 460.4000 282.2000 461.2000 286.2000 ;
	    RECT 463.6000 282.2000 464.4000 293.7000 ;
	    RECT 465.2000 293.6000 466.0000 293.7000 ;
	    RECT 468.2000 293.6000 470.8000 294.4000 ;
	    RECT 466.8000 291.6000 467.6000 293.2000 ;
	    RECT 468.2000 290.2000 468.8000 293.6000 ;
	    RECT 471.6000 291.4000 472.4000 294.8000 ;
	    RECT 478.6000 294.2000 479.4000 294.4000 ;
	    RECT 484.4000 294.2000 485.0000 296.4000 ;
	    RECT 489.2000 295.0000 490.0000 299.8000 ;
	    RECT 487.6000 294.2000 489.2000 294.4000 ;
	    RECT 478.2000 293.6000 489.2000 294.2000 ;
	    RECT 494.4000 294.2000 495.2000 299.8000 ;
	    RECT 500.8000 294.2000 501.6000 299.8000 ;
	    RECT 507.2000 294.2000 508.0000 299.8000 ;
	    RECT 494.4000 293.8000 496.2000 294.2000 ;
	    RECT 500.8000 293.8000 502.6000 294.2000 ;
	    RECT 507.2000 293.8000 509.0000 294.2000 ;
	    RECT 494.6000 293.6000 496.2000 293.8000 ;
	    RECT 501.0000 293.6000 502.6000 293.8000 ;
	    RECT 507.4000 293.6000 509.0000 293.8000 ;
	    RECT 476.4000 292.8000 477.2000 293.0000 ;
	    RECT 473.4000 292.2000 477.2000 292.8000 ;
	    RECT 478.2000 292.3000 478.8000 293.6000 ;
	    RECT 485.4000 293.4000 486.2000 293.6000 ;
	    RECT 487.0000 292.4000 487.8000 292.6000 ;
	    RECT 479.6000 292.3000 480.4000 292.4000 ;
	    RECT 473.4000 292.0000 474.2000 292.2000 ;
	    RECT 478.1000 291.7000 480.4000 292.3000 ;
	    RECT 475.0000 291.4000 475.8000 291.6000 ;
	    RECT 471.6000 290.8000 475.8000 291.4000 ;
	    RECT 470.0000 290.2000 470.8000 290.4000 ;
	    RECT 467.8000 289.6000 468.8000 290.2000 ;
	    RECT 469.4000 289.6000 470.8000 290.2000 ;
	    RECT 467.8000 282.2000 468.6000 289.6000 ;
	    RECT 469.4000 288.4000 470.0000 289.6000 ;
	    RECT 469.2000 287.6000 470.0000 288.4000 ;
	    RECT 471.6000 282.2000 472.4000 290.8000 ;
	    RECT 478.2000 290.4000 478.8000 291.7000 ;
	    RECT 479.6000 291.6000 480.4000 291.7000 ;
	    RECT 482.8000 291.8000 487.8000 292.4000 ;
	    RECT 482.8000 291.6000 483.6000 291.8000 ;
	    RECT 492.4000 291.6000 494.0000 292.4000 ;
	    RECT 484.4000 291.0000 490.0000 291.2000 ;
	    RECT 484.2000 290.8000 490.0000 291.0000 ;
	    RECT 476.4000 289.8000 478.8000 290.4000 ;
	    RECT 480.2000 290.6000 490.0000 290.8000 ;
	    RECT 480.2000 290.2000 485.0000 290.6000 ;
	    RECT 476.4000 288.8000 477.0000 289.8000 ;
	    RECT 475.6000 288.4000 477.0000 288.8000 ;
	    RECT 478.6000 289.0000 479.4000 289.2000 ;
	    RECT 480.2000 289.0000 480.8000 290.2000 ;
	    RECT 478.6000 288.4000 480.8000 289.0000 ;
	    RECT 481.4000 289.0000 486.8000 289.6000 ;
	    RECT 481.4000 288.8000 482.2000 289.0000 ;
	    RECT 486.0000 288.8000 486.8000 289.0000 ;
	    RECT 474.8000 288.0000 477.0000 288.4000 ;
	    RECT 474.8000 287.6000 476.2000 288.0000 ;
	    RECT 479.8000 287.4000 480.6000 287.6000 ;
	    RECT 482.6000 287.4000 483.4000 287.6000 ;
	    RECT 476.4000 286.2000 477.2000 287.0000 ;
	    RECT 479.8000 286.8000 483.4000 287.4000 ;
	    RECT 480.6000 286.2000 481.2000 286.8000 ;
	    RECT 486.0000 286.2000 486.8000 287.0000 ;
	    RECT 475.8000 282.2000 477.0000 286.2000 ;
	    RECT 480.4000 282.2000 481.2000 286.2000 ;
	    RECT 484.8000 285.6000 486.8000 286.2000 ;
	    RECT 484.8000 282.2000 485.6000 285.6000 ;
	    RECT 489.2000 282.2000 490.0000 290.6000 ;
	    RECT 495.6000 290.4000 496.2000 293.6000 ;
	    RECT 498.8000 291.6000 500.4000 292.4000 ;
	    RECT 502.0000 290.4000 502.6000 293.6000 ;
	    RECT 505.2000 291.6000 506.8000 292.4000 ;
	    RECT 508.4000 290.4000 509.0000 293.6000 ;
	    RECT 495.6000 289.6000 496.4000 290.4000 ;
	    RECT 502.0000 289.6000 502.8000 290.4000 ;
	    RECT 508.4000 289.6000 509.2000 290.4000 ;
	    RECT 494.0000 287.6000 494.8000 289.2000 ;
	    RECT 495.6000 287.0000 496.2000 289.6000 ;
	    RECT 497.2000 288.3000 498.0000 288.4000 ;
	    RECT 500.4000 288.3000 501.2000 289.2000 ;
	    RECT 497.2000 287.7000 501.2000 288.3000 ;
	    RECT 497.2000 287.6000 498.0000 287.7000 ;
	    RECT 500.4000 287.6000 501.2000 287.7000 ;
	    RECT 502.0000 287.0000 502.6000 289.6000 ;
	    RECT 506.8000 287.6000 507.6000 289.2000 ;
	    RECT 508.4000 287.0000 509.0000 289.6000 ;
	    RECT 492.6000 286.4000 496.2000 287.0000 ;
	    RECT 492.6000 286.2000 493.2000 286.4000 ;
	    RECT 492.4000 282.2000 493.2000 286.2000 ;
	    RECT 495.6000 286.2000 496.2000 286.4000 ;
	    RECT 499.0000 286.4000 502.6000 287.0000 ;
	    RECT 499.0000 286.2000 499.6000 286.4000 ;
	    RECT 495.6000 282.2000 496.4000 286.2000 ;
	    RECT 498.8000 282.2000 499.6000 286.2000 ;
	    RECT 502.0000 286.2000 502.6000 286.4000 ;
	    RECT 505.4000 286.4000 509.0000 287.0000 ;
	    RECT 505.4000 286.2000 506.0000 286.4000 ;
	    RECT 502.0000 282.2000 502.8000 286.2000 ;
	    RECT 505.2000 282.2000 506.0000 286.2000 ;
	    RECT 508.4000 286.2000 509.0000 286.4000 ;
	    RECT 508.4000 282.2000 509.2000 286.2000 ;
	    RECT 4.4000 272.4000 5.2000 279.8000 ;
	    RECT 6.8000 273.6000 7.6000 274.4000 ;
	    RECT 6.8000 272.4000 7.4000 273.6000 ;
	    RECT 8.2000 272.4000 9.0000 279.8000 ;
	    RECT 3.0000 271.8000 5.2000 272.4000 ;
	    RECT 6.0000 271.8000 7.4000 272.4000 ;
	    RECT 8.0000 271.8000 9.0000 272.4000 ;
	    RECT 15.0000 272.4000 15.8000 279.8000 ;
	    RECT 16.4000 274.3000 17.2000 274.4000 ;
	    RECT 18.8000 274.3000 19.6000 279.8000 ;
	    RECT 23.0000 275.8000 24.2000 279.8000 ;
	    RECT 27.6000 275.8000 28.4000 279.8000 ;
	    RECT 32.0000 276.4000 32.8000 279.8000 ;
	    RECT 32.0000 275.8000 34.0000 276.4000 ;
	    RECT 23.6000 275.0000 24.4000 275.8000 ;
	    RECT 27.8000 275.2000 28.4000 275.8000 ;
	    RECT 27.0000 274.6000 30.6000 275.2000 ;
	    RECT 33.2000 275.0000 34.0000 275.8000 ;
	    RECT 27.0000 274.4000 27.8000 274.6000 ;
	    RECT 29.8000 274.4000 30.6000 274.6000 ;
	    RECT 16.4000 273.7000 19.6000 274.3000 ;
	    RECT 16.4000 273.6000 17.2000 273.7000 ;
	    RECT 16.6000 272.4000 17.2000 273.6000 ;
	    RECT 15.0000 271.8000 16.0000 272.4000 ;
	    RECT 16.6000 271.8000 18.0000 272.4000 ;
	    RECT 3.0000 271.2000 3.6000 271.8000 ;
	    RECT 6.0000 271.6000 6.8000 271.8000 ;
	    RECT 2.4000 270.4000 3.6000 271.2000 ;
	    RECT 3.0000 267.4000 3.6000 270.4000 ;
	    RECT 4.4000 268.8000 5.2000 270.4000 ;
	    RECT 8.0000 268.4000 8.6000 271.8000 ;
	    RECT 9.2000 270.3000 10.0000 270.4000 ;
	    RECT 14.0000 270.3000 14.8000 270.4000 ;
	    RECT 9.2000 269.7000 14.8000 270.3000 ;
	    RECT 9.2000 268.8000 10.0000 269.7000 ;
	    RECT 14.0000 268.8000 14.8000 269.7000 ;
	    RECT 15.4000 270.3000 16.0000 271.8000 ;
	    RECT 17.2000 271.6000 18.0000 271.8000 ;
	    RECT 18.8000 271.2000 19.6000 273.7000 ;
	    RECT 22.8000 273.2000 24.2000 274.0000 ;
	    RECT 23.6000 272.2000 24.2000 273.2000 ;
	    RECT 25.8000 273.0000 28.0000 273.6000 ;
	    RECT 25.8000 272.8000 26.6000 273.0000 ;
	    RECT 23.6000 271.6000 26.0000 272.2000 ;
	    RECT 18.8000 270.6000 23.0000 271.2000 ;
	    RECT 17.2000 270.3000 18.0000 270.4000 ;
	    RECT 15.4000 269.7000 18.0000 270.3000 ;
	    RECT 15.4000 268.4000 16.0000 269.7000 ;
	    RECT 17.2000 269.6000 18.0000 269.7000 ;
	    RECT 6.0000 267.6000 8.6000 268.4000 ;
	    RECT 10.8000 268.3000 11.6000 268.4000 ;
	    RECT 12.4000 268.3000 13.2000 268.4000 ;
	    RECT 10.8000 268.2000 13.2000 268.3000 ;
	    RECT 10.0000 267.7000 14.0000 268.2000 ;
	    RECT 10.0000 267.6000 11.6000 267.7000 ;
	    RECT 12.4000 267.6000 14.0000 267.7000 ;
	    RECT 15.4000 267.6000 18.0000 268.4000 ;
	    RECT 3.0000 266.8000 5.2000 267.4000 ;
	    RECT 4.4000 262.2000 5.2000 266.8000 ;
	    RECT 6.2000 266.2000 6.8000 267.6000 ;
	    RECT 10.0000 267.2000 10.8000 267.6000 ;
	    RECT 13.2000 267.2000 14.0000 267.6000 ;
	    RECT 7.8000 266.2000 11.4000 266.6000 ;
	    RECT 12.6000 266.2000 16.2000 266.6000 ;
	    RECT 17.2000 266.2000 17.8000 267.6000 ;
	    RECT 18.8000 267.2000 19.6000 270.6000 ;
	    RECT 22.2000 270.4000 23.0000 270.6000 ;
	    RECT 25.4000 270.3000 26.0000 271.6000 ;
	    RECT 27.4000 271.8000 28.0000 273.0000 ;
	    RECT 28.6000 273.0000 29.4000 273.2000 ;
	    RECT 33.2000 273.0000 34.0000 273.2000 ;
	    RECT 28.6000 272.4000 34.0000 273.0000 ;
	    RECT 27.4000 271.4000 32.2000 271.8000 ;
	    RECT 36.4000 271.4000 37.2000 279.8000 ;
	    RECT 38.8000 273.6000 39.6000 274.4000 ;
	    RECT 38.8000 272.4000 39.4000 273.6000 ;
	    RECT 40.2000 272.4000 41.0000 279.8000 ;
	    RECT 46.6000 276.4000 47.4000 279.8000 ;
	    RECT 46.6000 275.6000 48.4000 276.4000 ;
	    RECT 45.2000 273.6000 46.0000 274.4000 ;
	    RECT 45.2000 272.4000 45.8000 273.6000 ;
	    RECT 46.6000 272.4000 47.4000 275.6000 ;
	    RECT 38.0000 271.8000 39.4000 272.4000 ;
	    RECT 40.0000 271.8000 41.0000 272.4000 ;
	    RECT 44.4000 271.8000 45.8000 272.4000 ;
	    RECT 46.4000 271.8000 47.4000 272.4000 ;
	    RECT 53.4000 272.4000 54.2000 279.8000 ;
	    RECT 54.8000 273.6000 55.6000 274.4000 ;
	    RECT 55.0000 272.4000 55.6000 273.6000 ;
	    RECT 58.0000 273.6000 58.8000 274.4000 ;
	    RECT 58.0000 272.4000 58.6000 273.6000 ;
	    RECT 59.4000 272.4000 60.2000 279.8000 ;
	    RECT 64.4000 273.6000 65.2000 274.4000 ;
	    RECT 64.4000 272.4000 65.0000 273.6000 ;
	    RECT 65.8000 272.4000 66.6000 279.8000 ;
	    RECT 70.8000 273.6000 71.6000 274.4000 ;
	    RECT 70.8000 272.4000 71.4000 273.6000 ;
	    RECT 72.2000 272.4000 73.0000 279.8000 ;
	    RECT 78.6000 274.4000 79.4000 279.8000 ;
	    RECT 77.2000 273.6000 78.0000 274.4000 ;
	    RECT 78.6000 273.6000 80.4000 274.4000 ;
	    RECT 83.6000 273.6000 84.4000 274.4000 ;
	    RECT 77.2000 272.4000 77.8000 273.6000 ;
	    RECT 78.6000 272.4000 79.4000 273.6000 ;
	    RECT 83.6000 272.4000 84.2000 273.6000 ;
	    RECT 85.0000 272.4000 85.8000 279.8000 ;
	    RECT 90.0000 273.6000 90.8000 274.4000 ;
	    RECT 90.0000 272.4000 90.6000 273.6000 ;
	    RECT 91.4000 272.4000 92.2000 279.8000 ;
	    RECT 53.4000 271.8000 54.4000 272.4000 ;
	    RECT 55.0000 271.8000 56.4000 272.4000 ;
	    RECT 38.0000 271.6000 38.8000 271.8000 ;
	    RECT 27.4000 271.2000 37.2000 271.4000 ;
	    RECT 31.4000 271.0000 37.2000 271.2000 ;
	    RECT 31.6000 270.8000 37.2000 271.0000 ;
	    RECT 26.8000 270.3000 27.6000 270.4000 ;
	    RECT 20.6000 269.8000 21.4000 270.0000 ;
	    RECT 20.6000 269.2000 24.4000 269.8000 ;
	    RECT 25.3000 269.7000 27.6000 270.3000 ;
	    RECT 23.6000 269.0000 24.4000 269.2000 ;
	    RECT 25.4000 268.4000 26.0000 269.7000 ;
	    RECT 26.8000 269.6000 27.6000 269.7000 ;
	    RECT 30.0000 270.2000 30.8000 270.4000 ;
	    RECT 30.0000 269.6000 35.0000 270.2000 ;
	    RECT 31.6000 269.4000 32.4000 269.6000 ;
	    RECT 34.2000 269.4000 35.0000 269.6000 ;
	    RECT 32.6000 268.4000 33.4000 268.6000 ;
	    RECT 40.0000 268.4000 40.6000 271.8000 ;
	    RECT 44.4000 271.6000 45.2000 271.8000 ;
	    RECT 41.2000 268.8000 42.0000 270.4000 ;
	    RECT 46.4000 268.4000 47.0000 271.8000 ;
	    RECT 53.8000 270.4000 54.4000 271.8000 ;
	    RECT 55.6000 271.6000 56.4000 271.8000 ;
	    RECT 57.2000 271.8000 58.6000 272.4000 ;
	    RECT 59.2000 271.8000 60.2000 272.4000 ;
	    RECT 63.6000 271.8000 65.0000 272.4000 ;
	    RECT 65.6000 271.8000 66.6000 272.4000 ;
	    RECT 70.0000 271.8000 71.4000 272.4000 ;
	    RECT 72.0000 271.8000 73.0000 272.4000 ;
	    RECT 76.4000 271.8000 77.8000 272.4000 ;
	    RECT 78.4000 271.8000 79.4000 272.4000 ;
	    RECT 82.8000 271.8000 84.2000 272.4000 ;
	    RECT 84.8000 271.8000 85.8000 272.4000 ;
	    RECT 89.2000 271.8000 90.6000 272.4000 ;
	    RECT 91.2000 271.8000 92.2000 272.4000 ;
	    RECT 57.2000 271.6000 58.0000 271.8000 ;
	    RECT 59.2000 270.4000 59.8000 271.8000 ;
	    RECT 63.6000 271.6000 64.4000 271.8000 ;
	    RECT 65.6000 270.4000 66.2000 271.8000 ;
	    RECT 70.0000 271.6000 70.8000 271.8000 ;
	    RECT 72.0000 270.4000 72.6000 271.8000 ;
	    RECT 76.4000 271.6000 77.2000 271.8000 ;
	    RECT 47.6000 270.3000 48.4000 270.4000 ;
	    RECT 52.4000 270.3000 53.2000 270.4000 ;
	    RECT 47.6000 269.7000 53.2000 270.3000 ;
	    RECT 47.6000 268.8000 48.4000 269.7000 ;
	    RECT 52.4000 268.8000 53.2000 269.7000 ;
	    RECT 53.8000 269.6000 54.8000 270.4000 ;
	    RECT 58.8000 269.6000 59.8000 270.4000 ;
	    RECT 53.8000 268.4000 54.4000 269.6000 ;
	    RECT 59.2000 268.4000 59.8000 269.6000 ;
	    RECT 60.4000 268.8000 61.2000 270.4000 ;
	    RECT 65.2000 269.6000 66.2000 270.4000 ;
	    RECT 65.6000 268.4000 66.2000 269.6000 ;
	    RECT 66.8000 268.8000 67.6000 270.4000 ;
	    RECT 71.6000 269.6000 72.6000 270.4000 ;
	    RECT 72.0000 268.4000 72.6000 269.6000 ;
	    RECT 73.2000 268.8000 74.0000 270.4000 ;
	    RECT 78.4000 268.4000 79.0000 271.8000 ;
	    RECT 82.8000 271.6000 83.6000 271.8000 ;
	    RECT 79.6000 270.3000 80.4000 270.4000 ;
	    RECT 82.8000 270.3000 83.6000 270.4000 ;
	    RECT 79.6000 269.7000 83.6000 270.3000 ;
	    RECT 79.6000 268.8000 80.4000 269.7000 ;
	    RECT 82.8000 269.6000 83.6000 269.7000 ;
	    RECT 84.8000 268.4000 85.4000 271.8000 ;
	    RECT 89.2000 271.6000 90.0000 271.8000 ;
	    RECT 86.0000 268.8000 86.8000 270.4000 ;
	    RECT 87.6000 270.3000 88.4000 270.4000 ;
	    RECT 91.2000 270.3000 91.8000 271.8000 ;
	    RECT 95.6000 271.4000 96.4000 279.8000 ;
	    RECT 100.0000 276.4000 100.8000 279.8000 ;
	    RECT 98.8000 275.8000 100.8000 276.4000 ;
	    RECT 104.4000 275.8000 105.2000 279.8000 ;
	    RECT 108.6000 275.8000 109.8000 279.8000 ;
	    RECT 98.8000 275.0000 99.6000 275.8000 ;
	    RECT 104.4000 275.2000 105.0000 275.8000 ;
	    RECT 102.2000 274.6000 105.8000 275.2000 ;
	    RECT 108.4000 275.0000 109.2000 275.8000 ;
	    RECT 102.2000 274.4000 103.0000 274.6000 ;
	    RECT 105.0000 274.4000 105.8000 274.6000 ;
	    RECT 98.8000 273.0000 99.6000 273.2000 ;
	    RECT 103.4000 273.0000 104.2000 273.2000 ;
	    RECT 98.8000 272.4000 104.2000 273.0000 ;
	    RECT 104.8000 273.0000 107.0000 273.6000 ;
	    RECT 104.8000 271.8000 105.4000 273.0000 ;
	    RECT 106.2000 272.8000 107.0000 273.0000 ;
	    RECT 108.6000 273.2000 110.0000 274.0000 ;
	    RECT 108.6000 272.2000 109.2000 273.2000 ;
	    RECT 100.6000 271.4000 105.4000 271.8000 ;
	    RECT 95.6000 271.2000 105.4000 271.4000 ;
	    RECT 106.8000 271.6000 109.2000 272.2000 ;
	    RECT 95.6000 271.0000 101.4000 271.2000 ;
	    RECT 95.6000 270.8000 101.2000 271.0000 ;
	    RECT 87.6000 269.7000 91.8000 270.3000 ;
	    RECT 87.6000 269.6000 88.4000 269.7000 ;
	    RECT 91.2000 268.4000 91.8000 269.7000 ;
	    RECT 92.4000 268.8000 93.2000 270.4000 ;
	    RECT 102.0000 270.2000 102.8000 270.4000 ;
	    RECT 97.8000 269.6000 102.8000 270.2000 ;
	    RECT 97.8000 269.4000 98.6000 269.6000 ;
	    RECT 100.4000 269.4000 101.2000 269.6000 ;
	    RECT 99.4000 268.4000 100.2000 268.6000 ;
	    RECT 106.8000 268.4000 107.4000 271.6000 ;
	    RECT 113.2000 271.2000 114.0000 279.8000 ;
	    RECT 123.8000 272.4000 124.6000 279.8000 ;
	    RECT 130.2000 278.4000 132.2000 279.8000 ;
	    RECT 129.2000 277.6000 132.2000 278.4000 ;
	    RECT 125.2000 273.6000 126.0000 274.4000 ;
	    RECT 125.4000 272.4000 126.0000 273.6000 ;
	    RECT 123.8000 271.8000 124.8000 272.4000 ;
	    RECT 125.4000 271.8000 126.8000 272.4000 ;
	    RECT 130.2000 271.8000 132.2000 277.6000 ;
	    RECT 138.2000 272.6000 139.0000 279.8000 ;
	    RECT 143.0000 272.6000 143.8000 279.8000 ;
	    RECT 147.8000 272.6000 148.6000 279.8000 ;
	    RECT 137.2000 271.8000 139.0000 272.6000 ;
	    RECT 142.0000 271.8000 143.8000 272.6000 ;
	    RECT 146.8000 271.8000 148.6000 272.6000 ;
	    RECT 150.0000 271.8000 150.8000 279.8000 ;
	    RECT 153.2000 272.4000 154.0000 279.8000 ;
	    RECT 151.8000 271.8000 154.0000 272.4000 ;
	    RECT 109.8000 270.6000 114.0000 271.2000 ;
	    RECT 109.8000 270.4000 110.6000 270.6000 ;
	    RECT 113.2000 270.3000 114.0000 270.6000 ;
	    RECT 122.8000 270.3000 123.6000 270.4000 ;
	    RECT 111.4000 269.8000 112.2000 270.0000 ;
	    RECT 108.4000 269.2000 112.2000 269.8000 ;
	    RECT 113.2000 269.7000 123.6000 270.3000 ;
	    RECT 108.4000 269.0000 109.2000 269.2000 ;
	    RECT 25.4000 267.8000 36.4000 268.4000 ;
	    RECT 25.8000 267.6000 26.6000 267.8000 ;
	    RECT 18.8000 266.6000 22.6000 267.2000 ;
	    RECT 6.0000 262.2000 6.8000 266.2000 ;
	    RECT 7.6000 266.0000 11.6000 266.2000 ;
	    RECT 7.6000 262.2000 8.4000 266.0000 ;
	    RECT 10.8000 262.2000 11.6000 266.0000 ;
	    RECT 12.4000 266.0000 16.4000 266.2000 ;
	    RECT 12.4000 262.2000 13.2000 266.0000 ;
	    RECT 15.6000 262.2000 16.4000 266.0000 ;
	    RECT 17.2000 262.2000 18.0000 266.2000 ;
	    RECT 18.8000 262.2000 19.6000 266.6000 ;
	    RECT 21.8000 266.4000 22.6000 266.6000 ;
	    RECT 31.6000 265.6000 32.2000 267.8000 ;
	    RECT 34.8000 267.6000 36.4000 267.8000 ;
	    RECT 38.0000 267.6000 40.6000 268.4000 ;
	    RECT 42.8000 268.2000 43.6000 268.4000 ;
	    RECT 42.0000 267.6000 43.6000 268.2000 ;
	    RECT 44.4000 267.6000 47.0000 268.4000 ;
	    RECT 49.2000 268.3000 50.0000 268.4000 ;
	    RECT 50.8000 268.3000 51.6000 268.4000 ;
	    RECT 49.2000 268.2000 51.6000 268.3000 ;
	    RECT 48.4000 267.7000 52.4000 268.2000 ;
	    RECT 48.4000 267.6000 50.0000 267.7000 ;
	    RECT 50.8000 267.6000 52.4000 267.7000 ;
	    RECT 53.8000 267.6000 56.4000 268.4000 ;
	    RECT 57.2000 267.6000 59.8000 268.4000 ;
	    RECT 62.0000 268.2000 62.8000 268.4000 ;
	    RECT 61.2000 267.6000 62.8000 268.2000 ;
	    RECT 63.6000 267.6000 66.2000 268.4000 ;
	    RECT 68.4000 268.2000 69.2000 268.4000 ;
	    RECT 67.6000 267.6000 69.2000 268.2000 ;
	    RECT 70.0000 267.6000 72.6000 268.4000 ;
	    RECT 74.8000 268.2000 75.6000 268.4000 ;
	    RECT 74.0000 267.6000 75.6000 268.2000 ;
	    RECT 76.4000 267.6000 79.0000 268.4000 ;
	    RECT 81.2000 268.2000 82.0000 268.4000 ;
	    RECT 80.4000 267.6000 82.0000 268.2000 ;
	    RECT 82.8000 267.6000 85.4000 268.4000 ;
	    RECT 87.6000 268.2000 88.4000 268.4000 ;
	    RECT 86.8000 267.6000 88.4000 268.2000 ;
	    RECT 89.2000 267.6000 91.8000 268.4000 ;
	    RECT 94.0000 268.2000 94.8000 268.4000 ;
	    RECT 93.2000 267.6000 94.8000 268.2000 ;
	    RECT 96.4000 267.8000 107.4000 268.4000 ;
	    RECT 96.4000 267.6000 98.0000 267.8000 ;
	    RECT 29.8000 265.4000 30.6000 265.6000 ;
	    RECT 23.6000 264.2000 24.4000 265.0000 ;
	    RECT 27.8000 264.8000 30.6000 265.4000 ;
	    RECT 31.6000 264.8000 32.4000 265.6000 ;
	    RECT 27.8000 264.2000 28.4000 264.8000 ;
	    RECT 33.2000 264.2000 34.0000 265.0000 ;
	    RECT 23.0000 263.6000 24.4000 264.2000 ;
	    RECT 23.0000 262.2000 24.2000 263.6000 ;
	    RECT 27.6000 262.2000 28.4000 264.2000 ;
	    RECT 32.0000 263.6000 34.0000 264.2000 ;
	    RECT 32.0000 262.2000 32.8000 263.6000 ;
	    RECT 36.4000 262.2000 37.2000 267.0000 ;
	    RECT 38.2000 266.2000 38.8000 267.6000 ;
	    RECT 42.0000 267.2000 42.8000 267.6000 ;
	    RECT 39.8000 266.2000 43.4000 266.6000 ;
	    RECT 44.6000 266.2000 45.2000 267.6000 ;
	    RECT 48.4000 267.2000 49.2000 267.6000 ;
	    RECT 51.6000 267.2000 52.4000 267.6000 ;
	    RECT 46.2000 266.2000 49.8000 266.6000 ;
	    RECT 51.0000 266.2000 54.6000 266.6000 ;
	    RECT 55.6000 266.2000 56.2000 267.6000 ;
	    RECT 57.4000 266.2000 58.0000 267.6000 ;
	    RECT 61.2000 267.2000 62.0000 267.6000 ;
	    RECT 59.0000 266.2000 62.6000 266.6000 ;
	    RECT 63.8000 266.2000 64.4000 267.6000 ;
	    RECT 67.6000 267.2000 68.4000 267.6000 ;
	    RECT 65.4000 266.2000 69.0000 266.6000 ;
	    RECT 70.2000 266.2000 70.8000 267.6000 ;
	    RECT 74.0000 267.2000 74.8000 267.6000 ;
	    RECT 71.8000 266.2000 75.4000 266.6000 ;
	    RECT 76.6000 266.2000 77.2000 267.6000 ;
	    RECT 80.4000 267.2000 81.2000 267.6000 ;
	    RECT 78.2000 266.2000 81.8000 266.6000 ;
	    RECT 83.0000 266.4000 83.6000 267.6000 ;
	    RECT 86.8000 267.2000 87.6000 267.6000 ;
	    RECT 38.0000 262.2000 38.8000 266.2000 ;
	    RECT 39.6000 266.0000 43.6000 266.2000 ;
	    RECT 39.6000 262.2000 40.4000 266.0000 ;
	    RECT 42.8000 262.2000 43.6000 266.0000 ;
	    RECT 44.4000 262.2000 45.2000 266.2000 ;
	    RECT 46.0000 266.0000 50.0000 266.2000 ;
	    RECT 46.0000 262.2000 46.8000 266.0000 ;
	    RECT 49.2000 262.2000 50.0000 266.0000 ;
	    RECT 50.8000 266.0000 54.8000 266.2000 ;
	    RECT 50.8000 262.2000 51.6000 266.0000 ;
	    RECT 54.0000 262.2000 54.8000 266.0000 ;
	    RECT 55.6000 262.2000 56.4000 266.2000 ;
	    RECT 57.2000 262.2000 58.0000 266.2000 ;
	    RECT 58.8000 266.0000 62.8000 266.2000 ;
	    RECT 58.8000 262.2000 59.6000 266.0000 ;
	    RECT 62.0000 262.2000 62.8000 266.0000 ;
	    RECT 63.6000 262.2000 64.4000 266.2000 ;
	    RECT 65.2000 266.0000 69.2000 266.2000 ;
	    RECT 65.2000 262.2000 66.0000 266.0000 ;
	    RECT 68.4000 262.2000 69.2000 266.0000 ;
	    RECT 70.0000 262.2000 70.8000 266.2000 ;
	    RECT 71.6000 266.0000 75.6000 266.2000 ;
	    RECT 71.6000 262.2000 72.4000 266.0000 ;
	    RECT 74.8000 262.2000 75.6000 266.0000 ;
	    RECT 76.4000 262.2000 77.2000 266.2000 ;
	    RECT 78.0000 266.0000 82.0000 266.2000 ;
	    RECT 78.0000 262.2000 78.8000 266.0000 ;
	    RECT 81.2000 262.2000 82.0000 266.0000 ;
	    RECT 82.8000 262.2000 83.6000 266.4000 ;
	    RECT 84.6000 266.2000 88.2000 266.6000 ;
	    RECT 89.4000 266.2000 90.0000 267.6000 ;
	    RECT 93.2000 267.2000 94.0000 267.6000 ;
	    RECT 91.0000 266.2000 94.6000 266.6000 ;
	    RECT 84.4000 266.0000 88.4000 266.2000 ;
	    RECT 84.4000 262.2000 85.2000 266.0000 ;
	    RECT 87.6000 262.2000 88.4000 266.0000 ;
	    RECT 89.2000 262.2000 90.0000 266.2000 ;
	    RECT 90.8000 266.0000 94.8000 266.2000 ;
	    RECT 90.8000 262.2000 91.6000 266.0000 ;
	    RECT 94.0000 262.2000 94.8000 266.0000 ;
	    RECT 95.6000 262.2000 96.4000 267.0000 ;
	    RECT 100.6000 265.6000 101.2000 267.8000 ;
	    RECT 102.0000 267.6000 102.8000 267.8000 ;
	    RECT 106.2000 267.6000 107.0000 267.8000 ;
	    RECT 113.2000 267.2000 114.0000 269.7000 ;
	    RECT 122.8000 268.8000 123.6000 269.7000 ;
	    RECT 124.2000 268.4000 124.8000 271.8000 ;
	    RECT 126.0000 271.6000 126.8000 271.8000 ;
	    RECT 121.2000 268.2000 122.0000 268.4000 ;
	    RECT 121.2000 267.6000 122.8000 268.2000 ;
	    RECT 124.2000 267.6000 126.8000 268.4000 ;
	    RECT 127.6000 267.6000 128.4000 269.2000 ;
	    RECT 129.2000 268.8000 130.0000 270.4000 ;
	    RECT 131.0000 268.4000 131.6000 271.8000 ;
	    RECT 132.4000 270.3000 133.2000 270.4000 ;
	    RECT 134.0000 270.3000 134.8000 270.4000 ;
	    RECT 132.4000 269.7000 134.8000 270.3000 ;
	    RECT 132.4000 268.8000 133.2000 269.7000 ;
	    RECT 134.0000 269.6000 134.8000 269.7000 ;
	    RECT 137.4000 268.4000 138.0000 271.8000 ;
	    RECT 142.0000 271.6000 142.8000 271.8000 ;
	    RECT 138.8000 269.6000 139.6000 271.2000 ;
	    RECT 142.2000 268.4000 142.8000 271.6000 ;
	    RECT 143.6000 269.6000 144.4000 271.2000 ;
	    RECT 147.0000 270.4000 147.6000 271.8000 ;
	    RECT 146.8000 269.6000 147.6000 270.4000 ;
	    RECT 148.4000 269.6000 149.2000 271.2000 ;
	    RECT 150.0000 269.6000 150.6000 271.8000 ;
	    RECT 151.8000 271.2000 152.4000 271.8000 ;
	    RECT 151.2000 270.4000 152.4000 271.2000 ;
	    RECT 154.8000 271.4000 155.6000 279.8000 ;
	    RECT 159.2000 276.4000 160.0000 279.8000 ;
	    RECT 158.0000 275.8000 160.0000 276.4000 ;
	    RECT 163.6000 275.8000 164.4000 279.8000 ;
	    RECT 167.8000 275.8000 169.0000 279.8000 ;
	    RECT 158.0000 275.0000 158.8000 275.8000 ;
	    RECT 163.6000 275.2000 164.2000 275.8000 ;
	    RECT 161.4000 274.6000 165.0000 275.2000 ;
	    RECT 167.6000 275.0000 168.4000 275.8000 ;
	    RECT 161.4000 274.4000 162.2000 274.6000 ;
	    RECT 164.2000 274.4000 165.0000 274.6000 ;
	    RECT 158.0000 273.0000 158.8000 273.2000 ;
	    RECT 162.6000 273.0000 163.4000 273.2000 ;
	    RECT 158.0000 272.4000 163.4000 273.0000 ;
	    RECT 164.0000 273.0000 166.2000 273.6000 ;
	    RECT 164.0000 271.8000 164.6000 273.0000 ;
	    RECT 165.4000 272.8000 166.2000 273.0000 ;
	    RECT 167.8000 273.2000 169.2000 274.0000 ;
	    RECT 167.8000 272.2000 168.4000 273.2000 ;
	    RECT 159.8000 271.4000 164.6000 271.8000 ;
	    RECT 154.8000 271.2000 164.6000 271.4000 ;
	    RECT 166.0000 271.6000 168.4000 272.2000 ;
	    RECT 154.8000 271.0000 160.6000 271.2000 ;
	    RECT 154.8000 270.8000 160.4000 271.0000 ;
	    RECT 147.0000 268.4000 147.6000 269.6000 ;
	    RECT 130.8000 268.2000 131.6000 268.4000 ;
	    RECT 134.0000 268.2000 134.8000 268.4000 ;
	    RECT 129.2000 267.6000 131.6000 268.2000 ;
	    RECT 133.2000 267.6000 134.8000 268.2000 ;
	    RECT 137.2000 267.6000 138.0000 268.4000 ;
	    RECT 142.0000 267.6000 142.8000 268.4000 ;
	    RECT 146.8000 267.6000 147.6000 268.4000 ;
	    RECT 122.0000 267.2000 122.8000 267.6000 ;
	    RECT 110.2000 266.6000 114.0000 267.2000 ;
	    RECT 110.2000 266.4000 111.0000 266.6000 ;
	    RECT 98.8000 264.2000 99.6000 265.0000 ;
	    RECT 100.4000 264.8000 101.2000 265.6000 ;
	    RECT 102.2000 265.4000 103.0000 265.6000 ;
	    RECT 102.2000 264.8000 105.0000 265.4000 ;
	    RECT 104.4000 264.2000 105.0000 264.8000 ;
	    RECT 108.4000 264.2000 109.2000 265.0000 ;
	    RECT 98.8000 263.6000 100.8000 264.2000 ;
	    RECT 100.0000 262.2000 100.8000 263.6000 ;
	    RECT 104.4000 262.2000 105.2000 264.2000 ;
	    RECT 108.4000 263.6000 109.8000 264.2000 ;
	    RECT 108.6000 262.2000 109.8000 263.6000 ;
	    RECT 113.2000 262.2000 114.0000 266.6000 ;
	    RECT 121.4000 266.2000 125.0000 266.6000 ;
	    RECT 126.0000 266.2000 126.6000 267.6000 ;
	    RECT 129.2000 266.2000 129.8000 267.6000 ;
	    RECT 133.2000 267.2000 134.0000 267.6000 ;
	    RECT 131.0000 266.2000 134.6000 266.6000 ;
	    RECT 121.2000 266.0000 125.2000 266.2000 ;
	    RECT 121.2000 262.2000 122.0000 266.0000 ;
	    RECT 124.4000 262.2000 125.2000 266.0000 ;
	    RECT 126.0000 262.2000 126.8000 266.2000 ;
	    RECT 127.6000 262.8000 128.4000 266.2000 ;
	    RECT 129.2000 263.4000 130.0000 266.2000 ;
	    RECT 130.8000 266.0000 134.8000 266.2000 ;
	    RECT 130.8000 262.8000 131.6000 266.0000 ;
	    RECT 127.6000 262.2000 131.6000 262.8000 ;
	    RECT 134.0000 262.2000 134.8000 266.0000 ;
	    RECT 135.6000 264.8000 136.4000 266.4000 ;
	    RECT 137.4000 264.4000 138.0000 267.6000 ;
	    RECT 140.4000 264.8000 141.2000 266.4000 ;
	    RECT 137.2000 262.2000 138.0000 264.4000 ;
	    RECT 142.2000 264.2000 142.8000 267.6000 ;
	    RECT 145.2000 264.8000 146.0000 266.4000 ;
	    RECT 147.0000 264.2000 147.6000 267.6000 ;
	    RECT 142.0000 262.2000 142.8000 264.2000 ;
	    RECT 146.8000 262.2000 147.6000 264.2000 ;
	    RECT 150.0000 262.2000 150.8000 269.6000 ;
	    RECT 151.8000 267.4000 152.4000 270.4000 ;
	    RECT 161.2000 270.2000 162.0000 270.4000 ;
	    RECT 157.0000 269.6000 162.0000 270.2000 ;
	    RECT 157.0000 269.4000 157.8000 269.6000 ;
	    RECT 158.6000 268.4000 159.4000 268.6000 ;
	    RECT 166.0000 268.4000 166.6000 271.6000 ;
	    RECT 172.4000 271.2000 173.2000 279.8000 ;
	    RECT 174.6000 272.6000 175.4000 279.8000 ;
	    RECT 174.6000 271.8000 176.4000 272.6000 ;
	    RECT 181.4000 272.4000 183.4000 279.8000 ;
	    RECT 187.6000 273.6000 188.4000 274.4000 ;
	    RECT 187.6000 272.4000 188.2000 273.6000 ;
	    RECT 189.0000 272.4000 189.8000 279.8000 ;
	    RECT 195.4000 274.4000 196.2000 279.8000 ;
	    RECT 194.0000 273.6000 194.8000 274.4000 ;
	    RECT 195.4000 273.6000 197.2000 274.4000 ;
	    RECT 194.0000 272.4000 194.6000 273.6000 ;
	    RECT 195.4000 272.4000 196.2000 273.6000 ;
	    RECT 202.2000 272.6000 203.0000 279.8000 ;
	    RECT 207.0000 278.4000 207.8000 279.8000 ;
	    RECT 206.0000 277.6000 207.8000 278.4000 ;
	    RECT 207.0000 272.6000 207.8000 277.6000 ;
	    RECT 180.4000 271.8000 183.4000 272.4000 ;
	    RECT 186.8000 271.8000 188.2000 272.4000 ;
	    RECT 188.8000 271.8000 189.8000 272.4000 ;
	    RECT 193.2000 271.8000 194.6000 272.4000 ;
	    RECT 195.2000 271.8000 196.2000 272.4000 ;
	    RECT 201.2000 271.8000 203.0000 272.6000 ;
	    RECT 206.0000 271.8000 207.8000 272.6000 ;
	    RECT 210.0000 273.6000 210.8000 274.4000 ;
	    RECT 210.0000 272.4000 210.6000 273.6000 ;
	    RECT 211.4000 272.4000 212.2000 279.8000 ;
	    RECT 209.2000 271.8000 210.6000 272.4000 ;
	    RECT 211.2000 271.8000 212.2000 272.4000 ;
	    RECT 218.2000 271.8000 220.2000 279.8000 ;
	    RECT 223.6000 275.0000 224.4000 279.0000 ;
	    RECT 227.8000 278.4000 228.6000 279.8000 ;
	    RECT 226.8000 277.6000 228.6000 278.4000 ;
	    RECT 169.0000 270.6000 173.2000 271.2000 ;
	    RECT 169.0000 270.4000 169.8000 270.6000 ;
	    RECT 170.6000 269.8000 171.4000 270.0000 ;
	    RECT 167.6000 269.2000 171.4000 269.8000 ;
	    RECT 167.6000 269.0000 168.4000 269.2000 ;
	    RECT 155.6000 267.8000 166.6000 268.4000 ;
	    RECT 155.6000 267.6000 157.2000 267.8000 ;
	    RECT 151.8000 266.8000 154.0000 267.4000 ;
	    RECT 153.2000 262.2000 154.0000 266.8000 ;
	    RECT 154.8000 262.2000 155.6000 267.0000 ;
	    RECT 159.8000 265.6000 160.4000 267.8000 ;
	    RECT 165.4000 267.6000 166.2000 267.8000 ;
	    RECT 172.4000 267.2000 173.2000 270.6000 ;
	    RECT 174.0000 269.6000 174.8000 271.2000 ;
	    RECT 175.6000 270.3000 176.2000 271.8000 ;
	    RECT 180.4000 271.6000 182.6000 271.8000 ;
	    RECT 186.8000 271.6000 187.6000 271.8000 ;
	    RECT 180.4000 270.3000 181.2000 270.4000 ;
	    RECT 175.6000 269.7000 181.2000 270.3000 ;
	    RECT 169.4000 266.6000 173.2000 267.2000 ;
	    RECT 169.4000 266.4000 170.2000 266.6000 ;
	    RECT 158.0000 264.2000 158.8000 265.0000 ;
	    RECT 159.6000 264.8000 160.4000 265.6000 ;
	    RECT 161.4000 265.4000 162.2000 265.6000 ;
	    RECT 161.4000 264.8000 164.2000 265.4000 ;
	    RECT 163.6000 264.2000 164.2000 264.8000 ;
	    RECT 167.6000 264.2000 168.4000 265.0000 ;
	    RECT 158.0000 263.6000 160.0000 264.2000 ;
	    RECT 159.2000 262.2000 160.0000 263.6000 ;
	    RECT 163.6000 262.2000 164.4000 264.2000 ;
	    RECT 167.6000 263.6000 169.0000 264.2000 ;
	    RECT 167.8000 262.2000 169.0000 263.6000 ;
	    RECT 172.4000 262.2000 173.2000 266.6000 ;
	    RECT 175.6000 268.4000 176.2000 269.7000 ;
	    RECT 180.4000 268.8000 181.2000 269.7000 ;
	    RECT 182.0000 268.4000 182.6000 271.6000 ;
	    RECT 183.6000 268.8000 184.4000 270.4000 ;
	    RECT 186.9000 270.3000 187.5000 271.6000 ;
	    RECT 185.2000 269.7000 187.5000 270.3000 ;
	    RECT 175.6000 267.6000 176.4000 268.4000 ;
	    RECT 178.8000 268.2000 179.6000 268.4000 ;
	    RECT 182.0000 268.2000 182.8000 268.4000 ;
	    RECT 178.8000 267.6000 180.4000 268.2000 ;
	    RECT 182.0000 267.6000 184.4000 268.2000 ;
	    RECT 185.2000 267.6000 186.0000 269.7000 ;
	    RECT 188.8000 268.4000 189.4000 271.8000 ;
	    RECT 193.2000 271.6000 194.0000 271.8000 ;
	    RECT 190.0000 268.8000 190.8000 270.4000 ;
	    RECT 195.2000 268.4000 195.8000 271.8000 ;
	    RECT 196.4000 268.8000 197.2000 270.4000 ;
	    RECT 201.4000 268.4000 202.0000 271.8000 ;
	    RECT 202.8000 269.6000 203.6000 271.2000 ;
	    RECT 206.2000 268.4000 206.8000 271.8000 ;
	    RECT 209.2000 271.6000 210.0000 271.8000 ;
	    RECT 207.6000 269.6000 208.4000 271.2000 ;
	    RECT 211.2000 268.4000 211.8000 271.8000 ;
	    RECT 212.4000 268.8000 213.2000 270.4000 ;
	    RECT 214.0000 270.3000 214.8000 270.4000 ;
	    RECT 217.2000 270.3000 218.0000 270.4000 ;
	    RECT 214.0000 269.7000 218.0000 270.3000 ;
	    RECT 214.0000 269.6000 214.8000 269.7000 ;
	    RECT 217.2000 268.8000 218.0000 269.7000 ;
	    RECT 218.8000 268.4000 219.4000 271.8000 ;
	    RECT 223.6000 271.6000 224.2000 275.0000 ;
	    RECT 227.8000 272.8000 228.6000 277.6000 ;
	    RECT 233.2000 275.0000 234.0000 279.0000 ;
	    RECT 227.8000 272.2000 229.4000 272.8000 ;
	    RECT 223.6000 271.0000 227.4000 271.6000 ;
	    RECT 220.4000 268.8000 221.2000 270.4000 ;
	    RECT 186.8000 267.6000 189.4000 268.4000 ;
	    RECT 191.6000 268.2000 192.4000 268.4000 ;
	    RECT 190.8000 267.6000 192.4000 268.2000 ;
	    RECT 193.2000 267.6000 195.8000 268.4000 ;
	    RECT 198.0000 268.3000 198.8000 268.4000 ;
	    RECT 199.6000 268.3000 200.4000 268.4000 ;
	    RECT 198.0000 268.2000 200.4000 268.3000 ;
	    RECT 197.2000 267.7000 200.4000 268.2000 ;
	    RECT 197.2000 267.6000 198.8000 267.7000 ;
	    RECT 199.6000 267.6000 200.4000 267.7000 ;
	    RECT 201.2000 268.3000 202.0000 268.4000 ;
	    RECT 204.4000 268.3000 205.2000 268.4000 ;
	    RECT 201.2000 267.7000 205.2000 268.3000 ;
	    RECT 201.2000 267.6000 202.0000 267.7000 ;
	    RECT 204.4000 267.6000 205.2000 267.7000 ;
	    RECT 206.0000 267.6000 206.8000 268.4000 ;
	    RECT 209.2000 267.6000 211.8000 268.4000 ;
	    RECT 214.0000 268.2000 214.8000 268.4000 ;
	    RECT 213.2000 267.6000 214.8000 268.2000 ;
	    RECT 215.6000 268.2000 216.4000 268.4000 ;
	    RECT 218.8000 268.2000 219.6000 268.4000 ;
	    RECT 215.6000 267.6000 217.2000 268.2000 ;
	    RECT 218.8000 267.6000 221.2000 268.2000 ;
	    RECT 222.0000 267.6000 222.8000 269.2000 ;
	    RECT 223.6000 268.8000 224.4000 270.4000 ;
	    RECT 225.2000 268.8000 226.0000 270.4000 ;
	    RECT 226.8000 269.0000 227.4000 271.0000 ;
	    RECT 226.8000 268.2000 228.2000 269.0000 ;
	    RECT 228.8000 268.4000 229.4000 272.2000 ;
	    RECT 233.2000 271.6000 233.8000 275.0000 ;
	    RECT 237.4000 272.8000 238.2000 279.8000 ;
	    RECT 242.8000 275.0000 243.6000 279.0000 ;
	    RECT 247.0000 278.4000 247.8000 279.8000 ;
	    RECT 246.0000 277.6000 247.8000 278.4000 ;
	    RECT 237.4000 272.2000 239.0000 272.8000 ;
	    RECT 238.0000 271.6000 239.0000 272.2000 ;
	    RECT 230.0000 269.6000 230.8000 271.2000 ;
	    RECT 233.2000 271.0000 237.0000 271.6000 ;
	    RECT 233.2000 268.8000 234.0000 270.4000 ;
	    RECT 234.8000 268.8000 235.6000 270.4000 ;
	    RECT 236.4000 269.0000 237.0000 271.0000 ;
	    RECT 226.8000 267.8000 227.8000 268.2000 ;
	    RECT 175.6000 264.2000 176.2000 267.6000 ;
	    RECT 179.6000 267.2000 180.4000 267.6000 ;
	    RECT 177.2000 264.8000 178.0000 266.4000 ;
	    RECT 179.0000 266.2000 182.6000 266.6000 ;
	    RECT 183.8000 266.2000 184.4000 267.6000 ;
	    RECT 187.0000 266.2000 187.6000 267.6000 ;
	    RECT 190.8000 267.2000 191.6000 267.6000 ;
	    RECT 188.6000 266.2000 192.2000 266.6000 ;
	    RECT 193.4000 266.2000 194.0000 267.6000 ;
	    RECT 197.2000 267.2000 198.0000 267.6000 ;
	    RECT 195.0000 266.2000 198.6000 266.6000 ;
	    RECT 178.8000 266.0000 182.8000 266.2000 ;
	    RECT 175.6000 262.2000 176.4000 264.2000 ;
	    RECT 178.8000 262.2000 179.6000 266.0000 ;
	    RECT 182.0000 262.8000 182.8000 266.0000 ;
	    RECT 183.6000 263.4000 184.4000 266.2000 ;
	    RECT 185.2000 262.8000 186.0000 266.2000 ;
	    RECT 182.0000 262.2000 186.0000 262.8000 ;
	    RECT 186.8000 262.2000 187.6000 266.2000 ;
	    RECT 188.4000 266.0000 192.4000 266.2000 ;
	    RECT 188.4000 262.2000 189.2000 266.0000 ;
	    RECT 191.6000 262.2000 192.4000 266.0000 ;
	    RECT 193.2000 262.2000 194.0000 266.2000 ;
	    RECT 194.8000 266.0000 198.8000 266.2000 ;
	    RECT 194.8000 262.2000 195.6000 266.0000 ;
	    RECT 198.0000 262.2000 198.8000 266.0000 ;
	    RECT 199.6000 264.8000 200.4000 266.4000 ;
	    RECT 201.4000 264.2000 202.0000 267.6000 ;
	    RECT 204.4000 264.8000 205.2000 266.4000 ;
	    RECT 206.2000 264.2000 206.8000 267.6000 ;
	    RECT 209.4000 266.2000 210.0000 267.6000 ;
	    RECT 213.2000 267.2000 214.0000 267.6000 ;
	    RECT 216.4000 267.2000 217.2000 267.6000 ;
	    RECT 211.0000 266.2000 214.6000 266.6000 ;
	    RECT 215.8000 266.2000 219.4000 266.6000 ;
	    RECT 220.6000 266.2000 221.2000 267.6000 ;
	    RECT 223.6000 267.2000 227.8000 267.8000 ;
	    RECT 228.8000 267.6000 230.8000 268.4000 ;
	    RECT 236.4000 268.2000 237.8000 269.0000 ;
	    RECT 238.4000 268.4000 239.0000 271.6000 ;
	    RECT 242.8000 271.6000 243.4000 275.0000 ;
	    RECT 247.0000 272.8000 247.8000 277.6000 ;
	    RECT 247.0000 272.2000 248.6000 272.8000 ;
	    RECT 239.6000 269.6000 240.4000 271.2000 ;
	    RECT 242.8000 271.0000 246.6000 271.6000 ;
	    RECT 241.2000 270.3000 242.0000 270.4000 ;
	    RECT 242.8000 270.3000 243.6000 270.4000 ;
	    RECT 241.2000 269.7000 243.6000 270.3000 ;
	    RECT 241.2000 269.6000 242.0000 269.7000 ;
	    RECT 242.8000 268.8000 243.6000 269.7000 ;
	    RECT 244.4000 268.8000 245.2000 270.4000 ;
	    RECT 246.0000 269.0000 246.6000 271.0000 ;
	    RECT 236.4000 267.8000 237.4000 268.2000 ;
	    RECT 201.2000 262.2000 202.0000 264.2000 ;
	    RECT 206.0000 262.2000 206.8000 264.2000 ;
	    RECT 209.2000 262.2000 210.0000 266.2000 ;
	    RECT 210.8000 266.0000 214.8000 266.2000 ;
	    RECT 210.8000 262.2000 211.6000 266.0000 ;
	    RECT 214.0000 262.2000 214.8000 266.0000 ;
	    RECT 215.6000 266.0000 219.6000 266.2000 ;
	    RECT 215.6000 262.2000 216.4000 266.0000 ;
	    RECT 218.8000 262.8000 219.6000 266.0000 ;
	    RECT 220.4000 263.4000 221.2000 266.2000 ;
	    RECT 222.0000 262.8000 222.8000 266.2000 ;
	    RECT 223.6000 265.0000 224.2000 267.2000 ;
	    RECT 228.8000 267.0000 229.4000 267.6000 ;
	    RECT 228.6000 266.6000 229.4000 267.0000 ;
	    RECT 227.8000 266.0000 229.4000 266.6000 ;
	    RECT 233.2000 267.2000 237.4000 267.8000 ;
	    RECT 238.4000 267.6000 240.4000 268.4000 ;
	    RECT 246.0000 268.2000 247.4000 269.0000 ;
	    RECT 248.0000 268.4000 248.6000 272.2000 ;
	    RECT 252.4000 272.4000 253.2000 279.8000 ;
	    RECT 255.6000 278.3000 256.4000 279.8000 ;
	    RECT 257.2000 278.3000 258.0000 278.4000 ;
	    RECT 255.6000 277.7000 258.0000 278.3000 ;
	    RECT 252.4000 271.8000 254.6000 272.4000 ;
	    RECT 255.6000 271.8000 256.4000 277.7000 ;
	    RECT 257.2000 277.6000 258.0000 277.7000 ;
	    RECT 254.0000 271.2000 254.6000 271.8000 ;
	    RECT 249.2000 269.6000 250.0000 271.2000 ;
	    RECT 254.0000 270.4000 255.2000 271.2000 ;
	    RECT 246.0000 267.8000 247.0000 268.2000 ;
	    RECT 223.6000 263.0000 224.4000 265.0000 ;
	    RECT 227.8000 263.0000 228.6000 266.0000 ;
	    RECT 233.2000 265.0000 233.8000 267.2000 ;
	    RECT 238.4000 267.0000 239.0000 267.6000 ;
	    RECT 238.2000 266.6000 239.0000 267.0000 ;
	    RECT 237.4000 266.0000 239.0000 266.6000 ;
	    RECT 242.8000 267.2000 247.0000 267.8000 ;
	    RECT 248.0000 267.6000 250.0000 268.4000 ;
	    RECT 233.2000 263.0000 234.0000 265.0000 ;
	    RECT 237.4000 263.0000 238.2000 266.0000 ;
	    RECT 242.8000 265.0000 243.4000 267.2000 ;
	    RECT 248.0000 267.0000 248.6000 267.6000 ;
	    RECT 254.0000 267.4000 254.6000 270.4000 ;
	    RECT 255.8000 269.6000 256.4000 271.8000 ;
	    RECT 247.8000 266.6000 248.6000 267.0000 ;
	    RECT 247.0000 266.0000 248.6000 266.6000 ;
	    RECT 252.4000 266.8000 254.6000 267.4000 ;
	    RECT 242.8000 263.0000 243.6000 265.0000 ;
	    RECT 247.0000 263.0000 247.8000 266.0000 ;
	    RECT 218.8000 262.2000 222.8000 262.8000 ;
	    RECT 252.4000 262.2000 253.2000 266.8000 ;
	    RECT 255.6000 262.2000 256.4000 269.6000 ;
	    RECT 263.6000 271.2000 264.4000 279.8000 ;
	    RECT 267.8000 275.8000 269.0000 279.8000 ;
	    RECT 272.4000 275.8000 273.2000 279.8000 ;
	    RECT 276.8000 276.4000 277.6000 279.8000 ;
	    RECT 276.8000 275.8000 278.8000 276.4000 ;
	    RECT 268.4000 275.0000 269.2000 275.8000 ;
	    RECT 272.6000 275.2000 273.2000 275.8000 ;
	    RECT 271.8000 274.6000 275.4000 275.2000 ;
	    RECT 278.0000 275.0000 278.8000 275.8000 ;
	    RECT 271.8000 274.4000 272.6000 274.6000 ;
	    RECT 274.6000 274.4000 275.4000 274.6000 ;
	    RECT 267.6000 273.2000 269.0000 274.0000 ;
	    RECT 268.4000 272.2000 269.0000 273.2000 ;
	    RECT 270.6000 273.0000 272.8000 273.6000 ;
	    RECT 270.6000 272.8000 271.4000 273.0000 ;
	    RECT 268.4000 271.6000 270.8000 272.2000 ;
	    RECT 263.6000 270.6000 267.8000 271.2000 ;
	    RECT 263.6000 267.2000 264.4000 270.6000 ;
	    RECT 267.0000 270.4000 267.8000 270.6000 ;
	    RECT 270.2000 270.4000 270.8000 271.6000 ;
	    RECT 272.2000 271.8000 272.8000 273.0000 ;
	    RECT 273.4000 273.0000 274.2000 273.2000 ;
	    RECT 278.0000 273.0000 278.8000 273.2000 ;
	    RECT 273.4000 272.4000 278.8000 273.0000 ;
	    RECT 272.2000 271.4000 277.0000 271.8000 ;
	    RECT 281.2000 271.4000 282.0000 279.8000 ;
	    RECT 272.2000 271.2000 282.0000 271.4000 ;
	    RECT 276.2000 271.0000 282.0000 271.2000 ;
	    RECT 276.4000 270.8000 282.0000 271.0000 ;
	    RECT 265.4000 269.8000 266.2000 270.0000 ;
	    RECT 265.4000 269.2000 269.2000 269.8000 ;
	    RECT 270.0000 269.6000 270.8000 270.4000 ;
	    RECT 274.8000 270.2000 275.6000 270.4000 ;
	    RECT 284.4000 270.3000 285.2000 279.8000 ;
	    RECT 289.8000 274.4000 290.6000 279.8000 ;
	    RECT 296.6000 278.4000 298.6000 279.8000 ;
	    RECT 295.6000 277.6000 298.6000 278.4000 ;
	    RECT 288.4000 273.6000 289.2000 274.4000 ;
	    RECT 289.8000 273.6000 291.6000 274.4000 ;
	    RECT 286.0000 271.6000 286.8000 273.2000 ;
	    RECT 288.4000 272.4000 289.0000 273.6000 ;
	    RECT 289.8000 272.4000 290.6000 273.6000 ;
	    RECT 287.6000 271.8000 289.0000 272.4000 ;
	    RECT 289.6000 271.8000 290.6000 272.4000 ;
	    RECT 296.6000 271.8000 298.6000 277.6000 ;
	    RECT 304.6000 272.4000 305.4000 279.8000 ;
	    RECT 309.0000 278.4000 309.8000 279.8000 ;
	    RECT 309.0000 277.6000 310.8000 278.4000 ;
	    RECT 306.0000 273.6000 306.8000 274.4000 ;
	    RECT 306.2000 272.4000 306.8000 273.6000 ;
	    RECT 309.0000 272.6000 309.8000 277.6000 ;
	    RECT 313.8000 272.6000 314.6000 279.8000 ;
	    RECT 320.6000 274.4000 322.6000 279.8000 ;
	    RECT 319.6000 273.6000 322.6000 274.4000 ;
	    RECT 287.6000 271.6000 288.4000 271.8000 ;
	    RECT 287.7000 270.3000 288.3000 271.6000 ;
	    RECT 274.8000 269.6000 279.8000 270.2000 ;
	    RECT 268.4000 269.0000 269.2000 269.2000 ;
	    RECT 270.2000 268.4000 270.8000 269.6000 ;
	    RECT 276.4000 269.4000 277.2000 269.6000 ;
	    RECT 279.0000 269.4000 279.8000 269.6000 ;
	    RECT 284.4000 269.7000 288.3000 270.3000 ;
	    RECT 277.4000 268.4000 278.2000 268.6000 ;
	    RECT 270.2000 267.8000 281.2000 268.4000 ;
	    RECT 270.6000 267.6000 271.4000 267.8000 ;
	    RECT 263.6000 266.6000 267.4000 267.2000 ;
	    RECT 263.6000 262.2000 264.4000 266.6000 ;
	    RECT 266.6000 266.4000 267.4000 266.6000 ;
	    RECT 276.4000 265.6000 277.0000 267.8000 ;
	    RECT 279.6000 267.6000 281.2000 267.8000 ;
	    RECT 274.6000 265.4000 275.4000 265.6000 ;
	    RECT 268.4000 264.2000 269.2000 265.0000 ;
	    RECT 272.6000 264.8000 275.4000 265.4000 ;
	    RECT 276.4000 264.8000 277.2000 265.6000 ;
	    RECT 272.6000 264.2000 273.2000 264.8000 ;
	    RECT 278.0000 264.2000 278.8000 265.0000 ;
	    RECT 267.8000 263.6000 269.2000 264.2000 ;
	    RECT 267.8000 262.2000 269.0000 263.6000 ;
	    RECT 272.4000 262.2000 273.2000 264.2000 ;
	    RECT 276.8000 263.6000 278.8000 264.2000 ;
	    RECT 276.8000 262.2000 277.6000 263.6000 ;
	    RECT 281.2000 262.2000 282.0000 267.0000 ;
	    RECT 282.8000 266.8000 283.6000 268.4000 ;
	    RECT 284.4000 266.2000 285.2000 269.7000 ;
	    RECT 289.6000 268.4000 290.2000 271.8000 ;
	    RECT 290.8000 268.8000 291.6000 270.4000 ;
	    RECT 287.6000 267.6000 290.2000 268.4000 ;
	    RECT 292.4000 268.2000 293.2000 268.4000 ;
	    RECT 291.6000 267.6000 293.2000 268.2000 ;
	    RECT 294.0000 267.6000 294.8000 269.2000 ;
	    RECT 295.6000 268.8000 296.4000 270.4000 ;
	    RECT 297.4000 268.4000 298.0000 271.8000 ;
	    RECT 303.6000 271.6000 305.6000 272.4000 ;
	    RECT 306.2000 271.8000 307.6000 272.4000 ;
	    RECT 309.0000 271.8000 310.8000 272.6000 ;
	    RECT 313.8000 271.8000 315.6000 272.6000 ;
	    RECT 320.6000 271.8000 322.6000 273.6000 ;
	    RECT 326.8000 273.6000 327.6000 274.4000 ;
	    RECT 326.8000 272.4000 327.4000 273.6000 ;
	    RECT 328.2000 272.4000 329.0000 279.8000 ;
	    RECT 326.0000 271.8000 327.4000 272.4000 ;
	    RECT 328.0000 271.8000 329.0000 272.4000 ;
	    RECT 306.8000 271.6000 307.6000 271.8000 ;
	    RECT 298.8000 268.8000 299.6000 270.4000 ;
	    RECT 302.0000 270.3000 302.8000 270.4000 ;
	    RECT 300.5000 269.7000 302.8000 270.3000 ;
	    RECT 300.5000 268.4000 301.1000 269.7000 ;
	    RECT 302.0000 269.6000 302.8000 269.7000 ;
	    RECT 303.6000 268.8000 304.4000 270.4000 ;
	    RECT 305.0000 268.4000 305.6000 271.6000 ;
	    RECT 308.4000 269.6000 309.2000 271.2000 ;
	    RECT 310.0000 268.4000 310.6000 271.8000 ;
	    RECT 313.2000 269.6000 314.0000 271.2000 ;
	    RECT 314.8000 270.3000 315.4000 271.8000 ;
	    RECT 319.6000 270.3000 320.4000 270.4000 ;
	    RECT 314.8000 269.7000 320.4000 270.3000 ;
	    RECT 314.8000 268.4000 315.4000 269.7000 ;
	    RECT 319.6000 268.8000 320.4000 269.7000 ;
	    RECT 321.2000 268.4000 321.8000 271.8000 ;
	    RECT 326.0000 271.6000 326.8000 271.8000 ;
	    RECT 322.8000 268.8000 323.6000 270.4000 ;
	    RECT 326.1000 270.3000 326.7000 271.6000 ;
	    RECT 324.4000 269.7000 326.7000 270.3000 ;
	    RECT 297.2000 268.2000 298.0000 268.4000 ;
	    RECT 300.4000 268.2000 301.2000 268.4000 ;
	    RECT 295.6000 267.6000 298.0000 268.2000 ;
	    RECT 299.6000 267.6000 301.2000 268.2000 ;
	    RECT 302.0000 268.2000 302.8000 268.4000 ;
	    RECT 302.0000 267.6000 303.6000 268.2000 ;
	    RECT 305.0000 267.6000 307.6000 268.4000 ;
	    RECT 310.0000 267.6000 310.8000 268.4000 ;
	    RECT 314.8000 267.6000 315.6000 268.4000 ;
	    RECT 318.0000 268.2000 318.8000 268.4000 ;
	    RECT 321.2000 268.2000 322.0000 268.4000 ;
	    RECT 318.0000 267.6000 319.6000 268.2000 ;
	    RECT 321.2000 267.6000 323.6000 268.2000 ;
	    RECT 324.4000 267.6000 325.2000 269.7000 ;
	    RECT 328.0000 268.4000 328.6000 271.8000 ;
	    RECT 332.4000 271.2000 333.2000 279.8000 ;
	    RECT 336.6000 275.8000 337.8000 279.8000 ;
	    RECT 341.2000 275.8000 342.0000 279.8000 ;
	    RECT 345.6000 276.4000 346.4000 279.8000 ;
	    RECT 345.6000 275.8000 347.6000 276.4000 ;
	    RECT 337.2000 275.0000 338.0000 275.8000 ;
	    RECT 341.4000 275.2000 342.0000 275.8000 ;
	    RECT 340.6000 274.6000 344.2000 275.2000 ;
	    RECT 346.8000 275.0000 347.6000 275.8000 ;
	    RECT 340.6000 274.4000 341.4000 274.6000 ;
	    RECT 343.4000 274.4000 344.2000 274.6000 ;
	    RECT 336.4000 273.2000 337.8000 274.0000 ;
	    RECT 337.2000 272.2000 337.8000 273.2000 ;
	    RECT 339.4000 273.0000 341.6000 273.6000 ;
	    RECT 339.4000 272.8000 340.2000 273.0000 ;
	    RECT 337.2000 271.6000 339.6000 272.2000 ;
	    RECT 332.4000 270.6000 336.6000 271.2000 ;
	    RECT 329.2000 268.8000 330.0000 270.4000 ;
	    RECT 326.0000 267.6000 328.6000 268.4000 ;
	    RECT 330.8000 268.2000 331.6000 268.4000 ;
	    RECT 330.0000 267.6000 331.6000 268.2000 ;
	    RECT 287.8000 266.2000 288.4000 267.6000 ;
	    RECT 291.6000 267.2000 292.4000 267.6000 ;
	    RECT 289.4000 266.2000 293.0000 266.6000 ;
	    RECT 295.6000 266.2000 296.2000 267.6000 ;
	    RECT 299.6000 267.2000 300.4000 267.6000 ;
	    RECT 302.8000 267.2000 303.6000 267.6000 ;
	    RECT 297.4000 266.2000 301.0000 266.6000 ;
	    RECT 302.2000 266.2000 305.8000 266.6000 ;
	    RECT 306.8000 266.2000 307.4000 267.6000 ;
	    RECT 284.4000 265.6000 286.2000 266.2000 ;
	    RECT 285.4000 262.2000 286.2000 265.6000 ;
	    RECT 287.6000 262.2000 288.4000 266.2000 ;
	    RECT 289.2000 266.0000 293.2000 266.2000 ;
	    RECT 289.2000 262.2000 290.0000 266.0000 ;
	    RECT 292.4000 262.2000 293.2000 266.0000 ;
	    RECT 294.0000 262.8000 294.8000 266.2000 ;
	    RECT 295.6000 263.4000 296.4000 266.2000 ;
	    RECT 297.2000 266.0000 301.2000 266.2000 ;
	    RECT 297.2000 262.8000 298.0000 266.0000 ;
	    RECT 294.0000 262.2000 298.0000 262.8000 ;
	    RECT 300.4000 262.2000 301.2000 266.0000 ;
	    RECT 302.0000 266.0000 306.0000 266.2000 ;
	    RECT 302.0000 262.2000 302.8000 266.0000 ;
	    RECT 305.2000 262.2000 306.0000 266.0000 ;
	    RECT 306.8000 262.2000 307.6000 266.2000 ;
	    RECT 310.0000 264.2000 310.6000 267.6000 ;
	    RECT 311.6000 264.8000 312.4000 266.4000 ;
	    RECT 314.8000 264.2000 315.4000 267.6000 ;
	    RECT 318.8000 267.2000 319.6000 267.6000 ;
	    RECT 316.4000 264.8000 317.2000 266.4000 ;
	    RECT 318.2000 266.2000 321.8000 266.6000 ;
	    RECT 323.0000 266.2000 323.6000 267.6000 ;
	    RECT 326.2000 266.2000 326.8000 267.6000 ;
	    RECT 330.0000 267.2000 330.8000 267.6000 ;
	    RECT 332.4000 267.2000 333.2000 270.6000 ;
	    RECT 335.8000 270.4000 336.6000 270.6000 ;
	    RECT 339.0000 270.4000 339.6000 271.6000 ;
	    RECT 341.0000 271.8000 341.6000 273.0000 ;
	    RECT 342.2000 273.0000 343.0000 273.2000 ;
	    RECT 346.8000 273.0000 347.6000 273.2000 ;
	    RECT 342.2000 272.4000 347.6000 273.0000 ;
	    RECT 341.0000 271.4000 345.8000 271.8000 ;
	    RECT 350.0000 271.4000 350.8000 279.8000 ;
	    RECT 352.4000 273.6000 353.2000 274.4000 ;
	    RECT 352.4000 272.4000 353.0000 273.6000 ;
	    RECT 353.8000 272.4000 354.6000 279.8000 ;
	    RECT 358.8000 273.6000 359.6000 274.4000 ;
	    RECT 358.8000 272.4000 359.4000 273.6000 ;
	    RECT 360.2000 272.4000 361.0000 279.8000 ;
	    RECT 351.6000 271.8000 353.0000 272.4000 ;
	    RECT 353.6000 271.8000 354.6000 272.4000 ;
	    RECT 358.0000 271.8000 359.4000 272.4000 ;
	    RECT 360.0000 271.8000 361.0000 272.4000 ;
	    RECT 351.6000 271.6000 352.4000 271.8000 ;
	    RECT 341.0000 271.2000 350.8000 271.4000 ;
	    RECT 345.0000 271.0000 350.8000 271.2000 ;
	    RECT 345.2000 270.8000 350.8000 271.0000 ;
	    RECT 353.6000 270.4000 354.2000 271.8000 ;
	    RECT 358.0000 271.6000 358.8000 271.8000 ;
	    RECT 360.0000 270.4000 360.6000 271.8000 ;
	    RECT 334.2000 269.8000 335.0000 270.0000 ;
	    RECT 334.2000 269.2000 338.0000 269.8000 ;
	    RECT 338.8000 269.6000 339.6000 270.4000 ;
	    RECT 343.6000 270.2000 344.4000 270.4000 ;
	    RECT 343.6000 269.6000 348.6000 270.2000 ;
	    RECT 353.2000 269.6000 354.2000 270.4000 ;
	    RECT 337.2000 269.0000 338.0000 269.2000 ;
	    RECT 339.0000 268.4000 339.6000 269.6000 ;
	    RECT 345.2000 269.4000 346.0000 269.6000 ;
	    RECT 347.8000 269.4000 348.6000 269.6000 ;
	    RECT 346.2000 268.4000 347.0000 268.6000 ;
	    RECT 353.6000 268.4000 354.2000 269.6000 ;
	    RECT 354.8000 270.3000 355.6000 270.4000 ;
	    RECT 356.4000 270.3000 357.2000 270.4000 ;
	    RECT 354.8000 269.7000 357.2000 270.3000 ;
	    RECT 354.8000 268.8000 355.6000 269.7000 ;
	    RECT 356.4000 269.6000 357.2000 269.7000 ;
	    RECT 359.6000 269.6000 360.6000 270.4000 ;
	    RECT 360.0000 268.4000 360.6000 269.6000 ;
	    RECT 361.2000 268.8000 362.0000 270.4000 ;
	    RECT 366.0000 270.3000 366.8000 279.8000 ;
	    RECT 370.0000 273.6000 370.8000 274.4000 ;
	    RECT 367.6000 271.6000 368.4000 273.2000 ;
	    RECT 370.0000 272.4000 370.6000 273.6000 ;
	    RECT 371.4000 272.4000 372.2000 279.8000 ;
	    RECT 369.2000 271.8000 370.6000 272.4000 ;
	    RECT 371.2000 271.8000 372.2000 272.4000 ;
	    RECT 375.6000 271.8000 376.4000 279.8000 ;
	    RECT 378.8000 272.4000 379.6000 279.8000 ;
	    RECT 381.0000 272.4000 381.8000 279.8000 ;
	    RECT 377.4000 271.8000 379.6000 272.4000 ;
	    RECT 380.4000 271.8000 381.8000 272.4000 ;
	    RECT 369.2000 271.6000 370.0000 271.8000 ;
	    RECT 369.3000 270.3000 369.9000 271.6000 ;
	    RECT 366.0000 269.7000 369.9000 270.3000 ;
	    RECT 339.0000 267.8000 350.0000 268.4000 ;
	    RECT 339.4000 267.6000 340.2000 267.8000 ;
	    RECT 332.4000 266.6000 336.2000 267.2000 ;
	    RECT 327.8000 266.2000 331.4000 266.6000 ;
	    RECT 318.0000 266.0000 322.0000 266.2000 ;
	    RECT 310.0000 262.2000 310.8000 264.2000 ;
	    RECT 314.8000 262.2000 315.6000 264.2000 ;
	    RECT 318.0000 262.2000 318.8000 266.0000 ;
	    RECT 321.2000 262.8000 322.0000 266.0000 ;
	    RECT 322.8000 263.4000 323.6000 266.2000 ;
	    RECT 324.4000 262.8000 325.2000 266.2000 ;
	    RECT 321.2000 262.2000 325.2000 262.8000 ;
	    RECT 326.0000 262.2000 326.8000 266.2000 ;
	    RECT 327.6000 266.0000 331.6000 266.2000 ;
	    RECT 327.6000 262.2000 328.4000 266.0000 ;
	    RECT 330.8000 262.2000 331.6000 266.0000 ;
	    RECT 332.4000 262.2000 333.2000 266.6000 ;
	    RECT 335.4000 266.4000 336.2000 266.6000 ;
	    RECT 345.2000 265.6000 345.8000 267.8000 ;
	    RECT 348.4000 267.6000 350.0000 267.8000 ;
	    RECT 351.6000 267.6000 354.2000 268.4000 ;
	    RECT 356.4000 268.2000 357.2000 268.4000 ;
	    RECT 355.6000 267.6000 357.2000 268.2000 ;
	    RECT 358.0000 267.6000 360.6000 268.4000 ;
	    RECT 362.8000 268.2000 363.6000 268.4000 ;
	    RECT 362.0000 267.6000 363.6000 268.2000 ;
	    RECT 343.4000 265.4000 344.2000 265.6000 ;
	    RECT 337.2000 264.2000 338.0000 265.0000 ;
	    RECT 341.4000 264.8000 344.2000 265.4000 ;
	    RECT 345.2000 264.8000 346.0000 265.6000 ;
	    RECT 341.4000 264.2000 342.0000 264.8000 ;
	    RECT 346.8000 264.2000 347.6000 265.0000 ;
	    RECT 336.6000 263.6000 338.0000 264.2000 ;
	    RECT 336.6000 262.2000 337.8000 263.6000 ;
	    RECT 341.2000 262.2000 342.0000 264.2000 ;
	    RECT 345.6000 263.6000 347.6000 264.2000 ;
	    RECT 345.6000 262.2000 346.4000 263.6000 ;
	    RECT 350.0000 262.2000 350.8000 267.0000 ;
	    RECT 351.8000 266.2000 352.4000 267.6000 ;
	    RECT 355.6000 267.2000 356.4000 267.6000 ;
	    RECT 353.4000 266.2000 357.0000 266.6000 ;
	    RECT 358.2000 266.2000 358.8000 267.6000 ;
	    RECT 362.0000 267.2000 362.8000 267.6000 ;
	    RECT 364.4000 266.8000 365.2000 268.4000 ;
	    RECT 359.8000 266.2000 363.4000 266.6000 ;
	    RECT 366.0000 266.2000 366.8000 269.7000 ;
	    RECT 371.2000 268.4000 371.8000 271.8000 ;
	    RECT 372.4000 268.8000 373.2000 270.4000 ;
	    RECT 375.6000 269.6000 376.2000 271.8000 ;
	    RECT 377.4000 271.2000 378.0000 271.8000 ;
	    RECT 376.8000 270.4000 378.0000 271.2000 ;
	    RECT 380.4000 270.4000 381.0000 271.8000 ;
	    RECT 385.2000 271.2000 386.0000 279.8000 ;
	    RECT 389.4000 272.4000 390.2000 279.8000 ;
	    RECT 395.4000 278.4000 396.2000 279.8000 ;
	    RECT 395.4000 277.6000 397.2000 278.4000 ;
	    RECT 390.8000 273.6000 392.4000 274.4000 ;
	    RECT 394.0000 273.6000 394.8000 274.4000 ;
	    RECT 391.0000 272.4000 391.6000 273.6000 ;
	    RECT 394.0000 272.4000 394.6000 273.6000 ;
	    RECT 395.4000 272.4000 396.2000 277.6000 ;
	    RECT 389.4000 271.8000 390.4000 272.4000 ;
	    RECT 391.0000 271.8000 392.4000 272.4000 ;
	    RECT 382.0000 270.8000 386.0000 271.2000 ;
	    RECT 381.8000 270.6000 386.0000 270.8000 ;
	    RECT 369.2000 267.6000 371.8000 268.4000 ;
	    RECT 374.0000 268.2000 374.8000 268.4000 ;
	    RECT 373.2000 267.6000 374.8000 268.2000 ;
	    RECT 369.4000 266.2000 370.0000 267.6000 ;
	    RECT 373.2000 267.2000 374.0000 267.6000 ;
	    RECT 371.0000 266.2000 374.6000 266.6000 ;
	    RECT 351.6000 262.2000 352.4000 266.2000 ;
	    RECT 353.2000 266.0000 357.2000 266.2000 ;
	    RECT 353.2000 262.2000 354.0000 266.0000 ;
	    RECT 356.4000 262.2000 357.2000 266.0000 ;
	    RECT 358.0000 262.2000 358.8000 266.2000 ;
	    RECT 359.6000 266.0000 363.6000 266.2000 ;
	    RECT 359.6000 262.2000 360.4000 266.0000 ;
	    RECT 362.8000 262.2000 363.6000 266.0000 ;
	    RECT 366.0000 265.6000 367.8000 266.2000 ;
	    RECT 367.0000 262.2000 367.8000 265.6000 ;
	    RECT 369.2000 262.2000 370.0000 266.2000 ;
	    RECT 370.8000 266.0000 374.8000 266.2000 ;
	    RECT 370.8000 262.2000 371.6000 266.0000 ;
	    RECT 374.0000 262.2000 374.8000 266.0000 ;
	    RECT 375.6000 262.2000 376.4000 269.6000 ;
	    RECT 377.4000 267.4000 378.0000 270.4000 ;
	    RECT 378.8000 268.8000 379.6000 270.4000 ;
	    RECT 380.4000 269.6000 381.2000 270.4000 ;
	    RECT 381.8000 270.0000 382.6000 270.6000 ;
	    RECT 377.4000 266.8000 379.6000 267.4000 ;
	    RECT 378.8000 262.2000 379.6000 266.8000 ;
	    RECT 380.4000 266.2000 381.0000 269.6000 ;
	    RECT 381.8000 267.0000 382.4000 270.0000 ;
	    RECT 383.2000 268.4000 384.0000 269.2000 ;
	    RECT 388.4000 268.8000 389.2000 270.4000 ;
	    RECT 389.8000 270.3000 390.4000 271.8000 ;
	    RECT 391.6000 271.6000 392.4000 271.8000 ;
	    RECT 393.2000 271.8000 394.6000 272.4000 ;
	    RECT 395.2000 271.8000 396.2000 272.4000 ;
	    RECT 393.2000 271.6000 394.0000 271.8000 ;
	    RECT 393.3000 270.3000 393.9000 271.6000 ;
	    RECT 389.8000 269.7000 393.9000 270.3000 ;
	    RECT 389.8000 268.4000 390.4000 269.7000 ;
	    RECT 395.2000 268.4000 395.8000 271.8000 ;
	    RECT 396.4000 268.8000 397.2000 270.4000 ;
	    RECT 399.6000 270.3000 400.4000 270.4000 ;
	    RECT 398.1000 269.7000 400.4000 270.3000 ;
	    RECT 398.1000 268.4000 398.7000 269.7000 ;
	    RECT 399.6000 269.6000 400.4000 269.7000 ;
	    RECT 401.2000 270.3000 402.0000 279.8000 ;
	    RECT 411.6000 273.6000 412.4000 274.4000 ;
	    RECT 402.8000 271.6000 403.6000 273.2000 ;
	    RECT 411.6000 272.4000 412.2000 273.6000 ;
	    RECT 413.0000 272.4000 413.8000 279.8000 ;
	    RECT 410.8000 271.8000 412.2000 272.4000 ;
	    RECT 412.8000 271.8000 413.8000 272.4000 ;
	    RECT 410.8000 271.6000 411.6000 271.8000 ;
	    RECT 410.9000 270.3000 411.5000 271.6000 ;
	    RECT 401.2000 269.7000 411.5000 270.3000 ;
	    RECT 383.4000 268.3000 384.4000 268.4000 ;
	    RECT 386.8000 268.3000 387.6000 268.4000 ;
	    RECT 383.4000 268.2000 387.6000 268.3000 ;
	    RECT 383.4000 267.7000 388.4000 268.2000 ;
	    RECT 383.4000 267.6000 384.4000 267.7000 ;
	    RECT 386.8000 267.6000 388.4000 267.7000 ;
	    RECT 389.8000 267.6000 392.4000 268.4000 ;
	    RECT 393.2000 267.6000 395.8000 268.4000 ;
	    RECT 398.0000 268.2000 398.8000 268.4000 ;
	    RECT 397.2000 267.6000 398.8000 268.2000 ;
	    RECT 387.6000 267.2000 388.4000 267.6000 ;
	    RECT 381.8000 266.4000 384.2000 267.0000 ;
	    RECT 380.4000 262.2000 381.2000 266.2000 ;
	    RECT 383.6000 264.2000 384.2000 266.4000 ;
	    RECT 385.2000 264.8000 386.0000 266.4000 ;
	    RECT 387.0000 266.2000 390.6000 266.6000 ;
	    RECT 391.6000 266.2000 392.2000 267.6000 ;
	    RECT 393.4000 266.2000 394.0000 267.6000 ;
	    RECT 397.2000 267.2000 398.0000 267.6000 ;
	    RECT 399.6000 266.8000 400.4000 268.4000 ;
	    RECT 395.0000 266.2000 398.6000 266.6000 ;
	    RECT 401.2000 266.2000 402.0000 269.7000 ;
	    RECT 412.8000 268.4000 413.4000 271.8000 ;
	    RECT 414.0000 268.8000 414.8000 270.4000 ;
	    RECT 410.8000 267.6000 413.4000 268.4000 ;
	    RECT 415.6000 268.2000 416.4000 268.4000 ;
	    RECT 414.8000 267.6000 416.4000 268.2000 ;
	    RECT 411.0000 266.2000 411.6000 267.6000 ;
	    RECT 414.8000 267.2000 415.6000 267.6000 ;
	    RECT 417.2000 266.8000 418.0000 268.4000 ;
	    RECT 412.6000 266.2000 416.2000 266.6000 ;
	    RECT 418.8000 266.2000 419.6000 279.8000 ;
	    RECT 422.8000 273.6000 423.6000 274.4000 ;
	    RECT 420.4000 271.6000 421.2000 273.2000 ;
	    RECT 422.8000 272.4000 423.4000 273.6000 ;
	    RECT 424.2000 272.4000 425.0000 279.8000 ;
	    RECT 429.2000 273.6000 430.0000 274.4000 ;
	    RECT 429.2000 272.4000 429.8000 273.6000 ;
	    RECT 430.6000 272.4000 431.4000 279.8000 ;
	    RECT 422.0000 271.8000 423.4000 272.4000 ;
	    RECT 424.0000 271.8000 425.0000 272.4000 ;
	    RECT 428.4000 271.8000 429.8000 272.4000 ;
	    RECT 430.4000 271.8000 431.4000 272.4000 ;
	    RECT 422.0000 271.6000 422.8000 271.8000 ;
	    RECT 422.0000 270.3000 422.8000 270.4000 ;
	    RECT 424.0000 270.3000 424.6000 271.8000 ;
	    RECT 428.4000 271.6000 429.2000 271.8000 ;
	    RECT 430.4000 270.4000 431.0000 271.8000 ;
	    RECT 436.4000 271.2000 437.2000 279.8000 ;
	    RECT 439.6000 271.2000 440.4000 279.8000 ;
	    RECT 442.8000 271.2000 443.6000 279.8000 ;
	    RECT 446.0000 271.2000 446.8000 279.8000 ;
	    RECT 451.8000 272.4000 452.6000 279.8000 ;
	    RECT 457.2000 275.6000 458.0000 279.8000 ;
	    RECT 460.4000 275.8000 461.2000 279.8000 ;
	    RECT 460.4000 275.6000 461.0000 275.8000 ;
	    RECT 457.4000 275.0000 461.0000 275.6000 ;
	    RECT 453.2000 273.6000 454.0000 274.4000 ;
	    RECT 453.4000 272.4000 454.0000 273.6000 ;
	    RECT 458.8000 272.8000 459.6000 274.4000 ;
	    RECT 460.4000 272.4000 461.0000 275.0000 ;
	    RECT 451.8000 271.8000 452.8000 272.4000 ;
	    RECT 453.4000 271.8000 454.8000 272.4000 ;
	    RECT 434.8000 270.4000 437.2000 271.2000 ;
	    RECT 438.2000 270.4000 440.4000 271.2000 ;
	    RECT 441.4000 270.4000 443.6000 271.2000 ;
	    RECT 445.0000 270.4000 446.8000 271.2000 ;
	    RECT 422.0000 269.7000 424.6000 270.3000 ;
	    RECT 422.0000 269.6000 422.8000 269.7000 ;
	    RECT 424.0000 268.4000 424.6000 269.7000 ;
	    RECT 425.2000 268.8000 426.0000 270.4000 ;
	    RECT 430.0000 269.6000 431.0000 270.4000 ;
	    RECT 430.4000 268.4000 431.0000 269.6000 ;
	    RECT 431.6000 268.8000 432.4000 270.4000 ;
	    RECT 422.0000 267.6000 424.6000 268.4000 ;
	    RECT 426.8000 268.2000 427.6000 268.4000 ;
	    RECT 426.0000 267.6000 427.6000 268.2000 ;
	    RECT 428.4000 267.6000 431.0000 268.4000 ;
	    RECT 433.2000 268.2000 434.0000 268.4000 ;
	    RECT 432.4000 267.6000 434.0000 268.2000 ;
	    RECT 434.8000 267.6000 435.6000 270.4000 ;
	    RECT 438.2000 269.0000 439.0000 270.4000 ;
	    RECT 441.4000 269.0000 442.2000 270.4000 ;
	    RECT 445.0000 269.0000 445.8000 270.4000 ;
	    RECT 436.4000 268.2000 439.0000 269.0000 ;
	    RECT 439.8000 268.2000 442.2000 269.0000 ;
	    RECT 443.2000 268.2000 445.8000 269.0000 ;
	    RECT 450.8000 268.8000 451.6000 270.4000 ;
	    RECT 452.2000 268.4000 452.8000 271.8000 ;
	    RECT 454.0000 271.6000 454.8000 271.8000 ;
	    RECT 460.4000 271.6000 461.2000 272.4000 ;
	    RECT 462.0000 271.8000 462.8000 279.8000 ;
	    RECT 465.2000 272.4000 466.0000 279.8000 ;
	    RECT 463.8000 271.8000 466.0000 272.4000 ;
	    RECT 466.8000 272.4000 467.6000 279.8000 ;
	    RECT 466.8000 271.8000 469.0000 272.4000 ;
	    RECT 470.0000 271.8000 470.8000 279.8000 ;
	    RECT 457.2000 269.6000 458.8000 270.4000 ;
	    RECT 460.4000 268.4000 461.0000 271.6000 ;
	    RECT 438.2000 267.6000 439.0000 268.2000 ;
	    RECT 441.4000 267.6000 442.2000 268.2000 ;
	    RECT 445.0000 267.6000 445.8000 268.2000 ;
	    RECT 449.2000 268.2000 450.0000 268.4000 ;
	    RECT 449.2000 267.6000 450.8000 268.2000 ;
	    RECT 452.2000 267.6000 454.8000 268.4000 ;
	    RECT 459.4000 268.2000 461.0000 268.4000 ;
	    RECT 459.2000 267.8000 461.0000 268.2000 ;
	    RECT 462.0000 269.6000 462.6000 271.8000 ;
	    RECT 463.8000 271.2000 464.4000 271.8000 ;
	    RECT 463.2000 270.4000 464.4000 271.2000 ;
	    RECT 468.4000 271.2000 469.0000 271.8000 ;
	    RECT 468.4000 270.4000 469.6000 271.2000 ;
	    RECT 422.2000 266.2000 422.8000 267.6000 ;
	    RECT 426.0000 267.2000 426.8000 267.6000 ;
	    RECT 423.8000 266.2000 427.4000 266.6000 ;
	    RECT 428.6000 266.2000 429.2000 267.6000 ;
	    RECT 432.4000 267.2000 433.2000 267.6000 ;
	    RECT 434.8000 266.8000 437.2000 267.6000 ;
	    RECT 438.2000 266.8000 440.4000 267.6000 ;
	    RECT 441.4000 266.8000 443.6000 267.6000 ;
	    RECT 445.0000 266.8000 446.8000 267.6000 ;
	    RECT 450.0000 267.2000 450.8000 267.6000 ;
	    RECT 430.2000 266.2000 433.8000 266.6000 ;
	    RECT 386.8000 266.0000 390.8000 266.2000 ;
	    RECT 383.6000 262.2000 384.4000 264.2000 ;
	    RECT 386.8000 262.2000 387.6000 266.0000 ;
	    RECT 390.0000 262.2000 390.8000 266.0000 ;
	    RECT 391.6000 262.2000 392.4000 266.2000 ;
	    RECT 393.2000 262.2000 394.0000 266.2000 ;
	    RECT 394.8000 266.0000 398.8000 266.2000 ;
	    RECT 394.8000 262.2000 395.6000 266.0000 ;
	    RECT 398.0000 262.2000 398.8000 266.0000 ;
	    RECT 401.2000 265.6000 403.0000 266.2000 ;
	    RECT 402.2000 262.2000 403.0000 265.6000 ;
	    RECT 404.4000 264.3000 405.2000 264.4000 ;
	    RECT 410.8000 264.3000 411.6000 266.2000 ;
	    RECT 404.4000 263.7000 411.6000 264.3000 ;
	    RECT 404.4000 263.6000 405.2000 263.7000 ;
	    RECT 410.8000 262.2000 411.6000 263.7000 ;
	    RECT 412.4000 266.0000 416.4000 266.2000 ;
	    RECT 412.4000 262.2000 413.2000 266.0000 ;
	    RECT 415.6000 262.2000 416.4000 266.0000 ;
	    RECT 418.8000 265.6000 420.6000 266.2000 ;
	    RECT 419.8000 264.4000 420.6000 265.6000 ;
	    RECT 418.8000 263.6000 420.6000 264.4000 ;
	    RECT 419.8000 262.2000 420.6000 263.6000 ;
	    RECT 422.0000 262.2000 422.8000 266.2000 ;
	    RECT 423.6000 266.0000 427.6000 266.2000 ;
	    RECT 423.6000 262.2000 424.4000 266.0000 ;
	    RECT 426.8000 262.2000 427.6000 266.0000 ;
	    RECT 428.4000 262.2000 429.2000 266.2000 ;
	    RECT 430.0000 266.0000 434.0000 266.2000 ;
	    RECT 430.0000 262.2000 430.8000 266.0000 ;
	    RECT 433.2000 262.2000 434.0000 266.0000 ;
	    RECT 436.4000 262.2000 437.2000 266.8000 ;
	    RECT 439.6000 262.2000 440.4000 266.8000 ;
	    RECT 442.8000 262.2000 443.6000 266.8000 ;
	    RECT 446.0000 262.2000 446.8000 266.8000 ;
	    RECT 449.4000 266.2000 453.0000 266.6000 ;
	    RECT 454.0000 266.2000 454.6000 267.6000 ;
	    RECT 449.2000 266.0000 453.2000 266.2000 ;
	    RECT 449.2000 262.2000 450.0000 266.0000 ;
	    RECT 452.4000 262.2000 453.2000 266.0000 ;
	    RECT 454.0000 262.2000 454.8000 266.2000 ;
	    RECT 459.2000 262.2000 460.0000 267.8000 ;
	    RECT 462.0000 262.2000 462.8000 269.6000 ;
	    RECT 463.8000 267.4000 464.4000 270.4000 ;
	    RECT 465.2000 270.3000 466.0000 270.4000 ;
	    RECT 466.8000 270.3000 467.6000 270.4000 ;
	    RECT 465.2000 269.7000 467.6000 270.3000 ;
	    RECT 465.2000 268.8000 466.0000 269.7000 ;
	    RECT 466.8000 268.8000 467.6000 269.7000 ;
	    RECT 468.4000 267.4000 469.0000 270.4000 ;
	    RECT 470.2000 269.6000 470.8000 271.8000 ;
	    RECT 463.8000 266.8000 466.0000 267.4000 ;
	    RECT 465.2000 262.2000 466.0000 266.8000 ;
	    RECT 466.8000 266.8000 469.0000 267.4000 ;
	    RECT 466.8000 262.2000 467.6000 266.8000 ;
	    RECT 470.0000 262.2000 470.8000 269.6000 ;
	    RECT 471.6000 271.2000 472.4000 279.8000 ;
	    RECT 475.8000 275.8000 477.0000 279.8000 ;
	    RECT 480.4000 275.8000 481.2000 279.8000 ;
	    RECT 484.8000 276.4000 485.6000 279.8000 ;
	    RECT 484.8000 275.8000 486.8000 276.4000 ;
	    RECT 476.4000 275.0000 477.2000 275.8000 ;
	    RECT 480.6000 275.2000 481.2000 275.8000 ;
	    RECT 479.8000 274.6000 483.4000 275.2000 ;
	    RECT 486.0000 275.0000 486.8000 275.8000 ;
	    RECT 479.8000 274.4000 480.6000 274.6000 ;
	    RECT 482.6000 274.4000 483.4000 274.6000 ;
	    RECT 475.6000 273.2000 477.0000 274.0000 ;
	    RECT 476.4000 272.2000 477.0000 273.2000 ;
	    RECT 478.6000 273.0000 480.8000 273.6000 ;
	    RECT 478.6000 272.8000 479.4000 273.0000 ;
	    RECT 476.4000 271.6000 478.8000 272.2000 ;
	    RECT 471.6000 270.6000 475.8000 271.2000 ;
	    RECT 471.6000 267.2000 472.4000 270.6000 ;
	    RECT 475.0000 270.4000 475.8000 270.6000 ;
	    RECT 478.2000 270.3000 478.8000 271.6000 ;
	    RECT 480.2000 271.8000 480.8000 273.0000 ;
	    RECT 481.4000 273.0000 482.2000 273.2000 ;
	    RECT 486.0000 273.0000 486.8000 273.2000 ;
	    RECT 481.4000 272.4000 486.8000 273.0000 ;
	    RECT 480.2000 271.4000 485.0000 271.8000 ;
	    RECT 489.2000 271.4000 490.0000 279.8000 ;
	    RECT 480.2000 271.2000 490.0000 271.4000 ;
	    RECT 484.2000 271.0000 490.0000 271.2000 ;
	    RECT 484.4000 270.8000 490.0000 271.0000 ;
	    RECT 479.6000 270.3000 480.4000 270.4000 ;
	    RECT 473.4000 269.8000 474.2000 270.0000 ;
	    RECT 473.4000 269.2000 477.2000 269.8000 ;
	    RECT 478.1000 269.7000 480.4000 270.3000 ;
	    RECT 476.4000 269.0000 477.2000 269.2000 ;
	    RECT 478.2000 268.4000 478.8000 269.7000 ;
	    RECT 479.6000 269.6000 480.4000 269.7000 ;
	    RECT 482.8000 270.2000 483.6000 270.4000 ;
	    RECT 482.8000 269.6000 487.8000 270.2000 ;
	    RECT 484.4000 269.4000 485.2000 269.6000 ;
	    RECT 487.0000 269.4000 487.8000 269.6000 ;
	    RECT 485.4000 268.4000 486.2000 268.6000 ;
	    RECT 478.2000 267.8000 489.2000 268.4000 ;
	    RECT 478.6000 267.6000 479.4000 267.8000 ;
	    RECT 471.6000 266.6000 475.4000 267.2000 ;
	    RECT 471.6000 262.2000 472.4000 266.6000 ;
	    RECT 474.6000 266.4000 475.4000 266.6000 ;
	    RECT 484.4000 265.6000 485.0000 267.8000 ;
	    RECT 487.6000 267.6000 489.2000 267.8000 ;
	    RECT 492.4000 268.3000 493.2000 279.8000 ;
	    RECT 496.6000 272.4000 497.4000 279.8000 ;
	    RECT 498.0000 273.6000 498.8000 274.4000 ;
	    RECT 498.2000 272.4000 498.8000 273.6000 ;
	    RECT 496.6000 271.8000 497.6000 272.4000 ;
	    RECT 498.2000 271.8000 499.6000 272.4000 ;
	    RECT 495.6000 268.8000 496.4000 270.4000 ;
	    RECT 497.0000 268.4000 497.6000 271.8000 ;
	    RECT 498.8000 271.6000 499.6000 271.8000 ;
	    RECT 500.4000 271.8000 501.2000 279.8000 ;
	    RECT 503.6000 272.4000 504.4000 279.8000 ;
	    RECT 502.2000 271.8000 504.4000 272.4000 ;
	    RECT 505.2000 272.4000 506.0000 279.8000 ;
	    RECT 508.4000 278.3000 509.2000 279.8000 ;
	    RECT 510.0000 278.3000 510.8000 278.4000 ;
	    RECT 508.4000 277.7000 510.8000 278.3000 ;
	    RECT 505.2000 271.8000 507.4000 272.4000 ;
	    RECT 508.4000 271.8000 509.2000 277.7000 ;
	    RECT 510.0000 277.6000 510.8000 277.7000 ;
	    RECT 500.4000 269.6000 501.0000 271.8000 ;
	    RECT 502.2000 271.2000 502.8000 271.8000 ;
	    RECT 501.6000 270.4000 502.8000 271.2000 ;
	    RECT 506.8000 271.2000 507.4000 271.8000 ;
	    RECT 506.8000 270.4000 508.0000 271.2000 ;
	    RECT 494.0000 268.3000 494.8000 268.4000 ;
	    RECT 492.4000 268.2000 494.8000 268.3000 ;
	    RECT 492.4000 267.7000 495.6000 268.2000 ;
	    RECT 482.6000 265.4000 483.4000 265.6000 ;
	    RECT 476.4000 264.2000 477.2000 265.0000 ;
	    RECT 480.6000 264.8000 483.4000 265.4000 ;
	    RECT 484.4000 264.8000 485.2000 265.6000 ;
	    RECT 480.6000 264.2000 481.2000 264.8000 ;
	    RECT 486.0000 264.2000 486.8000 265.0000 ;
	    RECT 475.8000 263.6000 477.2000 264.2000 ;
	    RECT 475.8000 262.2000 477.0000 263.6000 ;
	    RECT 480.4000 262.2000 481.2000 264.2000 ;
	    RECT 484.8000 263.6000 486.8000 264.2000 ;
	    RECT 484.8000 262.2000 485.6000 263.6000 ;
	    RECT 489.2000 262.2000 490.0000 267.0000 ;
	    RECT 490.8000 264.8000 491.6000 266.4000 ;
	    RECT 492.4000 262.2000 493.2000 267.7000 ;
	    RECT 494.0000 267.6000 495.6000 267.7000 ;
	    RECT 497.0000 267.6000 499.6000 268.4000 ;
	    RECT 494.8000 267.2000 495.6000 267.6000 ;
	    RECT 494.2000 266.2000 497.8000 266.6000 ;
	    RECT 498.8000 266.2000 499.4000 267.6000 ;
	    RECT 494.0000 266.0000 498.0000 266.2000 ;
	    RECT 494.0000 262.2000 494.8000 266.0000 ;
	    RECT 497.2000 262.2000 498.0000 266.0000 ;
	    RECT 498.8000 262.2000 499.6000 266.2000 ;
	    RECT 500.4000 262.2000 501.2000 269.6000 ;
	    RECT 502.2000 267.4000 502.8000 270.4000 ;
	    RECT 503.6000 270.3000 504.4000 270.4000 ;
	    RECT 505.2000 270.3000 506.0000 270.4000 ;
	    RECT 503.6000 269.7000 506.0000 270.3000 ;
	    RECT 503.6000 268.8000 504.4000 269.7000 ;
	    RECT 505.2000 268.8000 506.0000 269.7000 ;
	    RECT 506.8000 267.4000 507.4000 270.4000 ;
	    RECT 508.6000 269.6000 509.2000 271.8000 ;
	    RECT 502.2000 266.8000 504.4000 267.4000 ;
	    RECT 503.6000 262.2000 504.4000 266.8000 ;
	    RECT 505.2000 266.8000 507.4000 267.4000 ;
	    RECT 505.2000 262.2000 506.0000 266.8000 ;
	    RECT 508.4000 262.2000 509.2000 269.6000 ;
	    RECT 4.4000 255.2000 5.2000 259.8000 ;
	    RECT 9.2000 255.2000 10.0000 259.8000 ;
	    RECT 3.0000 254.6000 5.2000 255.2000 ;
	    RECT 7.8000 254.6000 10.0000 255.2000 ;
	    RECT 10.8000 255.4000 11.6000 259.8000 ;
	    RECT 15.0000 258.4000 16.2000 259.8000 ;
	    RECT 15.0000 257.8000 16.4000 258.4000 ;
	    RECT 19.6000 257.8000 20.4000 259.8000 ;
	    RECT 24.0000 258.4000 24.8000 259.8000 ;
	    RECT 24.0000 257.8000 26.0000 258.4000 ;
	    RECT 15.6000 257.0000 16.4000 257.8000 ;
	    RECT 19.8000 257.2000 20.4000 257.8000 ;
	    RECT 19.8000 256.6000 22.6000 257.2000 ;
	    RECT 21.8000 256.4000 22.6000 256.6000 ;
	    RECT 23.6000 256.4000 24.4000 257.2000 ;
	    RECT 25.2000 257.0000 26.0000 257.8000 ;
	    RECT 13.8000 255.4000 14.6000 255.6000 ;
	    RECT 10.8000 254.8000 14.6000 255.4000 ;
	    RECT 3.0000 251.6000 3.6000 254.6000 ;
	    RECT 4.4000 251.6000 5.2000 253.2000 ;
	    RECT 7.8000 251.6000 8.4000 254.6000 ;
	    RECT 9.2000 252.3000 10.0000 253.2000 ;
	    RECT 10.8000 252.3000 11.6000 254.8000 ;
	    RECT 17.8000 254.2000 18.6000 254.4000 ;
	    RECT 23.6000 254.2000 24.2000 256.4000 ;
	    RECT 28.4000 255.0000 29.2000 259.8000 ;
	    RECT 30.0000 255.8000 30.8000 259.8000 ;
	    RECT 31.6000 256.0000 32.4000 259.8000 ;
	    RECT 34.8000 256.0000 35.6000 259.8000 ;
	    RECT 31.6000 255.8000 35.6000 256.0000 ;
	    RECT 30.2000 254.4000 30.8000 255.8000 ;
	    RECT 31.8000 255.4000 35.4000 255.8000 ;
	    RECT 38.0000 255.2000 38.8000 259.8000 ;
	    RECT 41.2000 255.2000 42.0000 259.8000 ;
	    RECT 44.4000 255.2000 45.2000 259.8000 ;
	    RECT 47.6000 255.2000 48.4000 259.8000 ;
	    RECT 50.8000 255.8000 51.6000 259.8000 ;
	    RECT 52.4000 256.0000 53.2000 259.8000 ;
	    RECT 55.6000 256.0000 56.4000 259.8000 ;
	    RECT 52.4000 255.8000 56.4000 256.0000 ;
	    RECT 57.2000 255.8000 58.0000 259.8000 ;
	    RECT 58.8000 256.0000 59.6000 259.8000 ;
	    RECT 62.0000 256.0000 62.8000 259.8000 ;
	    RECT 65.2000 257.8000 66.0000 259.8000 ;
	    RECT 58.8000 255.8000 62.8000 256.0000 ;
	    RECT 34.0000 254.4000 34.8000 254.8000 ;
	    RECT 36.4000 254.4000 38.8000 255.2000 ;
	    RECT 39.8000 254.4000 42.0000 255.2000 ;
	    RECT 43.0000 254.4000 45.2000 255.2000 ;
	    RECT 46.6000 254.4000 48.4000 255.2000 ;
	    RECT 51.0000 254.4000 51.6000 255.8000 ;
	    RECT 52.6000 255.4000 56.2000 255.8000 ;
	    RECT 54.8000 254.4000 55.6000 254.8000 ;
	    RECT 57.4000 254.4000 58.0000 255.8000 ;
	    RECT 59.0000 255.4000 62.6000 255.8000 ;
	    RECT 63.6000 255.6000 64.4000 257.2000 ;
	    RECT 61.2000 254.4000 62.0000 254.8000 ;
	    RECT 65.4000 254.4000 66.0000 257.8000 ;
	    RECT 68.4000 255.0000 69.2000 259.8000 ;
	    RECT 72.8000 258.4000 73.6000 259.8000 ;
	    RECT 71.6000 257.8000 73.6000 258.4000 ;
	    RECT 77.2000 257.8000 78.0000 259.8000 ;
	    RECT 81.4000 258.4000 82.6000 259.8000 ;
	    RECT 81.2000 257.8000 82.6000 258.4000 ;
	    RECT 71.6000 257.0000 72.4000 257.8000 ;
	    RECT 77.2000 257.2000 77.8000 257.8000 ;
	    RECT 73.2000 255.6000 74.0000 257.2000 ;
	    RECT 75.0000 256.6000 77.8000 257.2000 ;
	    RECT 81.2000 257.0000 82.0000 257.8000 ;
	    RECT 75.0000 256.4000 75.8000 256.6000 ;
	    RECT 26.8000 254.2000 28.4000 254.4000 ;
	    RECT 17.4000 253.6000 28.4000 254.2000 ;
	    RECT 30.0000 253.6000 32.6000 254.4000 ;
	    RECT 34.0000 253.8000 35.6000 254.4000 ;
	    RECT 34.8000 253.6000 35.6000 253.8000 ;
	    RECT 15.6000 252.8000 16.4000 253.0000 ;
	    RECT 9.2000 251.7000 11.6000 252.3000 ;
	    RECT 12.6000 252.2000 16.4000 252.8000 ;
	    RECT 12.6000 252.0000 13.4000 252.2000 ;
	    RECT 9.2000 251.6000 10.0000 251.7000 ;
	    RECT 2.4000 250.8000 3.6000 251.6000 ;
	    RECT 7.2000 250.8000 8.4000 251.6000 ;
	    RECT 3.0000 250.2000 3.6000 250.8000 ;
	    RECT 7.8000 250.2000 8.4000 250.8000 ;
	    RECT 10.8000 251.4000 11.6000 251.7000 ;
	    RECT 14.2000 251.4000 15.0000 251.6000 ;
	    RECT 10.8000 250.8000 15.0000 251.4000 ;
	    RECT 3.0000 249.6000 5.2000 250.2000 ;
	    RECT 7.8000 249.6000 10.0000 250.2000 ;
	    RECT 4.4000 242.2000 5.2000 249.6000 ;
	    RECT 9.2000 242.2000 10.0000 249.6000 ;
	    RECT 10.8000 242.2000 11.6000 250.8000 ;
	    RECT 17.4000 250.4000 18.0000 253.6000 ;
	    RECT 24.6000 253.4000 25.4000 253.6000 ;
	    RECT 23.6000 252.4000 24.4000 252.6000 ;
	    RECT 26.2000 252.4000 27.0000 252.6000 ;
	    RECT 22.0000 251.8000 27.0000 252.4000 ;
	    RECT 30.0000 252.3000 30.8000 252.4000 ;
	    RECT 32.0000 252.3000 32.6000 253.6000 ;
	    RECT 22.0000 251.6000 22.8000 251.8000 ;
	    RECT 30.0000 251.7000 32.6000 252.3000 ;
	    RECT 30.0000 251.6000 30.8000 251.7000 ;
	    RECT 23.6000 251.0000 29.2000 251.2000 ;
	    RECT 23.4000 250.8000 29.2000 251.0000 ;
	    RECT 15.6000 249.8000 18.0000 250.4000 ;
	    RECT 19.4000 250.6000 29.2000 250.8000 ;
	    RECT 19.4000 250.2000 24.2000 250.6000 ;
	    RECT 15.6000 248.8000 16.2000 249.8000 ;
	    RECT 14.8000 248.0000 16.2000 248.8000 ;
	    RECT 17.8000 249.0000 18.6000 249.2000 ;
	    RECT 19.4000 249.0000 20.0000 250.2000 ;
	    RECT 17.8000 248.4000 20.0000 249.0000 ;
	    RECT 20.6000 249.0000 26.0000 249.6000 ;
	    RECT 20.6000 248.8000 21.4000 249.0000 ;
	    RECT 25.2000 248.8000 26.0000 249.0000 ;
	    RECT 19.0000 247.4000 19.8000 247.6000 ;
	    RECT 21.8000 247.4000 22.6000 247.6000 ;
	    RECT 15.6000 246.2000 16.4000 247.0000 ;
	    RECT 19.0000 246.8000 22.6000 247.4000 ;
	    RECT 19.8000 246.2000 20.4000 246.8000 ;
	    RECT 25.2000 246.2000 26.0000 247.0000 ;
	    RECT 15.0000 242.2000 16.2000 246.2000 ;
	    RECT 19.6000 242.2000 20.4000 246.2000 ;
	    RECT 24.0000 245.6000 26.0000 246.2000 ;
	    RECT 24.0000 242.2000 24.8000 245.6000 ;
	    RECT 28.4000 242.2000 29.2000 250.6000 ;
	    RECT 30.0000 250.2000 30.8000 250.4000 ;
	    RECT 32.0000 250.2000 32.6000 251.7000 ;
	    RECT 33.2000 251.6000 34.0000 253.2000 ;
	    RECT 36.4000 251.6000 37.2000 254.4000 ;
	    RECT 39.8000 253.8000 40.6000 254.4000 ;
	    RECT 43.0000 253.8000 43.8000 254.4000 ;
	    RECT 46.6000 253.8000 47.4000 254.4000 ;
	    RECT 38.0000 253.0000 40.6000 253.8000 ;
	    RECT 41.4000 253.0000 43.8000 253.8000 ;
	    RECT 44.8000 253.0000 47.4000 253.8000 ;
	    RECT 50.8000 253.6000 53.4000 254.4000 ;
	    RECT 54.8000 253.8000 56.4000 254.4000 ;
	    RECT 55.6000 253.6000 56.4000 253.8000 ;
	    RECT 57.2000 253.6000 59.8000 254.4000 ;
	    RECT 61.2000 254.3000 62.8000 254.4000 ;
	    RECT 63.6000 254.3000 64.4000 254.4000 ;
	    RECT 61.2000 253.8000 64.4000 254.3000 ;
	    RECT 62.0000 253.7000 64.4000 253.8000 ;
	    RECT 62.0000 253.6000 62.8000 253.7000 ;
	    RECT 63.6000 253.6000 64.4000 253.7000 ;
	    RECT 65.2000 253.6000 66.0000 254.4000 ;
	    RECT 69.2000 254.2000 70.8000 254.4000 ;
	    RECT 73.4000 254.2000 74.0000 255.6000 ;
	    RECT 83.0000 255.4000 83.8000 255.6000 ;
	    RECT 86.0000 255.4000 86.8000 259.8000 ;
	    RECT 90.2000 256.4000 91.0000 259.8000 ;
	    RECT 83.0000 254.8000 86.8000 255.4000 ;
	    RECT 89.2000 255.8000 91.0000 256.4000 ;
	    RECT 92.4000 255.8000 93.2000 259.8000 ;
	    RECT 94.0000 256.0000 94.8000 259.8000 ;
	    RECT 97.2000 256.0000 98.0000 259.8000 ;
	    RECT 114.8000 259.2000 118.8000 259.8000 ;
	    RECT 94.0000 255.8000 98.0000 256.0000 ;
	    RECT 98.8000 257.0000 99.6000 259.0000 ;
	    RECT 79.0000 254.2000 79.8000 254.4000 ;
	    RECT 69.2000 253.6000 80.2000 254.2000 ;
	    RECT 39.8000 251.6000 40.6000 253.0000 ;
	    RECT 43.0000 251.6000 43.8000 253.0000 ;
	    RECT 46.6000 251.6000 47.4000 253.0000 ;
	    RECT 36.4000 250.8000 38.8000 251.6000 ;
	    RECT 39.8000 250.8000 42.0000 251.6000 ;
	    RECT 43.0000 250.8000 45.2000 251.6000 ;
	    RECT 46.6000 250.8000 48.4000 251.6000 ;
	    RECT 30.0000 249.6000 31.4000 250.2000 ;
	    RECT 32.0000 249.6000 33.0000 250.2000 ;
	    RECT 30.8000 248.4000 31.4000 249.6000 ;
	    RECT 30.8000 247.6000 31.6000 248.4000 ;
	    RECT 32.2000 242.2000 33.0000 249.6000 ;
	    RECT 38.0000 242.2000 38.8000 250.8000 ;
	    RECT 41.2000 242.2000 42.0000 250.8000 ;
	    RECT 44.4000 242.2000 45.2000 250.8000 ;
	    RECT 47.6000 242.2000 48.4000 250.8000 ;
	    RECT 50.8000 250.2000 51.6000 250.4000 ;
	    RECT 52.8000 250.2000 53.4000 253.6000 ;
	    RECT 54.0000 251.6000 54.8000 253.2000 ;
	    RECT 57.2000 250.2000 58.0000 250.4000 ;
	    RECT 59.2000 250.2000 59.8000 253.6000 ;
	    RECT 60.4000 251.6000 61.2000 253.2000 ;
	    RECT 62.0000 252.3000 62.8000 252.4000 ;
	    RECT 65.4000 252.3000 66.0000 253.6000 ;
	    RECT 72.2000 253.4000 73.0000 253.6000 ;
	    RECT 70.6000 252.4000 71.4000 252.6000 ;
	    RECT 62.0000 251.7000 66.0000 252.3000 ;
	    RECT 62.0000 251.6000 62.8000 251.7000 ;
	    RECT 65.4000 250.2000 66.0000 251.7000 ;
	    RECT 66.8000 250.8000 67.6000 252.4000 ;
	    RECT 70.6000 252.3000 75.6000 252.4000 ;
	    RECT 76.4000 252.3000 77.2000 252.4000 ;
	    RECT 70.6000 251.8000 77.2000 252.3000 ;
	    RECT 74.8000 251.7000 77.2000 251.8000 ;
	    RECT 74.8000 251.6000 75.6000 251.7000 ;
	    RECT 76.4000 251.6000 77.2000 251.7000 ;
	    RECT 78.0000 252.3000 78.8000 252.4000 ;
	    RECT 79.6000 252.3000 80.2000 253.6000 ;
	    RECT 81.2000 252.8000 82.0000 253.0000 ;
	    RECT 78.0000 251.7000 80.3000 252.3000 ;
	    RECT 81.2000 252.2000 85.0000 252.8000 ;
	    RECT 84.2000 252.0000 85.0000 252.2000 ;
	    RECT 78.0000 251.6000 78.8000 251.7000 ;
	    RECT 68.4000 251.0000 74.0000 251.2000 ;
	    RECT 68.4000 250.8000 74.2000 251.0000 ;
	    RECT 68.4000 250.6000 78.2000 250.8000 ;
	    RECT 50.8000 249.6000 52.2000 250.2000 ;
	    RECT 52.8000 249.6000 53.8000 250.2000 ;
	    RECT 57.2000 249.6000 58.6000 250.2000 ;
	    RECT 59.2000 249.6000 60.2000 250.2000 ;
	    RECT 51.6000 248.4000 52.2000 249.6000 ;
	    RECT 51.6000 247.6000 52.4000 248.4000 ;
	    RECT 53.0000 242.2000 53.8000 249.6000 ;
	    RECT 58.0000 248.4000 58.6000 249.6000 ;
	    RECT 58.0000 247.6000 58.8000 248.4000 ;
	    RECT 59.4000 242.2000 60.2000 249.6000 ;
	    RECT 65.2000 249.4000 67.0000 250.2000 ;
	    RECT 66.2000 242.2000 67.0000 249.4000 ;
	    RECT 68.4000 242.2000 69.2000 250.6000 ;
	    RECT 73.4000 250.2000 78.2000 250.6000 ;
	    RECT 71.6000 249.0000 77.0000 249.6000 ;
	    RECT 71.6000 248.8000 72.4000 249.0000 ;
	    RECT 76.2000 248.8000 77.0000 249.0000 ;
	    RECT 77.6000 249.0000 78.2000 250.2000 ;
	    RECT 79.6000 250.4000 80.2000 251.7000 ;
	    RECT 82.6000 251.4000 83.4000 251.6000 ;
	    RECT 86.0000 251.4000 86.8000 254.8000 ;
	    RECT 87.6000 253.6000 88.4000 255.2000 ;
	    RECT 82.6000 250.8000 86.8000 251.4000 ;
	    RECT 79.6000 249.8000 82.0000 250.4000 ;
	    RECT 79.0000 249.0000 79.8000 249.2000 ;
	    RECT 77.6000 248.4000 79.8000 249.0000 ;
	    RECT 81.4000 248.8000 82.0000 249.8000 ;
	    RECT 81.4000 248.0000 82.8000 248.8000 ;
	    RECT 75.0000 247.4000 75.8000 247.6000 ;
	    RECT 77.8000 247.4000 78.6000 247.6000 ;
	    RECT 71.6000 246.2000 72.4000 247.0000 ;
	    RECT 75.0000 246.8000 78.6000 247.4000 ;
	    RECT 77.2000 246.2000 77.8000 246.8000 ;
	    RECT 81.2000 246.2000 82.0000 247.0000 ;
	    RECT 71.6000 245.6000 73.6000 246.2000 ;
	    RECT 72.8000 242.2000 73.6000 245.6000 ;
	    RECT 77.2000 242.2000 78.0000 246.2000 ;
	    RECT 81.4000 242.2000 82.6000 246.2000 ;
	    RECT 86.0000 242.2000 86.8000 250.8000 ;
	    RECT 89.2000 252.3000 90.0000 255.8000 ;
	    RECT 92.6000 254.4000 93.2000 255.8000 ;
	    RECT 94.2000 255.4000 97.8000 255.8000 ;
	    RECT 98.8000 254.8000 99.4000 257.0000 ;
	    RECT 103.0000 256.0000 103.8000 259.0000 ;
	    RECT 103.0000 255.4000 104.6000 256.0000 ;
	    RECT 114.8000 255.8000 115.6000 259.2000 ;
	    RECT 116.4000 255.8000 117.2000 258.6000 ;
	    RECT 118.0000 256.0000 118.8000 259.2000 ;
	    RECT 121.2000 256.0000 122.0000 259.8000 ;
	    RECT 118.0000 255.8000 122.0000 256.0000 ;
	    RECT 122.8000 257.0000 123.6000 259.0000 ;
	    RECT 103.8000 255.0000 104.6000 255.4000 ;
	    RECT 96.4000 254.4000 97.2000 254.8000 ;
	    RECT 90.8000 254.3000 91.6000 254.4000 ;
	    RECT 92.4000 254.3000 95.0000 254.4000 ;
	    RECT 90.8000 253.7000 95.0000 254.3000 ;
	    RECT 96.4000 253.8000 98.0000 254.4000 ;
	    RECT 98.8000 254.2000 103.0000 254.8000 ;
	    RECT 90.8000 253.6000 91.6000 253.7000 ;
	    RECT 92.4000 253.6000 95.0000 253.7000 ;
	    RECT 97.2000 253.6000 98.0000 253.8000 ;
	    RECT 102.0000 253.8000 103.0000 254.2000 ;
	    RECT 104.0000 254.4000 104.6000 255.0000 ;
	    RECT 116.4000 254.4000 117.0000 255.8000 ;
	    RECT 118.2000 255.4000 121.8000 255.8000 ;
	    RECT 122.8000 254.8000 123.4000 257.0000 ;
	    RECT 127.0000 256.0000 127.8000 259.0000 ;
	    RECT 134.0000 257.8000 134.8000 259.8000 ;
	    RECT 127.0000 255.4000 128.6000 256.0000 ;
	    RECT 132.4000 255.6000 133.2000 257.2000 ;
	    RECT 127.8000 255.0000 128.6000 255.4000 ;
	    RECT 120.4000 254.4000 121.2000 254.8000 ;
	    RECT 104.0000 254.3000 106.0000 254.4000 ;
	    RECT 113.2000 254.3000 114.0000 254.4000 ;
	    RECT 89.2000 251.7000 93.1000 252.3000 ;
	    RECT 89.2000 242.2000 90.0000 251.7000 ;
	    RECT 92.5000 250.4000 93.1000 251.7000 ;
	    RECT 90.8000 248.8000 91.6000 250.4000 ;
	    RECT 92.4000 250.2000 93.2000 250.4000 ;
	    RECT 94.4000 250.2000 95.0000 253.6000 ;
	    RECT 95.6000 251.6000 96.4000 253.2000 ;
	    RECT 98.8000 251.6000 99.6000 253.2000 ;
	    RECT 100.4000 251.6000 101.2000 253.2000 ;
	    RECT 102.0000 253.0000 103.4000 253.8000 ;
	    RECT 104.0000 253.7000 114.0000 254.3000 ;
	    RECT 104.0000 253.6000 106.0000 253.7000 ;
	    RECT 113.2000 253.6000 114.0000 253.7000 ;
	    RECT 102.0000 251.0000 102.6000 253.0000 ;
	    RECT 98.8000 250.4000 102.6000 251.0000 ;
	    RECT 92.4000 249.6000 93.8000 250.2000 ;
	    RECT 94.4000 249.6000 95.4000 250.2000 ;
	    RECT 93.2000 248.4000 93.8000 249.6000 ;
	    RECT 93.2000 247.6000 94.0000 248.4000 ;
	    RECT 94.6000 242.2000 95.4000 249.6000 ;
	    RECT 98.8000 247.0000 99.4000 250.4000 ;
	    RECT 104.0000 249.8000 104.6000 253.6000 ;
	    RECT 114.8000 252.8000 115.6000 254.4000 ;
	    RECT 116.4000 253.8000 118.8000 254.4000 ;
	    RECT 120.4000 253.8000 122.0000 254.4000 ;
	    RECT 122.8000 254.2000 127.0000 254.8000 ;
	    RECT 118.0000 253.6000 118.8000 253.8000 ;
	    RECT 121.2000 253.6000 122.0000 253.8000 ;
	    RECT 126.0000 253.8000 127.0000 254.2000 ;
	    RECT 128.0000 254.4000 128.6000 255.0000 ;
	    RECT 134.2000 254.4000 134.8000 257.8000 ;
	    RECT 105.2000 252.3000 106.0000 252.4000 ;
	    RECT 113.2000 252.3000 114.0000 252.4000 ;
	    RECT 105.2000 251.7000 114.0000 252.3000 ;
	    RECT 105.2000 250.8000 106.0000 251.7000 ;
	    RECT 113.2000 251.6000 114.0000 251.7000 ;
	    RECT 116.4000 251.6000 117.2000 253.2000 ;
	    RECT 118.2000 250.2000 118.8000 253.6000 ;
	    RECT 119.6000 251.6000 120.4000 253.2000 ;
	    RECT 122.8000 251.6000 123.6000 253.2000 ;
	    RECT 124.4000 251.6000 125.2000 253.2000 ;
	    RECT 126.0000 253.0000 127.4000 253.8000 ;
	    RECT 128.0000 253.6000 130.0000 254.4000 ;
	    RECT 134.0000 253.6000 134.8000 254.4000 ;
	    RECT 126.0000 251.0000 126.6000 253.0000 ;
	    RECT 122.8000 250.4000 126.6000 251.0000 ;
	    RECT 103.0000 249.2000 104.6000 249.8000 ;
	    RECT 98.8000 243.0000 99.6000 247.0000 ;
	    RECT 103.0000 242.2000 103.8000 249.2000 ;
	    RECT 117.4000 248.4000 119.4000 250.2000 ;
	    RECT 116.4000 247.6000 119.4000 248.4000 ;
	    RECT 117.4000 242.2000 119.4000 247.6000 ;
	    RECT 122.8000 247.0000 123.4000 250.4000 ;
	    RECT 128.0000 249.8000 128.6000 253.6000 ;
	    RECT 129.2000 250.8000 130.0000 252.4000 ;
	    RECT 134.2000 250.4000 134.8000 253.6000 ;
	    RECT 138.8000 257.8000 139.6000 259.8000 ;
	    RECT 138.8000 254.4000 139.4000 257.8000 ;
	    RECT 140.4000 255.6000 141.2000 257.2000 ;
	    RECT 142.0000 255.4000 142.8000 259.8000 ;
	    RECT 146.2000 258.4000 147.4000 259.8000 ;
	    RECT 146.2000 257.8000 147.6000 258.4000 ;
	    RECT 150.8000 257.8000 151.6000 259.8000 ;
	    RECT 155.2000 258.4000 156.0000 259.8000 ;
	    RECT 155.2000 257.8000 157.2000 258.4000 ;
	    RECT 146.8000 257.0000 147.6000 257.8000 ;
	    RECT 151.0000 257.2000 151.6000 257.8000 ;
	    RECT 151.0000 256.6000 153.8000 257.2000 ;
	    RECT 153.0000 256.4000 153.8000 256.6000 ;
	    RECT 154.8000 256.4000 155.6000 257.2000 ;
	    RECT 156.4000 257.0000 157.2000 257.8000 ;
	    RECT 145.0000 255.4000 145.8000 255.6000 ;
	    RECT 142.0000 254.8000 145.8000 255.4000 ;
	    RECT 138.8000 253.6000 139.6000 254.4000 ;
	    RECT 135.6000 250.8000 136.4000 252.4000 ;
	    RECT 137.2000 250.8000 138.0000 252.4000 ;
	    RECT 127.0000 249.2000 128.6000 249.8000 ;
	    RECT 134.0000 250.2000 134.8000 250.4000 ;
	    RECT 138.8000 250.2000 139.4000 253.6000 ;
	    RECT 142.0000 251.4000 142.8000 254.8000 ;
	    RECT 149.0000 254.2000 149.8000 254.4000 ;
	    RECT 154.8000 254.2000 155.4000 256.4000 ;
	    RECT 159.6000 255.0000 160.4000 259.8000 ;
	    RECT 161.2000 256.0000 162.0000 259.8000 ;
	    RECT 164.4000 256.0000 165.2000 259.8000 ;
	    RECT 161.2000 255.8000 165.2000 256.0000 ;
	    RECT 166.0000 255.8000 166.8000 259.8000 ;
	    RECT 167.6000 255.8000 168.4000 259.8000 ;
	    RECT 169.2000 256.0000 170.0000 259.8000 ;
	    RECT 172.4000 256.0000 173.2000 259.8000 ;
	    RECT 169.2000 255.8000 173.2000 256.0000 ;
	    RECT 161.4000 255.4000 165.0000 255.8000 ;
	    RECT 162.0000 254.4000 162.8000 254.8000 ;
	    RECT 166.0000 254.4000 166.6000 255.8000 ;
	    RECT 167.8000 254.4000 168.4000 255.8000 ;
	    RECT 169.4000 255.4000 173.0000 255.8000 ;
	    RECT 174.0000 255.2000 174.8000 259.8000 ;
	    RECT 171.6000 254.4000 172.4000 254.8000 ;
	    RECT 174.0000 254.6000 176.2000 255.2000 ;
	    RECT 158.0000 254.2000 159.6000 254.4000 ;
	    RECT 148.6000 253.6000 159.6000 254.2000 ;
	    RECT 161.2000 253.8000 162.8000 254.4000 ;
	    RECT 161.2000 253.6000 162.0000 253.8000 ;
	    RECT 164.2000 253.6000 166.8000 254.4000 ;
	    RECT 167.6000 253.6000 170.2000 254.4000 ;
	    RECT 171.6000 253.8000 173.2000 254.4000 ;
	    RECT 172.4000 253.6000 173.2000 253.8000 ;
	    RECT 146.8000 252.8000 147.6000 253.0000 ;
	    RECT 143.8000 252.2000 147.6000 252.8000 ;
	    RECT 143.8000 252.0000 144.6000 252.2000 ;
	    RECT 145.4000 251.4000 146.2000 251.6000 ;
	    RECT 142.0000 250.8000 146.2000 251.4000 ;
	    RECT 134.0000 249.4000 135.8000 250.2000 ;
	    RECT 122.8000 243.0000 123.6000 247.0000 ;
	    RECT 127.0000 244.4000 127.8000 249.2000 ;
	    RECT 127.0000 243.6000 128.4000 244.4000 ;
	    RECT 127.0000 242.2000 127.8000 243.6000 ;
	    RECT 135.0000 242.2000 135.8000 249.4000 ;
	    RECT 137.8000 249.4000 139.6000 250.2000 ;
	    RECT 137.8000 244.4000 138.6000 249.4000 ;
	    RECT 137.2000 243.6000 138.6000 244.4000 ;
	    RECT 137.8000 242.2000 138.6000 243.6000 ;
	    RECT 142.0000 242.2000 142.8000 250.8000 ;
	    RECT 148.6000 250.4000 149.2000 253.6000 ;
	    RECT 155.8000 253.4000 156.6000 253.6000 ;
	    RECT 154.8000 252.4000 155.6000 252.6000 ;
	    RECT 157.4000 252.4000 158.2000 252.6000 ;
	    RECT 153.2000 251.8000 158.2000 252.4000 ;
	    RECT 153.2000 251.6000 154.0000 251.8000 ;
	    RECT 162.8000 251.6000 163.6000 253.2000 ;
	    RECT 154.8000 251.0000 160.4000 251.2000 ;
	    RECT 154.6000 250.8000 160.4000 251.0000 ;
	    RECT 146.8000 249.8000 149.2000 250.4000 ;
	    RECT 150.6000 250.6000 160.4000 250.8000 ;
	    RECT 150.6000 250.2000 155.4000 250.6000 ;
	    RECT 146.8000 248.8000 147.4000 249.8000 ;
	    RECT 146.0000 248.0000 147.4000 248.8000 ;
	    RECT 149.0000 249.0000 149.8000 249.2000 ;
	    RECT 150.6000 249.0000 151.2000 250.2000 ;
	    RECT 149.0000 248.4000 151.2000 249.0000 ;
	    RECT 151.8000 249.0000 157.2000 249.6000 ;
	    RECT 151.8000 248.8000 152.6000 249.0000 ;
	    RECT 156.4000 248.8000 157.2000 249.0000 ;
	    RECT 150.2000 247.4000 151.0000 247.6000 ;
	    RECT 153.0000 247.4000 153.8000 247.6000 ;
	    RECT 146.8000 246.2000 147.6000 247.0000 ;
	    RECT 150.2000 246.8000 153.8000 247.4000 ;
	    RECT 151.0000 246.2000 151.6000 246.8000 ;
	    RECT 156.4000 246.2000 157.2000 247.0000 ;
	    RECT 146.2000 242.2000 147.4000 246.2000 ;
	    RECT 150.8000 242.2000 151.6000 246.2000 ;
	    RECT 155.2000 245.6000 157.2000 246.2000 ;
	    RECT 155.2000 242.2000 156.0000 245.6000 ;
	    RECT 159.6000 242.2000 160.4000 250.6000 ;
	    RECT 164.2000 250.2000 164.8000 253.6000 ;
	    RECT 169.6000 252.3000 170.2000 253.6000 ;
	    RECT 166.1000 251.7000 170.2000 252.3000 ;
	    RECT 166.1000 250.4000 166.7000 251.7000 ;
	    RECT 166.0000 250.2000 166.8000 250.4000 ;
	    RECT 163.8000 249.6000 164.8000 250.2000 ;
	    RECT 165.4000 249.6000 166.8000 250.2000 ;
	    RECT 167.6000 250.2000 168.4000 250.4000 ;
	    RECT 169.6000 250.2000 170.2000 251.7000 ;
	    RECT 170.8000 251.6000 171.6000 253.2000 ;
	    RECT 175.6000 251.6000 176.2000 254.6000 ;
	    RECT 177.2000 252.4000 178.0000 259.8000 ;
	    RECT 178.8000 255.2000 179.6000 259.8000 ;
	    RECT 178.8000 254.6000 181.0000 255.2000 ;
	    RECT 175.6000 250.8000 176.8000 251.6000 ;
	    RECT 175.6000 250.2000 176.2000 250.8000 ;
	    RECT 177.4000 250.2000 178.0000 252.4000 ;
	    RECT 180.4000 251.6000 181.0000 254.6000 ;
	    RECT 182.0000 252.4000 182.8000 259.8000 ;
	    RECT 180.4000 250.8000 181.6000 251.6000 ;
	    RECT 180.4000 250.2000 181.0000 250.8000 ;
	    RECT 182.2000 250.2000 182.8000 252.4000 ;
	    RECT 167.6000 249.6000 169.0000 250.2000 ;
	    RECT 169.6000 249.6000 170.6000 250.2000 ;
	    RECT 163.8000 242.2000 164.6000 249.6000 ;
	    RECT 165.4000 248.4000 166.0000 249.6000 ;
	    RECT 165.2000 247.6000 166.0000 248.4000 ;
	    RECT 168.4000 248.4000 169.0000 249.6000 ;
	    RECT 168.4000 247.6000 169.2000 248.4000 ;
	    RECT 169.8000 242.2000 170.6000 249.6000 ;
	    RECT 174.0000 249.6000 176.2000 250.2000 ;
	    RECT 174.0000 242.2000 174.8000 249.6000 ;
	    RECT 177.2000 242.2000 178.0000 250.2000 ;
	    RECT 178.8000 249.6000 181.0000 250.2000 ;
	    RECT 178.8000 242.2000 179.6000 249.6000 ;
	    RECT 182.0000 242.2000 182.8000 250.2000 ;
	    RECT 183.6000 252.4000 184.4000 259.8000 ;
	    RECT 186.8000 255.2000 187.6000 259.8000 ;
	    RECT 185.4000 254.6000 187.6000 255.2000 ;
	    RECT 183.6000 250.2000 184.2000 252.4000 ;
	    RECT 185.4000 251.6000 186.0000 254.6000 ;
	    RECT 186.8000 251.6000 187.6000 253.2000 ;
	    RECT 188.4000 252.4000 189.2000 259.8000 ;
	    RECT 191.6000 255.2000 192.4000 259.8000 ;
	    RECT 193.2000 255.8000 194.0000 259.8000 ;
	    RECT 194.8000 256.0000 195.6000 259.8000 ;
	    RECT 198.0000 256.0000 198.8000 259.8000 ;
	    RECT 194.8000 255.8000 198.8000 256.0000 ;
	    RECT 190.2000 254.6000 192.4000 255.2000 ;
	    RECT 184.8000 250.8000 186.0000 251.6000 ;
	    RECT 185.4000 250.2000 186.0000 250.8000 ;
	    RECT 188.4000 250.2000 189.0000 252.4000 ;
	    RECT 190.2000 251.6000 190.8000 254.6000 ;
	    RECT 193.4000 254.4000 194.0000 255.8000 ;
	    RECT 195.0000 255.4000 198.6000 255.8000 ;
	    RECT 199.6000 255.2000 200.4000 259.8000 ;
	    RECT 197.2000 254.4000 198.0000 254.8000 ;
	    RECT 199.6000 254.6000 201.8000 255.2000 ;
	    RECT 193.2000 253.6000 195.8000 254.4000 ;
	    RECT 197.2000 253.8000 198.8000 254.4000 ;
	    RECT 198.0000 253.6000 198.8000 253.8000 ;
	    RECT 189.6000 250.8000 190.8000 251.6000 ;
	    RECT 190.2000 250.2000 190.8000 250.8000 ;
	    RECT 195.2000 250.4000 195.8000 253.6000 ;
	    RECT 196.4000 251.6000 197.2000 253.2000 ;
	    RECT 199.6000 251.6000 200.4000 253.2000 ;
	    RECT 201.2000 251.6000 201.8000 254.6000 ;
	    RECT 202.8000 252.4000 203.6000 259.8000 ;
	    RECT 223.6000 259.2000 227.6000 259.8000 ;
	    RECT 208.2000 256.0000 209.0000 259.0000 ;
	    RECT 212.4000 257.0000 213.2000 259.0000 ;
	    RECT 207.4000 255.4000 209.0000 256.0000 ;
	    RECT 207.4000 255.0000 208.2000 255.4000 ;
	    RECT 207.4000 254.4000 208.0000 255.0000 ;
	    RECT 212.6000 254.8000 213.2000 257.0000 ;
	    RECT 206.0000 253.6000 208.0000 254.4000 ;
	    RECT 209.0000 254.2000 213.2000 254.8000 ;
	    RECT 214.0000 257.0000 214.8000 259.0000 ;
	    RECT 214.0000 254.8000 214.6000 257.0000 ;
	    RECT 218.2000 256.0000 219.0000 259.0000 ;
	    RECT 218.2000 255.4000 219.8000 256.0000 ;
	    RECT 223.6000 255.8000 224.4000 259.2000 ;
	    RECT 225.2000 255.8000 226.0000 258.6000 ;
	    RECT 226.8000 256.0000 227.6000 259.2000 ;
	    RECT 230.0000 256.0000 230.8000 259.8000 ;
	    RECT 226.8000 255.8000 230.8000 256.0000 ;
	    RECT 231.6000 255.8000 232.4000 259.8000 ;
	    RECT 233.2000 256.0000 234.0000 259.8000 ;
	    RECT 236.4000 256.0000 237.2000 259.8000 ;
	    RECT 233.2000 255.8000 237.2000 256.0000 ;
	    RECT 238.0000 256.0000 238.8000 259.8000 ;
	    RECT 241.2000 256.0000 242.0000 259.8000 ;
	    RECT 238.0000 255.8000 242.0000 256.0000 ;
	    RECT 242.8000 255.8000 243.6000 259.8000 ;
	    RECT 244.4000 259.2000 248.4000 259.8000 ;
	    RECT 244.4000 255.8000 245.2000 259.2000 ;
	    RECT 246.0000 255.8000 246.8000 258.6000 ;
	    RECT 247.6000 256.0000 248.4000 259.2000 ;
	    RECT 250.8000 256.0000 251.6000 259.8000 ;
	    RECT 247.6000 255.8000 251.6000 256.0000 ;
	    RECT 254.0000 257.8000 254.8000 259.8000 ;
	    RECT 219.0000 255.0000 219.8000 255.4000 ;
	    RECT 214.0000 254.2000 218.2000 254.8000 ;
	    RECT 209.0000 253.8000 210.0000 254.2000 ;
	    RECT 201.2000 250.8000 202.4000 251.6000 ;
	    RECT 193.2000 250.2000 194.0000 250.4000 ;
	    RECT 183.6000 242.2000 184.4000 250.2000 ;
	    RECT 185.4000 249.6000 187.6000 250.2000 ;
	    RECT 186.8000 242.2000 187.6000 249.6000 ;
	    RECT 188.4000 242.2000 189.2000 250.2000 ;
	    RECT 190.2000 249.6000 192.4000 250.2000 ;
	    RECT 193.2000 249.6000 194.6000 250.2000 ;
	    RECT 195.2000 249.6000 197.2000 250.4000 ;
	    RECT 201.2000 250.2000 201.8000 250.8000 ;
	    RECT 203.0000 250.2000 203.6000 252.4000 ;
	    RECT 206.0000 250.8000 206.8000 252.4000 ;
	    RECT 199.6000 249.6000 201.8000 250.2000 ;
	    RECT 191.6000 242.2000 192.4000 249.6000 ;
	    RECT 194.0000 248.4000 194.6000 249.6000 ;
	    RECT 194.0000 247.6000 194.8000 248.4000 ;
	    RECT 195.4000 242.2000 196.2000 249.6000 ;
	    RECT 199.6000 242.2000 200.4000 249.6000 ;
	    RECT 202.8000 242.2000 203.6000 250.2000 ;
	    RECT 207.4000 249.8000 208.0000 253.6000 ;
	    RECT 208.6000 253.0000 210.0000 253.8000 ;
	    RECT 217.2000 253.8000 218.2000 254.2000 ;
	    RECT 219.2000 254.4000 219.8000 255.0000 ;
	    RECT 225.2000 254.4000 225.8000 255.8000 ;
	    RECT 227.0000 255.4000 230.6000 255.8000 ;
	    RECT 229.2000 254.4000 230.0000 254.8000 ;
	    RECT 231.8000 254.4000 232.4000 255.8000 ;
	    RECT 233.4000 255.4000 237.0000 255.8000 ;
	    RECT 238.2000 255.4000 241.8000 255.8000 ;
	    RECT 235.6000 254.4000 236.4000 254.8000 ;
	    RECT 238.8000 254.4000 239.6000 254.8000 ;
	    RECT 242.8000 254.4000 243.4000 255.8000 ;
	    RECT 246.0000 254.4000 246.6000 255.8000 ;
	    RECT 247.8000 255.4000 251.4000 255.8000 ;
	    RECT 250.0000 254.4000 250.8000 254.8000 ;
	    RECT 254.0000 254.4000 254.6000 257.8000 ;
	    RECT 265.2000 257.6000 266.0000 259.8000 ;
	    RECT 255.6000 256.3000 256.4000 257.2000 ;
	    RECT 263.6000 256.3000 264.4000 256.4000 ;
	    RECT 255.6000 255.7000 264.4000 256.3000 ;
	    RECT 255.6000 255.6000 256.4000 255.7000 ;
	    RECT 263.6000 255.6000 264.4000 255.7000 ;
	    RECT 265.2000 254.4000 265.8000 257.6000 ;
	    RECT 266.8000 255.6000 267.6000 257.2000 ;
	    RECT 268.4000 255.2000 269.2000 259.8000 ;
	    RECT 268.4000 254.6000 270.6000 255.2000 ;
	    RECT 209.4000 251.0000 210.0000 253.0000 ;
	    RECT 210.8000 251.6000 211.6000 253.2000 ;
	    RECT 212.4000 251.6000 213.2000 253.2000 ;
	    RECT 214.0000 251.6000 214.8000 253.2000 ;
	    RECT 215.6000 251.6000 216.4000 253.2000 ;
	    RECT 217.2000 253.0000 218.6000 253.8000 ;
	    RECT 219.2000 253.6000 221.2000 254.4000 ;
	    RECT 217.2000 251.0000 217.8000 253.0000 ;
	    RECT 209.4000 250.4000 213.2000 251.0000 ;
	    RECT 207.4000 249.2000 209.0000 249.8000 ;
	    RECT 208.2000 244.4000 209.0000 249.2000 ;
	    RECT 212.6000 247.0000 213.2000 250.4000 ;
	    RECT 207.6000 243.6000 209.0000 244.4000 ;
	    RECT 208.2000 242.2000 209.0000 243.6000 ;
	    RECT 212.4000 243.0000 213.2000 247.0000 ;
	    RECT 214.0000 250.4000 217.8000 251.0000 ;
	    RECT 214.0000 247.0000 214.6000 250.4000 ;
	    RECT 219.2000 249.8000 219.8000 253.6000 ;
	    RECT 223.6000 252.8000 224.4000 254.4000 ;
	    RECT 225.2000 253.8000 227.6000 254.4000 ;
	    RECT 229.2000 254.3000 230.8000 254.4000 ;
	    RECT 231.6000 254.3000 234.2000 254.4000 ;
	    RECT 229.2000 253.8000 234.2000 254.3000 ;
	    RECT 235.6000 253.8000 237.2000 254.4000 ;
	    RECT 226.8000 253.6000 227.6000 253.8000 ;
	    RECT 230.0000 253.7000 234.2000 253.8000 ;
	    RECT 230.0000 253.6000 230.8000 253.7000 ;
	    RECT 231.6000 253.6000 234.2000 253.7000 ;
	    RECT 236.4000 253.6000 237.2000 253.8000 ;
	    RECT 238.0000 253.8000 239.6000 254.4000 ;
	    RECT 238.0000 253.6000 238.8000 253.8000 ;
	    RECT 241.0000 253.6000 243.6000 254.4000 ;
	    RECT 220.4000 250.8000 221.2000 252.4000 ;
	    RECT 225.2000 251.6000 226.0000 253.2000 ;
	    RECT 227.0000 250.2000 227.6000 253.6000 ;
	    RECT 228.4000 251.6000 229.2000 253.2000 ;
	    RECT 231.6000 250.2000 232.4000 250.4000 ;
	    RECT 233.6000 250.2000 234.2000 253.6000 ;
	    RECT 234.8000 251.6000 235.6000 253.2000 ;
	    RECT 236.5000 252.3000 237.1000 253.6000 ;
	    RECT 239.6000 252.3000 240.4000 253.2000 ;
	    RECT 236.5000 251.7000 240.4000 252.3000 ;
	    RECT 239.6000 251.6000 240.4000 251.7000 ;
	    RECT 241.0000 250.2000 241.6000 253.6000 ;
	    RECT 244.4000 252.3000 245.2000 254.4000 ;
	    RECT 246.0000 253.8000 248.4000 254.4000 ;
	    RECT 250.0000 253.8000 251.6000 254.4000 ;
	    RECT 247.6000 253.6000 248.4000 253.8000 ;
	    RECT 250.8000 253.6000 251.6000 253.8000 ;
	    RECT 254.0000 253.6000 254.8000 254.4000 ;
	    RECT 265.2000 253.6000 266.0000 254.4000 ;
	    RECT 242.9000 251.7000 245.2000 252.3000 ;
	    RECT 242.9000 250.4000 243.5000 251.7000 ;
	    RECT 246.0000 251.6000 246.8000 253.2000 ;
	    RECT 242.8000 250.2000 243.6000 250.4000 ;
	    RECT 247.8000 250.2000 248.4000 253.6000 ;
	    RECT 249.2000 252.3000 250.0000 253.2000 ;
	    RECT 250.8000 252.3000 251.6000 252.4000 ;
	    RECT 249.2000 251.7000 251.6000 252.3000 ;
	    RECT 249.2000 251.6000 250.0000 251.7000 ;
	    RECT 250.8000 251.6000 251.6000 251.7000 ;
	    RECT 252.4000 250.8000 253.2000 252.4000 ;
	    RECT 254.0000 250.2000 254.6000 253.6000 ;
	    RECT 255.6000 252.3000 256.4000 252.4000 ;
	    RECT 260.4000 252.3000 261.2000 252.4000 ;
	    RECT 255.6000 251.7000 261.2000 252.3000 ;
	    RECT 255.6000 251.6000 256.4000 251.7000 ;
	    RECT 260.4000 251.6000 261.2000 251.7000 ;
	    RECT 262.0000 252.3000 262.8000 252.4000 ;
	    RECT 263.6000 252.3000 264.4000 252.4000 ;
	    RECT 262.0000 251.7000 264.4000 252.3000 ;
	    RECT 262.0000 251.6000 262.8000 251.7000 ;
	    RECT 263.6000 250.8000 264.4000 251.7000 ;
	    RECT 265.2000 250.2000 265.8000 253.6000 ;
	    RECT 270.0000 251.6000 270.6000 254.6000 ;
	    RECT 271.6000 252.4000 272.4000 259.8000 ;
	    RECT 270.0000 250.8000 271.2000 251.6000 ;
	    RECT 270.0000 250.2000 270.6000 250.8000 ;
	    RECT 271.8000 250.2000 272.4000 252.4000 ;
	    RECT 218.2000 249.2000 219.8000 249.8000 ;
	    RECT 214.0000 243.0000 214.8000 247.0000 ;
	    RECT 218.2000 244.4000 219.0000 249.2000 ;
	    RECT 226.2000 248.4000 228.2000 250.2000 ;
	    RECT 231.6000 249.6000 233.0000 250.2000 ;
	    RECT 233.6000 249.6000 234.6000 250.2000 ;
	    RECT 232.4000 248.4000 233.0000 249.6000 ;
	    RECT 225.2000 247.6000 228.2000 248.4000 ;
	    RECT 231.6000 247.6000 233.2000 248.4000 ;
	    RECT 218.2000 243.6000 219.6000 244.4000 ;
	    RECT 218.2000 242.2000 219.0000 243.6000 ;
	    RECT 226.2000 242.2000 228.2000 247.6000 ;
	    RECT 233.8000 242.2000 234.6000 249.6000 ;
	    RECT 240.6000 249.6000 241.6000 250.2000 ;
	    RECT 242.2000 249.6000 243.6000 250.2000 ;
	    RECT 240.6000 248.4000 241.4000 249.6000 ;
	    RECT 242.2000 248.4000 242.8000 249.6000 ;
	    RECT 239.6000 247.6000 241.4000 248.4000 ;
	    RECT 242.0000 247.6000 242.8000 248.4000 ;
	    RECT 240.6000 242.2000 241.4000 247.6000 ;
	    RECT 247.0000 242.2000 249.0000 250.2000 ;
	    RECT 253.0000 249.4000 254.8000 250.2000 ;
	    RECT 264.2000 249.4000 266.0000 250.2000 ;
	    RECT 268.4000 249.6000 270.6000 250.2000 ;
	    RECT 253.0000 248.4000 253.8000 249.4000 ;
	    RECT 252.4000 247.6000 253.8000 248.4000 ;
	    RECT 253.0000 242.2000 253.8000 247.6000 ;
	    RECT 264.2000 242.2000 265.0000 249.4000 ;
	    RECT 268.4000 242.2000 269.2000 249.6000 ;
	    RECT 271.6000 242.2000 272.4000 250.2000 ;
	    RECT 273.2000 255.4000 274.0000 259.8000 ;
	    RECT 277.4000 258.4000 278.6000 259.8000 ;
	    RECT 277.4000 257.8000 278.8000 258.4000 ;
	    RECT 282.0000 257.8000 282.8000 259.8000 ;
	    RECT 286.4000 258.4000 287.2000 259.8000 ;
	    RECT 286.4000 257.8000 288.4000 258.4000 ;
	    RECT 278.0000 257.0000 278.8000 257.8000 ;
	    RECT 282.2000 257.2000 282.8000 257.8000 ;
	    RECT 282.2000 256.6000 285.0000 257.2000 ;
	    RECT 284.2000 256.4000 285.0000 256.6000 ;
	    RECT 286.0000 255.6000 286.8000 257.2000 ;
	    RECT 287.6000 257.0000 288.4000 257.8000 ;
	    RECT 276.2000 255.4000 277.0000 255.6000 ;
	    RECT 273.2000 254.8000 277.0000 255.4000 ;
	    RECT 273.2000 251.4000 274.0000 254.8000 ;
	    RECT 280.2000 254.2000 281.0000 254.4000 ;
	    RECT 286.0000 254.2000 286.6000 255.6000 ;
	    RECT 290.8000 255.0000 291.6000 259.8000 ;
	    RECT 295.0000 256.4000 295.8000 259.8000 ;
	    RECT 294.0000 255.8000 295.8000 256.4000 ;
	    RECT 297.2000 255.8000 298.0000 259.8000 ;
	    RECT 298.8000 256.0000 299.6000 259.8000 ;
	    RECT 302.0000 256.0000 302.8000 259.8000 ;
	    RECT 298.8000 255.8000 302.8000 256.0000 ;
	    RECT 289.2000 254.2000 290.8000 254.4000 ;
	    RECT 279.8000 253.6000 290.8000 254.2000 ;
	    RECT 292.4000 253.6000 293.2000 255.2000 ;
	    RECT 278.0000 252.8000 278.8000 253.0000 ;
	    RECT 275.0000 252.2000 278.8000 252.8000 ;
	    RECT 275.0000 252.0000 275.8000 252.2000 ;
	    RECT 276.6000 251.4000 277.4000 251.6000 ;
	    RECT 273.2000 250.8000 277.4000 251.4000 ;
	    RECT 273.2000 242.2000 274.0000 250.8000 ;
	    RECT 279.8000 250.4000 280.4000 253.6000 ;
	    RECT 287.0000 253.4000 287.8000 253.6000 ;
	    RECT 286.0000 252.4000 286.8000 252.6000 ;
	    RECT 288.6000 252.4000 289.4000 252.6000 ;
	    RECT 284.4000 251.8000 289.4000 252.4000 ;
	    RECT 294.0000 252.3000 294.8000 255.8000 ;
	    RECT 297.4000 254.4000 298.0000 255.8000 ;
	    RECT 299.0000 255.4000 302.6000 255.8000 ;
	    RECT 303.6000 255.2000 304.4000 259.8000 ;
	    RECT 301.2000 254.4000 302.0000 254.8000 ;
	    RECT 303.6000 254.6000 305.8000 255.2000 ;
	    RECT 295.6000 254.3000 296.4000 254.4000 ;
	    RECT 297.2000 254.3000 299.8000 254.4000 ;
	    RECT 295.6000 253.7000 299.8000 254.3000 ;
	    RECT 301.2000 253.8000 302.8000 254.4000 ;
	    RECT 295.6000 253.6000 296.4000 253.7000 ;
	    RECT 297.2000 253.6000 299.8000 253.7000 ;
	    RECT 302.0000 253.6000 302.8000 253.8000 ;
	    RECT 284.4000 251.6000 285.2000 251.8000 ;
	    RECT 294.0000 251.7000 297.9000 252.3000 ;
	    RECT 286.0000 251.0000 291.6000 251.2000 ;
	    RECT 285.8000 250.8000 291.6000 251.0000 ;
	    RECT 278.0000 249.8000 280.4000 250.4000 ;
	    RECT 281.8000 250.6000 291.6000 250.8000 ;
	    RECT 281.8000 250.2000 286.6000 250.6000 ;
	    RECT 278.0000 248.8000 278.6000 249.8000 ;
	    RECT 277.2000 248.0000 278.6000 248.8000 ;
	    RECT 280.2000 249.0000 281.0000 249.2000 ;
	    RECT 281.8000 249.0000 282.4000 250.2000 ;
	    RECT 280.2000 248.4000 282.4000 249.0000 ;
	    RECT 283.0000 249.0000 288.4000 249.6000 ;
	    RECT 283.0000 248.8000 283.8000 249.0000 ;
	    RECT 287.6000 248.8000 288.4000 249.0000 ;
	    RECT 281.4000 247.4000 282.2000 247.6000 ;
	    RECT 284.2000 247.4000 285.0000 247.6000 ;
	    RECT 278.0000 246.2000 278.8000 247.0000 ;
	    RECT 281.4000 246.8000 285.0000 247.4000 ;
	    RECT 282.2000 246.2000 282.8000 246.8000 ;
	    RECT 287.6000 246.2000 288.4000 247.0000 ;
	    RECT 277.4000 242.2000 278.6000 246.2000 ;
	    RECT 282.0000 242.2000 282.8000 246.2000 ;
	    RECT 286.4000 245.6000 288.4000 246.2000 ;
	    RECT 286.4000 242.2000 287.2000 245.6000 ;
	    RECT 290.8000 242.2000 291.6000 250.6000 ;
	    RECT 294.0000 242.2000 294.8000 251.7000 ;
	    RECT 297.3000 250.4000 297.9000 251.7000 ;
	    RECT 295.6000 248.8000 296.4000 250.4000 ;
	    RECT 297.2000 250.2000 298.0000 250.4000 ;
	    RECT 299.2000 250.2000 299.8000 253.6000 ;
	    RECT 300.4000 251.6000 301.2000 253.2000 ;
	    RECT 305.2000 251.6000 305.8000 254.6000 ;
	    RECT 306.8000 252.4000 307.6000 259.8000 ;
	    RECT 305.2000 250.8000 306.4000 251.6000 ;
	    RECT 305.2000 250.2000 305.8000 250.8000 ;
	    RECT 307.0000 250.2000 307.6000 252.4000 ;
	    RECT 297.2000 249.6000 298.6000 250.2000 ;
	    RECT 299.2000 249.6000 300.2000 250.2000 ;
	    RECT 298.0000 248.4000 298.6000 249.6000 ;
	    RECT 298.0000 247.6000 298.8000 248.4000 ;
	    RECT 299.4000 242.2000 300.2000 249.6000 ;
	    RECT 303.6000 249.6000 305.8000 250.2000 ;
	    RECT 303.6000 242.2000 304.4000 249.6000 ;
	    RECT 306.8000 242.2000 307.6000 250.2000 ;
	    RECT 308.4000 252.4000 309.2000 259.8000 ;
	    RECT 311.6000 255.2000 312.4000 259.8000 ;
	    RECT 310.2000 254.6000 312.4000 255.2000 ;
	    RECT 313.2000 255.4000 314.0000 259.8000 ;
	    RECT 317.4000 258.4000 318.6000 259.8000 ;
	    RECT 317.4000 257.8000 318.8000 258.4000 ;
	    RECT 322.0000 257.8000 322.8000 259.8000 ;
	    RECT 326.4000 258.4000 327.2000 259.8000 ;
	    RECT 326.4000 257.8000 328.4000 258.4000 ;
	    RECT 318.0000 257.0000 318.8000 257.8000 ;
	    RECT 322.2000 257.2000 322.8000 257.8000 ;
	    RECT 322.2000 256.6000 325.0000 257.2000 ;
	    RECT 324.2000 256.4000 325.0000 256.6000 ;
	    RECT 326.0000 256.4000 326.8000 257.2000 ;
	    RECT 327.6000 257.0000 328.4000 257.8000 ;
	    RECT 316.2000 255.4000 317.0000 255.6000 ;
	    RECT 313.2000 254.8000 317.0000 255.4000 ;
	    RECT 308.4000 250.2000 309.0000 252.4000 ;
	    RECT 310.2000 251.6000 310.8000 254.6000 ;
	    RECT 309.6000 250.8000 310.8000 251.6000 ;
	    RECT 310.2000 250.2000 310.8000 250.8000 ;
	    RECT 313.2000 251.4000 314.0000 254.8000 ;
	    RECT 320.2000 254.2000 321.0000 254.4000 ;
	    RECT 326.0000 254.2000 326.6000 256.4000 ;
	    RECT 330.8000 255.0000 331.6000 259.8000 ;
	    RECT 335.0000 256.4000 335.8000 259.8000 ;
	    RECT 334.0000 255.8000 335.8000 256.4000 ;
	    RECT 337.2000 255.8000 338.0000 259.8000 ;
	    RECT 338.8000 256.0000 339.6000 259.8000 ;
	    RECT 342.0000 256.0000 342.8000 259.8000 ;
	    RECT 338.8000 255.8000 342.8000 256.0000 ;
	    RECT 329.2000 254.2000 330.8000 254.4000 ;
	    RECT 319.8000 253.6000 330.8000 254.2000 ;
	    RECT 332.4000 253.6000 333.2000 255.2000 ;
	    RECT 318.0000 252.8000 318.8000 253.0000 ;
	    RECT 315.0000 252.2000 318.8000 252.8000 ;
	    RECT 319.8000 252.4000 320.4000 253.6000 ;
	    RECT 327.0000 253.4000 327.8000 253.6000 ;
	    RECT 326.0000 252.4000 326.8000 252.6000 ;
	    RECT 328.6000 252.4000 329.4000 252.6000 ;
	    RECT 315.0000 252.0000 315.8000 252.2000 ;
	    RECT 319.6000 251.6000 320.4000 252.4000 ;
	    RECT 324.4000 251.8000 329.4000 252.4000 ;
	    RECT 334.0000 252.3000 334.8000 255.8000 ;
	    RECT 337.4000 254.4000 338.0000 255.8000 ;
	    RECT 339.0000 255.4000 342.6000 255.8000 ;
	    RECT 343.6000 255.2000 344.4000 259.8000 ;
	    RECT 341.2000 254.4000 342.0000 254.8000 ;
	    RECT 343.6000 254.6000 345.8000 255.2000 ;
	    RECT 337.2000 253.6000 339.8000 254.4000 ;
	    RECT 341.2000 253.8000 342.8000 254.4000 ;
	    RECT 342.0000 253.6000 342.8000 253.8000 ;
	    RECT 324.4000 251.6000 325.2000 251.8000 ;
	    RECT 334.0000 251.7000 337.9000 252.3000 ;
	    RECT 316.6000 251.4000 317.4000 251.6000 ;
	    RECT 313.2000 250.8000 317.4000 251.4000 ;
	    RECT 308.4000 242.2000 309.2000 250.2000 ;
	    RECT 310.2000 249.6000 312.4000 250.2000 ;
	    RECT 311.6000 242.2000 312.4000 249.6000 ;
	    RECT 313.2000 242.2000 314.0000 250.8000 ;
	    RECT 319.8000 250.4000 320.4000 251.6000 ;
	    RECT 326.0000 251.0000 331.6000 251.2000 ;
	    RECT 325.8000 250.8000 331.6000 251.0000 ;
	    RECT 318.0000 249.8000 320.4000 250.4000 ;
	    RECT 321.8000 250.6000 331.6000 250.8000 ;
	    RECT 321.8000 250.2000 326.6000 250.6000 ;
	    RECT 318.0000 248.8000 318.6000 249.8000 ;
	    RECT 317.2000 248.0000 318.6000 248.8000 ;
	    RECT 320.2000 249.0000 321.0000 249.2000 ;
	    RECT 321.8000 249.0000 322.4000 250.2000 ;
	    RECT 320.2000 248.4000 322.4000 249.0000 ;
	    RECT 323.0000 249.0000 328.4000 249.6000 ;
	    RECT 323.0000 248.8000 323.8000 249.0000 ;
	    RECT 327.6000 248.8000 328.4000 249.0000 ;
	    RECT 321.4000 247.4000 322.2000 247.6000 ;
	    RECT 324.2000 247.4000 325.0000 247.6000 ;
	    RECT 318.0000 246.2000 318.8000 247.0000 ;
	    RECT 321.4000 246.8000 325.0000 247.4000 ;
	    RECT 322.2000 246.2000 322.8000 246.8000 ;
	    RECT 327.6000 246.2000 328.4000 247.0000 ;
	    RECT 317.4000 242.2000 318.6000 246.2000 ;
	    RECT 322.0000 242.2000 322.8000 246.2000 ;
	    RECT 326.4000 245.6000 328.4000 246.2000 ;
	    RECT 326.4000 242.2000 327.2000 245.6000 ;
	    RECT 330.8000 242.2000 331.6000 250.6000 ;
	    RECT 334.0000 242.2000 334.8000 251.7000 ;
	    RECT 337.3000 250.4000 337.9000 251.7000 ;
	    RECT 335.6000 248.8000 336.4000 250.4000 ;
	    RECT 337.2000 250.2000 338.0000 250.4000 ;
	    RECT 339.2000 250.2000 339.8000 253.6000 ;
	    RECT 340.4000 251.6000 341.2000 253.2000 ;
	    RECT 343.6000 251.6000 344.4000 253.2000 ;
	    RECT 345.2000 251.6000 345.8000 254.6000 ;
	    RECT 346.8000 252.4000 347.6000 259.8000 ;
	    RECT 345.2000 250.8000 346.4000 251.6000 ;
	    RECT 345.2000 250.2000 345.8000 250.8000 ;
	    RECT 347.0000 250.2000 347.6000 252.4000 ;
	    RECT 337.2000 249.6000 338.6000 250.2000 ;
	    RECT 339.2000 249.6000 340.2000 250.2000 ;
	    RECT 338.0000 248.4000 338.6000 249.6000 ;
	    RECT 338.0000 247.6000 338.8000 248.4000 ;
	    RECT 339.4000 242.2000 340.2000 249.6000 ;
	    RECT 343.6000 249.6000 345.8000 250.2000 ;
	    RECT 343.6000 242.2000 344.4000 249.6000 ;
	    RECT 346.8000 242.2000 347.6000 250.2000 ;
	    RECT 348.4000 255.8000 349.2000 259.8000 ;
	    RECT 351.6000 257.8000 352.4000 259.8000 ;
	    RECT 348.4000 254.4000 349.0000 255.8000 ;
	    RECT 351.6000 255.6000 352.2000 257.8000 ;
	    RECT 353.2000 255.6000 354.0000 257.2000 ;
	    RECT 349.8000 255.0000 352.2000 255.6000 ;
	    RECT 354.8000 255.4000 355.6000 259.8000 ;
	    RECT 359.0000 258.4000 360.2000 259.8000 ;
	    RECT 359.0000 257.8000 360.4000 258.4000 ;
	    RECT 363.6000 257.8000 364.4000 259.8000 ;
	    RECT 368.0000 258.4000 368.8000 259.8000 ;
	    RECT 368.0000 257.8000 370.0000 258.4000 ;
	    RECT 359.6000 257.0000 360.4000 257.8000 ;
	    RECT 363.8000 257.2000 364.4000 257.8000 ;
	    RECT 363.8000 256.6000 366.6000 257.2000 ;
	    RECT 365.8000 256.4000 366.6000 256.6000 ;
	    RECT 367.6000 256.4000 368.4000 257.2000 ;
	    RECT 369.2000 257.0000 370.0000 257.8000 ;
	    RECT 357.8000 255.4000 358.6000 255.6000 ;
	    RECT 348.4000 253.6000 349.2000 254.4000 ;
	    RECT 348.4000 252.4000 349.0000 253.6000 ;
	    RECT 348.4000 251.6000 349.2000 252.4000 ;
	    RECT 349.8000 252.0000 350.4000 255.0000 ;
	    RECT 354.8000 254.8000 358.6000 255.4000 ;
	    RECT 351.4000 253.6000 352.4000 254.4000 ;
	    RECT 351.2000 252.8000 352.0000 253.6000 ;
	    RECT 348.4000 250.2000 349.0000 251.6000 ;
	    RECT 349.8000 251.4000 350.6000 252.0000 ;
	    RECT 354.8000 251.4000 355.6000 254.8000 ;
	    RECT 361.8000 254.2000 362.6000 254.4000 ;
	    RECT 366.0000 254.2000 366.8000 254.4000 ;
	    RECT 367.6000 254.2000 368.2000 256.4000 ;
	    RECT 372.4000 255.0000 373.2000 259.8000 ;
	    RECT 374.0000 255.4000 374.8000 259.8000 ;
	    RECT 378.2000 258.4000 379.4000 259.8000 ;
	    RECT 378.2000 257.8000 379.6000 258.4000 ;
	    RECT 382.8000 257.8000 383.6000 259.8000 ;
	    RECT 387.2000 258.4000 388.0000 259.8000 ;
	    RECT 387.2000 257.8000 389.2000 258.4000 ;
	    RECT 378.8000 257.0000 379.6000 257.8000 ;
	    RECT 383.0000 257.2000 383.6000 257.8000 ;
	    RECT 383.0000 256.6000 385.8000 257.2000 ;
	    RECT 385.0000 256.4000 385.8000 256.6000 ;
	    RECT 386.8000 256.4000 387.6000 257.2000 ;
	    RECT 388.4000 257.0000 389.2000 257.8000 ;
	    RECT 377.0000 255.4000 377.8000 255.6000 ;
	    RECT 374.0000 254.8000 377.8000 255.4000 ;
	    RECT 370.8000 254.2000 372.4000 254.4000 ;
	    RECT 361.4000 253.6000 372.4000 254.2000 ;
	    RECT 359.6000 252.8000 360.4000 253.0000 ;
	    RECT 356.6000 252.2000 360.4000 252.8000 ;
	    RECT 356.6000 252.0000 357.4000 252.2000 ;
	    RECT 358.2000 251.4000 359.0000 251.6000 ;
	    RECT 349.8000 251.2000 354.0000 251.4000 ;
	    RECT 350.0000 250.8000 354.0000 251.2000 ;
	    RECT 348.4000 249.6000 349.8000 250.2000 ;
	    RECT 349.0000 242.2000 349.8000 249.6000 ;
	    RECT 353.2000 242.2000 354.0000 250.8000 ;
	    RECT 354.8000 250.8000 359.0000 251.4000 ;
	    RECT 354.8000 242.2000 355.6000 250.8000 ;
	    RECT 361.4000 250.4000 362.0000 253.6000 ;
	    RECT 368.6000 253.4000 369.4000 253.6000 ;
	    RECT 367.6000 252.4000 368.4000 252.6000 ;
	    RECT 370.2000 252.4000 371.0000 252.6000 ;
	    RECT 366.0000 251.8000 371.0000 252.4000 ;
	    RECT 366.0000 251.6000 366.8000 251.8000 ;
	    RECT 374.0000 251.4000 374.8000 254.8000 ;
	    RECT 381.0000 254.2000 381.8000 254.4000 ;
	    RECT 383.6000 254.2000 384.4000 254.4000 ;
	    RECT 386.8000 254.2000 387.4000 256.4000 ;
	    RECT 391.6000 255.0000 392.4000 259.8000 ;
	    RECT 393.2000 255.4000 394.0000 259.8000 ;
	    RECT 397.4000 258.4000 398.6000 259.8000 ;
	    RECT 397.4000 257.8000 398.8000 258.4000 ;
	    RECT 402.0000 257.8000 402.8000 259.8000 ;
	    RECT 406.4000 258.4000 407.2000 259.8000 ;
	    RECT 406.4000 257.8000 408.4000 258.4000 ;
	    RECT 398.0000 257.0000 398.8000 257.8000 ;
	    RECT 402.2000 257.2000 402.8000 257.8000 ;
	    RECT 402.2000 256.6000 405.0000 257.2000 ;
	    RECT 404.2000 256.4000 405.0000 256.6000 ;
	    RECT 406.0000 256.4000 406.8000 257.2000 ;
	    RECT 407.6000 257.0000 408.4000 257.8000 ;
	    RECT 396.2000 255.4000 397.0000 255.6000 ;
	    RECT 393.2000 254.8000 397.0000 255.4000 ;
	    RECT 390.0000 254.2000 391.6000 254.4000 ;
	    RECT 380.6000 253.6000 391.6000 254.2000 ;
	    RECT 378.8000 252.8000 379.6000 253.0000 ;
	    RECT 375.8000 252.2000 379.6000 252.8000 ;
	    RECT 375.8000 252.0000 376.6000 252.2000 ;
	    RECT 377.4000 251.4000 378.2000 251.6000 ;
	    RECT 367.6000 251.0000 373.2000 251.2000 ;
	    RECT 367.4000 250.8000 373.2000 251.0000 ;
	    RECT 359.6000 249.8000 362.0000 250.4000 ;
	    RECT 363.4000 250.6000 373.2000 250.8000 ;
	    RECT 363.4000 250.2000 368.2000 250.6000 ;
	    RECT 359.6000 248.8000 360.2000 249.8000 ;
	    RECT 358.8000 248.0000 360.2000 248.8000 ;
	    RECT 361.8000 249.0000 362.6000 249.2000 ;
	    RECT 363.4000 249.0000 364.0000 250.2000 ;
	    RECT 361.8000 248.4000 364.0000 249.0000 ;
	    RECT 364.6000 249.0000 370.0000 249.6000 ;
	    RECT 364.6000 248.8000 365.4000 249.0000 ;
	    RECT 369.2000 248.8000 370.0000 249.0000 ;
	    RECT 363.0000 247.4000 363.8000 247.6000 ;
	    RECT 365.8000 247.4000 366.6000 247.6000 ;
	    RECT 359.6000 246.2000 360.4000 247.0000 ;
	    RECT 363.0000 246.8000 366.6000 247.4000 ;
	    RECT 363.8000 246.2000 364.4000 246.8000 ;
	    RECT 369.2000 246.2000 370.0000 247.0000 ;
	    RECT 359.0000 242.2000 360.2000 246.2000 ;
	    RECT 363.6000 242.2000 364.4000 246.2000 ;
	    RECT 368.0000 245.6000 370.0000 246.2000 ;
	    RECT 368.0000 242.2000 368.8000 245.6000 ;
	    RECT 372.4000 242.2000 373.2000 250.6000 ;
	    RECT 374.0000 250.8000 378.2000 251.4000 ;
	    RECT 374.0000 242.2000 374.8000 250.8000 ;
	    RECT 380.6000 250.4000 381.2000 253.6000 ;
	    RECT 387.8000 253.4000 388.6000 253.6000 ;
	    RECT 386.8000 252.4000 387.6000 252.6000 ;
	    RECT 389.4000 252.4000 390.2000 252.6000 ;
	    RECT 385.2000 251.8000 390.2000 252.4000 ;
	    RECT 385.2000 251.6000 386.0000 251.8000 ;
	    RECT 393.2000 251.4000 394.0000 254.8000 ;
	    RECT 400.2000 254.2000 401.0000 254.4000 ;
	    RECT 406.0000 254.2000 406.6000 256.4000 ;
	    RECT 410.8000 255.0000 411.6000 259.8000 ;
	    RECT 418.8000 255.8000 419.6000 259.8000 ;
	    RECT 420.4000 256.0000 421.2000 259.8000 ;
	    RECT 423.6000 256.0000 424.4000 259.8000 ;
	    RECT 420.4000 255.8000 424.4000 256.0000 ;
	    RECT 419.0000 254.4000 419.6000 255.8000 ;
	    RECT 420.6000 255.4000 424.2000 255.8000 ;
	    RECT 422.8000 254.4000 423.6000 254.8000 ;
	    RECT 409.2000 254.2000 410.8000 254.4000 ;
	    RECT 399.8000 253.6000 410.8000 254.2000 ;
	    RECT 418.8000 253.6000 421.4000 254.4000 ;
	    RECT 422.8000 253.8000 424.4000 254.4000 ;
	    RECT 423.6000 253.6000 424.4000 253.8000 ;
	    RECT 398.0000 252.8000 398.8000 253.0000 ;
	    RECT 395.0000 252.2000 398.8000 252.8000 ;
	    RECT 395.0000 252.0000 395.8000 252.2000 ;
	    RECT 396.6000 251.4000 397.4000 251.6000 ;
	    RECT 386.8000 251.0000 392.4000 251.2000 ;
	    RECT 386.6000 250.8000 392.4000 251.0000 ;
	    RECT 378.8000 249.8000 381.2000 250.4000 ;
	    RECT 382.6000 250.6000 392.4000 250.8000 ;
	    RECT 382.6000 250.2000 387.4000 250.6000 ;
	    RECT 378.8000 248.8000 379.4000 249.8000 ;
	    RECT 378.0000 248.0000 379.4000 248.8000 ;
	    RECT 381.0000 249.0000 381.8000 249.2000 ;
	    RECT 382.6000 249.0000 383.2000 250.2000 ;
	    RECT 381.0000 248.4000 383.2000 249.0000 ;
	    RECT 383.8000 249.0000 389.2000 249.6000 ;
	    RECT 383.8000 248.8000 384.6000 249.0000 ;
	    RECT 388.4000 248.8000 389.2000 249.0000 ;
	    RECT 382.2000 247.4000 383.0000 247.6000 ;
	    RECT 385.0000 247.4000 385.8000 247.6000 ;
	    RECT 378.8000 246.2000 379.6000 247.0000 ;
	    RECT 382.2000 246.8000 385.8000 247.4000 ;
	    RECT 383.0000 246.2000 383.6000 246.8000 ;
	    RECT 388.4000 246.2000 389.2000 247.0000 ;
	    RECT 378.2000 242.2000 379.4000 246.2000 ;
	    RECT 382.8000 242.2000 383.6000 246.2000 ;
	    RECT 387.2000 245.6000 389.2000 246.2000 ;
	    RECT 387.2000 242.2000 388.0000 245.6000 ;
	    RECT 391.6000 242.2000 392.4000 250.6000 ;
	    RECT 393.2000 250.8000 397.4000 251.4000 ;
	    RECT 393.2000 242.2000 394.0000 250.8000 ;
	    RECT 399.8000 250.4000 400.4000 253.6000 ;
	    RECT 407.0000 253.4000 407.8000 253.6000 ;
	    RECT 406.0000 252.4000 406.8000 252.6000 ;
	    RECT 408.6000 252.4000 409.4000 252.6000 ;
	    RECT 404.4000 251.8000 409.4000 252.4000 ;
	    RECT 404.4000 251.6000 405.2000 251.8000 ;
	    RECT 406.0000 251.0000 411.6000 251.2000 ;
	    RECT 405.8000 250.8000 411.6000 251.0000 ;
	    RECT 398.0000 249.8000 400.4000 250.4000 ;
	    RECT 401.8000 250.6000 411.6000 250.8000 ;
	    RECT 401.8000 250.2000 406.6000 250.6000 ;
	    RECT 398.0000 248.8000 398.6000 249.8000 ;
	    RECT 397.2000 248.0000 398.6000 248.8000 ;
	    RECT 400.2000 249.0000 401.0000 249.2000 ;
	    RECT 401.8000 249.0000 402.4000 250.2000 ;
	    RECT 400.2000 248.4000 402.4000 249.0000 ;
	    RECT 403.0000 249.0000 408.4000 249.6000 ;
	    RECT 403.0000 248.8000 403.8000 249.0000 ;
	    RECT 407.6000 248.8000 408.4000 249.0000 ;
	    RECT 401.4000 247.4000 402.2000 247.6000 ;
	    RECT 404.2000 247.4000 405.0000 247.6000 ;
	    RECT 398.0000 246.2000 398.8000 247.0000 ;
	    RECT 401.4000 246.8000 405.0000 247.4000 ;
	    RECT 402.2000 246.2000 402.8000 246.8000 ;
	    RECT 407.6000 246.2000 408.4000 247.0000 ;
	    RECT 397.4000 242.2000 398.6000 246.2000 ;
	    RECT 402.0000 242.2000 402.8000 246.2000 ;
	    RECT 406.4000 245.6000 408.4000 246.2000 ;
	    RECT 406.4000 242.2000 407.2000 245.6000 ;
	    RECT 410.8000 242.2000 411.6000 250.6000 ;
	    RECT 417.2000 250.3000 418.0000 250.4000 ;
	    RECT 418.8000 250.3000 419.6000 250.4000 ;
	    RECT 417.2000 250.2000 419.6000 250.3000 ;
	    RECT 420.8000 250.2000 421.4000 253.6000 ;
	    RECT 422.0000 251.6000 422.8000 253.2000 ;
	    RECT 417.2000 249.7000 420.2000 250.2000 ;
	    RECT 417.2000 249.6000 418.0000 249.7000 ;
	    RECT 418.8000 249.6000 420.2000 249.7000 ;
	    RECT 420.8000 249.6000 421.8000 250.2000 ;
	    RECT 419.6000 248.4000 420.2000 249.6000 ;
	    RECT 419.6000 247.6000 420.4000 248.4000 ;
	    RECT 421.0000 242.2000 421.8000 249.6000 ;
	    RECT 425.2000 242.2000 426.0000 259.8000 ;
	    RECT 428.4000 255.4000 429.2000 259.8000 ;
	    RECT 432.6000 258.4000 433.8000 259.8000 ;
	    RECT 432.6000 257.8000 434.0000 258.4000 ;
	    RECT 437.2000 257.8000 438.0000 259.8000 ;
	    RECT 441.6000 258.4000 442.4000 259.8000 ;
	    RECT 441.6000 257.8000 443.6000 258.4000 ;
	    RECT 433.2000 257.0000 434.0000 257.8000 ;
	    RECT 437.4000 257.2000 438.0000 257.8000 ;
	    RECT 437.4000 256.6000 440.2000 257.2000 ;
	    RECT 439.4000 256.4000 440.2000 256.6000 ;
	    RECT 441.2000 256.4000 442.0000 257.2000 ;
	    RECT 442.8000 257.0000 443.6000 257.8000 ;
	    RECT 431.4000 255.4000 432.2000 255.6000 ;
	    RECT 428.4000 254.8000 432.2000 255.4000 ;
	    RECT 428.4000 251.4000 429.2000 254.8000 ;
	    RECT 441.2000 254.4000 441.8000 256.4000 ;
	    RECT 446.0000 255.0000 446.8000 259.8000 ;
	    RECT 447.6000 255.6000 448.4000 257.2000 ;
	    RECT 435.4000 254.2000 436.2000 254.4000 ;
	    RECT 441.2000 254.2000 442.0000 254.4000 ;
	    RECT 444.4000 254.2000 446.0000 254.4000 ;
	    RECT 435.0000 253.6000 446.0000 254.2000 ;
	    RECT 433.2000 252.8000 434.0000 253.0000 ;
	    RECT 430.2000 252.2000 434.0000 252.8000 ;
	    RECT 430.2000 252.0000 431.0000 252.2000 ;
	    RECT 431.8000 251.4000 432.6000 251.6000 ;
	    RECT 428.4000 250.8000 432.6000 251.4000 ;
	    RECT 428.4000 242.2000 429.2000 250.8000 ;
	    RECT 435.0000 250.4000 435.6000 253.6000 ;
	    RECT 442.2000 253.4000 443.0000 253.6000 ;
	    RECT 443.8000 252.4000 444.6000 252.6000 ;
	    RECT 439.6000 251.8000 444.6000 252.4000 ;
	    RECT 439.6000 251.6000 440.4000 251.8000 ;
	    RECT 441.2000 251.0000 446.8000 251.2000 ;
	    RECT 441.0000 250.8000 446.8000 251.0000 ;
	    RECT 433.2000 249.8000 435.6000 250.4000 ;
	    RECT 437.0000 250.6000 446.8000 250.8000 ;
	    RECT 437.0000 250.2000 441.8000 250.6000 ;
	    RECT 433.2000 248.8000 433.8000 249.8000 ;
	    RECT 432.4000 248.0000 433.8000 248.8000 ;
	    RECT 435.4000 249.0000 436.2000 249.2000 ;
	    RECT 437.0000 249.0000 437.6000 250.2000 ;
	    RECT 435.4000 248.4000 437.6000 249.0000 ;
	    RECT 438.2000 249.0000 443.6000 249.6000 ;
	    RECT 438.2000 248.8000 439.0000 249.0000 ;
	    RECT 442.8000 248.8000 443.6000 249.0000 ;
	    RECT 436.6000 247.4000 437.4000 247.6000 ;
	    RECT 439.4000 247.4000 440.2000 247.6000 ;
	    RECT 433.2000 246.2000 434.0000 247.0000 ;
	    RECT 436.6000 246.8000 440.2000 247.4000 ;
	    RECT 437.4000 246.2000 438.0000 246.8000 ;
	    RECT 442.8000 246.2000 443.6000 247.0000 ;
	    RECT 432.6000 242.2000 433.8000 246.2000 ;
	    RECT 437.2000 242.2000 438.0000 246.2000 ;
	    RECT 441.6000 245.6000 443.6000 246.2000 ;
	    RECT 441.6000 242.2000 442.4000 245.6000 ;
	    RECT 446.0000 242.2000 446.8000 250.6000 ;
	    RECT 449.2000 242.2000 450.0000 259.8000 ;
	    RECT 450.8000 255.4000 451.6000 259.8000 ;
	    RECT 455.0000 258.4000 456.2000 259.8000 ;
	    RECT 455.0000 257.8000 456.4000 258.4000 ;
	    RECT 459.6000 257.8000 460.4000 259.8000 ;
	    RECT 464.0000 258.4000 464.8000 259.8000 ;
	    RECT 464.0000 257.8000 466.0000 258.4000 ;
	    RECT 455.6000 257.0000 456.4000 257.8000 ;
	    RECT 459.8000 257.2000 460.4000 257.8000 ;
	    RECT 459.8000 256.6000 462.6000 257.2000 ;
	    RECT 461.8000 256.4000 462.6000 256.6000 ;
	    RECT 463.6000 255.6000 464.4000 257.2000 ;
	    RECT 465.2000 257.0000 466.0000 257.8000 ;
	    RECT 453.8000 255.4000 454.6000 255.6000 ;
	    RECT 450.8000 254.8000 454.6000 255.4000 ;
	    RECT 450.8000 251.4000 451.6000 254.8000 ;
	    RECT 457.8000 254.2000 458.6000 254.4000 ;
	    RECT 463.6000 254.2000 464.2000 255.6000 ;
	    RECT 468.4000 255.0000 469.2000 259.8000 ;
	    RECT 470.0000 255.6000 470.8000 257.2000 ;
	    RECT 466.8000 254.2000 468.4000 254.4000 ;
	    RECT 457.4000 253.6000 468.4000 254.2000 ;
	    RECT 471.6000 254.3000 472.4000 259.8000 ;
	    RECT 473.2000 256.0000 474.0000 259.8000 ;
	    RECT 476.4000 256.0000 477.2000 259.8000 ;
	    RECT 473.2000 255.8000 477.2000 256.0000 ;
	    RECT 478.0000 255.8000 478.8000 259.8000 ;
	    RECT 473.4000 255.4000 477.0000 255.8000 ;
	    RECT 474.0000 254.4000 474.8000 254.8000 ;
	    RECT 478.0000 254.4000 478.6000 255.8000 ;
	    RECT 479.6000 255.4000 480.4000 259.8000 ;
	    RECT 483.8000 258.4000 485.0000 259.8000 ;
	    RECT 483.8000 257.8000 485.2000 258.4000 ;
	    RECT 488.4000 257.8000 489.2000 259.8000 ;
	    RECT 492.8000 258.4000 493.6000 259.8000 ;
	    RECT 492.8000 257.8000 494.8000 258.4000 ;
	    RECT 484.4000 257.0000 485.2000 257.8000 ;
	    RECT 488.6000 257.2000 489.2000 257.8000 ;
	    RECT 488.6000 256.6000 491.4000 257.2000 ;
	    RECT 490.6000 256.4000 491.4000 256.6000 ;
	    RECT 492.4000 256.4000 493.2000 257.2000 ;
	    RECT 494.0000 257.0000 494.8000 257.8000 ;
	    RECT 482.6000 255.4000 483.4000 255.6000 ;
	    RECT 479.6000 254.8000 483.4000 255.4000 ;
	    RECT 473.2000 254.3000 474.8000 254.4000 ;
	    RECT 471.6000 253.8000 474.8000 254.3000 ;
	    RECT 471.6000 253.7000 474.0000 253.8000 ;
	    RECT 455.6000 252.8000 456.4000 253.0000 ;
	    RECT 452.6000 252.2000 456.4000 252.8000 ;
	    RECT 457.4000 252.4000 458.0000 253.6000 ;
	    RECT 464.6000 253.4000 465.4000 253.6000 ;
	    RECT 463.6000 252.4000 464.4000 252.6000 ;
	    RECT 466.2000 252.4000 467.0000 252.6000 ;
	    RECT 452.6000 252.0000 453.4000 252.2000 ;
	    RECT 457.2000 251.6000 458.0000 252.4000 ;
	    RECT 462.0000 251.8000 467.0000 252.4000 ;
	    RECT 462.0000 251.6000 462.8000 251.8000 ;
	    RECT 454.2000 251.4000 455.0000 251.6000 ;
	    RECT 450.8000 250.8000 455.0000 251.4000 ;
	    RECT 450.8000 242.2000 451.6000 250.8000 ;
	    RECT 457.4000 250.4000 458.0000 251.6000 ;
	    RECT 463.6000 251.0000 469.2000 251.2000 ;
	    RECT 463.4000 250.8000 469.2000 251.0000 ;
	    RECT 455.6000 249.8000 458.0000 250.4000 ;
	    RECT 459.4000 250.6000 469.2000 250.8000 ;
	    RECT 459.4000 250.2000 464.2000 250.6000 ;
	    RECT 455.6000 248.8000 456.2000 249.8000 ;
	    RECT 454.8000 248.0000 456.2000 248.8000 ;
	    RECT 457.8000 249.0000 458.6000 249.2000 ;
	    RECT 459.4000 249.0000 460.0000 250.2000 ;
	    RECT 457.8000 248.4000 460.0000 249.0000 ;
	    RECT 460.6000 249.0000 466.0000 249.6000 ;
	    RECT 460.6000 248.8000 461.4000 249.0000 ;
	    RECT 465.2000 248.8000 466.0000 249.0000 ;
	    RECT 459.0000 247.4000 459.8000 247.6000 ;
	    RECT 461.8000 247.4000 462.6000 247.6000 ;
	    RECT 455.6000 246.2000 456.4000 247.0000 ;
	    RECT 459.0000 246.8000 462.6000 247.4000 ;
	    RECT 459.8000 246.2000 460.4000 246.8000 ;
	    RECT 465.2000 246.2000 466.0000 247.0000 ;
	    RECT 455.0000 242.2000 456.2000 246.2000 ;
	    RECT 459.6000 242.2000 460.4000 246.2000 ;
	    RECT 464.0000 245.6000 466.0000 246.2000 ;
	    RECT 464.0000 242.2000 464.8000 245.6000 ;
	    RECT 468.4000 242.2000 469.2000 250.6000 ;
	    RECT 471.6000 242.2000 472.4000 253.7000 ;
	    RECT 473.2000 253.6000 474.0000 253.7000 ;
	    RECT 476.2000 253.6000 478.8000 254.4000 ;
	    RECT 474.8000 251.6000 475.6000 253.2000 ;
	    RECT 476.2000 250.4000 476.8000 253.6000 ;
	    RECT 479.6000 251.4000 480.4000 254.8000 ;
	    RECT 486.6000 254.2000 487.4000 254.4000 ;
	    RECT 492.4000 254.2000 493.0000 256.4000 ;
	    RECT 497.2000 255.0000 498.0000 259.8000 ;
	    RECT 495.6000 254.2000 497.2000 254.4000 ;
	    RECT 500.0000 254.2000 500.8000 259.8000 ;
	    RECT 505.2000 255.8000 506.0000 259.8000 ;
	    RECT 506.8000 256.0000 507.6000 259.8000 ;
	    RECT 510.0000 256.0000 510.8000 259.8000 ;
	    RECT 506.8000 255.8000 510.8000 256.0000 ;
	    RECT 505.4000 254.4000 506.0000 255.8000 ;
	    RECT 507.0000 255.4000 510.6000 255.8000 ;
	    RECT 509.2000 254.4000 510.0000 254.8000 ;
	    RECT 486.2000 253.6000 497.2000 254.2000 ;
	    RECT 499.0000 253.8000 500.8000 254.2000 ;
	    RECT 499.0000 253.6000 500.6000 253.8000 ;
	    RECT 505.2000 253.6000 507.8000 254.4000 ;
	    RECT 509.2000 254.3000 510.8000 254.4000 ;
	    RECT 511.6000 254.3000 512.4000 259.8000 ;
	    RECT 513.2000 255.6000 514.0000 257.2000 ;
	    RECT 509.2000 253.8000 512.4000 254.3000 ;
	    RECT 510.0000 253.7000 512.4000 253.8000 ;
	    RECT 510.0000 253.6000 510.8000 253.7000 ;
	    RECT 484.4000 252.8000 485.2000 253.0000 ;
	    RECT 481.4000 252.2000 485.2000 252.8000 ;
	    RECT 486.2000 252.4000 486.8000 253.6000 ;
	    RECT 493.4000 253.4000 494.2000 253.6000 ;
	    RECT 495.0000 252.4000 495.8000 252.6000 ;
	    RECT 481.4000 252.0000 482.2000 252.2000 ;
	    RECT 486.0000 251.6000 486.8000 252.4000 ;
	    RECT 490.8000 251.8000 495.8000 252.4000 ;
	    RECT 490.8000 251.6000 491.6000 251.8000 ;
	    RECT 483.0000 251.4000 483.8000 251.6000 ;
	    RECT 479.6000 250.8000 483.8000 251.4000 ;
	    RECT 474.8000 249.6000 476.8000 250.4000 ;
	    RECT 478.0000 250.2000 478.8000 250.4000 ;
	    RECT 477.4000 249.6000 478.8000 250.2000 ;
	    RECT 475.8000 242.2000 476.6000 249.6000 ;
	    RECT 477.4000 248.4000 478.0000 249.6000 ;
	    RECT 477.2000 247.6000 478.0000 248.4000 ;
	    RECT 479.6000 242.2000 480.4000 250.8000 ;
	    RECT 486.2000 250.4000 486.8000 251.6000 ;
	    RECT 492.4000 251.0000 498.0000 251.2000 ;
	    RECT 492.2000 250.8000 498.0000 251.0000 ;
	    RECT 484.4000 249.8000 486.8000 250.4000 ;
	    RECT 488.2000 250.6000 498.0000 250.8000 ;
	    RECT 488.2000 250.2000 493.0000 250.6000 ;
	    RECT 484.4000 248.8000 485.0000 249.8000 ;
	    RECT 483.6000 248.0000 485.0000 248.8000 ;
	    RECT 486.6000 249.0000 487.4000 249.2000 ;
	    RECT 488.2000 249.0000 488.8000 250.2000 ;
	    RECT 486.6000 248.4000 488.8000 249.0000 ;
	    RECT 489.4000 249.0000 494.8000 249.6000 ;
	    RECT 489.4000 248.8000 490.2000 249.0000 ;
	    RECT 494.0000 248.8000 494.8000 249.0000 ;
	    RECT 487.8000 247.4000 488.6000 247.6000 ;
	    RECT 490.6000 247.4000 491.4000 247.6000 ;
	    RECT 484.4000 246.2000 485.2000 247.0000 ;
	    RECT 487.8000 246.8000 491.4000 247.4000 ;
	    RECT 488.6000 246.2000 489.2000 246.8000 ;
	    RECT 494.0000 246.2000 494.8000 247.0000 ;
	    RECT 483.8000 242.2000 485.0000 246.2000 ;
	    RECT 488.4000 242.2000 489.2000 246.2000 ;
	    RECT 492.8000 245.6000 494.8000 246.2000 ;
	    RECT 492.8000 242.2000 493.6000 245.6000 ;
	    RECT 497.2000 242.2000 498.0000 250.6000 ;
	    RECT 499.0000 250.4000 499.6000 253.6000 ;
	    RECT 501.2000 251.6000 502.8000 252.4000 ;
	    RECT 498.8000 249.6000 499.6000 250.4000 ;
	    RECT 505.2000 250.2000 506.0000 250.4000 ;
	    RECT 507.2000 250.2000 507.8000 253.6000 ;
	    RECT 508.4000 252.3000 509.2000 253.2000 ;
	    RECT 510.0000 252.3000 510.8000 252.4000 ;
	    RECT 508.4000 251.7000 510.8000 252.3000 ;
	    RECT 508.4000 251.6000 509.2000 251.7000 ;
	    RECT 510.0000 251.6000 510.8000 251.7000 ;
	    RECT 505.2000 249.6000 506.6000 250.2000 ;
	    RECT 507.2000 249.6000 508.2000 250.2000 ;
	    RECT 499.0000 247.0000 499.6000 249.6000 ;
	    RECT 500.4000 247.6000 501.2000 249.2000 ;
	    RECT 506.0000 248.4000 506.6000 249.6000 ;
	    RECT 506.0000 247.6000 506.8000 248.4000 ;
	    RECT 499.0000 246.4000 502.6000 247.0000 ;
	    RECT 499.0000 246.2000 499.6000 246.4000 ;
	    RECT 498.8000 242.2000 499.6000 246.2000 ;
	    RECT 502.0000 242.2000 502.8000 246.4000 ;
	    RECT 507.4000 242.2000 508.2000 249.6000 ;
	    RECT 511.6000 242.2000 512.4000 253.7000 ;
	    RECT 4.4000 232.4000 5.2000 239.8000 ;
	    RECT 9.2000 232.4000 10.0000 239.8000 ;
	    RECT 13.4000 238.4000 14.2000 239.8000 ;
	    RECT 12.4000 237.6000 14.2000 238.4000 ;
	    RECT 3.0000 231.8000 5.2000 232.4000 ;
	    RECT 7.8000 231.8000 10.0000 232.4000 ;
	    RECT 13.4000 232.4000 14.2000 237.6000 ;
	    RECT 19.8000 234.4000 20.6000 239.8000 ;
	    RECT 14.8000 233.6000 16.4000 234.4000 ;
	    RECT 18.8000 233.6000 20.6000 234.4000 ;
	    RECT 21.2000 234.3000 22.0000 234.4000 ;
	    RECT 23.6000 234.3000 24.4000 239.8000 ;
	    RECT 27.8000 235.8000 29.0000 239.8000 ;
	    RECT 32.4000 235.8000 33.2000 239.8000 ;
	    RECT 36.8000 236.4000 37.6000 239.8000 ;
	    RECT 36.8000 235.8000 38.8000 236.4000 ;
	    RECT 28.4000 235.0000 29.2000 235.8000 ;
	    RECT 32.6000 235.2000 33.2000 235.8000 ;
	    RECT 31.8000 234.6000 35.4000 235.2000 ;
	    RECT 38.0000 235.0000 38.8000 235.8000 ;
	    RECT 31.8000 234.4000 32.6000 234.6000 ;
	    RECT 34.6000 234.4000 35.4000 234.6000 ;
	    RECT 21.2000 233.7000 24.4000 234.3000 ;
	    RECT 21.2000 233.6000 22.0000 233.7000 ;
	    RECT 15.0000 232.4000 15.6000 233.6000 ;
	    RECT 19.8000 232.4000 20.6000 233.6000 ;
	    RECT 21.4000 232.4000 22.0000 233.6000 ;
	    RECT 13.4000 231.8000 14.4000 232.4000 ;
	    RECT 15.0000 231.8000 16.4000 232.4000 ;
	    RECT 19.8000 231.8000 20.8000 232.4000 ;
	    RECT 21.4000 231.8000 22.8000 232.4000 ;
	    RECT 3.0000 231.2000 3.6000 231.8000 ;
	    RECT 7.8000 231.2000 8.4000 231.8000 ;
	    RECT 2.4000 230.4000 3.6000 231.2000 ;
	    RECT 7.2000 230.4000 8.4000 231.2000 ;
	    RECT 3.0000 227.4000 3.6000 230.4000 ;
	    RECT 4.4000 228.8000 5.2000 230.4000 ;
	    RECT 7.8000 227.4000 8.4000 230.4000 ;
	    RECT 9.2000 230.3000 10.0000 230.4000 ;
	    RECT 10.8000 230.3000 11.6000 230.4000 ;
	    RECT 9.2000 229.7000 11.6000 230.3000 ;
	    RECT 9.2000 228.8000 10.0000 229.7000 ;
	    RECT 10.8000 229.6000 11.6000 229.7000 ;
	    RECT 12.4000 228.8000 13.2000 230.4000 ;
	    RECT 13.8000 228.4000 14.4000 231.8000 ;
	    RECT 15.6000 231.6000 16.4000 231.8000 ;
	    RECT 18.8000 228.8000 19.6000 230.4000 ;
	    RECT 20.2000 228.4000 20.8000 231.8000 ;
	    RECT 22.0000 231.6000 22.8000 231.8000 ;
	    RECT 23.6000 231.2000 24.4000 233.7000 ;
	    RECT 27.6000 233.2000 29.0000 234.0000 ;
	    RECT 28.4000 232.2000 29.0000 233.2000 ;
	    RECT 30.6000 233.0000 32.8000 233.6000 ;
	    RECT 30.6000 232.8000 31.4000 233.0000 ;
	    RECT 28.4000 231.6000 30.8000 232.2000 ;
	    RECT 23.6000 230.6000 27.8000 231.2000 ;
	    RECT 10.8000 228.2000 11.6000 228.4000 ;
	    RECT 10.8000 227.6000 12.4000 228.2000 ;
	    RECT 13.8000 227.6000 16.4000 228.4000 ;
	    RECT 17.2000 228.2000 18.0000 228.4000 ;
	    RECT 17.2000 227.6000 18.8000 228.2000 ;
	    RECT 20.2000 227.6000 22.8000 228.4000 ;
	    RECT 3.0000 226.8000 5.2000 227.4000 ;
	    RECT 7.8000 226.8000 10.0000 227.4000 ;
	    RECT 11.6000 227.2000 12.4000 227.6000 ;
	    RECT 4.4000 222.2000 5.2000 226.8000 ;
	    RECT 9.2000 222.2000 10.0000 226.8000 ;
	    RECT 11.0000 226.2000 14.6000 226.6000 ;
	    RECT 15.6000 226.2000 16.2000 227.6000 ;
	    RECT 18.0000 227.2000 18.8000 227.6000 ;
	    RECT 17.4000 226.2000 21.0000 226.6000 ;
	    RECT 22.0000 226.2000 22.6000 227.6000 ;
	    RECT 23.6000 227.2000 24.4000 230.6000 ;
	    RECT 27.0000 230.4000 27.8000 230.6000 ;
	    RECT 30.2000 230.3000 30.8000 231.6000 ;
	    RECT 32.2000 231.8000 32.8000 233.0000 ;
	    RECT 33.4000 233.0000 34.2000 233.2000 ;
	    RECT 38.0000 233.0000 38.8000 233.2000 ;
	    RECT 33.4000 232.4000 38.8000 233.0000 ;
	    RECT 32.2000 231.4000 37.0000 231.8000 ;
	    RECT 41.2000 231.4000 42.0000 239.8000 ;
	    RECT 45.4000 232.4000 46.2000 239.8000 ;
	    RECT 46.8000 233.6000 47.6000 234.4000 ;
	    RECT 47.0000 232.4000 47.6000 233.6000 ;
	    RECT 50.0000 233.6000 50.8000 234.4000 ;
	    RECT 50.0000 232.4000 50.6000 233.6000 ;
	    RECT 51.4000 232.4000 52.2000 239.8000 ;
	    RECT 56.4000 233.6000 57.2000 234.4000 ;
	    RECT 56.4000 232.4000 57.0000 233.6000 ;
	    RECT 57.8000 232.4000 58.6000 239.8000 ;
	    RECT 45.4000 231.8000 46.4000 232.4000 ;
	    RECT 47.0000 231.8000 48.4000 232.4000 ;
	    RECT 32.2000 231.2000 42.0000 231.4000 ;
	    RECT 36.2000 231.0000 42.0000 231.2000 ;
	    RECT 36.4000 230.8000 42.0000 231.0000 ;
	    RECT 31.6000 230.3000 32.4000 230.4000 ;
	    RECT 25.4000 229.8000 26.2000 230.0000 ;
	    RECT 25.4000 229.2000 29.2000 229.8000 ;
	    RECT 30.1000 229.7000 32.4000 230.3000 ;
	    RECT 28.4000 229.0000 29.2000 229.2000 ;
	    RECT 30.2000 228.4000 30.8000 229.7000 ;
	    RECT 31.6000 229.6000 32.4000 229.7000 ;
	    RECT 34.8000 230.2000 35.6000 230.4000 ;
	    RECT 34.8000 229.6000 39.8000 230.2000 ;
	    RECT 36.4000 229.4000 37.2000 229.6000 ;
	    RECT 39.0000 229.4000 39.8000 229.6000 ;
	    RECT 44.4000 228.8000 45.2000 230.4000 ;
	    RECT 37.4000 228.4000 38.2000 228.6000 ;
	    RECT 45.8000 228.4000 46.4000 231.8000 ;
	    RECT 47.6000 231.6000 48.4000 231.8000 ;
	    RECT 49.2000 231.8000 50.6000 232.4000 ;
	    RECT 51.2000 231.8000 52.2000 232.4000 ;
	    RECT 55.6000 231.8000 57.0000 232.4000 ;
	    RECT 57.6000 231.8000 58.6000 232.4000 ;
	    RECT 49.2000 231.6000 50.0000 231.8000 ;
	    RECT 47.6000 230.3000 48.4000 230.4000 ;
	    RECT 51.2000 230.3000 51.8000 231.8000 ;
	    RECT 55.6000 231.6000 56.4000 231.8000 ;
	    RECT 47.6000 229.7000 51.8000 230.3000 ;
	    RECT 47.6000 229.6000 48.4000 229.7000 ;
	    RECT 51.2000 228.4000 51.8000 229.7000 ;
	    RECT 52.4000 230.3000 53.2000 230.4000 ;
	    RECT 57.6000 230.3000 58.2000 231.8000 ;
	    RECT 62.0000 231.2000 62.8000 239.8000 ;
	    RECT 66.2000 235.8000 67.4000 239.8000 ;
	    RECT 70.8000 235.8000 71.6000 239.8000 ;
	    RECT 75.2000 236.4000 76.0000 239.8000 ;
	    RECT 75.2000 235.8000 77.2000 236.4000 ;
	    RECT 66.8000 235.0000 67.6000 235.8000 ;
	    RECT 71.0000 235.2000 71.6000 235.8000 ;
	    RECT 70.2000 234.6000 73.8000 235.2000 ;
	    RECT 76.4000 235.0000 77.2000 235.8000 ;
	    RECT 70.2000 234.4000 71.0000 234.6000 ;
	    RECT 73.0000 234.4000 73.8000 234.6000 ;
	    RECT 66.0000 233.2000 67.4000 234.0000 ;
	    RECT 66.8000 232.2000 67.4000 233.2000 ;
	    RECT 69.0000 233.0000 71.2000 233.6000 ;
	    RECT 69.0000 232.8000 69.8000 233.0000 ;
	    RECT 66.8000 231.6000 69.2000 232.2000 ;
	    RECT 62.0000 230.6000 66.2000 231.2000 ;
	    RECT 52.4000 229.7000 58.2000 230.3000 ;
	    RECT 52.4000 228.8000 53.2000 229.7000 ;
	    RECT 57.6000 228.4000 58.2000 229.7000 ;
	    RECT 58.8000 230.3000 59.6000 230.4000 ;
	    RECT 60.4000 230.3000 61.2000 230.4000 ;
	    RECT 58.8000 229.7000 61.2000 230.3000 ;
	    RECT 58.8000 228.8000 59.6000 229.7000 ;
	    RECT 60.4000 229.6000 61.2000 229.7000 ;
	    RECT 30.0000 227.8000 41.2000 228.4000 ;
	    RECT 30.0000 227.6000 31.4000 227.8000 ;
	    RECT 23.6000 226.6000 27.4000 227.2000 ;
	    RECT 10.8000 226.0000 14.8000 226.2000 ;
	    RECT 10.8000 222.2000 11.6000 226.0000 ;
	    RECT 14.0000 222.2000 14.8000 226.0000 ;
	    RECT 15.6000 222.2000 16.4000 226.2000 ;
	    RECT 17.2000 226.0000 21.2000 226.2000 ;
	    RECT 17.2000 222.2000 18.0000 226.0000 ;
	    RECT 20.4000 222.2000 21.2000 226.0000 ;
	    RECT 22.0000 222.2000 22.8000 226.2000 ;
	    RECT 23.6000 222.2000 24.4000 226.6000 ;
	    RECT 26.6000 226.4000 27.4000 226.6000 ;
	    RECT 36.4000 225.6000 37.0000 227.8000 ;
	    RECT 39.6000 227.6000 41.2000 227.8000 ;
	    RECT 42.8000 228.2000 43.6000 228.4000 ;
	    RECT 42.8000 227.6000 44.4000 228.2000 ;
	    RECT 45.8000 227.6000 48.4000 228.4000 ;
	    RECT 49.2000 227.6000 51.8000 228.4000 ;
	    RECT 54.0000 228.2000 54.8000 228.4000 ;
	    RECT 53.2000 227.6000 54.8000 228.2000 ;
	    RECT 55.6000 227.6000 58.2000 228.4000 ;
	    RECT 60.4000 228.2000 61.2000 228.4000 ;
	    RECT 59.6000 227.6000 61.2000 228.2000 ;
	    RECT 43.6000 227.2000 44.4000 227.6000 ;
	    RECT 34.6000 225.4000 35.4000 225.6000 ;
	    RECT 28.4000 224.2000 29.2000 225.0000 ;
	    RECT 32.6000 224.8000 35.4000 225.4000 ;
	    RECT 36.4000 224.8000 37.2000 225.6000 ;
	    RECT 32.6000 224.2000 33.2000 224.8000 ;
	    RECT 38.0000 224.2000 38.8000 225.0000 ;
	    RECT 27.8000 223.6000 29.2000 224.2000 ;
	    RECT 27.8000 222.2000 29.0000 223.6000 ;
	    RECT 32.4000 222.2000 33.2000 224.2000 ;
	    RECT 36.8000 223.6000 38.8000 224.2000 ;
	    RECT 36.8000 222.2000 37.6000 223.6000 ;
	    RECT 41.2000 222.2000 42.0000 227.0000 ;
	    RECT 43.0000 226.2000 46.6000 226.6000 ;
	    RECT 47.6000 226.2000 48.2000 227.6000 ;
	    RECT 49.4000 226.2000 50.0000 227.6000 ;
	    RECT 53.2000 227.2000 54.0000 227.6000 ;
	    RECT 51.0000 226.2000 54.6000 226.6000 ;
	    RECT 55.8000 226.2000 56.4000 227.6000 ;
	    RECT 59.6000 227.2000 60.4000 227.6000 ;
	    RECT 62.0000 227.2000 62.8000 230.6000 ;
	    RECT 65.4000 230.4000 66.2000 230.6000 ;
	    RECT 68.6000 230.4000 69.2000 231.6000 ;
	    RECT 70.6000 231.8000 71.2000 233.0000 ;
	    RECT 71.8000 233.0000 72.6000 233.2000 ;
	    RECT 76.4000 233.0000 77.2000 233.2000 ;
	    RECT 71.8000 232.4000 77.2000 233.0000 ;
	    RECT 70.6000 231.4000 75.4000 231.8000 ;
	    RECT 79.6000 231.4000 80.4000 239.8000 ;
	    RECT 82.0000 233.6000 82.8000 234.4000 ;
	    RECT 82.0000 232.4000 82.6000 233.6000 ;
	    RECT 83.4000 232.4000 84.2000 239.8000 ;
	    RECT 88.4000 233.6000 89.2000 234.4000 ;
	    RECT 88.4000 232.4000 89.0000 233.6000 ;
	    RECT 89.8000 232.4000 90.6000 239.8000 ;
	    RECT 94.8000 233.6000 95.6000 234.4000 ;
	    RECT 94.8000 232.4000 95.4000 233.6000 ;
	    RECT 96.2000 232.4000 97.0000 239.8000 ;
	    RECT 81.2000 231.8000 82.6000 232.4000 ;
	    RECT 83.2000 231.8000 84.2000 232.4000 ;
	    RECT 87.6000 231.8000 89.0000 232.4000 ;
	    RECT 89.6000 231.8000 90.6000 232.4000 ;
	    RECT 94.0000 231.8000 95.4000 232.4000 ;
	    RECT 96.0000 231.8000 97.0000 232.4000 ;
	    RECT 81.2000 231.6000 82.0000 231.8000 ;
	    RECT 70.6000 231.2000 80.4000 231.4000 ;
	    RECT 74.6000 231.0000 80.4000 231.2000 ;
	    RECT 74.8000 230.8000 80.4000 231.0000 ;
	    RECT 83.2000 230.4000 83.8000 231.8000 ;
	    RECT 87.6000 231.6000 88.4000 231.8000 ;
	    RECT 63.8000 229.8000 64.6000 230.0000 ;
	    RECT 63.8000 229.2000 67.6000 229.8000 ;
	    RECT 68.4000 229.6000 69.2000 230.4000 ;
	    RECT 73.2000 230.2000 74.0000 230.4000 ;
	    RECT 73.2000 229.6000 78.2000 230.2000 ;
	    RECT 82.8000 229.6000 83.8000 230.4000 ;
	    RECT 66.8000 229.0000 67.6000 229.2000 ;
	    RECT 68.6000 228.4000 69.2000 229.6000 ;
	    RECT 74.8000 229.4000 75.6000 229.6000 ;
	    RECT 77.4000 229.4000 78.2000 229.6000 ;
	    RECT 75.8000 228.4000 76.6000 228.6000 ;
	    RECT 83.2000 228.4000 83.8000 229.6000 ;
	    RECT 84.4000 230.3000 85.2000 230.4000 ;
	    RECT 89.6000 230.3000 90.2000 231.8000 ;
	    RECT 94.0000 231.6000 94.8000 231.8000 ;
	    RECT 96.0000 230.4000 96.6000 231.8000 ;
	    RECT 106.8000 231.4000 107.6000 239.8000 ;
	    RECT 111.2000 236.4000 112.0000 239.8000 ;
	    RECT 110.0000 235.8000 112.0000 236.4000 ;
	    RECT 115.6000 235.8000 116.4000 239.8000 ;
	    RECT 119.8000 235.8000 121.0000 239.8000 ;
	    RECT 110.0000 235.0000 110.8000 235.8000 ;
	    RECT 115.6000 235.2000 116.2000 235.8000 ;
	    RECT 113.4000 234.6000 117.0000 235.2000 ;
	    RECT 119.6000 235.0000 120.4000 235.8000 ;
	    RECT 113.4000 234.4000 114.2000 234.6000 ;
	    RECT 116.2000 234.4000 117.0000 234.6000 ;
	    RECT 110.0000 233.0000 110.8000 233.2000 ;
	    RECT 114.6000 233.0000 115.4000 233.2000 ;
	    RECT 110.0000 232.4000 115.4000 233.0000 ;
	    RECT 116.0000 233.0000 118.2000 233.6000 ;
	    RECT 116.0000 231.8000 116.6000 233.0000 ;
	    RECT 117.4000 232.8000 118.2000 233.0000 ;
	    RECT 119.8000 233.2000 121.2000 234.0000 ;
	    RECT 119.8000 232.2000 120.4000 233.2000 ;
	    RECT 111.8000 231.4000 116.6000 231.8000 ;
	    RECT 106.8000 231.2000 116.6000 231.4000 ;
	    RECT 118.0000 231.6000 120.4000 232.2000 ;
	    RECT 106.8000 231.0000 112.6000 231.2000 ;
	    RECT 106.8000 230.8000 112.4000 231.0000 ;
	    RECT 84.4000 229.7000 90.2000 230.3000 ;
	    RECT 84.4000 228.8000 85.2000 229.7000 ;
	    RECT 89.6000 228.4000 90.2000 229.7000 ;
	    RECT 90.8000 228.8000 91.6000 230.4000 ;
	    RECT 95.6000 229.6000 96.6000 230.4000 ;
	    RECT 96.0000 228.4000 96.6000 229.6000 ;
	    RECT 97.2000 228.8000 98.0000 230.4000 ;
	    RECT 113.2000 230.2000 114.0000 230.4000 ;
	    RECT 109.0000 229.6000 114.0000 230.2000 ;
	    RECT 109.0000 229.4000 109.8000 229.6000 ;
	    RECT 111.6000 229.4000 112.4000 229.6000 ;
	    RECT 110.6000 228.4000 111.4000 228.6000 ;
	    RECT 118.0000 228.4000 118.6000 231.6000 ;
	    RECT 124.4000 231.2000 125.2000 239.8000 ;
	    RECT 128.6000 231.8000 130.6000 239.8000 ;
	    RECT 134.8000 233.6000 135.6000 234.4000 ;
	    RECT 134.8000 232.4000 135.4000 233.6000 ;
	    RECT 136.2000 232.4000 137.0000 239.8000 ;
	    RECT 143.0000 238.4000 143.8000 239.8000 ;
	    RECT 142.0000 237.6000 143.8000 238.4000 ;
	    RECT 134.0000 231.8000 135.4000 232.4000 ;
	    RECT 136.0000 231.8000 137.0000 232.4000 ;
	    RECT 143.0000 232.4000 143.8000 237.6000 ;
	    RECT 144.4000 233.6000 145.2000 234.4000 ;
	    RECT 144.6000 232.4000 145.2000 233.6000 ;
	    RECT 147.4000 232.6000 148.2000 239.8000 ;
	    RECT 154.2000 238.4000 155.0000 239.8000 ;
	    RECT 153.2000 237.6000 155.0000 238.4000 ;
	    RECT 154.2000 232.6000 155.0000 237.6000 ;
	    RECT 160.2000 232.8000 161.0000 239.8000 ;
	    RECT 164.4000 235.0000 165.2000 239.0000 ;
	    RECT 143.0000 231.8000 144.0000 232.4000 ;
	    RECT 144.6000 231.8000 146.0000 232.4000 ;
	    RECT 147.4000 231.8000 149.2000 232.6000 ;
	    RECT 153.2000 231.8000 155.0000 232.6000 ;
	    RECT 159.4000 232.2000 161.0000 232.8000 ;
	    RECT 121.0000 230.6000 125.2000 231.2000 ;
	    RECT 121.0000 230.4000 121.8000 230.6000 ;
	    RECT 122.6000 229.8000 123.4000 230.0000 ;
	    RECT 119.6000 229.2000 123.4000 229.8000 ;
	    RECT 119.6000 229.0000 120.4000 229.2000 ;
	    RECT 68.6000 227.8000 79.6000 228.4000 ;
	    RECT 69.0000 227.6000 69.8000 227.8000 ;
	    RECT 62.0000 226.6000 65.8000 227.2000 ;
	    RECT 57.4000 226.2000 61.0000 226.6000 ;
	    RECT 42.8000 226.0000 46.8000 226.2000 ;
	    RECT 42.8000 222.2000 43.6000 226.0000 ;
	    RECT 46.0000 222.2000 46.8000 226.0000 ;
	    RECT 47.6000 222.2000 48.4000 226.2000 ;
	    RECT 49.2000 222.2000 50.0000 226.2000 ;
	    RECT 50.8000 226.0000 54.8000 226.2000 ;
	    RECT 50.8000 222.2000 51.6000 226.0000 ;
	    RECT 54.0000 222.2000 54.8000 226.0000 ;
	    RECT 55.6000 222.2000 56.4000 226.2000 ;
	    RECT 57.2000 226.0000 61.2000 226.2000 ;
	    RECT 57.2000 222.2000 58.0000 226.0000 ;
	    RECT 60.4000 222.2000 61.2000 226.0000 ;
	    RECT 62.0000 222.2000 62.8000 226.6000 ;
	    RECT 65.0000 226.4000 65.8000 226.6000 ;
	    RECT 74.8000 225.6000 75.4000 227.8000 ;
	    RECT 78.0000 227.6000 79.6000 227.8000 ;
	    RECT 81.2000 227.6000 83.8000 228.4000 ;
	    RECT 86.0000 228.2000 86.8000 228.4000 ;
	    RECT 85.2000 227.6000 86.8000 228.2000 ;
	    RECT 87.6000 227.6000 90.2000 228.4000 ;
	    RECT 92.4000 228.2000 93.2000 228.4000 ;
	    RECT 91.6000 227.6000 93.2000 228.2000 ;
	    RECT 94.0000 227.6000 96.6000 228.4000 ;
	    RECT 98.8000 228.2000 99.6000 228.4000 ;
	    RECT 98.0000 227.6000 99.6000 228.2000 ;
	    RECT 107.6000 227.8000 118.6000 228.4000 ;
	    RECT 107.6000 227.6000 109.2000 227.8000 ;
	    RECT 73.0000 225.4000 73.8000 225.6000 ;
	    RECT 66.8000 224.2000 67.6000 225.0000 ;
	    RECT 71.0000 224.8000 73.8000 225.4000 ;
	    RECT 74.8000 224.8000 75.6000 225.6000 ;
	    RECT 71.0000 224.2000 71.6000 224.8000 ;
	    RECT 76.4000 224.2000 77.2000 225.0000 ;
	    RECT 66.2000 223.6000 67.6000 224.2000 ;
	    RECT 66.2000 222.2000 67.4000 223.6000 ;
	    RECT 70.8000 222.2000 71.6000 224.2000 ;
	    RECT 75.2000 223.6000 77.2000 224.2000 ;
	    RECT 75.2000 222.2000 76.0000 223.6000 ;
	    RECT 79.6000 222.2000 80.4000 227.0000 ;
	    RECT 81.4000 226.2000 82.0000 227.6000 ;
	    RECT 85.2000 227.2000 86.0000 227.6000 ;
	    RECT 83.0000 226.2000 86.6000 226.6000 ;
	    RECT 87.8000 226.2000 88.4000 227.6000 ;
	    RECT 91.6000 227.2000 92.4000 227.6000 ;
	    RECT 89.4000 226.2000 93.0000 226.6000 ;
	    RECT 94.2000 226.2000 94.8000 227.6000 ;
	    RECT 98.0000 227.2000 98.8000 227.6000 ;
	    RECT 95.8000 226.2000 99.4000 226.6000 ;
	    RECT 81.2000 222.2000 82.0000 226.2000 ;
	    RECT 82.8000 226.0000 86.8000 226.2000 ;
	    RECT 82.8000 222.2000 83.6000 226.0000 ;
	    RECT 86.0000 222.2000 86.8000 226.0000 ;
	    RECT 87.6000 222.2000 88.4000 226.2000 ;
	    RECT 89.2000 226.0000 93.2000 226.2000 ;
	    RECT 89.2000 222.2000 90.0000 226.0000 ;
	    RECT 92.4000 222.2000 93.2000 226.0000 ;
	    RECT 94.0000 222.2000 94.8000 226.2000 ;
	    RECT 95.6000 226.0000 99.6000 226.2000 ;
	    RECT 95.6000 222.2000 96.4000 226.0000 ;
	    RECT 98.8000 222.2000 99.6000 226.0000 ;
	    RECT 106.8000 222.2000 107.6000 227.0000 ;
	    RECT 111.8000 226.4000 112.4000 227.8000 ;
	    RECT 117.4000 227.6000 118.2000 227.8000 ;
	    RECT 124.4000 227.2000 125.2000 230.6000 ;
	    RECT 126.0000 227.6000 126.8000 229.2000 ;
	    RECT 127.6000 228.8000 128.4000 230.4000 ;
	    RECT 129.4000 228.4000 130.0000 231.8000 ;
	    RECT 134.0000 231.6000 134.8000 231.8000 ;
	    RECT 130.8000 228.8000 131.6000 230.4000 ;
	    RECT 136.0000 228.4000 136.6000 231.8000 ;
	    RECT 137.2000 230.3000 138.0000 230.4000 ;
	    RECT 137.2000 229.7000 141.1000 230.3000 ;
	    RECT 137.2000 228.8000 138.0000 229.7000 ;
	    RECT 140.5000 228.4000 141.1000 229.7000 ;
	    RECT 142.0000 228.8000 142.8000 230.4000 ;
	    RECT 143.4000 228.4000 144.0000 231.8000 ;
	    RECT 145.2000 231.6000 146.0000 231.8000 ;
	    RECT 146.8000 229.6000 147.6000 231.2000 ;
	    RECT 148.4000 228.4000 149.0000 231.8000 ;
	    RECT 153.4000 228.4000 154.0000 231.8000 ;
	    RECT 154.8000 229.6000 155.6000 231.2000 ;
	    RECT 158.0000 229.6000 158.8000 231.2000 ;
	    RECT 159.4000 230.4000 160.0000 232.2000 ;
	    RECT 164.6000 231.6000 165.2000 235.0000 ;
	    RECT 168.6000 231.8000 170.6000 239.8000 ;
	    RECT 176.6000 232.6000 177.4000 239.8000 ;
	    RECT 175.6000 231.8000 177.4000 232.6000 ;
	    RECT 179.6000 233.6000 180.4000 234.4000 ;
	    RECT 179.6000 232.4000 180.2000 233.6000 ;
	    RECT 181.0000 232.4000 181.8000 239.8000 ;
	    RECT 178.8000 231.8000 180.2000 232.4000 ;
	    RECT 180.8000 231.8000 181.8000 232.4000 ;
	    RECT 161.4000 231.0000 165.2000 231.6000 ;
	    RECT 159.4000 229.6000 160.4000 230.4000 ;
	    RECT 159.4000 228.4000 160.0000 229.6000 ;
	    RECT 161.4000 229.0000 162.0000 231.0000 ;
	    RECT 129.2000 228.2000 130.0000 228.4000 ;
	    RECT 132.4000 228.3000 133.2000 228.4000 ;
	    RECT 134.0000 228.3000 136.6000 228.4000 ;
	    RECT 132.4000 228.2000 136.6000 228.3000 ;
	    RECT 138.8000 228.2000 139.6000 228.4000 ;
	    RECT 127.6000 227.6000 130.0000 228.2000 ;
	    RECT 131.6000 227.7000 136.6000 228.2000 ;
	    RECT 131.6000 227.6000 133.2000 227.7000 ;
	    RECT 134.0000 227.6000 136.6000 227.7000 ;
	    RECT 138.0000 227.6000 139.6000 228.2000 ;
	    RECT 140.4000 228.2000 141.2000 228.4000 ;
	    RECT 140.4000 227.6000 142.0000 228.2000 ;
	    RECT 143.4000 227.6000 146.0000 228.4000 ;
	    RECT 148.4000 227.6000 149.2000 228.4000 ;
	    RECT 151.6000 228.3000 152.4000 228.4000 ;
	    RECT 150.1000 227.7000 152.4000 228.3000 ;
	    RECT 121.4000 226.6000 125.2000 227.2000 ;
	    RECT 121.4000 226.4000 122.2000 226.6000 ;
	    RECT 110.0000 224.2000 110.8000 225.0000 ;
	    RECT 111.6000 224.8000 112.4000 226.4000 ;
	    RECT 113.4000 225.4000 114.2000 225.6000 ;
	    RECT 113.4000 224.8000 116.2000 225.4000 ;
	    RECT 115.6000 224.2000 116.2000 224.8000 ;
	    RECT 119.6000 224.2000 120.4000 225.0000 ;
	    RECT 110.0000 223.6000 112.0000 224.2000 ;
	    RECT 111.2000 222.2000 112.0000 223.6000 ;
	    RECT 115.6000 222.2000 116.4000 224.2000 ;
	    RECT 119.6000 223.6000 121.0000 224.2000 ;
	    RECT 119.8000 222.2000 121.0000 223.6000 ;
	    RECT 124.4000 222.2000 125.2000 226.6000 ;
	    RECT 127.6000 226.2000 128.2000 227.6000 ;
	    RECT 131.6000 227.2000 132.4000 227.6000 ;
	    RECT 129.4000 226.2000 133.0000 226.6000 ;
	    RECT 134.2000 226.2000 134.8000 227.6000 ;
	    RECT 138.0000 227.2000 138.8000 227.6000 ;
	    RECT 141.2000 227.2000 142.0000 227.6000 ;
	    RECT 135.8000 226.2000 139.4000 226.6000 ;
	    RECT 140.6000 226.2000 144.2000 226.6000 ;
	    RECT 145.2000 226.2000 145.8000 227.6000 ;
	    RECT 146.8000 226.3000 147.6000 226.4000 ;
	    RECT 148.4000 226.3000 149.0000 227.6000 ;
	    RECT 150.1000 226.4000 150.7000 227.7000 ;
	    RECT 151.6000 227.6000 152.4000 227.7000 ;
	    RECT 153.2000 227.6000 154.0000 228.4000 ;
	    RECT 158.0000 227.6000 160.0000 228.4000 ;
	    RECT 160.6000 228.2000 162.0000 229.0000 ;
	    RECT 162.8000 228.8000 163.6000 230.4000 ;
	    RECT 164.4000 228.8000 165.2000 230.4000 ;
	    RECT 126.0000 222.8000 126.8000 226.2000 ;
	    RECT 127.6000 223.4000 128.4000 226.2000 ;
	    RECT 129.2000 226.0000 133.2000 226.2000 ;
	    RECT 129.2000 222.8000 130.0000 226.0000 ;
	    RECT 126.0000 222.2000 130.0000 222.8000 ;
	    RECT 132.4000 222.2000 133.2000 226.0000 ;
	    RECT 134.0000 222.2000 134.8000 226.2000 ;
	    RECT 135.6000 226.0000 139.6000 226.2000 ;
	    RECT 135.6000 222.2000 136.4000 226.0000 ;
	    RECT 138.8000 222.2000 139.6000 226.0000 ;
	    RECT 140.4000 226.0000 144.4000 226.2000 ;
	    RECT 140.4000 222.2000 141.2000 226.0000 ;
	    RECT 143.6000 222.2000 144.4000 226.0000 ;
	    RECT 145.2000 222.2000 146.0000 226.2000 ;
	    RECT 146.8000 225.7000 149.1000 226.3000 ;
	    RECT 146.8000 225.6000 147.6000 225.7000 ;
	    RECT 148.4000 224.2000 149.0000 225.7000 ;
	    RECT 150.0000 224.8000 150.8000 226.4000 ;
	    RECT 151.6000 224.8000 152.4000 226.4000 ;
	    RECT 153.4000 224.2000 154.0000 227.6000 ;
	    RECT 159.4000 227.0000 160.0000 227.6000 ;
	    RECT 161.0000 227.8000 162.0000 228.2000 ;
	    RECT 161.0000 227.2000 165.2000 227.8000 ;
	    RECT 166.0000 227.6000 166.8000 229.2000 ;
	    RECT 167.6000 228.8000 168.4000 230.4000 ;
	    RECT 169.4000 228.4000 170.0000 231.8000 ;
	    RECT 170.8000 230.3000 171.6000 230.4000 ;
	    RECT 175.8000 230.3000 176.4000 231.8000 ;
	    RECT 178.8000 231.6000 179.6000 231.8000 ;
	    RECT 170.8000 229.7000 176.4000 230.3000 ;
	    RECT 170.8000 228.8000 171.6000 229.7000 ;
	    RECT 175.8000 228.4000 176.4000 229.7000 ;
	    RECT 177.2000 229.6000 178.0000 231.2000 ;
	    RECT 180.8000 230.4000 181.4000 231.8000 ;
	    RECT 180.4000 229.6000 181.4000 230.4000 ;
	    RECT 180.8000 228.4000 181.4000 229.6000 ;
	    RECT 182.0000 228.8000 182.8000 230.4000 ;
	    RECT 186.8000 230.3000 187.6000 239.8000 ;
	    RECT 192.2000 236.4000 193.0000 239.8000 ;
	    RECT 192.2000 235.6000 194.0000 236.4000 ;
	    RECT 190.8000 233.6000 191.6000 234.4000 ;
	    RECT 188.4000 231.6000 189.2000 233.2000 ;
	    RECT 190.8000 232.4000 191.4000 233.6000 ;
	    RECT 192.2000 232.4000 193.0000 235.6000 ;
	    RECT 190.0000 231.8000 191.4000 232.4000 ;
	    RECT 192.0000 231.8000 193.0000 232.4000 ;
	    RECT 196.4000 231.8000 197.2000 239.8000 ;
	    RECT 199.6000 232.4000 200.4000 239.8000 ;
	    RECT 198.2000 231.8000 200.4000 232.4000 ;
	    RECT 201.8000 232.6000 202.6000 239.8000 ;
	    RECT 201.8000 231.8000 203.6000 232.6000 ;
	    RECT 208.6000 231.8000 210.6000 239.8000 ;
	    RECT 214.8000 233.6000 215.6000 234.4000 ;
	    RECT 214.8000 232.4000 215.4000 233.6000 ;
	    RECT 216.2000 232.4000 217.0000 239.8000 ;
	    RECT 214.0000 231.8000 215.4000 232.4000 ;
	    RECT 216.0000 231.8000 217.0000 232.4000 ;
	    RECT 223.0000 231.8000 225.0000 239.8000 ;
	    RECT 229.2000 233.6000 230.0000 234.4000 ;
	    RECT 229.2000 232.4000 229.8000 233.6000 ;
	    RECT 230.6000 232.4000 231.4000 239.8000 ;
	    RECT 237.4000 232.6000 238.2000 239.8000 ;
	    RECT 228.4000 231.8000 229.8000 232.4000 ;
	    RECT 230.4000 231.8000 231.4000 232.4000 ;
	    RECT 236.4000 231.8000 238.2000 232.6000 ;
	    RECT 239.6000 231.8000 240.4000 239.8000 ;
	    RECT 242.8000 232.4000 243.6000 239.8000 ;
	    RECT 241.4000 231.8000 243.6000 232.4000 ;
	    RECT 244.4000 231.8000 245.2000 239.8000 ;
	    RECT 247.6000 232.4000 248.4000 239.8000 ;
	    RECT 246.2000 231.8000 248.4000 232.4000 ;
	    RECT 249.2000 231.8000 250.0000 239.8000 ;
	    RECT 252.4000 232.4000 253.2000 239.8000 ;
	    RECT 251.0000 231.8000 253.2000 232.4000 ;
	    RECT 263.0000 231.8000 265.0000 239.8000 ;
	    RECT 269.2000 233.6000 270.0000 234.4000 ;
	    RECT 269.2000 232.4000 269.8000 233.6000 ;
	    RECT 270.6000 232.4000 271.4000 239.8000 ;
	    RECT 268.4000 231.8000 269.8000 232.4000 ;
	    RECT 270.4000 231.8000 271.4000 232.4000 ;
	    RECT 275.4000 232.6000 276.2000 239.8000 ;
	    RECT 275.4000 231.8000 277.2000 232.6000 ;
	    RECT 282.2000 232.4000 283.0000 239.8000 ;
	    RECT 283.6000 233.6000 284.4000 234.4000 ;
	    RECT 283.8000 232.4000 284.4000 233.6000 ;
	    RECT 282.2000 231.8000 283.2000 232.4000 ;
	    RECT 283.8000 231.8000 285.2000 232.4000 ;
	    RECT 288.6000 231.8000 290.6000 239.8000 ;
	    RECT 296.6000 232.6000 297.4000 239.8000 ;
	    RECT 295.6000 231.8000 297.4000 232.6000 ;
	    RECT 190.0000 231.6000 190.8000 231.8000 ;
	    RECT 190.1000 230.3000 190.7000 231.6000 ;
	    RECT 186.8000 229.7000 190.7000 230.3000 ;
	    RECT 169.2000 228.2000 170.0000 228.4000 ;
	    RECT 172.4000 228.3000 173.2000 228.4000 ;
	    RECT 174.0000 228.3000 174.8000 228.4000 ;
	    RECT 172.4000 228.2000 174.8000 228.3000 ;
	    RECT 167.6000 227.6000 170.0000 228.2000 ;
	    RECT 171.6000 227.7000 174.8000 228.2000 ;
	    RECT 171.6000 227.6000 173.2000 227.7000 ;
	    RECT 174.0000 227.6000 174.8000 227.7000 ;
	    RECT 175.6000 227.6000 176.4000 228.4000 ;
	    RECT 178.8000 227.6000 181.4000 228.4000 ;
	    RECT 183.6000 228.3000 184.4000 228.4000 ;
	    RECT 185.2000 228.3000 186.0000 228.4000 ;
	    RECT 183.6000 228.2000 186.0000 228.3000 ;
	    RECT 182.8000 227.7000 186.0000 228.2000 ;
	    RECT 182.8000 227.6000 184.4000 227.7000 ;
	    RECT 159.4000 226.6000 160.2000 227.0000 ;
	    RECT 159.4000 226.0000 161.0000 226.6000 ;
	    RECT 148.4000 222.2000 149.2000 224.2000 ;
	    RECT 153.2000 222.2000 154.0000 224.2000 ;
	    RECT 160.2000 223.0000 161.0000 226.0000 ;
	    RECT 164.6000 225.0000 165.2000 227.2000 ;
	    RECT 167.6000 226.2000 168.2000 227.6000 ;
	    RECT 171.6000 227.2000 172.4000 227.6000 ;
	    RECT 169.4000 226.2000 173.0000 226.6000 ;
	    RECT 164.4000 223.0000 165.2000 225.0000 ;
	    RECT 166.0000 222.8000 166.8000 226.2000 ;
	    RECT 167.6000 223.4000 168.4000 226.2000 ;
	    RECT 169.2000 226.0000 173.2000 226.2000 ;
	    RECT 169.2000 222.8000 170.0000 226.0000 ;
	    RECT 166.0000 222.2000 170.0000 222.8000 ;
	    RECT 172.4000 222.2000 173.2000 226.0000 ;
	    RECT 174.0000 224.8000 174.8000 226.4000 ;
	    RECT 175.8000 224.2000 176.4000 227.6000 ;
	    RECT 179.0000 226.2000 179.6000 227.6000 ;
	    RECT 182.8000 227.2000 183.6000 227.6000 ;
	    RECT 185.2000 226.8000 186.0000 227.7000 ;
	    RECT 180.6000 226.2000 184.2000 226.6000 ;
	    RECT 186.8000 226.2000 187.6000 229.7000 ;
	    RECT 192.0000 228.4000 192.6000 231.8000 ;
	    RECT 193.2000 230.3000 194.0000 230.4000 ;
	    RECT 194.8000 230.3000 195.6000 230.4000 ;
	    RECT 193.2000 229.7000 195.6000 230.3000 ;
	    RECT 193.2000 228.8000 194.0000 229.7000 ;
	    RECT 194.8000 229.6000 195.6000 229.7000 ;
	    RECT 196.4000 229.6000 197.0000 231.8000 ;
	    RECT 198.2000 231.2000 198.8000 231.8000 ;
	    RECT 197.6000 230.4000 198.8000 231.2000 ;
	    RECT 190.0000 227.6000 192.6000 228.4000 ;
	    RECT 194.8000 228.2000 195.6000 228.4000 ;
	    RECT 194.0000 227.6000 195.6000 228.2000 ;
	    RECT 190.2000 226.2000 190.8000 227.6000 ;
	    RECT 194.0000 227.2000 194.8000 227.6000 ;
	    RECT 191.8000 226.2000 195.4000 226.6000 ;
	    RECT 175.6000 222.2000 176.4000 224.2000 ;
	    RECT 178.8000 222.2000 179.6000 226.2000 ;
	    RECT 180.4000 226.0000 184.4000 226.2000 ;
	    RECT 180.4000 222.2000 181.2000 226.0000 ;
	    RECT 183.6000 222.2000 184.4000 226.0000 ;
	    RECT 186.8000 225.6000 188.6000 226.2000 ;
	    RECT 187.8000 222.2000 188.6000 225.6000 ;
	    RECT 190.0000 222.2000 190.8000 226.2000 ;
	    RECT 191.6000 226.0000 195.6000 226.2000 ;
	    RECT 191.6000 222.2000 192.4000 226.0000 ;
	    RECT 194.8000 222.2000 195.6000 226.0000 ;
	    RECT 196.4000 222.2000 197.2000 229.6000 ;
	    RECT 198.2000 227.4000 198.8000 230.4000 ;
	    RECT 199.6000 228.8000 200.4000 230.4000 ;
	    RECT 201.2000 229.6000 202.0000 231.2000 ;
	    RECT 202.8000 230.4000 203.4000 231.8000 ;
	    RECT 202.8000 229.6000 203.6000 230.4000 ;
	    RECT 202.8000 228.4000 203.4000 229.6000 ;
	    RECT 202.8000 227.6000 203.6000 228.4000 ;
	    RECT 206.0000 227.6000 206.8000 229.2000 ;
	    RECT 207.6000 228.8000 208.4000 230.4000 ;
	    RECT 209.4000 228.4000 210.0000 231.8000 ;
	    RECT 214.0000 231.6000 214.8000 231.8000 ;
	    RECT 210.8000 228.8000 211.6000 230.4000 ;
	    RECT 216.0000 228.4000 216.6000 231.8000 ;
	    RECT 217.2000 228.8000 218.0000 230.4000 ;
	    RECT 218.8000 229.6000 219.6000 230.4000 ;
	    RECT 218.9000 228.4000 219.5000 229.6000 ;
	    RECT 209.2000 228.2000 210.0000 228.4000 ;
	    RECT 212.4000 228.3000 213.2000 228.4000 ;
	    RECT 214.0000 228.3000 216.6000 228.4000 ;
	    RECT 212.4000 228.2000 216.6000 228.3000 ;
	    RECT 218.8000 228.2000 219.6000 228.4000 ;
	    RECT 207.6000 227.6000 210.0000 228.2000 ;
	    RECT 211.6000 227.7000 216.6000 228.2000 ;
	    RECT 211.6000 227.6000 213.2000 227.7000 ;
	    RECT 214.0000 227.6000 216.6000 227.7000 ;
	    RECT 218.0000 227.6000 219.6000 228.2000 ;
	    RECT 220.4000 227.6000 221.2000 229.2000 ;
	    RECT 222.0000 228.8000 222.8000 230.4000 ;
	    RECT 223.8000 228.4000 224.4000 231.8000 ;
	    RECT 228.4000 231.6000 229.2000 231.8000 ;
	    RECT 225.2000 228.8000 226.0000 230.4000 ;
	    RECT 230.4000 228.4000 231.0000 231.8000 ;
	    RECT 231.6000 230.3000 232.4000 230.4000 ;
	    RECT 233.2000 230.3000 234.0000 230.4000 ;
	    RECT 231.6000 229.7000 234.0000 230.3000 ;
	    RECT 231.6000 228.8000 232.4000 229.7000 ;
	    RECT 233.2000 229.6000 234.0000 229.7000 ;
	    RECT 236.6000 228.4000 237.2000 231.8000 ;
	    RECT 238.0000 229.6000 238.8000 231.2000 ;
	    RECT 239.6000 229.6000 240.2000 231.8000 ;
	    RECT 241.4000 231.2000 242.0000 231.8000 ;
	    RECT 240.8000 230.4000 242.0000 231.2000 ;
	    RECT 223.6000 228.2000 224.4000 228.4000 ;
	    RECT 226.8000 228.3000 227.6000 228.4000 ;
	    RECT 228.4000 228.3000 231.0000 228.4000 ;
	    RECT 226.8000 228.2000 231.0000 228.3000 ;
	    RECT 233.2000 228.2000 234.0000 228.4000 ;
	    RECT 222.0000 227.6000 224.4000 228.2000 ;
	    RECT 226.0000 227.7000 231.0000 228.2000 ;
	    RECT 226.0000 227.6000 227.6000 227.7000 ;
	    RECT 228.4000 227.6000 231.0000 227.7000 ;
	    RECT 232.4000 227.6000 234.0000 228.2000 ;
	    RECT 236.4000 227.6000 237.2000 228.4000 ;
	    RECT 198.2000 226.8000 200.4000 227.4000 ;
	    RECT 199.6000 222.2000 200.4000 226.8000 ;
	    RECT 202.8000 224.2000 203.4000 227.6000 ;
	    RECT 204.4000 224.8000 205.2000 226.4000 ;
	    RECT 207.6000 226.2000 208.2000 227.6000 ;
	    RECT 211.6000 227.2000 212.4000 227.6000 ;
	    RECT 209.4000 226.2000 213.0000 226.6000 ;
	    RECT 214.2000 226.2000 214.8000 227.6000 ;
	    RECT 218.0000 227.2000 218.8000 227.6000 ;
	    RECT 215.8000 226.2000 219.4000 226.6000 ;
	    RECT 222.0000 226.2000 222.6000 227.6000 ;
	    RECT 226.0000 227.2000 226.8000 227.6000 ;
	    RECT 223.8000 226.2000 227.4000 226.6000 ;
	    RECT 228.6000 226.2000 229.2000 227.6000 ;
	    RECT 232.4000 227.2000 233.2000 227.6000 ;
	    RECT 230.2000 226.2000 233.8000 226.6000 ;
	    RECT 202.8000 222.2000 203.6000 224.2000 ;
	    RECT 206.0000 222.8000 206.8000 226.2000 ;
	    RECT 207.6000 223.4000 208.4000 226.2000 ;
	    RECT 209.2000 226.0000 213.2000 226.2000 ;
	    RECT 209.2000 222.8000 210.0000 226.0000 ;
	    RECT 206.0000 222.2000 210.0000 222.8000 ;
	    RECT 212.4000 222.2000 213.2000 226.0000 ;
	    RECT 214.0000 222.2000 214.8000 226.2000 ;
	    RECT 215.6000 226.0000 219.6000 226.2000 ;
	    RECT 215.6000 222.2000 216.4000 226.0000 ;
	    RECT 218.8000 222.2000 219.6000 226.0000 ;
	    RECT 220.4000 222.8000 221.2000 226.2000 ;
	    RECT 222.0000 223.4000 222.8000 226.2000 ;
	    RECT 223.6000 226.0000 227.6000 226.2000 ;
	    RECT 223.6000 222.8000 224.4000 226.0000 ;
	    RECT 220.4000 222.2000 224.4000 222.8000 ;
	    RECT 226.8000 222.2000 227.6000 226.0000 ;
	    RECT 228.4000 222.2000 229.2000 226.2000 ;
	    RECT 230.0000 226.0000 234.0000 226.2000 ;
	    RECT 230.0000 222.2000 230.8000 226.0000 ;
	    RECT 233.2000 222.2000 234.0000 226.0000 ;
	    RECT 234.8000 224.8000 235.6000 226.4000 ;
	    RECT 236.6000 226.3000 237.2000 227.6000 ;
	    RECT 238.0000 226.3000 238.8000 226.4000 ;
	    RECT 236.5000 225.7000 238.8000 226.3000 ;
	    RECT 236.6000 224.2000 237.2000 225.7000 ;
	    RECT 238.0000 225.6000 238.8000 225.7000 ;
	    RECT 236.4000 222.2000 237.2000 224.2000 ;
	    RECT 239.6000 222.2000 240.4000 229.6000 ;
	    RECT 241.4000 227.4000 242.0000 230.4000 ;
	    RECT 242.8000 228.8000 243.6000 230.4000 ;
	    RECT 244.4000 229.6000 245.0000 231.8000 ;
	    RECT 246.2000 231.2000 246.8000 231.8000 ;
	    RECT 245.6000 230.4000 246.8000 231.2000 ;
	    RECT 241.4000 226.8000 243.6000 227.4000 ;
	    RECT 242.8000 222.2000 243.6000 226.8000 ;
	    RECT 244.4000 222.2000 245.2000 229.6000 ;
	    RECT 246.2000 227.4000 246.8000 230.4000 ;
	    RECT 247.6000 228.8000 248.4000 230.4000 ;
	    RECT 249.2000 229.6000 249.8000 231.8000 ;
	    RECT 251.0000 231.2000 251.6000 231.8000 ;
	    RECT 250.4000 230.4000 251.6000 231.2000 ;
	    RECT 246.2000 226.8000 248.4000 227.4000 ;
	    RECT 247.6000 222.2000 248.4000 226.8000 ;
	    RECT 249.2000 222.2000 250.0000 229.6000 ;
	    RECT 251.0000 227.4000 251.6000 230.4000 ;
	    RECT 252.4000 228.8000 253.2000 230.4000 ;
	    RECT 260.4000 227.6000 261.2000 229.2000 ;
	    RECT 262.0000 228.8000 262.8000 230.4000 ;
	    RECT 263.8000 228.4000 264.4000 231.8000 ;
	    RECT 268.4000 231.6000 269.2000 231.8000 ;
	    RECT 265.2000 228.8000 266.0000 230.4000 ;
	    RECT 270.4000 228.4000 271.0000 231.8000 ;
	    RECT 271.6000 228.8000 272.4000 230.4000 ;
	    RECT 274.8000 229.6000 275.6000 231.2000 ;
	    RECT 276.4000 228.4000 277.0000 231.8000 ;
	    RECT 281.2000 228.8000 282.0000 230.4000 ;
	    RECT 282.6000 228.4000 283.2000 231.8000 ;
	    RECT 284.4000 231.6000 285.2000 231.8000 ;
	    RECT 284.5000 230.3000 285.1000 231.6000 ;
	    RECT 284.5000 229.7000 286.8000 230.3000 ;
	    RECT 263.6000 228.2000 264.4000 228.4000 ;
	    RECT 266.8000 228.3000 267.6000 228.4000 ;
	    RECT 268.4000 228.3000 271.0000 228.4000 ;
	    RECT 266.8000 228.2000 271.0000 228.3000 ;
	    RECT 273.2000 228.2000 274.0000 228.4000 ;
	    RECT 262.0000 227.6000 264.4000 228.2000 ;
	    RECT 266.0000 227.7000 271.0000 228.2000 ;
	    RECT 266.0000 227.6000 267.6000 227.7000 ;
	    RECT 268.4000 227.6000 271.0000 227.7000 ;
	    RECT 272.4000 227.6000 274.0000 228.2000 ;
	    RECT 276.4000 227.6000 277.2000 228.4000 ;
	    RECT 279.6000 228.2000 280.4000 228.4000 ;
	    RECT 279.6000 227.6000 281.2000 228.2000 ;
	    RECT 282.6000 227.6000 285.2000 228.4000 ;
	    RECT 286.0000 227.6000 286.8000 229.7000 ;
	    RECT 287.6000 228.8000 288.4000 230.4000 ;
	    RECT 289.4000 228.4000 290.0000 231.8000 ;
	    RECT 290.8000 230.3000 291.6000 230.4000 ;
	    RECT 295.8000 230.3000 296.4000 231.8000 ;
	    RECT 290.8000 229.7000 296.4000 230.3000 ;
	    RECT 290.8000 228.8000 291.6000 229.7000 ;
	    RECT 295.8000 228.4000 296.4000 229.7000 ;
	    RECT 297.2000 229.6000 298.0000 231.2000 ;
	    RECT 289.2000 228.2000 290.0000 228.4000 ;
	    RECT 292.4000 228.2000 293.2000 228.4000 ;
	    RECT 287.6000 227.6000 290.0000 228.2000 ;
	    RECT 291.6000 227.6000 293.2000 228.2000 ;
	    RECT 295.6000 227.6000 296.4000 228.4000 ;
	    RECT 251.0000 226.8000 253.2000 227.4000 ;
	    RECT 252.4000 222.2000 253.2000 226.8000 ;
	    RECT 262.0000 226.2000 262.6000 227.6000 ;
	    RECT 266.0000 227.2000 266.8000 227.6000 ;
	    RECT 263.8000 226.2000 267.4000 226.6000 ;
	    RECT 268.6000 226.2000 269.2000 227.6000 ;
	    RECT 272.4000 227.2000 273.2000 227.6000 ;
	    RECT 270.2000 226.2000 273.8000 226.6000 ;
	    RECT 274.8000 226.3000 275.6000 226.4000 ;
	    RECT 276.4000 226.3000 277.0000 227.6000 ;
	    RECT 280.4000 227.2000 281.2000 227.6000 ;
	    RECT 260.4000 222.8000 261.2000 226.2000 ;
	    RECT 262.0000 223.4000 262.8000 226.2000 ;
	    RECT 263.6000 226.0000 267.6000 226.2000 ;
	    RECT 263.6000 222.8000 264.4000 226.0000 ;
	    RECT 260.4000 222.2000 264.4000 222.8000 ;
	    RECT 266.8000 222.2000 267.6000 226.0000 ;
	    RECT 268.4000 222.2000 269.2000 226.2000 ;
	    RECT 270.0000 226.0000 274.0000 226.2000 ;
	    RECT 270.0000 222.2000 270.8000 226.0000 ;
	    RECT 273.2000 222.2000 274.0000 226.0000 ;
	    RECT 274.8000 225.7000 277.1000 226.3000 ;
	    RECT 274.8000 225.6000 275.6000 225.7000 ;
	    RECT 276.4000 224.2000 277.0000 225.7000 ;
	    RECT 278.0000 224.8000 278.8000 226.4000 ;
	    RECT 279.8000 226.2000 283.4000 226.6000 ;
	    RECT 284.4000 226.2000 285.0000 227.6000 ;
	    RECT 287.6000 226.2000 288.2000 227.6000 ;
	    RECT 291.6000 227.2000 292.4000 227.6000 ;
	    RECT 289.4000 226.2000 293.0000 226.6000 ;
	    RECT 279.6000 226.0000 283.6000 226.2000 ;
	    RECT 276.4000 222.2000 277.2000 224.2000 ;
	    RECT 279.6000 222.2000 280.4000 226.0000 ;
	    RECT 282.8000 222.2000 283.6000 226.0000 ;
	    RECT 284.4000 222.2000 285.2000 226.2000 ;
	    RECT 286.0000 222.8000 286.8000 226.2000 ;
	    RECT 287.6000 223.4000 288.4000 226.2000 ;
	    RECT 289.2000 226.0000 293.2000 226.2000 ;
	    RECT 289.2000 222.8000 290.0000 226.0000 ;
	    RECT 286.0000 222.2000 290.0000 222.8000 ;
	    RECT 292.4000 222.2000 293.2000 226.0000 ;
	    RECT 294.0000 224.8000 294.8000 226.4000 ;
	    RECT 295.8000 224.2000 296.4000 227.6000 ;
	    RECT 295.6000 222.2000 296.4000 224.2000 ;
	    RECT 298.8000 222.2000 299.6000 239.8000 ;
	    RECT 302.0000 235.0000 302.8000 239.0000 ;
	    RECT 302.0000 231.6000 302.6000 235.0000 ;
	    RECT 306.2000 234.4000 307.0000 239.8000 ;
	    RECT 305.2000 233.6000 307.0000 234.4000 ;
	    RECT 306.2000 232.8000 307.0000 233.6000 ;
	    RECT 311.6000 235.0000 312.4000 239.0000 ;
	    RECT 306.2000 232.2000 307.8000 232.8000 ;
	    RECT 302.0000 231.0000 305.8000 231.6000 ;
	    RECT 302.0000 228.8000 302.8000 230.4000 ;
	    RECT 303.6000 228.8000 304.4000 230.4000 ;
	    RECT 305.2000 229.0000 305.8000 231.0000 ;
	    RECT 305.2000 228.2000 306.6000 229.0000 ;
	    RECT 307.2000 228.4000 307.8000 232.2000 ;
	    RECT 311.6000 231.6000 312.2000 235.0000 ;
	    RECT 315.8000 232.8000 316.6000 239.8000 ;
	    RECT 315.8000 232.2000 317.4000 232.8000 ;
	    RECT 308.4000 229.6000 309.2000 231.2000 ;
	    RECT 311.6000 231.0000 315.4000 231.6000 ;
	    RECT 311.6000 228.8000 312.4000 230.4000 ;
	    RECT 313.2000 228.8000 314.0000 230.4000 ;
	    RECT 314.8000 229.0000 315.4000 231.0000 ;
	    RECT 305.2000 227.8000 306.2000 228.2000 ;
	    RECT 302.0000 227.2000 306.2000 227.8000 ;
	    RECT 307.2000 227.6000 309.2000 228.4000 ;
	    RECT 314.8000 228.2000 316.2000 229.0000 ;
	    RECT 316.8000 228.4000 317.4000 232.2000 ;
	    RECT 321.2000 231.8000 322.0000 239.8000 ;
	    RECT 324.4000 232.4000 325.2000 239.8000 ;
	    RECT 323.0000 231.8000 325.2000 232.4000 ;
	    RECT 318.0000 229.6000 318.8000 231.2000 ;
	    RECT 321.2000 229.6000 321.8000 231.8000 ;
	    RECT 323.0000 231.2000 323.6000 231.8000 ;
	    RECT 322.4000 230.4000 323.6000 231.2000 ;
	    RECT 326.0000 231.2000 326.8000 239.8000 ;
	    RECT 330.2000 235.8000 331.4000 239.8000 ;
	    RECT 334.8000 235.8000 335.6000 239.8000 ;
	    RECT 339.2000 236.4000 340.0000 239.8000 ;
	    RECT 339.2000 235.8000 341.2000 236.4000 ;
	    RECT 330.8000 235.0000 331.6000 235.8000 ;
	    RECT 335.0000 235.2000 335.6000 235.8000 ;
	    RECT 334.2000 234.6000 337.8000 235.2000 ;
	    RECT 340.4000 235.0000 341.2000 235.8000 ;
	    RECT 334.2000 234.4000 335.0000 234.6000 ;
	    RECT 337.0000 234.4000 337.8000 234.6000 ;
	    RECT 330.0000 233.2000 331.4000 234.0000 ;
	    RECT 330.8000 232.2000 331.4000 233.2000 ;
	    RECT 333.0000 233.0000 335.2000 233.6000 ;
	    RECT 333.0000 232.8000 333.8000 233.0000 ;
	    RECT 330.8000 231.6000 333.2000 232.2000 ;
	    RECT 326.0000 230.6000 330.2000 231.2000 ;
	    RECT 314.8000 227.8000 315.8000 228.2000 ;
	    RECT 302.0000 225.0000 302.6000 227.2000 ;
	    RECT 307.2000 227.0000 307.8000 227.6000 ;
	    RECT 307.0000 226.6000 307.8000 227.0000 ;
	    RECT 306.2000 226.0000 307.8000 226.6000 ;
	    RECT 311.6000 227.2000 315.8000 227.8000 ;
	    RECT 316.8000 227.6000 318.8000 228.4000 ;
	    RECT 302.0000 223.0000 302.8000 225.0000 ;
	    RECT 306.2000 223.0000 307.0000 226.0000 ;
	    RECT 311.6000 225.0000 312.2000 227.2000 ;
	    RECT 316.8000 227.0000 317.4000 227.6000 ;
	    RECT 316.6000 226.6000 317.4000 227.0000 ;
	    RECT 315.8000 226.0000 317.4000 226.6000 ;
	    RECT 311.6000 223.0000 312.4000 225.0000 ;
	    RECT 315.8000 224.4000 316.6000 226.0000 ;
	    RECT 314.8000 223.6000 316.6000 224.4000 ;
	    RECT 315.8000 223.0000 316.6000 223.6000 ;
	    RECT 321.2000 222.2000 322.0000 229.6000 ;
	    RECT 323.0000 227.4000 323.6000 230.4000 ;
	    RECT 324.4000 228.8000 325.2000 230.4000 ;
	    RECT 323.0000 226.8000 325.2000 227.4000 ;
	    RECT 324.4000 222.2000 325.2000 226.8000 ;
	    RECT 326.0000 227.2000 326.8000 230.6000 ;
	    RECT 329.4000 230.4000 330.2000 230.6000 ;
	    RECT 327.8000 229.8000 328.6000 230.0000 ;
	    RECT 327.8000 229.2000 331.6000 229.8000 ;
	    RECT 330.8000 229.0000 331.6000 229.2000 ;
	    RECT 332.6000 228.4000 333.2000 231.6000 ;
	    RECT 334.6000 231.8000 335.2000 233.0000 ;
	    RECT 335.8000 233.0000 336.6000 233.2000 ;
	    RECT 340.4000 233.0000 341.2000 233.2000 ;
	    RECT 335.8000 232.4000 341.2000 233.0000 ;
	    RECT 334.6000 231.4000 339.4000 231.8000 ;
	    RECT 343.6000 231.4000 344.4000 239.8000 ;
	    RECT 347.8000 232.4000 348.6000 239.8000 ;
	    RECT 349.2000 233.6000 350.0000 234.4000 ;
	    RECT 349.4000 232.4000 350.0000 233.6000 ;
	    RECT 352.4000 233.6000 353.2000 234.4000 ;
	    RECT 352.4000 232.4000 353.0000 233.6000 ;
	    RECT 353.8000 232.4000 354.6000 239.8000 ;
	    RECT 347.8000 231.8000 348.8000 232.4000 ;
	    RECT 349.4000 231.8000 350.8000 232.4000 ;
	    RECT 334.6000 231.2000 344.4000 231.4000 ;
	    RECT 338.6000 231.0000 344.4000 231.2000 ;
	    RECT 338.8000 230.8000 344.4000 231.0000 ;
	    RECT 348.2000 230.4000 348.8000 231.8000 ;
	    RECT 350.0000 231.6000 350.8000 231.8000 ;
	    RECT 351.6000 231.8000 353.0000 232.4000 ;
	    RECT 353.6000 231.8000 354.6000 232.4000 ;
	    RECT 358.0000 232.4000 358.8000 239.8000 ;
	    RECT 358.0000 231.8000 360.2000 232.4000 ;
	    RECT 361.2000 231.8000 362.0000 239.8000 ;
	    RECT 351.6000 231.6000 352.4000 231.8000 ;
	    RECT 337.2000 230.2000 338.0000 230.4000 ;
	    RECT 337.2000 229.6000 342.2000 230.2000 ;
	    RECT 341.4000 229.4000 342.2000 229.6000 ;
	    RECT 346.8000 228.8000 347.6000 230.4000 ;
	    RECT 348.2000 229.6000 349.2000 230.4000 ;
	    RECT 350.1000 230.3000 350.7000 231.6000 ;
	    RECT 353.6000 230.3000 354.2000 231.8000 ;
	    RECT 359.6000 231.2000 360.2000 231.8000 ;
	    RECT 359.6000 230.4000 360.8000 231.2000 ;
	    RECT 350.1000 229.7000 354.2000 230.3000 ;
	    RECT 339.8000 228.4000 340.6000 228.6000 ;
	    RECT 348.2000 228.4000 348.8000 229.6000 ;
	    RECT 353.6000 228.4000 354.2000 229.7000 ;
	    RECT 354.8000 228.8000 355.6000 230.4000 ;
	    RECT 358.0000 228.8000 358.8000 230.4000 ;
	    RECT 332.6000 227.8000 343.6000 228.4000 ;
	    RECT 333.0000 227.6000 333.8000 227.8000 ;
	    RECT 338.8000 227.6000 339.6000 227.8000 ;
	    RECT 342.0000 227.6000 343.6000 227.8000 ;
	    RECT 345.2000 228.2000 346.0000 228.4000 ;
	    RECT 345.2000 227.6000 346.8000 228.2000 ;
	    RECT 348.2000 227.6000 350.8000 228.4000 ;
	    RECT 351.6000 227.6000 354.2000 228.4000 ;
	    RECT 356.4000 228.2000 357.2000 228.4000 ;
	    RECT 355.6000 227.6000 357.2000 228.2000 ;
	    RECT 326.0000 226.6000 329.8000 227.2000 ;
	    RECT 326.0000 222.2000 326.8000 226.6000 ;
	    RECT 329.0000 226.4000 329.8000 226.6000 ;
	    RECT 338.8000 225.6000 339.4000 227.6000 ;
	    RECT 346.0000 227.2000 346.8000 227.6000 ;
	    RECT 337.0000 225.4000 337.8000 225.6000 ;
	    RECT 330.8000 224.2000 331.6000 225.0000 ;
	    RECT 335.0000 224.8000 337.8000 225.4000 ;
	    RECT 338.8000 224.8000 339.6000 225.6000 ;
	    RECT 335.0000 224.2000 335.6000 224.8000 ;
	    RECT 340.4000 224.2000 341.2000 225.0000 ;
	    RECT 330.2000 223.6000 331.6000 224.2000 ;
	    RECT 330.2000 222.2000 331.4000 223.6000 ;
	    RECT 334.8000 222.2000 335.6000 224.2000 ;
	    RECT 339.2000 223.6000 341.2000 224.2000 ;
	    RECT 339.2000 222.2000 340.0000 223.6000 ;
	    RECT 343.6000 222.2000 344.4000 227.0000 ;
	    RECT 345.4000 226.2000 349.0000 226.6000 ;
	    RECT 350.0000 226.2000 350.6000 227.6000 ;
	    RECT 351.8000 226.2000 352.4000 227.6000 ;
	    RECT 355.6000 227.2000 356.4000 227.6000 ;
	    RECT 359.6000 227.4000 360.2000 230.4000 ;
	    RECT 361.4000 229.6000 362.0000 231.8000 ;
	    RECT 358.0000 226.8000 360.2000 227.4000 ;
	    RECT 353.4000 226.2000 357.0000 226.6000 ;
	    RECT 345.2000 226.0000 349.2000 226.2000 ;
	    RECT 345.2000 222.2000 346.0000 226.0000 ;
	    RECT 348.4000 222.2000 349.2000 226.0000 ;
	    RECT 350.0000 222.2000 350.8000 226.2000 ;
	    RECT 351.6000 222.2000 352.4000 226.2000 ;
	    RECT 353.2000 226.0000 357.2000 226.2000 ;
	    RECT 353.2000 222.2000 354.0000 226.0000 ;
	    RECT 356.4000 222.2000 357.2000 226.0000 ;
	    RECT 358.0000 222.2000 358.8000 226.8000 ;
	    RECT 361.2000 222.2000 362.0000 229.6000 ;
	    RECT 362.8000 231.2000 363.6000 239.8000 ;
	    RECT 367.0000 235.8000 368.2000 239.8000 ;
	    RECT 371.6000 235.8000 372.4000 239.8000 ;
	    RECT 376.0000 236.4000 376.8000 239.8000 ;
	    RECT 376.0000 235.8000 378.0000 236.4000 ;
	    RECT 367.6000 235.0000 368.4000 235.8000 ;
	    RECT 371.8000 235.2000 372.4000 235.8000 ;
	    RECT 371.0000 234.6000 374.6000 235.2000 ;
	    RECT 377.2000 235.0000 378.0000 235.8000 ;
	    RECT 371.0000 234.4000 371.8000 234.6000 ;
	    RECT 373.8000 234.4000 374.6000 234.6000 ;
	    RECT 366.8000 233.2000 368.2000 234.0000 ;
	    RECT 367.6000 232.2000 368.2000 233.2000 ;
	    RECT 369.8000 233.0000 372.0000 233.6000 ;
	    RECT 369.8000 232.8000 370.6000 233.0000 ;
	    RECT 367.6000 231.6000 370.0000 232.2000 ;
	    RECT 362.8000 230.6000 367.0000 231.2000 ;
	    RECT 362.8000 227.2000 363.6000 230.6000 ;
	    RECT 366.2000 230.4000 367.0000 230.6000 ;
	    RECT 369.4000 230.3000 370.0000 231.6000 ;
	    RECT 371.4000 231.8000 372.0000 233.0000 ;
	    RECT 372.6000 233.0000 373.4000 233.2000 ;
	    RECT 377.2000 233.0000 378.0000 233.2000 ;
	    RECT 372.6000 232.4000 378.0000 233.0000 ;
	    RECT 371.4000 231.4000 376.2000 231.8000 ;
	    RECT 380.4000 231.4000 381.2000 239.8000 ;
	    RECT 371.4000 231.2000 381.2000 231.4000 ;
	    RECT 375.4000 231.0000 381.2000 231.2000 ;
	    RECT 375.6000 230.8000 381.2000 231.0000 ;
	    RECT 370.8000 230.3000 371.6000 230.4000 ;
	    RECT 364.6000 229.8000 365.4000 230.0000 ;
	    RECT 364.6000 229.2000 368.4000 229.8000 ;
	    RECT 369.3000 229.7000 371.6000 230.3000 ;
	    RECT 367.6000 229.0000 368.4000 229.2000 ;
	    RECT 369.4000 228.4000 370.0000 229.7000 ;
	    RECT 370.8000 229.6000 371.6000 229.7000 ;
	    RECT 374.0000 230.2000 374.8000 230.4000 ;
	    RECT 374.0000 229.6000 379.0000 230.2000 ;
	    RECT 375.6000 229.4000 376.4000 229.6000 ;
	    RECT 378.2000 229.4000 379.0000 229.6000 ;
	    RECT 376.6000 228.4000 377.4000 228.6000 ;
	    RECT 369.4000 227.8000 380.4000 228.4000 ;
	    RECT 369.8000 227.6000 370.6000 227.8000 ;
	    RECT 362.8000 226.6000 366.6000 227.2000 ;
	    RECT 362.8000 222.2000 363.6000 226.6000 ;
	    RECT 365.8000 226.4000 366.6000 226.6000 ;
	    RECT 375.6000 225.6000 376.2000 227.8000 ;
	    RECT 378.8000 227.6000 380.4000 227.8000 ;
	    RECT 383.6000 228.3000 384.4000 239.8000 ;
	    RECT 387.8000 232.4000 388.6000 239.8000 ;
	    RECT 389.2000 233.6000 390.0000 234.4000 ;
	    RECT 389.4000 232.4000 390.0000 233.6000 ;
	    RECT 386.8000 231.6000 388.8000 232.4000 ;
	    RECT 389.4000 231.8000 390.8000 232.4000 ;
	    RECT 390.0000 231.6000 390.8000 231.8000 ;
	    RECT 391.6000 231.8000 392.4000 239.8000 ;
	    RECT 394.8000 232.4000 395.6000 239.8000 ;
	    RECT 393.4000 231.8000 395.6000 232.4000 ;
	    RECT 386.8000 228.8000 387.6000 230.4000 ;
	    RECT 388.2000 228.4000 388.8000 231.6000 ;
	    RECT 391.6000 229.6000 392.2000 231.8000 ;
	    RECT 393.4000 231.2000 394.0000 231.8000 ;
	    RECT 392.8000 230.4000 394.0000 231.2000 ;
	    RECT 385.2000 228.3000 386.0000 228.4000 ;
	    RECT 383.6000 228.2000 386.0000 228.3000 ;
	    RECT 383.6000 227.7000 386.8000 228.2000 ;
	    RECT 373.8000 225.4000 374.6000 225.6000 ;
	    RECT 367.6000 224.2000 368.4000 225.0000 ;
	    RECT 371.8000 224.8000 374.6000 225.4000 ;
	    RECT 375.6000 224.8000 376.4000 225.6000 ;
	    RECT 371.8000 224.2000 372.4000 224.8000 ;
	    RECT 377.2000 224.2000 378.0000 225.0000 ;
	    RECT 367.0000 223.6000 368.4000 224.2000 ;
	    RECT 367.0000 222.2000 368.2000 223.6000 ;
	    RECT 371.6000 222.2000 372.4000 224.2000 ;
	    RECT 376.0000 223.6000 378.0000 224.2000 ;
	    RECT 376.0000 222.2000 376.8000 223.6000 ;
	    RECT 380.4000 222.2000 381.2000 227.0000 ;
	    RECT 382.0000 224.8000 382.8000 226.4000 ;
	    RECT 383.6000 222.2000 384.4000 227.7000 ;
	    RECT 385.2000 227.6000 386.8000 227.7000 ;
	    RECT 388.2000 227.6000 390.8000 228.4000 ;
	    RECT 386.0000 227.2000 386.8000 227.6000 ;
	    RECT 385.4000 226.2000 389.0000 226.6000 ;
	    RECT 390.0000 226.2000 390.6000 227.6000 ;
	    RECT 385.2000 226.0000 389.2000 226.2000 ;
	    RECT 385.2000 222.2000 386.0000 226.0000 ;
	    RECT 388.4000 222.2000 389.2000 226.0000 ;
	    RECT 390.0000 222.2000 390.8000 226.2000 ;
	    RECT 391.6000 222.2000 392.4000 229.6000 ;
	    RECT 393.4000 227.4000 394.0000 230.4000 ;
	    RECT 394.8000 228.8000 395.6000 230.4000 ;
	    RECT 398.0000 230.3000 398.8000 239.8000 ;
	    RECT 402.0000 233.6000 402.8000 234.4000 ;
	    RECT 399.6000 231.6000 400.4000 233.2000 ;
	    RECT 402.0000 232.4000 402.6000 233.6000 ;
	    RECT 403.4000 232.4000 404.2000 239.8000 ;
	    RECT 401.2000 231.8000 402.6000 232.4000 ;
	    RECT 403.2000 231.8000 404.2000 232.4000 ;
	    RECT 401.2000 231.6000 402.0000 231.8000 ;
	    RECT 401.3000 230.3000 401.9000 231.6000 ;
	    RECT 403.2000 230.4000 403.8000 231.8000 ;
	    RECT 414.0000 231.2000 414.8000 239.8000 ;
	    RECT 418.2000 235.8000 419.4000 239.8000 ;
	    RECT 422.8000 235.8000 423.6000 239.8000 ;
	    RECT 427.2000 236.4000 428.0000 239.8000 ;
	    RECT 427.2000 235.8000 429.2000 236.4000 ;
	    RECT 418.8000 235.0000 419.6000 235.8000 ;
	    RECT 423.0000 235.2000 423.6000 235.8000 ;
	    RECT 422.2000 234.6000 425.8000 235.2000 ;
	    RECT 428.4000 235.0000 429.2000 235.8000 ;
	    RECT 422.2000 234.4000 423.0000 234.6000 ;
	    RECT 425.0000 234.4000 425.8000 234.6000 ;
	    RECT 418.0000 233.2000 419.4000 234.0000 ;
	    RECT 418.8000 232.2000 419.4000 233.2000 ;
	    RECT 421.0000 233.0000 423.2000 233.6000 ;
	    RECT 421.0000 232.8000 421.8000 233.0000 ;
	    RECT 418.8000 231.6000 421.2000 232.2000 ;
	    RECT 414.0000 230.6000 418.2000 231.2000 ;
	    RECT 398.0000 229.7000 401.9000 230.3000 ;
	    RECT 393.4000 226.8000 395.6000 227.4000 ;
	    RECT 396.4000 226.8000 397.2000 228.4000 ;
	    RECT 394.8000 222.2000 395.6000 226.8000 ;
	    RECT 398.0000 226.2000 398.8000 229.7000 ;
	    RECT 402.8000 229.6000 403.8000 230.4000 ;
	    RECT 403.2000 228.4000 403.8000 229.6000 ;
	    RECT 404.4000 228.8000 405.2000 230.4000 ;
	    RECT 401.2000 227.6000 403.8000 228.4000 ;
	    RECT 406.0000 228.3000 406.8000 228.4000 ;
	    RECT 412.4000 228.3000 413.2000 228.4000 ;
	    RECT 406.0000 228.2000 413.2000 228.3000 ;
	    RECT 405.2000 227.7000 413.2000 228.2000 ;
	    RECT 405.2000 227.6000 406.8000 227.7000 ;
	    RECT 412.4000 227.6000 413.2000 227.7000 ;
	    RECT 401.4000 226.2000 402.0000 227.6000 ;
	    RECT 405.2000 227.2000 406.0000 227.6000 ;
	    RECT 414.0000 227.2000 414.8000 230.6000 ;
	    RECT 417.4000 230.4000 418.2000 230.6000 ;
	    RECT 415.8000 229.8000 416.6000 230.0000 ;
	    RECT 415.8000 229.2000 419.6000 229.8000 ;
	    RECT 418.8000 229.0000 419.6000 229.2000 ;
	    RECT 420.6000 228.4000 421.2000 231.6000 ;
	    RECT 422.6000 231.8000 423.2000 233.0000 ;
	    RECT 423.8000 233.0000 424.6000 233.2000 ;
	    RECT 428.4000 233.0000 429.2000 233.2000 ;
	    RECT 423.8000 232.4000 429.2000 233.0000 ;
	    RECT 422.6000 231.4000 427.4000 231.8000 ;
	    RECT 431.6000 231.4000 432.4000 239.8000 ;
	    RECT 433.2000 235.8000 434.0000 239.8000 ;
	    RECT 433.4000 235.6000 434.0000 235.8000 ;
	    RECT 436.4000 235.8000 437.2000 239.8000 ;
	    RECT 439.6000 235.8000 440.4000 239.8000 ;
	    RECT 436.4000 235.6000 437.0000 235.8000 ;
	    RECT 433.4000 235.0000 437.0000 235.6000 ;
	    RECT 439.8000 235.6000 440.4000 235.8000 ;
	    RECT 442.8000 235.8000 443.6000 239.8000 ;
	    RECT 442.8000 235.6000 443.4000 235.8000 ;
	    RECT 439.8000 235.0000 443.4000 235.6000 ;
	    RECT 433.4000 232.4000 434.0000 235.0000 ;
	    RECT 434.8000 234.3000 435.6000 234.4000 ;
	    RECT 436.4000 234.3000 437.2000 234.4000 ;
	    RECT 434.8000 233.7000 437.2000 234.3000 ;
	    RECT 434.8000 232.8000 435.6000 233.7000 ;
	    RECT 436.4000 233.6000 437.2000 233.7000 ;
	    RECT 439.8000 232.4000 440.4000 235.0000 ;
	    RECT 441.2000 234.3000 442.0000 234.4000 ;
	    RECT 446.0000 234.3000 446.8000 239.8000 ;
	    RECT 441.2000 233.7000 446.8000 234.3000 ;
	    RECT 441.2000 232.8000 442.0000 233.7000 ;
	    RECT 433.2000 231.6000 434.0000 232.4000 ;
	    RECT 439.6000 231.6000 440.4000 232.4000 ;
	    RECT 422.6000 231.2000 432.4000 231.4000 ;
	    RECT 426.6000 231.0000 432.4000 231.2000 ;
	    RECT 426.8000 230.8000 432.4000 231.0000 ;
	    RECT 425.2000 230.2000 426.0000 230.4000 ;
	    RECT 425.2000 229.6000 430.2000 230.2000 ;
	    RECT 429.4000 229.4000 430.2000 229.6000 ;
	    RECT 427.8000 228.4000 428.6000 228.6000 ;
	    RECT 433.4000 228.4000 434.0000 231.6000 ;
	    RECT 435.6000 229.6000 437.2000 230.4000 ;
	    RECT 439.8000 228.4000 440.4000 231.6000 ;
	    RECT 446.0000 231.8000 446.8000 233.7000 ;
	    RECT 449.2000 232.4000 450.0000 239.8000 ;
	    RECT 451.6000 233.6000 452.4000 234.4000 ;
	    RECT 451.6000 232.4000 452.2000 233.6000 ;
	    RECT 453.0000 232.4000 453.8000 239.8000 ;
	    RECT 447.8000 231.8000 450.0000 232.4000 ;
	    RECT 450.8000 231.8000 452.2000 232.4000 ;
	    RECT 452.8000 231.8000 453.8000 232.4000 ;
	    RECT 442.0000 229.6000 443.6000 230.4000 ;
	    RECT 446.0000 229.6000 446.6000 231.8000 ;
	    RECT 447.8000 231.2000 448.4000 231.8000 ;
	    RECT 450.8000 231.6000 451.6000 231.8000 ;
	    RECT 447.2000 230.4000 448.4000 231.2000 ;
	    RECT 420.6000 227.8000 431.6000 228.4000 ;
	    RECT 433.4000 228.2000 435.0000 228.4000 ;
	    RECT 433.4000 227.8000 435.2000 228.2000 ;
	    RECT 439.8000 227.8000 442.0000 228.4000 ;
	    RECT 421.0000 227.6000 421.8000 227.8000 ;
	    RECT 414.0000 226.6000 417.8000 227.2000 ;
	    RECT 403.0000 226.2000 406.6000 226.6000 ;
	    RECT 398.0000 225.6000 399.8000 226.2000 ;
	    RECT 399.0000 222.2000 399.8000 225.6000 ;
	    RECT 401.2000 222.2000 402.0000 226.2000 ;
	    RECT 402.8000 226.0000 406.8000 226.2000 ;
	    RECT 402.8000 222.2000 403.6000 226.0000 ;
	    RECT 406.0000 222.2000 406.8000 226.0000 ;
	    RECT 414.0000 222.2000 414.8000 226.6000 ;
	    RECT 417.0000 226.4000 417.8000 226.6000 ;
	    RECT 426.8000 225.6000 427.4000 227.8000 ;
	    RECT 430.0000 227.6000 431.6000 227.8000 ;
	    RECT 425.0000 225.4000 425.8000 225.6000 ;
	    RECT 418.8000 224.2000 419.6000 225.0000 ;
	    RECT 423.0000 224.8000 425.8000 225.4000 ;
	    RECT 426.8000 224.8000 427.6000 225.6000 ;
	    RECT 423.0000 224.2000 423.6000 224.8000 ;
	    RECT 428.4000 224.2000 429.2000 225.0000 ;
	    RECT 418.2000 223.6000 419.6000 224.2000 ;
	    RECT 418.2000 222.2000 419.4000 223.6000 ;
	    RECT 422.8000 222.2000 423.6000 224.2000 ;
	    RECT 427.2000 223.6000 429.2000 224.2000 ;
	    RECT 427.2000 222.2000 428.0000 223.6000 ;
	    RECT 431.6000 222.2000 432.4000 227.0000 ;
	    RECT 434.4000 222.2000 435.2000 227.8000 ;
	    RECT 440.8000 227.6000 442.0000 227.8000 ;
	    RECT 440.8000 222.2000 441.6000 227.6000 ;
	    RECT 446.0000 222.2000 446.8000 229.6000 ;
	    RECT 447.8000 227.4000 448.4000 230.4000 ;
	    RECT 449.2000 228.8000 450.0000 230.4000 ;
	    RECT 452.8000 228.4000 453.4000 231.8000 ;
	    RECT 454.0000 228.8000 454.8000 230.4000 ;
	    RECT 450.8000 227.6000 453.4000 228.4000 ;
	    RECT 455.6000 228.3000 456.4000 228.4000 ;
	    RECT 457.2000 228.3000 458.0000 239.8000 ;
	    RECT 458.8000 234.3000 459.6000 234.4000 ;
	    RECT 460.4000 234.3000 461.2000 239.8000 ;
	    RECT 464.6000 235.8000 465.8000 239.8000 ;
	    RECT 469.2000 235.8000 470.0000 239.8000 ;
	    RECT 473.6000 236.4000 474.4000 239.8000 ;
	    RECT 473.6000 235.8000 475.6000 236.4000 ;
	    RECT 465.2000 235.0000 466.0000 235.8000 ;
	    RECT 469.4000 235.2000 470.0000 235.8000 ;
	    RECT 468.6000 234.6000 472.2000 235.2000 ;
	    RECT 474.8000 235.0000 475.6000 235.8000 ;
	    RECT 468.6000 234.4000 469.4000 234.6000 ;
	    RECT 471.4000 234.4000 472.2000 234.6000 ;
	    RECT 458.8000 233.7000 461.2000 234.3000 ;
	    RECT 458.8000 233.6000 459.6000 233.7000 ;
	    RECT 455.6000 228.2000 458.0000 228.3000 ;
	    RECT 454.8000 227.7000 458.0000 228.2000 ;
	    RECT 454.8000 227.6000 456.4000 227.7000 ;
	    RECT 447.8000 226.8000 450.0000 227.4000 ;
	    RECT 449.2000 222.2000 450.0000 226.8000 ;
	    RECT 451.0000 226.4000 451.6000 227.6000 ;
	    RECT 454.8000 227.2000 455.6000 227.6000 ;
	    RECT 450.8000 222.2000 451.6000 226.4000 ;
	    RECT 452.6000 226.2000 456.2000 226.6000 ;
	    RECT 452.4000 226.0000 456.4000 226.2000 ;
	    RECT 452.4000 222.2000 453.2000 226.0000 ;
	    RECT 455.6000 222.2000 456.4000 226.0000 ;
	    RECT 457.2000 222.2000 458.0000 227.7000 ;
	    RECT 460.4000 231.2000 461.2000 233.7000 ;
	    RECT 464.4000 233.2000 465.8000 234.0000 ;
	    RECT 465.2000 232.2000 465.8000 233.2000 ;
	    RECT 467.4000 233.0000 469.6000 233.6000 ;
	    RECT 467.4000 232.8000 468.2000 233.0000 ;
	    RECT 465.2000 231.6000 467.6000 232.2000 ;
	    RECT 460.4000 230.6000 464.6000 231.2000 ;
	    RECT 460.4000 227.2000 461.2000 230.6000 ;
	    RECT 463.8000 230.4000 464.6000 230.6000 ;
	    RECT 462.2000 229.8000 463.0000 230.0000 ;
	    RECT 462.2000 229.2000 466.0000 229.8000 ;
	    RECT 465.2000 229.0000 466.0000 229.2000 ;
	    RECT 467.0000 228.4000 467.6000 231.6000 ;
	    RECT 469.0000 231.8000 469.6000 233.0000 ;
	    RECT 470.2000 233.0000 471.0000 233.2000 ;
	    RECT 474.8000 233.0000 475.6000 233.2000 ;
	    RECT 470.2000 232.4000 475.6000 233.0000 ;
	    RECT 469.0000 231.4000 473.8000 231.8000 ;
	    RECT 478.0000 231.4000 478.8000 239.8000 ;
	    RECT 479.6000 235.8000 480.4000 239.8000 ;
	    RECT 479.8000 235.6000 480.4000 235.8000 ;
	    RECT 482.8000 235.6000 483.6000 239.8000 ;
	    RECT 479.8000 235.0000 483.4000 235.6000 ;
	    RECT 479.8000 232.4000 480.4000 235.0000 ;
	    RECT 481.2000 232.8000 482.0000 234.4000 ;
	    RECT 486.8000 233.6000 487.6000 234.4000 ;
	    RECT 486.8000 232.4000 487.4000 233.6000 ;
	    RECT 488.2000 232.4000 489.0000 239.8000 ;
	    RECT 479.6000 231.6000 480.4000 232.4000 ;
	    RECT 486.0000 231.8000 487.4000 232.4000 ;
	    RECT 488.0000 231.8000 489.0000 232.4000 ;
	    RECT 486.0000 231.6000 486.8000 231.8000 ;
	    RECT 469.0000 231.2000 478.8000 231.4000 ;
	    RECT 473.0000 231.0000 478.8000 231.2000 ;
	    RECT 473.2000 230.8000 478.8000 231.0000 ;
	    RECT 471.6000 230.2000 472.4000 230.4000 ;
	    RECT 471.6000 229.6000 476.6000 230.2000 ;
	    RECT 475.8000 229.4000 476.6000 229.6000 ;
	    RECT 474.2000 228.4000 475.0000 228.6000 ;
	    RECT 479.8000 228.4000 480.4000 231.6000 ;
	    RECT 482.0000 229.6000 483.6000 230.4000 ;
	    RECT 486.0000 230.3000 486.8000 230.4000 ;
	    RECT 488.0000 230.3000 488.6000 231.8000 ;
	    RECT 486.0000 229.7000 488.6000 230.3000 ;
	    RECT 486.0000 229.6000 486.8000 229.7000 ;
	    RECT 488.0000 228.4000 488.6000 229.7000 ;
	    RECT 489.2000 228.8000 490.0000 230.4000 ;
	    RECT 467.0000 227.8000 478.0000 228.4000 ;
	    RECT 479.8000 228.2000 481.4000 228.4000 ;
	    RECT 479.8000 227.8000 481.6000 228.2000 ;
	    RECT 467.4000 227.6000 468.2000 227.8000 ;
	    RECT 460.4000 226.6000 464.2000 227.2000 ;
	    RECT 458.8000 224.8000 459.6000 226.4000 ;
	    RECT 460.4000 222.2000 461.2000 226.6000 ;
	    RECT 463.4000 226.4000 464.2000 226.6000 ;
	    RECT 473.2000 225.6000 473.8000 227.8000 ;
	    RECT 476.4000 227.6000 478.0000 227.8000 ;
	    RECT 471.4000 225.4000 472.2000 225.6000 ;
	    RECT 465.2000 224.2000 466.0000 225.0000 ;
	    RECT 469.4000 224.8000 472.2000 225.4000 ;
	    RECT 473.2000 224.8000 474.0000 225.6000 ;
	    RECT 469.4000 224.2000 470.0000 224.8000 ;
	    RECT 474.8000 224.2000 475.6000 225.0000 ;
	    RECT 464.6000 223.6000 466.0000 224.2000 ;
	    RECT 464.6000 222.2000 465.8000 223.6000 ;
	    RECT 469.2000 222.2000 470.0000 224.2000 ;
	    RECT 473.6000 223.6000 475.6000 224.2000 ;
	    RECT 473.6000 222.2000 474.4000 223.6000 ;
	    RECT 478.0000 222.2000 478.8000 227.0000 ;
	    RECT 480.8000 222.2000 481.6000 227.8000 ;
	    RECT 486.0000 227.6000 488.6000 228.4000 ;
	    RECT 490.8000 228.3000 491.6000 228.4000 ;
	    RECT 492.4000 228.3000 493.2000 239.8000 ;
	    RECT 495.6000 231.4000 496.4000 239.8000 ;
	    RECT 500.0000 236.4000 500.8000 239.8000 ;
	    RECT 498.8000 235.8000 500.8000 236.4000 ;
	    RECT 504.4000 235.8000 505.2000 239.8000 ;
	    RECT 508.6000 235.8000 509.8000 239.8000 ;
	    RECT 498.8000 235.0000 499.6000 235.8000 ;
	    RECT 504.4000 235.2000 505.0000 235.8000 ;
	    RECT 502.2000 234.6000 505.8000 235.2000 ;
	    RECT 508.4000 235.0000 509.2000 235.8000 ;
	    RECT 502.2000 234.4000 503.0000 234.6000 ;
	    RECT 505.0000 234.4000 505.8000 234.6000 ;
	    RECT 498.8000 233.0000 499.6000 233.2000 ;
	    RECT 503.4000 233.0000 504.2000 233.2000 ;
	    RECT 498.8000 232.4000 504.2000 233.0000 ;
	    RECT 504.8000 233.0000 507.0000 233.6000 ;
	    RECT 504.8000 231.8000 505.4000 233.0000 ;
	    RECT 506.2000 232.8000 507.0000 233.0000 ;
	    RECT 508.6000 233.2000 510.0000 234.0000 ;
	    RECT 508.6000 232.2000 509.2000 233.2000 ;
	    RECT 500.6000 231.4000 505.4000 231.8000 ;
	    RECT 495.6000 231.2000 505.4000 231.4000 ;
	    RECT 506.8000 231.6000 509.2000 232.2000 ;
	    RECT 495.6000 231.0000 501.4000 231.2000 ;
	    RECT 495.6000 230.8000 501.2000 231.0000 ;
	    RECT 502.0000 230.2000 502.8000 230.4000 ;
	    RECT 497.8000 229.6000 502.8000 230.2000 ;
	    RECT 497.8000 229.4000 498.6000 229.6000 ;
	    RECT 500.4000 229.4000 501.2000 229.6000 ;
	    RECT 499.4000 228.4000 500.2000 228.6000 ;
	    RECT 506.8000 228.4000 507.4000 231.6000 ;
	    RECT 513.2000 231.2000 514.0000 239.8000 ;
	    RECT 509.8000 230.6000 514.0000 231.2000 ;
	    RECT 509.8000 230.4000 510.6000 230.6000 ;
	    RECT 511.4000 229.8000 512.2000 230.0000 ;
	    RECT 508.4000 229.2000 512.2000 229.8000 ;
	    RECT 508.4000 229.0000 509.2000 229.2000 ;
	    RECT 490.8000 228.2000 493.2000 228.3000 ;
	    RECT 490.0000 227.7000 493.2000 228.2000 ;
	    RECT 490.0000 227.6000 491.6000 227.7000 ;
	    RECT 486.2000 226.2000 486.8000 227.6000 ;
	    RECT 490.0000 227.2000 490.8000 227.6000 ;
	    RECT 487.8000 226.2000 491.4000 226.6000 ;
	    RECT 486.0000 222.2000 486.8000 226.2000 ;
	    RECT 487.6000 226.0000 491.6000 226.2000 ;
	    RECT 487.6000 222.2000 488.4000 226.0000 ;
	    RECT 490.8000 222.2000 491.6000 226.0000 ;
	    RECT 492.4000 222.2000 493.2000 227.7000 ;
	    RECT 496.4000 227.8000 507.4000 228.4000 ;
	    RECT 496.4000 227.6000 498.0000 227.8000 ;
	    RECT 494.0000 224.8000 494.8000 226.4000 ;
	    RECT 495.6000 222.2000 496.4000 227.0000 ;
	    RECT 500.6000 225.6000 501.2000 227.8000 ;
	    RECT 506.2000 227.6000 507.0000 227.8000 ;
	    RECT 513.2000 227.2000 514.0000 230.6000 ;
	    RECT 510.2000 226.6000 514.0000 227.2000 ;
	    RECT 510.2000 226.4000 511.0000 226.6000 ;
	    RECT 498.8000 224.2000 499.6000 225.0000 ;
	    RECT 500.4000 224.8000 501.2000 225.6000 ;
	    RECT 502.2000 225.4000 503.0000 225.6000 ;
	    RECT 502.2000 224.8000 505.0000 225.4000 ;
	    RECT 504.4000 224.2000 505.0000 224.8000 ;
	    RECT 508.4000 224.2000 509.2000 225.0000 ;
	    RECT 498.8000 223.6000 500.8000 224.2000 ;
	    RECT 500.0000 222.2000 500.8000 223.6000 ;
	    RECT 504.4000 222.2000 505.2000 224.2000 ;
	    RECT 508.4000 223.6000 509.8000 224.2000 ;
	    RECT 508.6000 222.2000 509.8000 223.6000 ;
	    RECT 513.2000 222.2000 514.0000 226.6000 ;
	    RECT 4.4000 215.2000 5.2000 219.8000 ;
	    RECT 3.0000 214.6000 5.2000 215.2000 ;
	    RECT 6.0000 215.2000 6.8000 219.8000 ;
	    RECT 6.0000 214.6000 8.2000 215.2000 ;
	    RECT 3.0000 211.6000 3.6000 214.6000 ;
	    RECT 4.4000 211.6000 5.2000 213.2000 ;
	    RECT 7.6000 211.6000 8.2000 214.6000 ;
	    RECT 9.2000 212.4000 10.0000 219.8000 ;
	    RECT 10.8000 216.0000 11.6000 219.8000 ;
	    RECT 14.0000 216.0000 14.8000 219.8000 ;
	    RECT 10.8000 215.8000 14.8000 216.0000 ;
	    RECT 15.6000 215.8000 16.4000 219.8000 ;
	    RECT 11.0000 215.4000 14.6000 215.8000 ;
	    RECT 11.6000 214.4000 12.4000 214.8000 ;
	    RECT 15.6000 214.4000 16.2000 215.8000 ;
	    RECT 17.2000 215.4000 18.0000 219.8000 ;
	    RECT 21.4000 218.4000 22.6000 219.8000 ;
	    RECT 21.4000 217.8000 22.8000 218.4000 ;
	    RECT 26.0000 217.8000 26.8000 219.8000 ;
	    RECT 30.4000 218.4000 31.2000 219.8000 ;
	    RECT 30.4000 217.8000 32.4000 218.4000 ;
	    RECT 22.0000 217.0000 22.8000 217.8000 ;
	    RECT 26.2000 217.2000 26.8000 217.8000 ;
	    RECT 26.2000 216.6000 29.0000 217.2000 ;
	    RECT 28.2000 216.4000 29.0000 216.6000 ;
	    RECT 30.0000 215.6000 30.8000 217.2000 ;
	    RECT 31.6000 217.0000 32.4000 217.8000 ;
	    RECT 20.2000 215.4000 21.0000 215.6000 ;
	    RECT 17.2000 214.8000 21.0000 215.4000 ;
	    RECT 10.8000 213.8000 12.4000 214.4000 ;
	    RECT 10.8000 213.6000 11.6000 213.8000 ;
	    RECT 13.8000 213.6000 16.4000 214.4000 ;
	    RECT 2.4000 210.8000 3.6000 211.6000 ;
	    RECT 3.0000 210.2000 3.6000 210.8000 ;
	    RECT 7.6000 210.8000 8.8000 211.6000 ;
	    RECT 7.6000 210.2000 8.2000 210.8000 ;
	    RECT 9.4000 210.2000 10.0000 212.4000 ;
	    RECT 12.4000 211.6000 13.2000 213.2000 ;
	    RECT 13.8000 212.4000 14.4000 213.6000 ;
	    RECT 13.8000 211.6000 14.8000 212.4000 ;
	    RECT 13.8000 210.2000 14.4000 211.6000 ;
	    RECT 17.2000 211.4000 18.0000 214.8000 ;
	    RECT 24.2000 214.2000 25.0000 214.4000 ;
	    RECT 30.0000 214.2000 30.6000 215.6000 ;
	    RECT 34.8000 215.0000 35.6000 219.8000 ;
	    RECT 36.4000 215.8000 37.2000 219.8000 ;
	    RECT 38.0000 216.0000 38.8000 219.8000 ;
	    RECT 41.2000 216.0000 42.0000 219.8000 ;
	    RECT 38.0000 215.8000 42.0000 216.0000 ;
	    RECT 36.6000 214.4000 37.2000 215.8000 ;
	    RECT 38.2000 215.4000 41.8000 215.8000 ;
	    RECT 42.8000 215.2000 43.6000 219.8000 ;
	    RECT 40.4000 214.4000 41.2000 214.8000 ;
	    RECT 42.8000 214.6000 45.0000 215.2000 ;
	    RECT 33.2000 214.2000 34.8000 214.4000 ;
	    RECT 23.8000 213.6000 34.8000 214.2000 ;
	    RECT 36.4000 213.6000 39.0000 214.4000 ;
	    RECT 40.4000 213.8000 42.0000 214.4000 ;
	    RECT 41.2000 213.6000 42.0000 213.8000 ;
	    RECT 22.0000 212.8000 22.8000 213.0000 ;
	    RECT 19.0000 212.2000 22.8000 212.8000 ;
	    RECT 19.0000 212.0000 19.8000 212.2000 ;
	    RECT 20.6000 211.4000 21.4000 211.6000 ;
	    RECT 17.2000 210.8000 21.4000 211.4000 ;
	    RECT 15.6000 210.2000 16.4000 210.4000 ;
	    RECT 3.0000 209.6000 5.2000 210.2000 ;
	    RECT 4.4000 202.2000 5.2000 209.6000 ;
	    RECT 6.0000 209.6000 8.2000 210.2000 ;
	    RECT 6.0000 202.2000 6.8000 209.6000 ;
	    RECT 9.2000 202.2000 10.0000 210.2000 ;
	    RECT 13.4000 209.6000 14.4000 210.2000 ;
	    RECT 15.0000 209.6000 16.4000 210.2000 ;
	    RECT 13.4000 202.2000 14.2000 209.6000 ;
	    RECT 15.0000 208.4000 15.6000 209.6000 ;
	    RECT 14.8000 208.3000 15.6000 208.4000 ;
	    RECT 17.2000 208.3000 18.0000 210.8000 ;
	    RECT 23.8000 210.4000 24.4000 213.6000 ;
	    RECT 31.0000 213.4000 31.8000 213.6000 ;
	    RECT 30.0000 212.4000 30.8000 212.6000 ;
	    RECT 32.6000 212.4000 33.4000 212.6000 ;
	    RECT 28.4000 211.8000 33.4000 212.4000 ;
	    RECT 36.4000 212.3000 37.2000 212.4000 ;
	    RECT 38.4000 212.3000 39.0000 213.6000 ;
	    RECT 28.4000 211.6000 29.2000 211.8000 ;
	    RECT 36.4000 211.7000 39.0000 212.3000 ;
	    RECT 36.4000 211.6000 37.2000 211.7000 ;
	    RECT 30.0000 211.0000 35.6000 211.2000 ;
	    RECT 29.8000 210.8000 35.6000 211.0000 ;
	    RECT 22.0000 209.8000 24.4000 210.4000 ;
	    RECT 25.8000 210.6000 35.6000 210.8000 ;
	    RECT 25.8000 210.2000 30.6000 210.6000 ;
	    RECT 22.0000 208.8000 22.6000 209.8000 ;
	    RECT 14.8000 207.7000 18.0000 208.3000 ;
	    RECT 21.2000 208.0000 22.6000 208.8000 ;
	    RECT 24.2000 209.0000 25.0000 209.2000 ;
	    RECT 25.8000 209.0000 26.4000 210.2000 ;
	    RECT 24.2000 208.4000 26.4000 209.0000 ;
	    RECT 27.0000 209.0000 32.4000 209.6000 ;
	    RECT 27.0000 208.8000 27.8000 209.0000 ;
	    RECT 31.6000 208.8000 32.4000 209.0000 ;
	    RECT 14.8000 207.6000 15.6000 207.7000 ;
	    RECT 17.2000 202.2000 18.0000 207.7000 ;
	    RECT 25.4000 207.4000 26.2000 207.6000 ;
	    RECT 28.2000 207.4000 29.0000 207.6000 ;
	    RECT 22.0000 206.2000 22.8000 207.0000 ;
	    RECT 25.4000 206.8000 29.0000 207.4000 ;
	    RECT 26.2000 206.2000 26.8000 206.8000 ;
	    RECT 31.6000 206.2000 32.4000 207.0000 ;
	    RECT 21.4000 202.2000 22.6000 206.2000 ;
	    RECT 26.0000 202.2000 26.8000 206.2000 ;
	    RECT 30.4000 205.6000 32.4000 206.2000 ;
	    RECT 30.4000 202.2000 31.2000 205.6000 ;
	    RECT 34.8000 202.2000 35.6000 210.6000 ;
	    RECT 36.4000 210.2000 37.2000 210.4000 ;
	    RECT 38.4000 210.2000 39.0000 211.7000 ;
	    RECT 39.6000 211.6000 40.4000 213.2000 ;
	    RECT 41.2000 212.3000 42.0000 212.4000 ;
	    RECT 42.8000 212.3000 43.6000 213.2000 ;
	    RECT 41.2000 211.7000 43.6000 212.3000 ;
	    RECT 41.2000 211.6000 42.0000 211.7000 ;
	    RECT 42.8000 211.6000 43.6000 211.7000 ;
	    RECT 44.4000 211.6000 45.0000 214.6000 ;
	    RECT 46.0000 212.4000 46.8000 219.8000 ;
	    RECT 47.6000 215.6000 48.4000 219.8000 ;
	    RECT 49.2000 216.0000 50.0000 219.8000 ;
	    RECT 52.4000 216.0000 53.2000 219.8000 ;
	    RECT 55.6000 217.8000 56.4000 219.8000 ;
	    RECT 60.4000 217.8000 61.2000 219.8000 ;
	    RECT 49.2000 215.8000 53.2000 216.0000 ;
	    RECT 54.0000 216.3000 54.8000 216.4000 ;
	    RECT 55.6000 216.3000 56.2000 217.8000 ;
	    RECT 57.2000 216.3000 58.0000 217.2000 ;
	    RECT 58.8000 216.3000 59.6000 217.2000 ;
	    RECT 47.8000 214.4000 48.4000 215.6000 ;
	    RECT 49.4000 215.4000 53.0000 215.8000 ;
	    RECT 54.0000 215.7000 56.3000 216.3000 ;
	    RECT 57.2000 215.7000 59.6000 216.3000 ;
	    RECT 54.0000 215.6000 54.8000 215.7000 ;
	    RECT 51.6000 214.4000 52.4000 214.8000 ;
	    RECT 55.6000 214.4000 56.2000 215.7000 ;
	    RECT 57.2000 215.6000 58.0000 215.7000 ;
	    RECT 58.8000 215.6000 59.6000 215.7000 ;
	    RECT 60.6000 214.4000 61.2000 217.8000 ;
	    RECT 62.0000 216.3000 62.8000 216.4000 ;
	    RECT 63.6000 216.3000 64.4000 219.8000 ;
	    RECT 62.0000 215.7000 64.4000 216.3000 ;
	    RECT 62.0000 215.6000 62.8000 215.7000 ;
	    RECT 47.6000 213.6000 50.2000 214.4000 ;
	    RECT 51.6000 213.8000 53.2000 214.4000 ;
	    RECT 52.4000 213.6000 53.2000 213.8000 ;
	    RECT 55.6000 213.6000 56.4000 214.4000 ;
	    RECT 57.2000 214.3000 58.0000 214.4000 ;
	    RECT 60.4000 214.3000 61.2000 214.4000 ;
	    RECT 57.2000 213.7000 61.2000 214.3000 ;
	    RECT 57.2000 213.6000 58.0000 213.7000 ;
	    RECT 60.4000 213.6000 61.2000 213.7000 ;
	    RECT 44.4000 210.8000 45.6000 211.6000 ;
	    RECT 44.4000 210.2000 45.0000 210.8000 ;
	    RECT 46.2000 210.2000 46.8000 212.4000 ;
	    RECT 36.4000 209.6000 37.8000 210.2000 ;
	    RECT 38.4000 209.6000 39.4000 210.2000 ;
	    RECT 37.2000 208.4000 37.8000 209.6000 ;
	    RECT 37.2000 207.6000 38.0000 208.4000 ;
	    RECT 38.6000 202.2000 39.4000 209.6000 ;
	    RECT 42.8000 209.6000 45.0000 210.2000 ;
	    RECT 42.8000 202.2000 43.6000 209.6000 ;
	    RECT 46.0000 208.3000 46.8000 210.2000 ;
	    RECT 47.6000 210.2000 48.4000 210.4000 ;
	    RECT 49.6000 210.2000 50.2000 213.6000 ;
	    RECT 50.8000 211.6000 51.6000 213.2000 ;
	    RECT 54.0000 210.8000 54.8000 212.4000 ;
	    RECT 55.6000 210.2000 56.2000 213.6000 ;
	    RECT 60.6000 210.2000 61.2000 213.6000 ;
	    RECT 63.6000 212.4000 64.4000 215.7000 ;
	    RECT 66.8000 215.2000 67.6000 219.8000 ;
	    RECT 65.4000 214.6000 67.6000 215.2000 ;
	    RECT 62.0000 210.8000 62.8000 212.4000 ;
	    RECT 63.6000 210.2000 64.2000 212.4000 ;
	    RECT 65.4000 211.6000 66.0000 214.6000 ;
	    RECT 64.8000 210.8000 66.0000 211.6000 ;
	    RECT 65.4000 210.2000 66.0000 210.8000 ;
	    RECT 68.4000 212.4000 69.2000 219.8000 ;
	    RECT 71.6000 215.2000 72.4000 219.8000 ;
	    RECT 70.2000 214.6000 72.4000 215.2000 ;
	    RECT 73.2000 215.0000 74.0000 219.8000 ;
	    RECT 77.6000 218.4000 78.4000 219.8000 ;
	    RECT 76.4000 217.8000 78.4000 218.4000 ;
	    RECT 82.0000 217.8000 82.8000 219.8000 ;
	    RECT 86.2000 218.4000 87.4000 219.8000 ;
	    RECT 86.0000 217.8000 87.4000 218.4000 ;
	    RECT 76.4000 217.0000 77.2000 217.8000 ;
	    RECT 82.0000 217.2000 82.6000 217.8000 ;
	    RECT 78.0000 215.6000 78.8000 217.2000 ;
	    RECT 79.8000 216.6000 82.6000 217.2000 ;
	    RECT 86.0000 217.0000 86.8000 217.8000 ;
	    RECT 79.8000 216.4000 80.6000 216.6000 ;
	    RECT 68.4000 210.2000 69.0000 212.4000 ;
	    RECT 70.2000 211.6000 70.8000 214.6000 ;
	    RECT 74.0000 214.2000 75.6000 214.4000 ;
	    RECT 78.2000 214.2000 78.8000 215.6000 ;
	    RECT 87.8000 215.4000 88.6000 215.6000 ;
	    RECT 90.8000 215.4000 91.6000 219.8000 ;
	    RECT 95.0000 218.4000 95.8000 219.8000 ;
	    RECT 94.0000 217.6000 95.8000 218.4000 ;
	    RECT 95.0000 216.4000 95.8000 217.6000 ;
	    RECT 99.8000 216.4000 100.6000 219.8000 ;
	    RECT 87.8000 214.8000 91.6000 215.4000 ;
	    RECT 94.0000 215.8000 95.8000 216.4000 ;
	    RECT 98.8000 215.8000 100.6000 216.4000 ;
	    RECT 102.0000 215.8000 102.8000 219.8000 ;
	    RECT 103.6000 216.0000 104.4000 219.8000 ;
	    RECT 106.8000 216.0000 107.6000 219.8000 ;
	    RECT 103.6000 215.8000 107.6000 216.0000 ;
	    RECT 114.8000 219.2000 118.8000 219.8000 ;
	    RECT 114.8000 215.8000 115.6000 219.2000 ;
	    RECT 116.4000 215.8000 117.2000 218.6000 ;
	    RECT 118.0000 216.0000 118.8000 219.2000 ;
	    RECT 121.2000 216.0000 122.0000 219.8000 ;
	    RECT 118.0000 215.8000 122.0000 216.0000 ;
	    RECT 122.8000 215.8000 123.6000 219.8000 ;
	    RECT 124.4000 216.0000 125.2000 219.8000 ;
	    RECT 127.6000 216.0000 128.4000 219.8000 ;
	    RECT 124.4000 215.8000 128.4000 216.0000 ;
	    RECT 79.6000 214.2000 80.4000 214.4000 ;
	    RECT 83.8000 214.2000 84.6000 214.4000 ;
	    RECT 74.0000 213.6000 85.0000 214.2000 ;
	    RECT 77.0000 213.4000 77.8000 213.6000 ;
	    RECT 71.6000 211.6000 72.4000 213.2000 ;
	    RECT 75.4000 212.4000 76.2000 212.6000 ;
	    RECT 75.4000 212.3000 80.4000 212.4000 ;
	    RECT 81.2000 212.3000 82.0000 212.4000 ;
	    RECT 75.4000 211.8000 82.0000 212.3000 ;
	    RECT 79.6000 211.7000 82.0000 211.8000 ;
	    RECT 79.6000 211.6000 80.4000 211.7000 ;
	    RECT 81.2000 211.6000 82.0000 211.7000 ;
	    RECT 69.6000 210.8000 70.8000 211.6000 ;
	    RECT 70.2000 210.2000 70.8000 210.8000 ;
	    RECT 73.2000 211.0000 78.8000 211.2000 ;
	    RECT 73.2000 210.8000 79.0000 211.0000 ;
	    RECT 73.2000 210.6000 83.0000 210.8000 ;
	    RECT 47.6000 209.6000 49.0000 210.2000 ;
	    RECT 49.6000 209.6000 50.6000 210.2000 ;
	    RECT 48.4000 208.4000 49.0000 209.6000 ;
	    RECT 48.4000 208.3000 49.2000 208.4000 ;
	    RECT 46.0000 207.7000 49.2000 208.3000 ;
	    RECT 46.0000 202.2000 46.8000 207.7000 ;
	    RECT 48.4000 207.6000 49.2000 207.7000 ;
	    RECT 49.8000 202.2000 50.6000 209.6000 ;
	    RECT 54.6000 209.4000 56.4000 210.2000 ;
	    RECT 60.4000 209.4000 62.2000 210.2000 ;
	    RECT 54.6000 202.2000 55.4000 209.4000 ;
	    RECT 61.4000 202.2000 62.2000 209.4000 ;
	    RECT 63.6000 202.2000 64.4000 210.2000 ;
	    RECT 65.4000 209.6000 67.6000 210.2000 ;
	    RECT 66.8000 202.2000 67.6000 209.6000 ;
	    RECT 68.4000 202.2000 69.2000 210.2000 ;
	    RECT 70.2000 209.6000 72.4000 210.2000 ;
	    RECT 71.6000 202.2000 72.4000 209.6000 ;
	    RECT 73.2000 202.2000 74.0000 210.6000 ;
	    RECT 78.2000 210.2000 83.0000 210.6000 ;
	    RECT 76.4000 209.0000 81.8000 209.6000 ;
	    RECT 76.4000 208.8000 77.2000 209.0000 ;
	    RECT 81.0000 208.8000 81.8000 209.0000 ;
	    RECT 82.4000 209.0000 83.0000 210.2000 ;
	    RECT 84.4000 210.4000 85.0000 213.6000 ;
	    RECT 86.0000 212.8000 86.8000 213.0000 ;
	    RECT 86.0000 212.2000 89.8000 212.8000 ;
	    RECT 89.0000 212.0000 89.8000 212.2000 ;
	    RECT 87.4000 211.4000 88.2000 211.6000 ;
	    RECT 90.8000 211.4000 91.6000 214.8000 ;
	    RECT 92.4000 213.6000 93.2000 215.2000 ;
	    RECT 87.4000 210.8000 91.6000 211.4000 ;
	    RECT 84.4000 209.8000 86.8000 210.4000 ;
	    RECT 83.8000 209.0000 84.6000 209.2000 ;
	    RECT 82.4000 208.4000 84.6000 209.0000 ;
	    RECT 86.2000 208.8000 86.8000 209.8000 ;
	    RECT 86.2000 208.0000 87.6000 208.8000 ;
	    RECT 79.8000 207.4000 80.6000 207.6000 ;
	    RECT 82.6000 207.4000 83.4000 207.6000 ;
	    RECT 76.4000 206.2000 77.2000 207.0000 ;
	    RECT 79.8000 206.8000 83.4000 207.4000 ;
	    RECT 82.0000 206.2000 82.6000 206.8000 ;
	    RECT 86.0000 206.2000 86.8000 207.0000 ;
	    RECT 76.4000 205.6000 78.4000 206.2000 ;
	    RECT 77.6000 202.2000 78.4000 205.6000 ;
	    RECT 82.0000 202.2000 82.8000 206.2000 ;
	    RECT 86.2000 202.2000 87.4000 206.2000 ;
	    RECT 90.8000 202.2000 91.6000 210.8000 ;
	    RECT 94.0000 202.2000 94.8000 215.8000 ;
	    RECT 97.2000 213.6000 98.0000 215.2000 ;
	    RECT 98.8000 212.3000 99.6000 215.8000 ;
	    RECT 102.2000 214.4000 102.8000 215.8000 ;
	    RECT 103.8000 215.4000 107.4000 215.8000 ;
	    RECT 106.0000 214.4000 106.8000 214.8000 ;
	    RECT 116.4000 214.4000 117.0000 215.8000 ;
	    RECT 118.2000 215.4000 121.8000 215.8000 ;
	    RECT 120.4000 214.4000 121.2000 214.8000 ;
	    RECT 123.0000 214.4000 123.6000 215.8000 ;
	    RECT 124.6000 215.4000 128.2000 215.8000 ;
	    RECT 129.2000 215.0000 130.0000 219.8000 ;
	    RECT 133.6000 218.4000 134.4000 219.8000 ;
	    RECT 132.4000 217.8000 134.4000 218.4000 ;
	    RECT 138.0000 217.8000 138.8000 219.8000 ;
	    RECT 142.2000 218.4000 143.4000 219.8000 ;
	    RECT 142.0000 217.8000 143.4000 218.4000 ;
	    RECT 132.4000 217.0000 133.2000 217.8000 ;
	    RECT 138.0000 217.2000 138.6000 217.8000 ;
	    RECT 134.0000 216.4000 134.8000 217.2000 ;
	    RECT 135.8000 216.6000 138.6000 217.2000 ;
	    RECT 142.0000 217.0000 142.8000 217.8000 ;
	    RECT 135.8000 216.4000 136.6000 216.6000 ;
	    RECT 126.8000 214.4000 127.6000 214.8000 ;
	    RECT 100.4000 214.3000 101.2000 214.4000 ;
	    RECT 102.0000 214.3000 104.6000 214.4000 ;
	    RECT 100.4000 213.7000 104.6000 214.3000 ;
	    RECT 106.0000 213.8000 107.6000 214.4000 ;
	    RECT 100.4000 213.6000 101.2000 213.7000 ;
	    RECT 102.0000 213.6000 104.6000 213.7000 ;
	    RECT 106.8000 213.6000 107.6000 213.8000 ;
	    RECT 98.8000 211.7000 102.7000 212.3000 ;
	    RECT 95.6000 208.8000 96.4000 210.4000 ;
	    RECT 98.8000 202.2000 99.6000 211.7000 ;
	    RECT 102.1000 210.4000 102.7000 211.7000 ;
	    RECT 100.4000 208.8000 101.2000 210.4000 ;
	    RECT 102.0000 210.2000 102.8000 210.4000 ;
	    RECT 104.0000 210.2000 104.6000 213.6000 ;
	    RECT 105.2000 211.6000 106.0000 213.2000 ;
	    RECT 114.8000 212.8000 115.6000 214.4000 ;
	    RECT 116.4000 213.8000 118.8000 214.4000 ;
	    RECT 120.4000 214.3000 122.0000 214.4000 ;
	    RECT 122.8000 214.3000 125.4000 214.4000 ;
	    RECT 120.4000 213.8000 125.4000 214.3000 ;
	    RECT 126.8000 213.8000 128.4000 214.4000 ;
	    RECT 118.0000 213.6000 118.8000 213.8000 ;
	    RECT 121.2000 213.7000 125.4000 213.8000 ;
	    RECT 121.2000 213.6000 122.0000 213.7000 ;
	    RECT 122.8000 213.6000 125.4000 213.7000 ;
	    RECT 127.6000 213.6000 128.4000 213.8000 ;
	    RECT 130.0000 214.2000 131.6000 214.4000 ;
	    RECT 134.2000 214.2000 134.8000 216.4000 ;
	    RECT 143.8000 215.4000 144.6000 215.6000 ;
	    RECT 146.8000 215.4000 147.6000 219.8000 ;
	    RECT 143.8000 214.8000 147.6000 215.4000 ;
	    RECT 139.8000 214.2000 140.6000 214.4000 ;
	    RECT 130.0000 213.6000 141.0000 214.2000 ;
	    RECT 116.4000 211.6000 117.2000 213.2000 ;
	    RECT 118.2000 210.2000 118.8000 213.6000 ;
	    RECT 119.6000 211.6000 120.4000 213.2000 ;
	    RECT 122.8000 210.2000 123.6000 210.4000 ;
	    RECT 124.8000 210.2000 125.4000 213.6000 ;
	    RECT 133.0000 213.4000 133.8000 213.6000 ;
	    RECT 126.0000 211.6000 126.8000 213.2000 ;
	    RECT 131.4000 212.4000 132.2000 212.6000 ;
	    RECT 131.4000 211.8000 136.4000 212.4000 ;
	    RECT 135.6000 211.6000 136.4000 211.8000 ;
	    RECT 129.2000 211.0000 134.8000 211.2000 ;
	    RECT 129.2000 210.8000 135.0000 211.0000 ;
	    RECT 129.2000 210.6000 139.0000 210.8000 ;
	    RECT 102.0000 209.6000 103.4000 210.2000 ;
	    RECT 104.0000 209.6000 105.0000 210.2000 ;
	    RECT 102.8000 208.4000 103.4000 209.6000 ;
	    RECT 102.8000 207.6000 103.6000 208.4000 ;
	    RECT 104.2000 202.2000 105.0000 209.6000 ;
	    RECT 117.4000 202.2000 119.4000 210.2000 ;
	    RECT 122.8000 209.6000 124.2000 210.2000 ;
	    RECT 124.8000 209.6000 125.8000 210.2000 ;
	    RECT 123.6000 208.4000 124.2000 209.6000 ;
	    RECT 123.6000 207.6000 124.4000 208.4000 ;
	    RECT 125.0000 202.2000 125.8000 209.6000 ;
	    RECT 129.2000 202.2000 130.0000 210.6000 ;
	    RECT 134.2000 210.2000 139.0000 210.6000 ;
	    RECT 132.4000 209.0000 137.8000 209.6000 ;
	    RECT 132.4000 208.8000 133.2000 209.0000 ;
	    RECT 137.0000 208.8000 137.8000 209.0000 ;
	    RECT 138.4000 209.0000 139.0000 210.2000 ;
	    RECT 140.4000 210.4000 141.0000 213.6000 ;
	    RECT 142.0000 212.8000 142.8000 213.0000 ;
	    RECT 142.0000 212.2000 145.8000 212.8000 ;
	    RECT 145.0000 212.0000 145.8000 212.2000 ;
	    RECT 143.4000 211.4000 144.2000 211.6000 ;
	    RECT 146.8000 211.4000 147.6000 214.8000 ;
	    RECT 150.0000 217.8000 150.8000 219.8000 ;
	    RECT 150.0000 214.4000 150.6000 217.8000 ;
	    RECT 151.6000 215.6000 152.4000 217.2000 ;
	    RECT 157.0000 216.0000 157.8000 219.0000 ;
	    RECT 161.2000 217.0000 162.0000 219.0000 ;
	    RECT 156.2000 215.4000 157.8000 216.0000 ;
	    RECT 156.2000 215.0000 157.0000 215.4000 ;
	    RECT 156.2000 214.4000 156.8000 215.0000 ;
	    RECT 161.4000 214.8000 162.0000 217.0000 ;
	    RECT 150.0000 213.6000 150.8000 214.4000 ;
	    RECT 154.8000 213.6000 156.8000 214.4000 ;
	    RECT 157.8000 214.2000 162.0000 214.8000 ;
	    RECT 157.8000 213.8000 158.8000 214.2000 ;
	    RECT 143.4000 210.8000 147.6000 211.4000 ;
	    RECT 148.4000 210.8000 149.2000 212.4000 ;
	    RECT 140.4000 209.8000 142.8000 210.4000 ;
	    RECT 139.8000 209.0000 140.6000 209.2000 ;
	    RECT 138.4000 208.4000 140.6000 209.0000 ;
	    RECT 142.2000 208.8000 142.8000 209.8000 ;
	    RECT 142.2000 208.0000 143.6000 208.8000 ;
	    RECT 135.8000 207.4000 136.6000 207.6000 ;
	    RECT 138.6000 207.4000 139.4000 207.6000 ;
	    RECT 132.4000 206.2000 133.2000 207.0000 ;
	    RECT 135.8000 206.8000 139.4000 207.4000 ;
	    RECT 138.0000 206.2000 138.6000 206.8000 ;
	    RECT 142.0000 206.2000 142.8000 207.0000 ;
	    RECT 132.4000 205.6000 134.4000 206.2000 ;
	    RECT 133.6000 202.2000 134.4000 205.6000 ;
	    RECT 138.0000 202.2000 138.8000 206.2000 ;
	    RECT 142.2000 202.2000 143.4000 206.2000 ;
	    RECT 146.8000 202.2000 147.6000 210.8000 ;
	    RECT 150.0000 210.2000 150.6000 213.6000 ;
	    RECT 154.8000 210.8000 155.6000 212.4000 ;
	    RECT 149.0000 209.4000 150.8000 210.2000 ;
	    RECT 156.2000 209.8000 156.8000 213.6000 ;
	    RECT 157.4000 213.0000 158.8000 213.8000 ;
	    RECT 158.2000 211.0000 158.8000 213.0000 ;
	    RECT 159.6000 211.6000 160.4000 213.2000 ;
	    RECT 161.2000 211.6000 162.0000 213.2000 ;
	    RECT 162.8000 212.4000 163.6000 219.8000 ;
	    RECT 166.0000 215.2000 166.8000 219.8000 ;
	    RECT 164.6000 214.6000 166.8000 215.2000 ;
	    RECT 167.6000 215.0000 168.4000 219.8000 ;
	    RECT 172.0000 218.4000 172.8000 219.8000 ;
	    RECT 170.8000 217.8000 172.8000 218.4000 ;
	    RECT 176.4000 217.8000 177.2000 219.8000 ;
	    RECT 180.6000 218.4000 181.8000 219.8000 ;
	    RECT 180.4000 217.8000 181.8000 218.4000 ;
	    RECT 170.8000 217.0000 171.6000 217.8000 ;
	    RECT 176.4000 217.2000 177.0000 217.8000 ;
	    RECT 172.4000 216.4000 173.2000 217.2000 ;
	    RECT 174.2000 216.6000 177.0000 217.2000 ;
	    RECT 180.4000 217.0000 181.2000 217.8000 ;
	    RECT 174.2000 216.4000 175.0000 216.6000 ;
	    RECT 158.2000 210.4000 162.0000 211.0000 ;
	    RECT 149.0000 208.4000 149.8000 209.4000 ;
	    RECT 156.2000 209.2000 157.8000 209.8000 ;
	    RECT 148.4000 207.6000 149.8000 208.4000 ;
	    RECT 149.0000 202.2000 149.8000 207.6000 ;
	    RECT 157.0000 204.4000 157.8000 209.2000 ;
	    RECT 161.4000 207.0000 162.0000 210.4000 ;
	    RECT 156.4000 203.6000 157.8000 204.4000 ;
	    RECT 157.0000 202.2000 157.8000 203.6000 ;
	    RECT 161.2000 203.0000 162.0000 207.0000 ;
	    RECT 162.8000 210.2000 163.4000 212.4000 ;
	    RECT 164.6000 211.6000 165.2000 214.6000 ;
	    RECT 168.4000 214.2000 170.0000 214.4000 ;
	    RECT 172.6000 214.2000 173.2000 216.4000 ;
	    RECT 182.2000 215.4000 183.0000 215.6000 ;
	    RECT 185.2000 215.4000 186.0000 219.8000 ;
	    RECT 182.2000 214.8000 186.0000 215.4000 ;
	    RECT 178.2000 214.2000 179.0000 214.4000 ;
	    RECT 168.4000 213.6000 179.4000 214.2000 ;
	    RECT 171.4000 213.4000 172.2000 213.6000 ;
	    RECT 169.8000 212.4000 170.6000 212.6000 ;
	    RECT 169.8000 211.8000 174.8000 212.4000 ;
	    RECT 174.0000 211.6000 174.8000 211.8000 ;
	    RECT 164.0000 210.8000 165.2000 211.6000 ;
	    RECT 164.6000 210.2000 165.2000 210.8000 ;
	    RECT 167.6000 211.0000 173.2000 211.2000 ;
	    RECT 167.6000 210.8000 173.4000 211.0000 ;
	    RECT 167.6000 210.6000 177.4000 210.8000 ;
	    RECT 162.8000 202.2000 163.6000 210.2000 ;
	    RECT 164.6000 209.6000 166.8000 210.2000 ;
	    RECT 166.0000 202.2000 166.8000 209.6000 ;
	    RECT 167.6000 202.2000 168.4000 210.6000 ;
	    RECT 172.6000 210.2000 177.4000 210.6000 ;
	    RECT 170.8000 209.0000 176.2000 209.6000 ;
	    RECT 170.8000 208.8000 171.6000 209.0000 ;
	    RECT 175.4000 208.8000 176.2000 209.0000 ;
	    RECT 176.8000 209.0000 177.4000 210.2000 ;
	    RECT 178.8000 210.4000 179.4000 213.6000 ;
	    RECT 180.4000 212.8000 181.2000 213.0000 ;
	    RECT 180.4000 212.2000 184.2000 212.8000 ;
	    RECT 183.4000 212.0000 184.2000 212.2000 ;
	    RECT 181.8000 211.4000 182.6000 211.6000 ;
	    RECT 185.2000 211.4000 186.0000 214.8000 ;
	    RECT 181.8000 210.8000 186.0000 211.4000 ;
	    RECT 178.8000 209.8000 181.2000 210.4000 ;
	    RECT 178.2000 209.0000 179.0000 209.2000 ;
	    RECT 176.8000 208.4000 179.0000 209.0000 ;
	    RECT 180.6000 208.8000 181.2000 209.8000 ;
	    RECT 180.6000 208.0000 182.0000 208.8000 ;
	    RECT 174.2000 207.4000 175.0000 207.6000 ;
	    RECT 177.0000 207.4000 177.8000 207.6000 ;
	    RECT 170.8000 206.2000 171.6000 207.0000 ;
	    RECT 174.2000 206.8000 177.8000 207.4000 ;
	    RECT 176.4000 206.2000 177.0000 206.8000 ;
	    RECT 180.4000 206.2000 181.2000 207.0000 ;
	    RECT 170.8000 205.6000 172.8000 206.2000 ;
	    RECT 172.0000 202.2000 172.8000 205.6000 ;
	    RECT 176.4000 202.2000 177.2000 206.2000 ;
	    RECT 180.6000 202.2000 181.8000 206.2000 ;
	    RECT 185.2000 202.2000 186.0000 210.8000 ;
	    RECT 186.8000 212.4000 187.6000 219.8000 ;
	    RECT 190.0000 215.2000 190.8000 219.8000 ;
	    RECT 188.6000 214.6000 190.8000 215.2000 ;
	    RECT 191.6000 215.2000 192.4000 219.8000 ;
	    RECT 191.6000 214.6000 193.8000 215.2000 ;
	    RECT 186.8000 210.2000 187.4000 212.4000 ;
	    RECT 188.6000 211.6000 189.2000 214.6000 ;
	    RECT 190.0000 211.6000 190.8000 213.2000 ;
	    RECT 193.2000 211.6000 193.8000 214.6000 ;
	    RECT 194.8000 212.4000 195.6000 219.8000 ;
	    RECT 199.0000 216.4000 199.8000 219.8000 ;
	    RECT 198.0000 215.8000 199.8000 216.4000 ;
	    RECT 201.2000 215.8000 202.0000 219.8000 ;
	    RECT 202.8000 216.0000 203.6000 219.8000 ;
	    RECT 206.0000 216.0000 206.8000 219.8000 ;
	    RECT 209.2000 217.6000 210.0000 219.8000 ;
	    RECT 202.8000 215.8000 206.8000 216.0000 ;
	    RECT 196.4000 213.6000 197.2000 215.2000 ;
	    RECT 188.0000 210.8000 189.2000 211.6000 ;
	    RECT 188.6000 210.2000 189.2000 210.8000 ;
	    RECT 193.2000 210.8000 194.4000 211.6000 ;
	    RECT 193.2000 210.2000 193.8000 210.8000 ;
	    RECT 195.0000 210.2000 195.6000 212.4000 ;
	    RECT 186.8000 202.2000 187.6000 210.2000 ;
	    RECT 188.6000 209.6000 190.8000 210.2000 ;
	    RECT 190.0000 202.2000 190.8000 209.6000 ;
	    RECT 191.6000 209.6000 193.8000 210.2000 ;
	    RECT 191.6000 202.2000 192.4000 209.6000 ;
	    RECT 194.8000 202.2000 195.6000 210.2000 ;
	    RECT 198.0000 212.3000 198.8000 215.8000 ;
	    RECT 201.4000 214.4000 202.0000 215.8000 ;
	    RECT 203.0000 215.4000 206.6000 215.8000 ;
	    RECT 207.6000 215.6000 208.4000 217.2000 ;
	    RECT 205.2000 214.4000 206.0000 214.8000 ;
	    RECT 209.4000 214.4000 210.0000 217.6000 ;
	    RECT 215.0000 216.4000 215.8000 219.8000 ;
	    RECT 214.0000 215.8000 215.8000 216.4000 ;
	    RECT 217.2000 215.8000 218.0000 219.8000 ;
	    RECT 218.8000 216.0000 219.6000 219.8000 ;
	    RECT 222.0000 216.0000 222.8000 219.8000 ;
	    RECT 218.8000 215.8000 222.8000 216.0000 ;
	    RECT 199.6000 214.3000 200.4000 214.4000 ;
	    RECT 201.2000 214.3000 203.8000 214.4000 ;
	    RECT 199.6000 213.7000 203.8000 214.3000 ;
	    RECT 205.2000 213.8000 206.8000 214.4000 ;
	    RECT 199.6000 213.6000 200.4000 213.7000 ;
	    RECT 201.2000 213.6000 203.8000 213.7000 ;
	    RECT 206.0000 213.6000 206.8000 213.8000 ;
	    RECT 209.2000 213.6000 210.0000 214.4000 ;
	    RECT 212.4000 213.6000 213.2000 215.2000 ;
	    RECT 198.0000 211.7000 201.9000 212.3000 ;
	    RECT 198.0000 202.2000 198.8000 211.7000 ;
	    RECT 201.3000 210.4000 201.9000 211.7000 ;
	    RECT 199.6000 208.8000 200.4000 210.4000 ;
	    RECT 201.2000 210.2000 202.0000 210.4000 ;
	    RECT 203.2000 210.2000 203.8000 213.6000 ;
	    RECT 204.4000 211.6000 205.2000 213.2000 ;
	    RECT 209.4000 210.2000 210.0000 213.6000 ;
	    RECT 210.8000 210.8000 211.6000 212.4000 ;
	    RECT 214.0000 212.3000 214.8000 215.8000 ;
	    RECT 217.4000 214.4000 218.0000 215.8000 ;
	    RECT 219.0000 215.4000 222.6000 215.8000 ;
	    RECT 223.6000 215.0000 224.4000 219.8000 ;
	    RECT 228.0000 218.4000 228.8000 219.8000 ;
	    RECT 226.8000 217.8000 228.8000 218.4000 ;
	    RECT 232.4000 217.8000 233.2000 219.8000 ;
	    RECT 236.6000 218.4000 237.8000 219.8000 ;
	    RECT 236.4000 217.8000 237.8000 218.4000 ;
	    RECT 226.8000 217.0000 227.6000 217.8000 ;
	    RECT 232.4000 217.2000 233.0000 217.8000 ;
	    RECT 228.4000 215.6000 229.2000 217.2000 ;
	    RECT 230.2000 216.6000 233.0000 217.2000 ;
	    RECT 236.4000 217.0000 237.2000 217.8000 ;
	    RECT 230.2000 216.4000 231.0000 216.6000 ;
	    RECT 221.2000 214.4000 222.0000 214.8000 ;
	    RECT 217.2000 213.6000 219.8000 214.4000 ;
	    RECT 221.2000 213.8000 222.8000 214.4000 ;
	    RECT 222.0000 213.6000 222.8000 213.8000 ;
	    RECT 224.4000 214.2000 226.0000 214.4000 ;
	    RECT 228.6000 214.2000 229.2000 215.6000 ;
	    RECT 238.2000 215.4000 239.0000 215.6000 ;
	    RECT 241.2000 215.4000 242.0000 219.8000 ;
	    RECT 246.6000 216.0000 247.4000 219.0000 ;
	    RECT 250.8000 217.0000 251.6000 219.0000 ;
	    RECT 238.2000 214.8000 242.0000 215.4000 ;
	    RECT 234.2000 214.2000 235.0000 214.4000 ;
	    RECT 224.4000 213.6000 235.4000 214.2000 ;
	    RECT 219.2000 212.4000 219.8000 213.6000 ;
	    RECT 227.4000 213.4000 228.2000 213.6000 ;
	    RECT 214.0000 211.7000 217.9000 212.3000 ;
	    RECT 201.2000 209.6000 202.6000 210.2000 ;
	    RECT 203.2000 209.6000 204.2000 210.2000 ;
	    RECT 202.0000 208.4000 202.6000 209.6000 ;
	    RECT 202.0000 207.6000 202.8000 208.4000 ;
	    RECT 203.4000 202.2000 204.2000 209.6000 ;
	    RECT 209.2000 209.4000 211.0000 210.2000 ;
	    RECT 210.2000 202.2000 211.0000 209.4000 ;
	    RECT 214.0000 202.2000 214.8000 211.7000 ;
	    RECT 217.3000 210.4000 217.9000 211.7000 ;
	    RECT 218.8000 211.6000 219.8000 212.4000 ;
	    RECT 220.4000 211.6000 221.2000 213.2000 ;
	    RECT 225.8000 212.4000 226.6000 212.6000 ;
	    RECT 228.4000 212.4000 229.2000 212.6000 ;
	    RECT 225.8000 211.8000 230.8000 212.4000 ;
	    RECT 230.0000 211.6000 230.8000 211.8000 ;
	    RECT 215.6000 208.8000 216.4000 210.4000 ;
	    RECT 217.2000 210.2000 218.0000 210.4000 ;
	    RECT 219.2000 210.2000 219.8000 211.6000 ;
	    RECT 223.6000 211.0000 229.2000 211.2000 ;
	    RECT 223.6000 210.8000 229.4000 211.0000 ;
	    RECT 223.6000 210.6000 233.4000 210.8000 ;
	    RECT 217.2000 209.6000 218.6000 210.2000 ;
	    RECT 219.2000 209.6000 220.2000 210.2000 ;
	    RECT 218.0000 208.4000 218.6000 209.6000 ;
	    RECT 218.0000 207.6000 218.8000 208.4000 ;
	    RECT 219.4000 202.2000 220.2000 209.6000 ;
	    RECT 223.6000 202.2000 224.4000 210.6000 ;
	    RECT 228.6000 210.2000 233.4000 210.6000 ;
	    RECT 226.8000 209.0000 232.2000 209.6000 ;
	    RECT 226.8000 208.8000 227.6000 209.0000 ;
	    RECT 231.4000 208.8000 232.2000 209.0000 ;
	    RECT 232.8000 209.0000 233.4000 210.2000 ;
	    RECT 234.8000 210.4000 235.4000 213.6000 ;
	    RECT 236.4000 212.8000 237.2000 213.0000 ;
	    RECT 236.4000 212.2000 240.2000 212.8000 ;
	    RECT 239.4000 212.0000 240.2000 212.2000 ;
	    RECT 237.8000 211.4000 238.6000 211.6000 ;
	    RECT 241.2000 211.4000 242.0000 214.8000 ;
	    RECT 245.8000 215.4000 247.4000 216.0000 ;
	    RECT 245.8000 215.0000 246.6000 215.4000 ;
	    RECT 245.8000 214.4000 246.4000 215.0000 ;
	    RECT 251.0000 214.8000 251.6000 217.0000 ;
	    RECT 262.6000 216.0000 263.4000 219.0000 ;
	    RECT 266.8000 217.0000 267.6000 219.0000 ;
	    RECT 244.4000 213.6000 246.4000 214.4000 ;
	    RECT 247.4000 214.2000 251.6000 214.8000 ;
	    RECT 261.8000 215.4000 263.4000 216.0000 ;
	    RECT 261.8000 215.0000 262.6000 215.4000 ;
	    RECT 261.8000 214.4000 262.4000 215.0000 ;
	    RECT 267.0000 214.8000 267.6000 217.0000 ;
	    RECT 247.4000 213.8000 248.4000 214.2000 ;
	    RECT 237.8000 210.8000 242.0000 211.4000 ;
	    RECT 244.4000 210.8000 245.2000 212.4000 ;
	    RECT 234.8000 209.8000 237.2000 210.4000 ;
	    RECT 234.2000 209.0000 235.0000 209.2000 ;
	    RECT 232.8000 208.4000 235.0000 209.0000 ;
	    RECT 236.6000 208.8000 237.2000 209.8000 ;
	    RECT 236.6000 208.0000 238.0000 208.8000 ;
	    RECT 230.2000 207.4000 231.0000 207.6000 ;
	    RECT 233.0000 207.4000 233.8000 207.6000 ;
	    RECT 226.8000 206.2000 227.6000 207.0000 ;
	    RECT 230.2000 206.8000 233.8000 207.4000 ;
	    RECT 232.4000 206.2000 233.0000 206.8000 ;
	    RECT 236.4000 206.2000 237.2000 207.0000 ;
	    RECT 226.8000 205.6000 228.8000 206.2000 ;
	    RECT 228.0000 202.2000 228.8000 205.6000 ;
	    RECT 232.4000 202.2000 233.2000 206.2000 ;
	    RECT 236.6000 202.2000 237.8000 206.2000 ;
	    RECT 241.2000 202.2000 242.0000 210.8000 ;
	    RECT 245.8000 209.8000 246.4000 213.6000 ;
	    RECT 247.0000 213.0000 248.4000 213.8000 ;
	    RECT 260.4000 213.6000 262.4000 214.4000 ;
	    RECT 263.4000 214.2000 267.6000 214.8000 ;
	    RECT 263.4000 213.8000 264.4000 214.2000 ;
	    RECT 247.8000 211.0000 248.4000 213.0000 ;
	    RECT 249.2000 211.6000 250.0000 213.2000 ;
	    RECT 250.8000 212.3000 251.6000 213.2000 ;
	    RECT 258.8000 212.3000 259.6000 212.4000 ;
	    RECT 250.8000 211.7000 259.6000 212.3000 ;
	    RECT 250.8000 211.6000 251.6000 211.7000 ;
	    RECT 258.8000 211.6000 259.6000 211.7000 ;
	    RECT 247.8000 210.4000 251.6000 211.0000 ;
	    RECT 260.4000 210.8000 261.2000 212.4000 ;
	    RECT 245.8000 209.2000 247.4000 209.8000 ;
	    RECT 246.6000 204.4000 247.4000 209.2000 ;
	    RECT 251.0000 207.0000 251.6000 210.4000 ;
	    RECT 252.4000 210.3000 253.2000 210.4000 ;
	    RECT 257.2000 210.3000 258.0000 210.4000 ;
	    RECT 252.4000 209.7000 258.0000 210.3000 ;
	    RECT 252.4000 209.6000 253.2000 209.7000 ;
	    RECT 257.2000 209.6000 258.0000 209.7000 ;
	    RECT 261.8000 209.8000 262.4000 213.6000 ;
	    RECT 263.0000 213.0000 264.4000 213.8000 ;
	    RECT 263.8000 211.0000 264.4000 213.0000 ;
	    RECT 265.2000 211.6000 266.0000 213.2000 ;
	    RECT 266.8000 211.6000 267.6000 213.2000 ;
	    RECT 268.4000 212.4000 269.2000 219.8000 ;
	    RECT 271.6000 215.2000 272.4000 219.8000 ;
	    RECT 270.2000 214.6000 272.4000 215.2000 ;
	    RECT 263.8000 210.4000 267.6000 211.0000 ;
	    RECT 261.8000 209.2000 263.4000 209.8000 ;
	    RECT 246.0000 203.6000 247.4000 204.4000 ;
	    RECT 246.6000 202.2000 247.4000 203.6000 ;
	    RECT 250.8000 203.0000 251.6000 207.0000 ;
	    RECT 262.6000 204.4000 263.4000 209.2000 ;
	    RECT 267.0000 207.0000 267.6000 210.4000 ;
	    RECT 262.6000 203.6000 264.4000 204.4000 ;
	    RECT 262.6000 202.2000 263.4000 203.6000 ;
	    RECT 266.8000 203.0000 267.6000 207.0000 ;
	    RECT 268.4000 210.2000 269.0000 212.4000 ;
	    RECT 270.2000 211.6000 270.8000 214.6000 ;
	    RECT 271.6000 211.6000 272.4000 213.2000 ;
	    RECT 273.2000 212.4000 274.0000 219.8000 ;
	    RECT 276.4000 215.2000 277.2000 219.8000 ;
	    RECT 280.6000 216.4000 281.4000 219.8000 ;
	    RECT 279.6000 215.8000 281.4000 216.4000 ;
	    RECT 282.8000 215.8000 283.6000 219.8000 ;
	    RECT 284.4000 216.0000 285.2000 219.8000 ;
	    RECT 287.6000 216.0000 288.4000 219.8000 ;
	    RECT 284.4000 215.8000 288.4000 216.0000 ;
	    RECT 275.0000 214.6000 277.2000 215.2000 ;
	    RECT 269.6000 210.8000 270.8000 211.6000 ;
	    RECT 270.2000 210.2000 270.8000 210.8000 ;
	    RECT 273.2000 210.2000 273.8000 212.4000 ;
	    RECT 275.0000 211.6000 275.6000 214.6000 ;
	    RECT 278.0000 213.6000 278.8000 215.2000 ;
	    RECT 274.4000 210.8000 275.6000 211.6000 ;
	    RECT 275.0000 210.2000 275.6000 210.8000 ;
	    RECT 279.6000 212.3000 280.4000 215.8000 ;
	    RECT 283.0000 214.4000 283.6000 215.8000 ;
	    RECT 284.6000 215.4000 288.2000 215.8000 ;
	    RECT 289.2000 215.4000 290.0000 219.8000 ;
	    RECT 293.4000 218.4000 294.6000 219.8000 ;
	    RECT 293.4000 217.8000 294.8000 218.4000 ;
	    RECT 298.0000 217.8000 298.8000 219.8000 ;
	    RECT 302.4000 218.4000 303.2000 219.8000 ;
	    RECT 302.4000 217.8000 304.4000 218.4000 ;
	    RECT 294.0000 217.0000 294.8000 217.8000 ;
	    RECT 298.2000 217.2000 298.8000 217.8000 ;
	    RECT 298.2000 216.6000 301.0000 217.2000 ;
	    RECT 300.2000 216.4000 301.0000 216.6000 ;
	    RECT 302.0000 216.4000 302.8000 217.2000 ;
	    RECT 303.6000 217.0000 304.4000 217.8000 ;
	    RECT 292.2000 215.4000 293.0000 215.6000 ;
	    RECT 289.2000 214.8000 293.0000 215.4000 ;
	    RECT 286.8000 214.4000 287.6000 214.8000 ;
	    RECT 282.8000 213.6000 285.4000 214.4000 ;
	    RECT 286.8000 213.8000 288.4000 214.4000 ;
	    RECT 287.6000 213.6000 288.4000 213.8000 ;
	    RECT 279.6000 211.7000 283.5000 212.3000 ;
	    RECT 268.4000 202.2000 269.2000 210.2000 ;
	    RECT 270.2000 209.6000 272.4000 210.2000 ;
	    RECT 271.6000 202.2000 272.4000 209.6000 ;
	    RECT 273.2000 202.2000 274.0000 210.2000 ;
	    RECT 275.0000 209.6000 277.2000 210.2000 ;
	    RECT 276.4000 202.2000 277.2000 209.6000 ;
	    RECT 279.6000 202.2000 280.4000 211.7000 ;
	    RECT 282.9000 210.4000 283.5000 211.7000 ;
	    RECT 284.8000 210.4000 285.4000 213.6000 ;
	    RECT 286.0000 212.3000 286.8000 213.2000 ;
	    RECT 287.6000 212.3000 288.4000 212.4000 ;
	    RECT 286.0000 211.7000 288.4000 212.3000 ;
	    RECT 286.0000 211.6000 286.8000 211.7000 ;
	    RECT 287.6000 211.6000 288.4000 211.7000 ;
	    RECT 289.2000 211.4000 290.0000 214.8000 ;
	    RECT 296.2000 214.2000 297.0000 214.4000 ;
	    RECT 302.0000 214.2000 302.6000 216.4000 ;
	    RECT 306.8000 215.0000 307.6000 219.8000 ;
	    RECT 308.4000 217.0000 309.2000 219.0000 ;
	    RECT 308.4000 214.8000 309.0000 217.0000 ;
	    RECT 312.6000 216.0000 313.4000 219.0000 ;
	    RECT 318.0000 217.0000 318.8000 219.0000 ;
	    RECT 312.6000 215.4000 314.2000 216.0000 ;
	    RECT 313.4000 215.0000 314.2000 215.4000 ;
	    RECT 305.2000 214.2000 306.8000 214.4000 ;
	    RECT 308.4000 214.2000 312.6000 214.8000 ;
	    RECT 295.8000 213.6000 306.8000 214.2000 ;
	    RECT 311.6000 213.8000 312.6000 214.2000 ;
	    RECT 313.6000 214.4000 314.2000 215.0000 ;
	    RECT 318.0000 214.8000 318.6000 217.0000 ;
	    RECT 322.2000 216.0000 323.0000 219.0000 ;
	    RECT 322.2000 215.4000 323.8000 216.0000 ;
	    RECT 323.0000 215.0000 323.8000 215.4000 ;
	    RECT 294.0000 212.8000 294.8000 213.0000 ;
	    RECT 291.0000 212.2000 294.8000 212.8000 ;
	    RECT 291.0000 212.0000 291.8000 212.2000 ;
	    RECT 292.6000 211.4000 293.4000 211.6000 ;
	    RECT 289.2000 210.8000 293.4000 211.4000 ;
	    RECT 281.2000 208.8000 282.0000 210.4000 ;
	    RECT 282.8000 210.2000 283.6000 210.4000 ;
	    RECT 282.8000 209.6000 284.2000 210.2000 ;
	    RECT 284.8000 209.6000 286.8000 210.4000 ;
	    RECT 283.6000 208.4000 284.2000 209.6000 ;
	    RECT 283.6000 207.6000 284.4000 208.4000 ;
	    RECT 285.0000 202.2000 285.8000 209.6000 ;
	    RECT 289.2000 202.2000 290.0000 210.8000 ;
	    RECT 295.8000 210.4000 296.4000 213.6000 ;
	    RECT 303.0000 213.4000 303.8000 213.6000 ;
	    RECT 304.6000 212.4000 305.4000 212.6000 ;
	    RECT 300.4000 211.8000 305.4000 212.4000 ;
	    RECT 300.4000 211.6000 301.2000 211.8000 ;
	    RECT 308.4000 211.6000 309.2000 213.2000 ;
	    RECT 310.0000 211.6000 310.8000 213.2000 ;
	    RECT 311.6000 213.0000 313.0000 213.8000 ;
	    RECT 313.6000 213.6000 315.6000 214.4000 ;
	    RECT 318.0000 214.2000 322.2000 214.8000 ;
	    RECT 321.2000 213.8000 322.2000 214.2000 ;
	    RECT 323.2000 214.4000 323.8000 215.0000 ;
	    RECT 327.6000 215.4000 328.4000 219.8000 ;
	    RECT 331.8000 218.4000 333.0000 219.8000 ;
	    RECT 331.8000 217.8000 333.2000 218.4000 ;
	    RECT 336.4000 217.8000 337.2000 219.8000 ;
	    RECT 340.8000 218.4000 341.6000 219.8000 ;
	    RECT 340.8000 217.8000 342.8000 218.4000 ;
	    RECT 332.4000 217.0000 333.2000 217.8000 ;
	    RECT 336.6000 217.2000 337.2000 217.8000 ;
	    RECT 336.6000 216.6000 339.4000 217.2000 ;
	    RECT 338.6000 216.4000 339.4000 216.6000 ;
	    RECT 340.4000 216.4000 341.2000 217.2000 ;
	    RECT 342.0000 217.0000 342.8000 217.8000 ;
	    RECT 330.6000 215.4000 331.4000 215.6000 ;
	    RECT 327.6000 214.8000 331.4000 215.4000 ;
	    RECT 302.0000 211.0000 307.6000 211.2000 ;
	    RECT 311.6000 211.0000 312.2000 213.0000 ;
	    RECT 301.8000 210.8000 307.6000 211.0000 ;
	    RECT 294.0000 209.8000 296.4000 210.4000 ;
	    RECT 297.8000 210.6000 307.6000 210.8000 ;
	    RECT 297.8000 210.2000 302.6000 210.6000 ;
	    RECT 294.0000 208.8000 294.6000 209.8000 ;
	    RECT 293.2000 208.0000 294.6000 208.8000 ;
	    RECT 296.2000 209.0000 297.0000 209.2000 ;
	    RECT 297.8000 209.0000 298.4000 210.2000 ;
	    RECT 296.2000 208.4000 298.4000 209.0000 ;
	    RECT 299.0000 209.0000 304.4000 209.6000 ;
	    RECT 299.0000 208.8000 299.8000 209.0000 ;
	    RECT 303.6000 208.8000 304.4000 209.0000 ;
	    RECT 297.4000 207.4000 298.2000 207.6000 ;
	    RECT 300.2000 207.4000 301.0000 207.6000 ;
	    RECT 294.0000 206.2000 294.8000 207.0000 ;
	    RECT 297.4000 206.8000 301.0000 207.4000 ;
	    RECT 298.2000 206.2000 298.8000 206.8000 ;
	    RECT 303.6000 206.2000 304.4000 207.0000 ;
	    RECT 293.4000 202.2000 294.6000 206.2000 ;
	    RECT 298.0000 202.2000 298.8000 206.2000 ;
	    RECT 302.4000 205.6000 304.4000 206.2000 ;
	    RECT 302.4000 202.2000 303.2000 205.6000 ;
	    RECT 306.8000 202.2000 307.6000 210.6000 ;
	    RECT 308.4000 210.4000 312.2000 211.0000 ;
	    RECT 308.4000 207.0000 309.0000 210.4000 ;
	    RECT 313.6000 209.8000 314.2000 213.6000 ;
	    RECT 314.8000 212.3000 315.6000 212.4000 ;
	    RECT 316.4000 212.3000 317.2000 212.4000 ;
	    RECT 314.8000 211.7000 317.2000 212.3000 ;
	    RECT 314.8000 210.8000 315.6000 211.7000 ;
	    RECT 316.4000 211.6000 317.2000 211.7000 ;
	    RECT 318.0000 211.6000 318.8000 213.2000 ;
	    RECT 319.6000 211.6000 320.4000 213.2000 ;
	    RECT 321.2000 213.0000 322.6000 213.8000 ;
	    RECT 323.2000 213.6000 325.2000 214.4000 ;
	    RECT 321.2000 211.0000 321.8000 213.0000 ;
	    RECT 312.6000 209.2000 314.2000 209.8000 ;
	    RECT 318.0000 210.4000 321.8000 211.0000 ;
	    RECT 308.4000 203.0000 309.2000 207.0000 ;
	    RECT 312.6000 206.4000 313.4000 209.2000 ;
	    RECT 311.6000 205.6000 313.4000 206.4000 ;
	    RECT 312.6000 202.2000 313.4000 205.6000 ;
	    RECT 318.0000 207.0000 318.6000 210.4000 ;
	    RECT 323.2000 209.8000 323.8000 213.6000 ;
	    RECT 324.4000 210.8000 325.2000 212.4000 ;
	    RECT 327.6000 211.4000 328.4000 214.8000 ;
	    RECT 334.6000 214.2000 335.4000 214.4000 ;
	    RECT 338.8000 214.2000 339.6000 214.4000 ;
	    RECT 340.4000 214.2000 341.0000 216.4000 ;
	    RECT 345.2000 215.0000 346.0000 219.8000 ;
	    RECT 346.8000 216.0000 347.6000 219.8000 ;
	    RECT 350.0000 216.0000 350.8000 219.8000 ;
	    RECT 346.8000 215.8000 350.8000 216.0000 ;
	    RECT 351.6000 215.8000 352.4000 219.8000 ;
	    RECT 353.2000 215.8000 354.0000 219.8000 ;
	    RECT 354.8000 216.0000 355.6000 219.8000 ;
	    RECT 358.0000 216.0000 358.8000 219.8000 ;
	    RECT 354.8000 215.8000 358.8000 216.0000 ;
	    RECT 347.0000 215.4000 350.6000 215.8000 ;
	    RECT 347.6000 214.4000 348.4000 214.8000 ;
	    RECT 351.6000 214.4000 352.2000 215.8000 ;
	    RECT 353.4000 214.4000 354.0000 215.8000 ;
	    RECT 355.0000 215.4000 358.6000 215.8000 ;
	    RECT 357.2000 214.4000 358.0000 214.8000 ;
	    RECT 343.6000 214.2000 345.2000 214.4000 ;
	    RECT 334.2000 213.6000 345.2000 214.2000 ;
	    RECT 346.8000 213.8000 348.4000 214.4000 ;
	    RECT 346.8000 213.6000 347.6000 213.8000 ;
	    RECT 349.8000 213.6000 352.4000 214.4000 ;
	    RECT 353.2000 213.6000 355.8000 214.4000 ;
	    RECT 357.2000 213.8000 358.8000 214.4000 ;
	    RECT 358.0000 213.6000 358.8000 213.8000 ;
	    RECT 332.4000 212.8000 333.2000 213.0000 ;
	    RECT 329.4000 212.2000 333.2000 212.8000 ;
	    RECT 329.4000 212.0000 330.2000 212.2000 ;
	    RECT 331.0000 211.4000 331.8000 211.6000 ;
	    RECT 327.6000 210.8000 331.8000 211.4000 ;
	    RECT 322.2000 209.2000 323.8000 209.8000 ;
	    RECT 322.2000 208.4000 323.0000 209.2000 ;
	    RECT 321.2000 207.6000 323.0000 208.4000 ;
	    RECT 318.0000 203.0000 318.8000 207.0000 ;
	    RECT 322.2000 202.2000 323.0000 207.6000 ;
	    RECT 327.6000 202.2000 328.4000 210.8000 ;
	    RECT 334.2000 210.4000 334.8000 213.6000 ;
	    RECT 341.4000 213.4000 342.2000 213.6000 ;
	    RECT 340.4000 212.4000 341.2000 212.6000 ;
	    RECT 343.0000 212.4000 343.8000 212.6000 ;
	    RECT 338.8000 211.8000 343.8000 212.4000 ;
	    RECT 338.8000 211.6000 339.6000 211.8000 ;
	    RECT 348.4000 211.6000 349.2000 213.2000 ;
	    RECT 340.4000 211.0000 346.0000 211.2000 ;
	    RECT 340.2000 210.8000 346.0000 211.0000 ;
	    RECT 332.4000 209.8000 334.8000 210.4000 ;
	    RECT 336.2000 210.6000 346.0000 210.8000 ;
	    RECT 336.2000 210.2000 341.0000 210.6000 ;
	    RECT 332.4000 208.8000 333.0000 209.8000 ;
	    RECT 331.6000 208.0000 333.0000 208.8000 ;
	    RECT 334.6000 209.0000 335.4000 209.2000 ;
	    RECT 336.2000 209.0000 336.8000 210.2000 ;
	    RECT 334.6000 208.4000 336.8000 209.0000 ;
	    RECT 337.4000 209.0000 342.8000 209.6000 ;
	    RECT 337.4000 208.8000 338.2000 209.0000 ;
	    RECT 342.0000 208.8000 342.8000 209.0000 ;
	    RECT 335.8000 207.4000 336.6000 207.6000 ;
	    RECT 338.6000 207.4000 339.4000 207.6000 ;
	    RECT 332.4000 206.2000 333.2000 207.0000 ;
	    RECT 335.8000 206.8000 339.4000 207.4000 ;
	    RECT 336.6000 206.2000 337.2000 206.8000 ;
	    RECT 342.0000 206.2000 342.8000 207.0000 ;
	    RECT 331.8000 202.2000 333.0000 206.2000 ;
	    RECT 336.4000 202.2000 337.2000 206.2000 ;
	    RECT 340.8000 205.6000 342.8000 206.2000 ;
	    RECT 340.8000 202.2000 341.6000 205.6000 ;
	    RECT 345.2000 202.2000 346.0000 210.6000 ;
	    RECT 349.8000 210.4000 350.4000 213.6000 ;
	    RECT 355.2000 212.3000 355.8000 213.6000 ;
	    RECT 351.7000 211.7000 355.8000 212.3000 ;
	    RECT 351.7000 210.4000 352.3000 211.7000 ;
	    RECT 348.4000 209.6000 350.4000 210.4000 ;
	    RECT 351.6000 210.2000 352.4000 210.4000 ;
	    RECT 351.0000 209.6000 352.4000 210.2000 ;
	    RECT 353.2000 210.2000 354.0000 210.4000 ;
	    RECT 355.2000 210.2000 355.8000 211.7000 ;
	    RECT 356.4000 211.6000 357.2000 213.2000 ;
	    RECT 359.6000 212.4000 360.4000 219.8000 ;
	    RECT 362.8000 215.2000 363.6000 219.8000 ;
	    RECT 361.4000 214.6000 363.6000 215.2000 ;
	    RECT 364.4000 215.4000 365.2000 219.8000 ;
	    RECT 368.6000 218.4000 369.8000 219.8000 ;
	    RECT 368.6000 217.8000 370.0000 218.4000 ;
	    RECT 373.2000 217.8000 374.0000 219.8000 ;
	    RECT 377.6000 218.4000 378.4000 219.8000 ;
	    RECT 377.6000 217.8000 379.6000 218.4000 ;
	    RECT 369.2000 217.0000 370.0000 217.8000 ;
	    RECT 373.4000 217.2000 374.0000 217.8000 ;
	    RECT 373.4000 216.6000 376.2000 217.2000 ;
	    RECT 375.4000 216.4000 376.2000 216.6000 ;
	    RECT 377.2000 216.4000 378.0000 217.2000 ;
	    RECT 378.8000 217.0000 379.6000 217.8000 ;
	    RECT 367.4000 215.4000 368.2000 215.6000 ;
	    RECT 364.4000 214.8000 368.2000 215.4000 ;
	    RECT 359.6000 210.2000 360.2000 212.4000 ;
	    RECT 361.4000 211.6000 362.0000 214.6000 ;
	    RECT 362.8000 211.6000 363.6000 213.2000 ;
	    RECT 360.8000 210.8000 362.0000 211.6000 ;
	    RECT 361.4000 210.2000 362.0000 210.8000 ;
	    RECT 364.4000 211.4000 365.2000 214.8000 ;
	    RECT 371.4000 214.2000 372.2000 214.4000 ;
	    RECT 377.2000 214.2000 377.8000 216.4000 ;
	    RECT 382.0000 215.0000 382.8000 219.8000 ;
	    RECT 386.2000 216.4000 387.0000 219.8000 ;
	    RECT 385.2000 215.8000 387.0000 216.4000 ;
	    RECT 388.4000 215.8000 389.2000 219.8000 ;
	    RECT 390.0000 216.0000 390.8000 219.8000 ;
	    RECT 393.2000 216.0000 394.0000 219.8000 ;
	    RECT 390.0000 215.8000 394.0000 216.0000 ;
	    RECT 380.4000 214.2000 382.0000 214.4000 ;
	    RECT 371.0000 213.6000 382.0000 214.2000 ;
	    RECT 383.6000 213.6000 384.4000 215.2000 ;
	    RECT 369.2000 212.8000 370.0000 213.0000 ;
	    RECT 366.2000 212.2000 370.0000 212.8000 ;
	    RECT 371.0000 212.4000 371.6000 213.6000 ;
	    RECT 378.2000 213.4000 379.0000 213.6000 ;
	    RECT 377.2000 212.4000 378.0000 212.6000 ;
	    RECT 379.8000 212.4000 380.6000 212.6000 ;
	    RECT 366.2000 212.0000 367.0000 212.2000 ;
	    RECT 370.8000 211.6000 371.6000 212.4000 ;
	    RECT 375.6000 211.8000 380.6000 212.4000 ;
	    RECT 385.2000 212.3000 386.0000 215.8000 ;
	    RECT 388.6000 214.4000 389.2000 215.8000 ;
	    RECT 390.2000 215.4000 393.8000 215.8000 ;
	    RECT 394.8000 215.2000 395.6000 219.8000 ;
	    RECT 392.4000 214.4000 393.2000 214.8000 ;
	    RECT 394.8000 214.6000 397.0000 215.2000 ;
	    RECT 388.4000 213.6000 391.0000 214.4000 ;
	    RECT 392.4000 213.8000 394.0000 214.4000 ;
	    RECT 393.2000 213.6000 394.0000 213.8000 ;
	    RECT 375.6000 211.6000 376.4000 211.8000 ;
	    RECT 385.2000 211.7000 389.1000 212.3000 ;
	    RECT 367.8000 211.4000 368.6000 211.6000 ;
	    RECT 364.4000 210.8000 368.6000 211.4000 ;
	    RECT 353.2000 209.6000 354.6000 210.2000 ;
	    RECT 355.2000 209.6000 356.2000 210.2000 ;
	    RECT 349.4000 202.2000 350.2000 209.6000 ;
	    RECT 351.0000 208.4000 351.6000 209.6000 ;
	    RECT 354.0000 208.4000 354.6000 209.6000 ;
	    RECT 350.8000 207.6000 351.6000 208.4000 ;
	    RECT 353.2000 207.6000 354.8000 208.4000 ;
	    RECT 355.4000 202.2000 356.2000 209.6000 ;
	    RECT 359.6000 202.2000 360.4000 210.2000 ;
	    RECT 361.4000 209.6000 363.6000 210.2000 ;
	    RECT 362.8000 202.2000 363.6000 209.6000 ;
	    RECT 364.4000 202.2000 365.2000 210.8000 ;
	    RECT 371.0000 210.4000 371.6000 211.6000 ;
	    RECT 377.2000 211.0000 382.8000 211.2000 ;
	    RECT 377.0000 210.8000 382.8000 211.0000 ;
	    RECT 369.2000 209.8000 371.6000 210.4000 ;
	    RECT 373.0000 210.6000 382.8000 210.8000 ;
	    RECT 373.0000 210.2000 377.8000 210.6000 ;
	    RECT 369.2000 208.8000 369.8000 209.8000 ;
	    RECT 368.4000 208.0000 369.8000 208.8000 ;
	    RECT 371.4000 209.0000 372.2000 209.2000 ;
	    RECT 373.0000 209.0000 373.6000 210.2000 ;
	    RECT 371.4000 208.4000 373.6000 209.0000 ;
	    RECT 374.2000 209.0000 379.6000 209.6000 ;
	    RECT 374.2000 208.8000 375.0000 209.0000 ;
	    RECT 378.8000 208.8000 379.6000 209.0000 ;
	    RECT 372.6000 207.4000 373.4000 207.6000 ;
	    RECT 375.4000 207.4000 376.2000 207.6000 ;
	    RECT 369.2000 206.2000 370.0000 207.0000 ;
	    RECT 372.6000 206.8000 376.2000 207.4000 ;
	    RECT 373.4000 206.2000 374.0000 206.8000 ;
	    RECT 378.8000 206.2000 379.6000 207.0000 ;
	    RECT 368.6000 202.2000 369.8000 206.2000 ;
	    RECT 373.2000 202.2000 374.0000 206.2000 ;
	    RECT 377.6000 205.6000 379.6000 206.2000 ;
	    RECT 377.6000 202.2000 378.4000 205.6000 ;
	    RECT 382.0000 202.2000 382.8000 210.6000 ;
	    RECT 385.2000 202.2000 386.0000 211.7000 ;
	    RECT 388.5000 210.4000 389.1000 211.7000 ;
	    RECT 386.8000 208.8000 387.6000 210.4000 ;
	    RECT 388.4000 210.2000 389.2000 210.4000 ;
	    RECT 390.4000 210.2000 391.0000 213.6000 ;
	    RECT 391.6000 211.6000 392.4000 213.2000 ;
	    RECT 394.8000 211.6000 395.6000 213.2000 ;
	    RECT 396.4000 211.6000 397.0000 214.6000 ;
	    RECT 398.0000 212.4000 398.8000 219.8000 ;
	    RECT 402.2000 216.4000 403.0000 219.8000 ;
	    RECT 401.2000 215.8000 403.0000 216.4000 ;
	    RECT 410.8000 215.8000 411.6000 219.8000 ;
	    RECT 412.4000 216.0000 413.2000 219.8000 ;
	    RECT 415.6000 216.0000 416.4000 219.8000 ;
	    RECT 412.4000 215.8000 416.4000 216.0000 ;
	    RECT 399.6000 213.6000 400.4000 215.2000 ;
	    RECT 396.4000 210.8000 397.6000 211.6000 ;
	    RECT 396.4000 210.2000 397.0000 210.8000 ;
	    RECT 398.2000 210.2000 398.8000 212.4000 ;
	    RECT 388.4000 209.6000 389.8000 210.2000 ;
	    RECT 390.4000 209.6000 391.4000 210.2000 ;
	    RECT 389.2000 208.4000 389.8000 209.6000 ;
	    RECT 389.2000 207.6000 390.0000 208.4000 ;
	    RECT 390.6000 202.2000 391.4000 209.6000 ;
	    RECT 394.8000 209.6000 397.0000 210.2000 ;
	    RECT 394.8000 202.2000 395.6000 209.6000 ;
	    RECT 398.0000 202.2000 398.8000 210.2000 ;
	    RECT 401.2000 212.3000 402.0000 215.8000 ;
	    RECT 411.0000 214.4000 411.6000 215.8000 ;
	    RECT 412.6000 215.4000 416.2000 215.8000 ;
	    RECT 417.2000 215.4000 418.0000 219.8000 ;
	    RECT 421.4000 218.4000 422.6000 219.8000 ;
	    RECT 421.4000 217.8000 422.8000 218.4000 ;
	    RECT 426.0000 217.8000 426.8000 219.8000 ;
	    RECT 430.4000 218.4000 431.2000 219.8000 ;
	    RECT 430.4000 217.8000 432.4000 218.4000 ;
	    RECT 422.0000 217.0000 422.8000 217.8000 ;
	    RECT 426.2000 217.2000 426.8000 217.8000 ;
	    RECT 426.2000 216.6000 429.0000 217.2000 ;
	    RECT 428.2000 216.4000 429.0000 216.6000 ;
	    RECT 430.0000 216.4000 430.8000 217.2000 ;
	    RECT 431.6000 217.0000 432.4000 217.8000 ;
	    RECT 420.2000 215.4000 421.0000 215.6000 ;
	    RECT 417.2000 214.8000 421.0000 215.4000 ;
	    RECT 414.8000 214.4000 415.6000 214.8000 ;
	    RECT 410.8000 213.6000 413.4000 214.4000 ;
	    RECT 414.8000 213.8000 416.4000 214.4000 ;
	    RECT 415.6000 213.6000 416.4000 213.8000 ;
	    RECT 401.2000 211.7000 411.5000 212.3000 ;
	    RECT 401.2000 202.2000 402.0000 211.7000 ;
	    RECT 410.9000 210.4000 411.5000 211.7000 ;
	    RECT 412.8000 210.4000 413.4000 213.6000 ;
	    RECT 414.0000 212.3000 414.8000 213.2000 ;
	    RECT 415.6000 212.3000 416.4000 212.4000 ;
	    RECT 414.0000 211.7000 416.4000 212.3000 ;
	    RECT 414.0000 211.6000 414.8000 211.7000 ;
	    RECT 415.6000 211.6000 416.4000 211.7000 ;
	    RECT 417.2000 211.4000 418.0000 214.8000 ;
	    RECT 424.2000 214.2000 425.0000 214.4000 ;
	    RECT 430.0000 214.2000 430.6000 216.4000 ;
	    RECT 434.8000 215.0000 435.6000 219.8000 ;
	    RECT 433.2000 214.2000 434.8000 214.4000 ;
	    RECT 423.8000 213.6000 434.8000 214.2000 ;
	    RECT 422.0000 212.8000 422.8000 213.0000 ;
	    RECT 419.0000 212.2000 422.8000 212.8000 ;
	    RECT 419.0000 212.0000 419.8000 212.2000 ;
	    RECT 420.6000 211.4000 421.4000 211.6000 ;
	    RECT 417.2000 210.8000 421.4000 211.4000 ;
	    RECT 402.8000 208.8000 403.6000 210.4000 ;
	    RECT 410.8000 210.2000 411.6000 210.4000 ;
	    RECT 410.8000 209.6000 412.2000 210.2000 ;
	    RECT 412.8000 209.6000 414.8000 210.4000 ;
	    RECT 411.6000 208.4000 412.2000 209.6000 ;
	    RECT 411.6000 207.6000 412.4000 208.4000 ;
	    RECT 413.0000 202.2000 413.8000 209.6000 ;
	    RECT 417.2000 202.2000 418.0000 210.8000 ;
	    RECT 423.8000 210.4000 424.4000 213.6000 ;
	    RECT 431.0000 213.4000 431.8000 213.6000 ;
	    RECT 432.6000 212.4000 433.4000 212.6000 ;
	    RECT 428.4000 211.8000 433.4000 212.4000 ;
	    RECT 428.4000 211.6000 429.2000 211.8000 ;
	    RECT 430.0000 211.0000 435.6000 211.2000 ;
	    RECT 429.8000 210.8000 435.6000 211.0000 ;
	    RECT 422.0000 209.8000 424.4000 210.4000 ;
	    RECT 425.8000 210.6000 435.6000 210.8000 ;
	    RECT 425.8000 210.2000 430.6000 210.6000 ;
	    RECT 422.0000 208.8000 422.6000 209.8000 ;
	    RECT 421.2000 208.0000 422.6000 208.8000 ;
	    RECT 424.2000 209.0000 425.0000 209.2000 ;
	    RECT 425.8000 209.0000 426.4000 210.2000 ;
	    RECT 424.2000 208.4000 426.4000 209.0000 ;
	    RECT 427.0000 209.0000 432.4000 209.6000 ;
	    RECT 427.0000 208.8000 427.8000 209.0000 ;
	    RECT 431.6000 208.8000 432.4000 209.0000 ;
	    RECT 425.4000 207.4000 426.2000 207.6000 ;
	    RECT 428.2000 207.4000 429.0000 207.6000 ;
	    RECT 422.0000 206.2000 422.8000 207.0000 ;
	    RECT 425.4000 206.8000 429.0000 207.4000 ;
	    RECT 426.2000 206.2000 426.8000 206.8000 ;
	    RECT 431.6000 206.2000 432.4000 207.0000 ;
	    RECT 421.4000 202.2000 422.6000 206.2000 ;
	    RECT 426.0000 202.2000 426.8000 206.2000 ;
	    RECT 430.4000 205.6000 432.4000 206.2000 ;
	    RECT 430.4000 202.2000 431.2000 205.6000 ;
	    RECT 434.8000 202.2000 435.6000 210.6000 ;
	    RECT 436.4000 202.2000 437.2000 219.8000 ;
	    RECT 440.2000 218.4000 441.0000 219.8000 ;
	    RECT 439.6000 217.6000 441.0000 218.4000 ;
	    RECT 440.2000 216.4000 441.0000 217.6000 ;
	    RECT 440.2000 215.8000 442.0000 216.4000 ;
	    RECT 439.6000 208.8000 440.4000 210.4000 ;
	    RECT 441.2000 202.2000 442.0000 215.8000 ;
	    RECT 442.8000 213.6000 443.6000 215.2000 ;
	    RECT 448.0000 214.2000 448.8000 219.8000 ;
	    RECT 452.4000 215.2000 453.2000 219.8000 ;
	    RECT 455.6000 215.2000 456.4000 219.8000 ;
	    RECT 448.0000 213.8000 449.8000 214.2000 ;
	    RECT 448.2000 213.6000 449.8000 213.8000 ;
	    RECT 450.8000 213.6000 451.6000 215.2000 ;
	    RECT 452.4000 214.4000 456.4000 215.2000 ;
	    RECT 446.0000 211.6000 448.4000 212.4000 ;
	    RECT 449.2000 210.4000 449.8000 213.6000 ;
	    RECT 455.6000 211.6000 456.4000 214.4000 ;
	    RECT 452.4000 210.8000 456.4000 211.6000 ;
	    RECT 449.2000 209.6000 450.0000 210.4000 ;
	    RECT 446.0000 208.3000 446.8000 208.4000 ;
	    RECT 447.6000 208.3000 448.4000 209.2000 ;
	    RECT 446.0000 207.7000 448.4000 208.3000 ;
	    RECT 446.0000 207.6000 446.8000 207.7000 ;
	    RECT 447.6000 207.6000 448.4000 207.7000 ;
	    RECT 449.2000 207.0000 449.8000 209.6000 ;
	    RECT 446.2000 206.4000 449.8000 207.0000 ;
	    RECT 446.2000 206.2000 446.8000 206.4000 ;
	    RECT 446.0000 202.2000 446.8000 206.2000 ;
	    RECT 449.2000 206.2000 449.8000 206.4000 ;
	    RECT 449.2000 202.2000 450.0000 206.2000 ;
	    RECT 452.4000 202.2000 453.2000 210.8000 ;
	    RECT 455.6000 202.2000 456.4000 210.8000 ;
	    RECT 458.8000 215.4000 459.6000 219.8000 ;
	    RECT 463.0000 218.4000 464.2000 219.8000 ;
	    RECT 463.0000 217.8000 464.4000 218.4000 ;
	    RECT 467.6000 217.8000 468.4000 219.8000 ;
	    RECT 472.0000 218.4000 472.8000 219.8000 ;
	    RECT 472.0000 217.8000 474.0000 218.4000 ;
	    RECT 463.6000 217.0000 464.4000 217.8000 ;
	    RECT 467.8000 217.2000 468.4000 217.8000 ;
	    RECT 467.8000 216.6000 470.6000 217.2000 ;
	    RECT 469.8000 216.4000 470.6000 216.6000 ;
	    RECT 471.6000 216.4000 472.4000 217.2000 ;
	    RECT 473.2000 217.0000 474.0000 217.8000 ;
	    RECT 461.8000 215.4000 462.6000 215.6000 ;
	    RECT 458.8000 214.8000 462.6000 215.4000 ;
	    RECT 458.8000 211.4000 459.6000 214.8000 ;
	    RECT 465.8000 214.2000 466.6000 214.4000 ;
	    RECT 471.6000 214.2000 472.2000 216.4000 ;
	    RECT 476.4000 215.0000 477.2000 219.8000 ;
	    RECT 478.0000 215.8000 478.8000 219.8000 ;
	    RECT 479.6000 216.0000 480.4000 219.8000 ;
	    RECT 482.8000 216.0000 483.6000 219.8000 ;
	    RECT 479.6000 215.8000 483.6000 216.0000 ;
	    RECT 478.2000 214.4000 478.8000 215.8000 ;
	    RECT 479.8000 215.4000 483.4000 215.8000 ;
	    RECT 484.4000 215.6000 485.2000 217.2000 ;
	    RECT 482.0000 214.4000 482.8000 214.8000 ;
	    RECT 474.8000 214.2000 476.4000 214.4000 ;
	    RECT 465.4000 213.6000 476.4000 214.2000 ;
	    RECT 478.0000 213.6000 480.6000 214.4000 ;
	    RECT 482.0000 214.3000 483.6000 214.4000 ;
	    RECT 486.0000 214.3000 486.8000 219.8000 ;
	    RECT 487.6000 216.0000 488.4000 219.8000 ;
	    RECT 490.8000 216.0000 491.6000 219.8000 ;
	    RECT 487.6000 215.8000 491.6000 216.0000 ;
	    RECT 492.4000 215.8000 493.2000 219.8000 ;
	    RECT 487.8000 215.4000 491.4000 215.8000 ;
	    RECT 488.4000 214.4000 489.2000 214.8000 ;
	    RECT 492.4000 214.4000 493.0000 215.8000 ;
	    RECT 494.0000 215.4000 494.8000 219.8000 ;
	    RECT 498.2000 218.4000 499.4000 219.8000 ;
	    RECT 498.2000 217.8000 499.6000 218.4000 ;
	    RECT 502.8000 217.8000 503.6000 219.8000 ;
	    RECT 507.2000 218.4000 508.0000 219.8000 ;
	    RECT 507.2000 217.8000 509.2000 218.4000 ;
	    RECT 498.8000 217.0000 499.6000 217.8000 ;
	    RECT 503.0000 217.2000 503.6000 217.8000 ;
	    RECT 503.0000 216.6000 505.8000 217.2000 ;
	    RECT 505.0000 216.4000 505.8000 216.6000 ;
	    RECT 506.8000 216.4000 507.6000 217.2000 ;
	    RECT 508.4000 217.0000 509.2000 217.8000 ;
	    RECT 497.0000 215.4000 497.8000 215.6000 ;
	    RECT 494.0000 214.8000 497.8000 215.4000 ;
	    RECT 482.0000 213.8000 486.8000 214.3000 ;
	    RECT 482.8000 213.7000 486.8000 213.8000 ;
	    RECT 482.8000 213.6000 483.6000 213.7000 ;
	    RECT 463.6000 212.8000 464.4000 213.0000 ;
	    RECT 460.6000 212.2000 464.4000 212.8000 ;
	    RECT 460.6000 212.0000 461.4000 212.2000 ;
	    RECT 462.2000 211.4000 463.0000 211.6000 ;
	    RECT 458.8000 210.8000 463.0000 211.4000 ;
	    RECT 458.8000 202.2000 459.6000 210.8000 ;
	    RECT 465.4000 210.4000 466.0000 213.6000 ;
	    RECT 472.6000 213.4000 473.4000 213.6000 ;
	    RECT 471.6000 212.4000 472.4000 212.6000 ;
	    RECT 474.2000 212.4000 475.0000 212.6000 ;
	    RECT 480.0000 212.4000 480.6000 213.6000 ;
	    RECT 470.0000 211.8000 475.0000 212.4000 ;
	    RECT 470.0000 211.6000 470.8000 211.8000 ;
	    RECT 479.6000 211.6000 480.6000 212.4000 ;
	    RECT 481.2000 211.6000 482.0000 213.2000 ;
	    RECT 471.6000 211.0000 477.2000 211.2000 ;
	    RECT 471.4000 210.8000 477.2000 211.0000 ;
	    RECT 463.6000 209.8000 466.0000 210.4000 ;
	    RECT 467.4000 210.6000 477.2000 210.8000 ;
	    RECT 467.4000 210.2000 472.2000 210.6000 ;
	    RECT 463.6000 208.8000 464.2000 209.8000 ;
	    RECT 462.8000 208.0000 464.2000 208.8000 ;
	    RECT 465.8000 209.0000 466.6000 209.2000 ;
	    RECT 467.4000 209.0000 468.0000 210.2000 ;
	    RECT 465.8000 208.4000 468.0000 209.0000 ;
	    RECT 468.6000 209.0000 474.0000 209.6000 ;
	    RECT 468.6000 208.8000 469.4000 209.0000 ;
	    RECT 473.2000 208.8000 474.0000 209.0000 ;
	    RECT 467.0000 207.4000 467.8000 207.6000 ;
	    RECT 469.8000 207.4000 470.6000 207.6000 ;
	    RECT 463.6000 206.2000 464.4000 207.0000 ;
	    RECT 467.0000 206.8000 470.6000 207.4000 ;
	    RECT 467.8000 206.2000 468.4000 206.8000 ;
	    RECT 473.2000 206.2000 474.0000 207.0000 ;
	    RECT 463.0000 202.2000 464.2000 206.2000 ;
	    RECT 467.6000 202.2000 468.4000 206.2000 ;
	    RECT 472.0000 205.6000 474.0000 206.2000 ;
	    RECT 472.0000 202.2000 472.8000 205.6000 ;
	    RECT 476.4000 202.2000 477.2000 210.6000 ;
	    RECT 478.0000 210.2000 478.8000 210.4000 ;
	    RECT 480.0000 210.2000 480.6000 211.6000 ;
	    RECT 478.0000 209.6000 479.4000 210.2000 ;
	    RECT 480.0000 209.6000 481.0000 210.2000 ;
	    RECT 478.8000 208.4000 479.4000 209.6000 ;
	    RECT 478.8000 207.6000 479.6000 208.4000 ;
	    RECT 480.2000 202.2000 481.0000 209.6000 ;
	    RECT 486.0000 202.2000 486.8000 213.7000 ;
	    RECT 487.6000 213.8000 489.2000 214.4000 ;
	    RECT 487.6000 213.6000 488.4000 213.8000 ;
	    RECT 490.6000 213.6000 493.2000 214.4000 ;
	    RECT 489.2000 211.6000 490.0000 213.2000 ;
	    RECT 490.6000 212.3000 491.2000 213.6000 ;
	    RECT 492.4000 212.3000 493.2000 212.4000 ;
	    RECT 490.6000 211.7000 493.2000 212.3000 ;
	    RECT 490.6000 210.2000 491.2000 211.7000 ;
	    RECT 492.4000 211.6000 493.2000 211.7000 ;
	    RECT 494.0000 211.4000 494.8000 214.8000 ;
	    RECT 501.0000 214.2000 501.8000 214.4000 ;
	    RECT 506.8000 214.2000 507.4000 216.4000 ;
	    RECT 511.6000 215.0000 512.4000 219.8000 ;
	    RECT 510.0000 214.2000 511.6000 214.4000 ;
	    RECT 500.6000 213.6000 511.6000 214.2000 ;
	    RECT 498.8000 212.8000 499.6000 213.0000 ;
	    RECT 495.8000 212.2000 499.6000 212.8000 ;
	    RECT 500.6000 212.4000 501.2000 213.6000 ;
	    RECT 507.8000 213.4000 508.6000 213.6000 ;
	    RECT 509.4000 212.4000 510.2000 212.6000 ;
	    RECT 495.8000 212.0000 496.6000 212.2000 ;
	    RECT 500.4000 211.6000 501.2000 212.4000 ;
	    RECT 505.2000 211.8000 510.2000 212.4000 ;
	    RECT 505.2000 211.6000 506.0000 211.8000 ;
	    RECT 497.4000 211.4000 498.2000 211.6000 ;
	    RECT 494.0000 210.8000 498.2000 211.4000 ;
	    RECT 492.4000 210.2000 493.2000 210.4000 ;
	    RECT 490.2000 209.6000 491.2000 210.2000 ;
	    RECT 491.8000 209.6000 493.2000 210.2000 ;
	    RECT 490.2000 202.2000 491.0000 209.6000 ;
	    RECT 491.8000 208.4000 492.4000 209.6000 ;
	    RECT 491.6000 207.6000 492.4000 208.4000 ;
	    RECT 494.0000 202.2000 494.8000 210.8000 ;
	    RECT 500.6000 210.4000 501.2000 211.6000 ;
	    RECT 506.8000 211.0000 512.4000 211.2000 ;
	    RECT 506.6000 210.8000 512.4000 211.0000 ;
	    RECT 498.8000 209.8000 501.2000 210.4000 ;
	    RECT 502.6000 210.6000 512.4000 210.8000 ;
	    RECT 502.6000 210.2000 507.4000 210.6000 ;
	    RECT 498.8000 208.8000 499.4000 209.8000 ;
	    RECT 498.0000 208.0000 499.4000 208.8000 ;
	    RECT 501.0000 209.0000 501.8000 209.2000 ;
	    RECT 502.6000 209.0000 503.2000 210.2000 ;
	    RECT 501.0000 208.4000 503.2000 209.0000 ;
	    RECT 503.8000 209.0000 509.2000 209.6000 ;
	    RECT 503.8000 208.8000 504.6000 209.0000 ;
	    RECT 508.4000 208.8000 509.2000 209.0000 ;
	    RECT 502.2000 207.4000 503.0000 207.6000 ;
	    RECT 505.0000 207.4000 505.8000 207.6000 ;
	    RECT 498.8000 206.2000 499.6000 207.0000 ;
	    RECT 502.2000 206.8000 505.8000 207.4000 ;
	    RECT 503.0000 206.2000 503.6000 206.8000 ;
	    RECT 508.4000 206.2000 509.2000 207.0000 ;
	    RECT 498.2000 202.2000 499.4000 206.2000 ;
	    RECT 502.8000 202.2000 503.6000 206.2000 ;
	    RECT 507.2000 205.6000 509.2000 206.2000 ;
	    RECT 507.2000 202.2000 508.0000 205.6000 ;
	    RECT 511.6000 202.2000 512.4000 210.6000 ;
	    RECT 4.4000 192.4000 5.2000 199.8000 ;
	    RECT 3.0000 191.8000 5.2000 192.4000 ;
	    RECT 6.0000 192.4000 6.8000 199.8000 ;
	    RECT 6.0000 191.8000 8.2000 192.4000 ;
	    RECT 9.2000 191.8000 10.0000 199.8000 ;
	    RECT 10.8000 192.4000 11.6000 199.8000 ;
	    RECT 10.8000 191.8000 13.0000 192.4000 ;
	    RECT 14.0000 191.8000 14.8000 199.8000 ;
	    RECT 18.2000 192.4000 19.0000 199.8000 ;
	    RECT 19.6000 194.3000 20.4000 194.4000 ;
	    RECT 22.0000 194.3000 22.8000 199.8000 ;
	    RECT 26.2000 195.8000 27.4000 199.8000 ;
	    RECT 30.8000 195.8000 31.6000 199.8000 ;
	    RECT 35.2000 196.4000 36.0000 199.8000 ;
	    RECT 35.2000 195.8000 37.2000 196.4000 ;
	    RECT 26.8000 195.0000 27.6000 195.8000 ;
	    RECT 31.0000 195.2000 31.6000 195.8000 ;
	    RECT 30.2000 194.6000 33.8000 195.2000 ;
	    RECT 36.4000 195.0000 37.2000 195.8000 ;
	    RECT 30.2000 194.4000 31.0000 194.6000 ;
	    RECT 33.0000 194.4000 33.8000 194.6000 ;
	    RECT 19.6000 193.7000 22.8000 194.3000 ;
	    RECT 19.6000 193.6000 20.4000 193.7000 ;
	    RECT 19.8000 192.4000 20.4000 193.6000 ;
	    RECT 18.2000 191.8000 19.2000 192.4000 ;
	    RECT 19.8000 191.8000 21.2000 192.4000 ;
	    RECT 3.0000 191.2000 3.6000 191.8000 ;
	    RECT 2.4000 190.4000 3.6000 191.2000 ;
	    RECT 7.6000 191.2000 8.2000 191.8000 ;
	    RECT 7.6000 190.4000 8.8000 191.2000 ;
	    RECT 3.0000 187.4000 3.6000 190.4000 ;
	    RECT 4.4000 188.8000 5.2000 190.4000 ;
	    RECT 6.0000 188.8000 6.8000 190.4000 ;
	    RECT 7.6000 187.4000 8.2000 190.4000 ;
	    RECT 9.4000 189.6000 10.0000 191.8000 ;
	    RECT 3.0000 186.8000 5.2000 187.4000 ;
	    RECT 4.4000 182.2000 5.2000 186.8000 ;
	    RECT 6.0000 186.8000 8.2000 187.4000 ;
	    RECT 6.0000 182.2000 6.8000 186.8000 ;
	    RECT 9.2000 182.2000 10.0000 189.6000 ;
	    RECT 12.4000 191.2000 13.0000 191.8000 ;
	    RECT 12.4000 190.4000 13.6000 191.2000 ;
	    RECT 12.4000 187.4000 13.0000 190.4000 ;
	    RECT 14.2000 189.6000 14.8000 191.8000 ;
	    RECT 10.8000 186.8000 13.0000 187.4000 ;
	    RECT 14.0000 188.3000 14.8000 189.6000 ;
	    RECT 17.2000 188.8000 18.0000 190.4000 ;
	    RECT 18.6000 188.4000 19.2000 191.8000 ;
	    RECT 20.4000 191.6000 21.2000 191.8000 ;
	    RECT 22.0000 191.2000 22.8000 193.7000 ;
	    RECT 26.0000 193.2000 27.4000 194.0000 ;
	    RECT 26.8000 192.2000 27.4000 193.2000 ;
	    RECT 29.0000 193.0000 31.2000 193.6000 ;
	    RECT 29.0000 192.8000 29.8000 193.0000 ;
	    RECT 26.8000 191.6000 29.2000 192.2000 ;
	    RECT 22.0000 190.6000 26.2000 191.2000 ;
	    RECT 15.6000 188.3000 16.4000 188.4000 ;
	    RECT 14.0000 188.2000 16.4000 188.3000 ;
	    RECT 14.0000 187.7000 17.2000 188.2000 ;
	    RECT 10.8000 182.2000 11.6000 186.8000 ;
	    RECT 14.0000 182.2000 14.8000 187.7000 ;
	    RECT 15.6000 187.6000 17.2000 187.7000 ;
	    RECT 18.6000 187.6000 21.2000 188.4000 ;
	    RECT 16.4000 187.2000 17.2000 187.6000 ;
	    RECT 15.8000 186.2000 19.4000 186.6000 ;
	    RECT 20.4000 186.2000 21.0000 187.6000 ;
	    RECT 22.0000 187.2000 22.8000 190.6000 ;
	    RECT 25.4000 190.4000 26.2000 190.6000 ;
	    RECT 23.8000 189.8000 24.6000 190.0000 ;
	    RECT 23.8000 189.2000 27.6000 189.8000 ;
	    RECT 26.8000 189.0000 27.6000 189.2000 ;
	    RECT 28.6000 188.4000 29.2000 191.6000 ;
	    RECT 30.6000 191.8000 31.2000 193.0000 ;
	    RECT 31.8000 193.0000 32.6000 193.2000 ;
	    RECT 36.4000 193.0000 37.2000 193.2000 ;
	    RECT 31.8000 192.4000 37.2000 193.0000 ;
	    RECT 30.6000 191.4000 35.4000 191.8000 ;
	    RECT 39.6000 191.4000 40.4000 199.8000 ;
	    RECT 41.2000 192.4000 42.0000 199.8000 ;
	    RECT 41.2000 191.8000 43.4000 192.4000 ;
	    RECT 44.4000 191.8000 45.2000 199.8000 ;
	    RECT 46.8000 193.6000 47.6000 194.4000 ;
	    RECT 46.8000 192.4000 47.4000 193.6000 ;
	    RECT 48.2000 192.4000 49.0000 199.8000 ;
	    RECT 53.2000 193.6000 54.0000 194.4000 ;
	    RECT 53.2000 192.4000 53.8000 193.6000 ;
	    RECT 54.6000 192.4000 55.4000 199.8000 ;
	    RECT 59.6000 193.6000 60.4000 194.4000 ;
	    RECT 59.6000 192.4000 60.2000 193.6000 ;
	    RECT 61.0000 192.4000 61.8000 199.8000 ;
	    RECT 67.8000 192.6000 68.6000 199.8000 ;
	    RECT 30.6000 191.2000 40.4000 191.4000 ;
	    RECT 34.6000 191.0000 40.4000 191.2000 ;
	    RECT 34.8000 190.8000 40.4000 191.0000 ;
	    RECT 42.8000 191.2000 43.4000 191.8000 ;
	    RECT 42.8000 190.4000 44.0000 191.2000 ;
	    RECT 33.2000 190.2000 34.0000 190.4000 ;
	    RECT 33.2000 189.6000 38.2000 190.2000 ;
	    RECT 34.8000 189.4000 35.6000 189.6000 ;
	    RECT 37.4000 189.4000 38.2000 189.6000 ;
	    RECT 41.2000 188.8000 42.0000 190.4000 ;
	    RECT 35.8000 188.4000 36.6000 188.6000 ;
	    RECT 28.6000 187.8000 39.6000 188.4000 ;
	    RECT 29.0000 187.6000 29.8000 187.8000 ;
	    RECT 33.2000 187.6000 34.0000 187.8000 ;
	    RECT 22.0000 186.6000 25.8000 187.2000 ;
	    RECT 15.6000 186.0000 19.6000 186.2000 ;
	    RECT 15.6000 182.2000 16.4000 186.0000 ;
	    RECT 18.8000 182.2000 19.6000 186.0000 ;
	    RECT 20.4000 182.2000 21.2000 186.2000 ;
	    RECT 22.0000 182.2000 22.8000 186.6000 ;
	    RECT 25.0000 186.4000 25.8000 186.6000 ;
	    RECT 34.8000 185.6000 35.4000 187.8000 ;
	    RECT 38.0000 187.6000 39.6000 187.8000 ;
	    RECT 42.8000 187.4000 43.4000 190.4000 ;
	    RECT 44.6000 189.6000 45.2000 191.8000 ;
	    RECT 46.0000 191.8000 47.4000 192.4000 ;
	    RECT 48.0000 191.8000 49.0000 192.4000 ;
	    RECT 52.4000 191.8000 53.8000 192.4000 ;
	    RECT 54.4000 191.8000 55.4000 192.4000 ;
	    RECT 58.8000 191.8000 60.2000 192.4000 ;
	    RECT 60.8000 191.8000 61.8000 192.4000 ;
	    RECT 66.8000 191.8000 68.6000 192.6000 ;
	    RECT 46.0000 191.6000 46.8000 191.8000 ;
	    RECT 48.0000 190.4000 48.6000 191.8000 ;
	    RECT 52.4000 191.6000 53.2000 191.8000 ;
	    RECT 47.6000 189.6000 48.6000 190.4000 ;
	    RECT 33.0000 185.4000 33.8000 185.6000 ;
	    RECT 26.8000 184.2000 27.6000 185.0000 ;
	    RECT 31.0000 184.8000 33.8000 185.4000 ;
	    RECT 34.8000 184.8000 35.6000 185.6000 ;
	    RECT 31.0000 184.2000 31.6000 184.8000 ;
	    RECT 36.4000 184.2000 37.2000 185.0000 ;
	    RECT 26.2000 183.6000 27.6000 184.2000 ;
	    RECT 26.2000 182.2000 27.4000 183.6000 ;
	    RECT 30.8000 182.2000 31.6000 184.2000 ;
	    RECT 35.2000 183.6000 37.2000 184.2000 ;
	    RECT 35.2000 182.2000 36.0000 183.6000 ;
	    RECT 39.6000 182.2000 40.4000 187.0000 ;
	    RECT 41.2000 186.8000 43.4000 187.4000 ;
	    RECT 41.2000 182.2000 42.0000 186.8000 ;
	    RECT 44.4000 182.2000 45.2000 189.6000 ;
	    RECT 48.0000 188.4000 48.6000 189.6000 ;
	    RECT 49.2000 190.3000 50.0000 190.4000 ;
	    RECT 54.4000 190.3000 55.0000 191.8000 ;
	    RECT 58.8000 191.6000 59.6000 191.8000 ;
	    RECT 49.2000 189.7000 55.0000 190.3000 ;
	    RECT 49.2000 188.8000 50.0000 189.7000 ;
	    RECT 54.4000 188.4000 55.0000 189.7000 ;
	    RECT 55.6000 188.8000 56.4000 190.4000 ;
	    RECT 60.8000 188.4000 61.4000 191.8000 ;
	    RECT 62.0000 188.8000 62.8000 190.4000 ;
	    RECT 63.6000 190.3000 64.4000 190.4000 ;
	    RECT 67.0000 190.3000 67.6000 191.8000 ;
	    RECT 70.0000 191.4000 70.8000 199.8000 ;
	    RECT 74.4000 196.4000 75.2000 199.8000 ;
	    RECT 73.2000 195.8000 75.2000 196.4000 ;
	    RECT 78.8000 195.8000 79.6000 199.8000 ;
	    RECT 83.0000 195.8000 84.2000 199.8000 ;
	    RECT 73.2000 195.0000 74.0000 195.8000 ;
	    RECT 78.8000 195.2000 79.4000 195.8000 ;
	    RECT 76.6000 194.6000 80.2000 195.2000 ;
	    RECT 82.8000 195.0000 83.6000 195.8000 ;
	    RECT 76.6000 194.4000 77.4000 194.6000 ;
	    RECT 79.4000 194.4000 80.2000 194.6000 ;
	    RECT 73.2000 193.0000 74.0000 193.2000 ;
	    RECT 77.8000 193.0000 78.6000 193.2000 ;
	    RECT 73.2000 192.4000 78.6000 193.0000 ;
	    RECT 79.2000 193.0000 81.4000 193.6000 ;
	    RECT 79.2000 191.8000 79.8000 193.0000 ;
	    RECT 80.6000 192.8000 81.4000 193.0000 ;
	    RECT 83.0000 193.2000 84.4000 194.0000 ;
	    RECT 83.0000 192.2000 83.6000 193.2000 ;
	    RECT 75.0000 191.4000 79.8000 191.8000 ;
	    RECT 70.0000 191.2000 79.8000 191.4000 ;
	    RECT 81.2000 191.6000 83.6000 192.2000 ;
	    RECT 63.6000 189.7000 67.6000 190.3000 ;
	    RECT 63.6000 189.6000 64.4000 189.7000 ;
	    RECT 67.0000 188.4000 67.6000 189.7000 ;
	    RECT 68.4000 189.6000 69.2000 191.2000 ;
	    RECT 70.0000 191.0000 75.8000 191.2000 ;
	    RECT 70.0000 190.8000 75.6000 191.0000 ;
	    RECT 76.4000 190.3000 77.2000 190.4000 ;
	    RECT 78.0000 190.3000 78.8000 190.4000 ;
	    RECT 76.4000 190.2000 78.8000 190.3000 ;
	    RECT 72.2000 189.7000 78.8000 190.2000 ;
	    RECT 72.2000 189.6000 77.2000 189.7000 ;
	    RECT 78.0000 189.6000 78.8000 189.7000 ;
	    RECT 79.6000 190.3000 80.4000 190.4000 ;
	    RECT 81.2000 190.3000 81.8000 191.6000 ;
	    RECT 87.6000 191.2000 88.4000 199.8000 ;
	    RECT 89.2000 192.4000 90.0000 199.8000 ;
	    RECT 89.2000 191.8000 91.4000 192.4000 ;
	    RECT 92.4000 191.8000 93.2000 199.8000 ;
	    RECT 96.6000 192.4000 97.4000 199.8000 ;
	    RECT 98.0000 193.6000 98.8000 194.4000 ;
	    RECT 98.2000 192.4000 98.8000 193.6000 ;
	    RECT 101.2000 193.6000 102.0000 194.4000 ;
	    RECT 101.2000 192.4000 101.8000 193.6000 ;
	    RECT 102.6000 192.4000 103.4000 199.8000 ;
	    RECT 117.0000 198.4000 117.8000 199.8000 ;
	    RECT 116.4000 197.6000 117.8000 198.4000 ;
	    RECT 117.0000 192.8000 117.8000 197.6000 ;
	    RECT 121.2000 195.0000 122.0000 199.0000 ;
	    RECT 96.6000 191.8000 97.6000 192.4000 ;
	    RECT 98.2000 191.8000 99.6000 192.4000 ;
	    RECT 84.2000 190.6000 88.4000 191.2000 ;
	    RECT 84.2000 190.4000 85.0000 190.6000 ;
	    RECT 79.6000 189.7000 81.9000 190.3000 ;
	    RECT 85.8000 189.8000 86.6000 190.0000 ;
	    RECT 79.6000 189.6000 80.4000 189.7000 ;
	    RECT 72.2000 189.4000 73.0000 189.6000 ;
	    RECT 73.8000 188.4000 74.6000 188.6000 ;
	    RECT 81.2000 188.4000 81.8000 189.7000 ;
	    RECT 82.8000 189.2000 86.6000 189.8000 ;
	    RECT 82.8000 189.0000 83.6000 189.2000 ;
	    RECT 46.0000 187.6000 48.6000 188.4000 ;
	    RECT 50.8000 188.2000 51.6000 188.4000 ;
	    RECT 50.0000 187.6000 51.6000 188.2000 ;
	    RECT 52.4000 187.6000 55.0000 188.4000 ;
	    RECT 57.2000 188.2000 58.0000 188.4000 ;
	    RECT 56.4000 187.6000 58.0000 188.2000 ;
	    RECT 58.8000 187.6000 61.4000 188.4000 ;
	    RECT 63.6000 188.2000 64.4000 188.4000 ;
	    RECT 62.8000 187.6000 64.4000 188.2000 ;
	    RECT 66.8000 187.6000 67.6000 188.4000 ;
	    RECT 70.8000 187.8000 81.8000 188.4000 ;
	    RECT 70.8000 187.6000 72.4000 187.8000 ;
	    RECT 46.2000 186.2000 46.8000 187.6000 ;
	    RECT 50.0000 187.2000 50.8000 187.6000 ;
	    RECT 47.8000 186.2000 51.4000 186.6000 ;
	    RECT 52.6000 186.2000 53.2000 187.6000 ;
	    RECT 56.4000 187.2000 57.2000 187.6000 ;
	    RECT 54.2000 186.2000 57.8000 186.6000 ;
	    RECT 59.0000 186.2000 59.6000 187.6000 ;
	    RECT 62.8000 187.2000 63.6000 187.6000 ;
	    RECT 60.6000 186.2000 64.2000 186.6000 ;
	    RECT 46.0000 182.2000 46.8000 186.2000 ;
	    RECT 47.6000 186.0000 51.6000 186.2000 ;
	    RECT 47.6000 182.2000 48.4000 186.0000 ;
	    RECT 50.8000 182.2000 51.6000 186.0000 ;
	    RECT 52.4000 182.2000 53.2000 186.2000 ;
	    RECT 54.0000 186.0000 58.0000 186.2000 ;
	    RECT 54.0000 182.2000 54.8000 186.0000 ;
	    RECT 57.2000 182.2000 58.0000 186.0000 ;
	    RECT 58.8000 182.2000 59.6000 186.2000 ;
	    RECT 60.4000 186.0000 64.4000 186.2000 ;
	    RECT 60.4000 182.2000 61.2000 186.0000 ;
	    RECT 63.6000 182.2000 64.4000 186.0000 ;
	    RECT 65.2000 184.8000 66.0000 186.4000 ;
	    RECT 67.0000 184.2000 67.6000 187.6000 ;
	    RECT 66.8000 182.2000 67.6000 184.2000 ;
	    RECT 70.0000 182.2000 70.8000 187.0000 ;
	    RECT 75.0000 185.6000 75.6000 187.8000 ;
	    RECT 80.6000 187.6000 81.4000 187.8000 ;
	    RECT 87.6000 187.2000 88.4000 190.6000 ;
	    RECT 90.8000 191.2000 91.4000 191.8000 ;
	    RECT 90.8000 190.4000 92.0000 191.2000 ;
	    RECT 90.8000 187.4000 91.4000 190.4000 ;
	    RECT 92.6000 189.6000 93.2000 191.8000 ;
	    RECT 97.0000 190.4000 97.6000 191.8000 ;
	    RECT 98.8000 191.6000 99.6000 191.8000 ;
	    RECT 100.4000 191.8000 101.8000 192.4000 ;
	    RECT 102.4000 191.8000 103.4000 192.4000 ;
	    RECT 116.2000 192.2000 117.8000 192.8000 ;
	    RECT 100.4000 191.6000 101.2000 191.8000 ;
	    RECT 84.6000 186.6000 88.4000 187.2000 ;
	    RECT 84.6000 186.4000 85.4000 186.6000 ;
	    RECT 73.2000 184.2000 74.0000 185.0000 ;
	    RECT 74.8000 184.8000 75.6000 185.6000 ;
	    RECT 76.6000 185.4000 77.4000 185.6000 ;
	    RECT 76.6000 184.8000 79.4000 185.4000 ;
	    RECT 78.8000 184.2000 79.4000 184.8000 ;
	    RECT 82.8000 184.2000 83.6000 185.0000 ;
	    RECT 73.2000 183.6000 75.2000 184.2000 ;
	    RECT 74.4000 182.2000 75.2000 183.6000 ;
	    RECT 78.8000 182.2000 79.6000 184.2000 ;
	    RECT 82.8000 183.6000 84.2000 184.2000 ;
	    RECT 83.0000 182.2000 84.2000 183.6000 ;
	    RECT 87.6000 182.2000 88.4000 186.6000 ;
	    RECT 89.2000 186.8000 91.4000 187.4000 ;
	    RECT 89.2000 182.2000 90.0000 186.8000 ;
	    RECT 92.4000 182.2000 93.2000 189.6000 ;
	    RECT 95.6000 188.8000 96.4000 190.4000 ;
	    RECT 97.0000 189.6000 98.0000 190.4000 ;
	    RECT 98.9000 190.3000 99.5000 191.6000 ;
	    RECT 102.4000 190.3000 103.0000 191.8000 ;
	    RECT 98.9000 189.7000 103.0000 190.3000 ;
	    RECT 97.0000 188.4000 97.6000 189.6000 ;
	    RECT 102.4000 188.4000 103.0000 189.7000 ;
	    RECT 103.6000 188.8000 104.4000 190.4000 ;
	    RECT 105.2000 190.3000 106.0000 190.4000 ;
	    RECT 114.8000 190.3000 115.6000 191.2000 ;
	    RECT 105.2000 189.7000 115.6000 190.3000 ;
	    RECT 105.2000 189.6000 106.0000 189.7000 ;
	    RECT 114.8000 189.6000 115.6000 189.7000 ;
	    RECT 116.2000 188.4000 116.8000 192.2000 ;
	    RECT 121.4000 191.6000 122.0000 195.0000 ;
	    RECT 118.2000 191.0000 122.0000 191.6000 ;
	    RECT 122.8000 195.0000 123.6000 199.0000 ;
	    RECT 122.8000 191.6000 123.4000 195.0000 ;
	    RECT 127.0000 192.8000 127.8000 199.8000 ;
	    RECT 127.0000 192.2000 128.6000 192.8000 ;
	    RECT 122.8000 191.0000 126.6000 191.6000 ;
	    RECT 118.2000 189.0000 118.8000 191.0000 ;
	    RECT 94.0000 188.2000 94.8000 188.4000 ;
	    RECT 94.0000 187.6000 95.6000 188.2000 ;
	    RECT 97.0000 187.6000 99.6000 188.4000 ;
	    RECT 100.4000 187.6000 103.0000 188.4000 ;
	    RECT 105.2000 188.2000 106.0000 188.4000 ;
	    RECT 104.4000 187.6000 106.0000 188.2000 ;
	    RECT 114.8000 187.6000 116.8000 188.4000 ;
	    RECT 117.4000 188.2000 118.8000 189.0000 ;
	    RECT 119.6000 188.8000 120.4000 190.4000 ;
	    RECT 121.2000 188.8000 122.0000 190.4000 ;
	    RECT 122.8000 188.8000 123.6000 190.4000 ;
	    RECT 124.4000 188.8000 125.2000 190.4000 ;
	    RECT 126.0000 189.0000 126.6000 191.0000 ;
	    RECT 94.8000 187.2000 95.6000 187.6000 ;
	    RECT 94.2000 186.2000 97.8000 186.6000 ;
	    RECT 98.8000 186.2000 99.4000 187.6000 ;
	    RECT 100.6000 186.2000 101.2000 187.6000 ;
	    RECT 104.4000 187.2000 105.2000 187.6000 ;
	    RECT 116.2000 187.0000 116.8000 187.6000 ;
	    RECT 117.8000 187.8000 118.8000 188.2000 ;
	    RECT 126.0000 188.2000 127.4000 189.0000 ;
	    RECT 128.0000 188.4000 128.6000 192.2000 ;
	    RECT 135.0000 191.8000 137.0000 199.8000 ;
	    RECT 143.0000 192.4000 143.8000 199.8000 ;
	    RECT 144.4000 193.6000 145.2000 194.4000 ;
	    RECT 144.6000 192.4000 145.2000 193.6000 ;
	    RECT 129.2000 189.6000 130.0000 191.2000 ;
	    RECT 128.0000 188.3000 130.0000 188.4000 ;
	    RECT 130.8000 188.3000 131.6000 188.4000 ;
	    RECT 126.0000 187.8000 127.0000 188.2000 ;
	    RECT 117.8000 187.2000 122.0000 187.8000 ;
	    RECT 116.2000 186.6000 117.0000 187.0000 ;
	    RECT 102.2000 186.2000 105.8000 186.6000 ;
	    RECT 94.0000 186.0000 98.0000 186.2000 ;
	    RECT 94.0000 182.2000 94.8000 186.0000 ;
	    RECT 97.2000 182.2000 98.0000 186.0000 ;
	    RECT 98.8000 182.2000 99.6000 186.2000 ;
	    RECT 100.4000 182.2000 101.2000 186.2000 ;
	    RECT 102.0000 186.0000 106.0000 186.2000 ;
	    RECT 116.2000 186.0000 117.8000 186.6000 ;
	    RECT 102.0000 182.2000 102.8000 186.0000 ;
	    RECT 105.2000 182.2000 106.0000 186.0000 ;
	    RECT 117.0000 183.0000 117.8000 186.0000 ;
	    RECT 121.4000 185.0000 122.0000 187.2000 ;
	    RECT 121.2000 183.0000 122.0000 185.0000 ;
	    RECT 122.8000 187.2000 127.0000 187.8000 ;
	    RECT 128.0000 187.7000 131.6000 188.3000 ;
	    RECT 128.0000 187.6000 130.0000 187.7000 ;
	    RECT 130.8000 187.6000 131.6000 187.7000 ;
	    RECT 132.4000 187.6000 133.2000 189.2000 ;
	    RECT 134.0000 188.8000 134.8000 190.4000 ;
	    RECT 135.8000 188.4000 136.4000 191.8000 ;
	    RECT 142.0000 191.6000 144.0000 192.4000 ;
	    RECT 144.6000 191.8000 146.0000 192.4000 ;
	    RECT 149.4000 191.8000 151.4000 199.8000 ;
	    RECT 155.6000 193.6000 156.4000 194.4000 ;
	    RECT 155.6000 192.4000 156.2000 193.6000 ;
	    RECT 157.0000 192.4000 157.8000 199.8000 ;
	    RECT 154.8000 191.8000 156.2000 192.4000 ;
	    RECT 156.8000 191.8000 157.8000 192.4000 ;
	    RECT 161.8000 192.6000 162.6000 199.8000 ;
	    RECT 168.6000 192.6000 169.4000 199.8000 ;
	    RECT 161.8000 191.8000 163.6000 192.6000 ;
	    RECT 167.6000 191.8000 169.4000 192.6000 ;
	    RECT 171.6000 193.6000 172.4000 194.4000 ;
	    RECT 171.6000 192.4000 172.2000 193.6000 ;
	    RECT 173.0000 192.4000 173.8000 199.8000 ;
	    RECT 179.4000 196.4000 180.2000 199.8000 ;
	    RECT 179.4000 195.6000 181.2000 196.4000 ;
	    RECT 178.0000 193.6000 178.8000 194.4000 ;
	    RECT 178.0000 192.4000 178.6000 193.6000 ;
	    RECT 179.4000 192.4000 180.2000 195.6000 ;
	    RECT 170.8000 191.8000 172.2000 192.4000 ;
	    RECT 172.8000 191.8000 173.8000 192.4000 ;
	    RECT 177.2000 191.8000 178.6000 192.4000 ;
	    RECT 179.2000 191.8000 180.2000 192.4000 ;
	    RECT 186.2000 192.4000 187.0000 199.8000 ;
	    RECT 192.6000 198.4000 194.6000 199.8000 ;
	    RECT 191.6000 197.6000 194.6000 198.4000 ;
	    RECT 187.6000 193.6000 188.4000 194.4000 ;
	    RECT 187.8000 192.4000 188.4000 193.6000 ;
	    RECT 186.2000 191.8000 187.2000 192.4000 ;
	    RECT 187.8000 191.8000 189.2000 192.4000 ;
	    RECT 192.6000 191.8000 194.6000 197.6000 ;
	    RECT 198.6000 196.4000 199.4000 199.8000 ;
	    RECT 198.0000 195.6000 199.4000 196.4000 ;
	    RECT 198.6000 192.6000 199.4000 195.6000 ;
	    RECT 198.6000 191.8000 200.4000 192.6000 ;
	    RECT 205.4000 192.4000 206.2000 199.8000 ;
	    RECT 206.8000 193.6000 207.6000 194.4000 ;
	    RECT 207.0000 192.4000 207.6000 193.6000 ;
	    RECT 205.4000 191.8000 206.4000 192.4000 ;
	    RECT 207.0000 191.8000 208.4000 192.4000 ;
	    RECT 211.8000 191.8000 213.8000 199.8000 ;
	    RECT 219.8000 196.4000 220.6000 199.8000 ;
	    RECT 218.8000 195.6000 220.6000 196.4000 ;
	    RECT 219.8000 192.6000 220.6000 195.6000 ;
	    RECT 218.8000 191.8000 220.6000 192.6000 ;
	    RECT 222.0000 192.4000 222.8000 199.8000 ;
	    RECT 222.0000 191.8000 224.2000 192.4000 ;
	    RECT 225.2000 191.8000 226.0000 199.8000 ;
	    RECT 145.2000 191.6000 146.0000 191.8000 ;
	    RECT 137.2000 188.8000 138.0000 190.4000 ;
	    RECT 138.8000 190.3000 139.6000 190.4000 ;
	    RECT 138.8000 189.7000 141.1000 190.3000 ;
	    RECT 138.8000 189.6000 139.6000 189.7000 ;
	    RECT 140.5000 188.4000 141.1000 189.7000 ;
	    RECT 142.0000 188.8000 142.8000 190.4000 ;
	    RECT 143.4000 188.4000 144.0000 191.6000 ;
	    RECT 135.6000 188.2000 136.4000 188.4000 ;
	    RECT 138.8000 188.2000 139.6000 188.4000 ;
	    RECT 134.0000 187.6000 136.4000 188.2000 ;
	    RECT 138.0000 187.6000 139.6000 188.2000 ;
	    RECT 140.4000 188.2000 141.2000 188.4000 ;
	    RECT 140.4000 187.6000 142.0000 188.2000 ;
	    RECT 143.4000 187.6000 146.0000 188.4000 ;
	    RECT 146.8000 187.6000 147.6000 189.2000 ;
	    RECT 148.4000 188.8000 149.2000 190.4000 ;
	    RECT 150.2000 188.4000 150.8000 191.8000 ;
	    RECT 154.8000 191.6000 155.6000 191.8000 ;
	    RECT 151.6000 188.8000 152.4000 190.4000 ;
	    RECT 156.8000 188.4000 157.4000 191.8000 ;
	    RECT 158.0000 188.8000 158.8000 190.4000 ;
	    RECT 161.2000 189.6000 162.0000 191.2000 ;
	    RECT 162.8000 188.4000 163.4000 191.8000 ;
	    RECT 167.8000 188.4000 168.4000 191.8000 ;
	    RECT 170.8000 191.6000 171.6000 191.8000 ;
	    RECT 169.2000 189.6000 170.0000 191.2000 ;
	    RECT 172.8000 188.4000 173.4000 191.8000 ;
	    RECT 177.2000 191.6000 178.0000 191.8000 ;
	    RECT 174.0000 188.8000 174.8000 190.4000 ;
	    RECT 179.2000 188.4000 179.8000 191.8000 ;
	    RECT 180.4000 188.8000 181.2000 190.4000 ;
	    RECT 185.2000 188.8000 186.0000 190.4000 ;
	    RECT 186.6000 188.4000 187.2000 191.8000 ;
	    RECT 188.4000 191.6000 189.2000 191.8000 ;
	    RECT 191.6000 188.8000 192.4000 190.4000 ;
	    RECT 193.2000 188.4000 193.8000 191.8000 ;
	    RECT 194.8000 188.8000 195.6000 190.4000 ;
	    RECT 198.0000 189.6000 198.8000 191.2000 ;
	    RECT 150.0000 188.2000 150.8000 188.4000 ;
	    RECT 153.2000 188.3000 154.0000 188.4000 ;
	    RECT 154.8000 188.3000 157.4000 188.4000 ;
	    RECT 153.2000 188.2000 157.4000 188.3000 ;
	    RECT 159.6000 188.2000 160.4000 188.4000 ;
	    RECT 148.4000 187.6000 150.8000 188.2000 ;
	    RECT 152.4000 187.7000 157.4000 188.2000 ;
	    RECT 152.4000 187.6000 154.0000 187.7000 ;
	    RECT 154.8000 187.6000 157.4000 187.7000 ;
	    RECT 158.8000 187.6000 160.4000 188.2000 ;
	    RECT 162.8000 187.6000 163.6000 188.4000 ;
	    RECT 167.6000 187.6000 168.4000 188.4000 ;
	    RECT 170.8000 187.6000 173.4000 188.4000 ;
	    RECT 175.6000 188.2000 176.4000 188.4000 ;
	    RECT 174.8000 187.6000 176.4000 188.2000 ;
	    RECT 177.2000 187.6000 179.8000 188.4000 ;
	    RECT 182.0000 188.2000 182.8000 188.4000 ;
	    RECT 181.2000 187.6000 182.8000 188.2000 ;
	    RECT 183.6000 188.2000 184.4000 188.4000 ;
	    RECT 186.6000 188.3000 189.2000 188.4000 ;
	    RECT 190.0000 188.3000 190.8000 188.4000 ;
	    RECT 186.6000 188.2000 190.8000 188.3000 ;
	    RECT 193.2000 188.2000 194.0000 188.4000 ;
	    RECT 183.6000 187.6000 185.2000 188.2000 ;
	    RECT 186.6000 187.7000 191.6000 188.2000 ;
	    RECT 186.6000 187.6000 189.2000 187.7000 ;
	    RECT 190.0000 187.6000 191.6000 187.7000 ;
	    RECT 193.2000 187.6000 195.6000 188.2000 ;
	    RECT 196.4000 187.6000 197.2000 189.2000 ;
	    RECT 199.6000 188.4000 200.2000 191.8000 ;
	    RECT 204.4000 188.8000 205.2000 190.4000 ;
	    RECT 205.8000 188.4000 206.4000 191.8000 ;
	    RECT 207.6000 191.6000 208.4000 191.8000 ;
	    RECT 210.8000 188.8000 211.6000 190.4000 ;
	    RECT 212.4000 188.4000 213.0000 191.8000 ;
	    RECT 214.0000 188.8000 214.8000 190.4000 ;
	    RECT 199.6000 187.6000 200.4000 188.4000 ;
	    RECT 202.8000 188.2000 203.6000 188.4000 ;
	    RECT 205.8000 188.3000 208.4000 188.4000 ;
	    RECT 209.2000 188.3000 210.0000 188.4000 ;
	    RECT 205.8000 188.2000 210.0000 188.3000 ;
	    RECT 212.4000 188.2000 213.2000 188.4000 ;
	    RECT 215.6000 188.3000 216.4000 189.2000 ;
	    RECT 219.0000 188.4000 219.6000 191.8000 ;
	    RECT 223.6000 191.2000 224.2000 191.8000 ;
	    RECT 220.4000 189.6000 221.2000 191.2000 ;
	    RECT 223.6000 190.4000 224.8000 191.2000 ;
	    RECT 217.2000 188.3000 218.0000 188.4000 ;
	    RECT 202.8000 187.6000 204.4000 188.2000 ;
	    RECT 205.8000 187.7000 210.8000 188.2000 ;
	    RECT 205.8000 187.6000 208.4000 187.7000 ;
	    RECT 209.2000 187.6000 210.8000 187.7000 ;
	    RECT 212.4000 187.6000 214.8000 188.2000 ;
	    RECT 215.6000 187.7000 218.0000 188.3000 ;
	    RECT 215.6000 187.6000 216.4000 187.7000 ;
	    RECT 217.2000 187.6000 218.0000 187.7000 ;
	    RECT 218.8000 187.6000 219.6000 188.4000 ;
	    RECT 122.8000 185.0000 123.4000 187.2000 ;
	    RECT 128.0000 187.0000 128.6000 187.6000 ;
	    RECT 127.8000 186.6000 128.6000 187.0000 ;
	    RECT 127.0000 186.0000 128.6000 186.6000 ;
	    RECT 134.0000 186.2000 134.6000 187.6000 ;
	    RECT 138.0000 187.2000 138.8000 187.6000 ;
	    RECT 141.2000 187.2000 142.0000 187.6000 ;
	    RECT 135.8000 186.2000 139.4000 186.6000 ;
	    RECT 140.6000 186.2000 144.2000 186.6000 ;
	    RECT 145.2000 186.2000 145.8000 187.6000 ;
	    RECT 148.4000 186.2000 149.0000 187.6000 ;
	    RECT 152.4000 187.2000 153.2000 187.6000 ;
	    RECT 150.2000 186.2000 153.8000 186.6000 ;
	    RECT 155.0000 186.2000 155.6000 187.6000 ;
	    RECT 158.8000 187.2000 159.6000 187.6000 ;
	    RECT 156.6000 186.2000 160.2000 186.6000 ;
	    RECT 122.8000 183.0000 123.6000 185.0000 ;
	    RECT 127.0000 183.0000 127.8000 186.0000 ;
	    RECT 132.4000 182.8000 133.2000 186.2000 ;
	    RECT 134.0000 183.4000 134.8000 186.2000 ;
	    RECT 135.6000 186.0000 139.6000 186.2000 ;
	    RECT 135.6000 182.8000 136.4000 186.0000 ;
	    RECT 132.4000 182.2000 136.4000 182.8000 ;
	    RECT 138.8000 182.2000 139.6000 186.0000 ;
	    RECT 140.4000 186.0000 144.4000 186.2000 ;
	    RECT 140.4000 182.2000 141.2000 186.0000 ;
	    RECT 143.6000 182.2000 144.4000 186.0000 ;
	    RECT 145.2000 182.2000 146.0000 186.2000 ;
	    RECT 146.8000 182.8000 147.6000 186.2000 ;
	    RECT 148.4000 183.4000 149.2000 186.2000 ;
	    RECT 150.0000 186.0000 154.0000 186.2000 ;
	    RECT 150.0000 182.8000 150.8000 186.0000 ;
	    RECT 146.8000 182.2000 150.8000 182.8000 ;
	    RECT 153.2000 182.2000 154.0000 186.0000 ;
	    RECT 154.8000 182.2000 155.6000 186.2000 ;
	    RECT 156.4000 186.0000 160.4000 186.2000 ;
	    RECT 156.4000 182.2000 157.2000 186.0000 ;
	    RECT 159.6000 182.2000 160.4000 186.0000 ;
	    RECT 162.8000 184.4000 163.4000 187.6000 ;
	    RECT 164.4000 184.8000 165.2000 186.4000 ;
	    RECT 166.0000 184.8000 166.8000 186.4000 ;
	    RECT 167.8000 184.4000 168.4000 187.6000 ;
	    RECT 171.0000 186.2000 171.6000 187.6000 ;
	    RECT 174.8000 187.2000 175.6000 187.6000 ;
	    RECT 172.6000 186.2000 176.2000 186.6000 ;
	    RECT 177.4000 186.2000 178.0000 187.6000 ;
	    RECT 181.2000 187.2000 182.0000 187.6000 ;
	    RECT 184.4000 187.2000 185.2000 187.6000 ;
	    RECT 179.0000 186.2000 182.6000 186.6000 ;
	    RECT 183.8000 186.2000 187.4000 186.6000 ;
	    RECT 188.4000 186.2000 189.0000 187.6000 ;
	    RECT 190.8000 187.2000 191.6000 187.6000 ;
	    RECT 190.2000 186.2000 193.8000 186.6000 ;
	    RECT 195.0000 186.2000 195.6000 187.6000 ;
	    RECT 162.8000 182.2000 163.6000 184.4000 ;
	    RECT 167.6000 182.2000 168.4000 184.4000 ;
	    RECT 170.8000 182.2000 171.6000 186.2000 ;
	    RECT 172.4000 186.0000 176.4000 186.2000 ;
	    RECT 172.4000 182.2000 173.2000 186.0000 ;
	    RECT 175.6000 182.2000 176.4000 186.0000 ;
	    RECT 177.2000 182.2000 178.0000 186.2000 ;
	    RECT 178.8000 186.0000 182.8000 186.2000 ;
	    RECT 178.8000 182.2000 179.6000 186.0000 ;
	    RECT 182.0000 182.2000 182.8000 186.0000 ;
	    RECT 183.6000 186.0000 187.6000 186.2000 ;
	    RECT 183.6000 182.2000 184.4000 186.0000 ;
	    RECT 186.8000 182.2000 187.6000 186.0000 ;
	    RECT 188.4000 182.2000 189.2000 186.2000 ;
	    RECT 190.0000 186.0000 194.0000 186.2000 ;
	    RECT 190.0000 182.2000 190.8000 186.0000 ;
	    RECT 193.2000 182.8000 194.0000 186.0000 ;
	    RECT 194.8000 183.4000 195.6000 186.2000 ;
	    RECT 196.4000 182.8000 197.2000 186.2000 ;
	    RECT 193.2000 182.2000 197.2000 182.8000 ;
	    RECT 199.6000 184.2000 200.2000 187.6000 ;
	    RECT 203.6000 187.2000 204.4000 187.6000 ;
	    RECT 201.2000 184.8000 202.0000 186.4000 ;
	    RECT 203.0000 186.2000 206.6000 186.6000 ;
	    RECT 207.6000 186.2000 208.2000 187.6000 ;
	    RECT 210.0000 187.2000 210.8000 187.6000 ;
	    RECT 209.4000 186.2000 213.0000 186.6000 ;
	    RECT 214.2000 186.2000 214.8000 187.6000 ;
	    RECT 202.8000 186.0000 206.8000 186.2000 ;
	    RECT 199.6000 182.2000 200.4000 184.2000 ;
	    RECT 202.8000 182.2000 203.6000 186.0000 ;
	    RECT 206.0000 182.2000 206.8000 186.0000 ;
	    RECT 207.6000 182.2000 208.4000 186.2000 ;
	    RECT 209.2000 186.0000 213.2000 186.2000 ;
	    RECT 209.2000 182.2000 210.0000 186.0000 ;
	    RECT 212.4000 182.8000 213.2000 186.0000 ;
	    RECT 214.0000 183.4000 214.8000 186.2000 ;
	    RECT 215.6000 182.8000 216.4000 186.2000 ;
	    RECT 217.2000 184.8000 218.0000 186.4000 ;
	    RECT 219.0000 184.2000 219.6000 187.6000 ;
	    RECT 223.6000 187.4000 224.2000 190.4000 ;
	    RECT 225.4000 189.6000 226.0000 191.8000 ;
	    RECT 212.4000 182.2000 216.4000 182.8000 ;
	    RECT 218.8000 182.2000 219.6000 184.2000 ;
	    RECT 222.0000 186.8000 224.2000 187.4000 ;
	    RECT 222.0000 182.2000 222.8000 186.8000 ;
	    RECT 225.2000 182.2000 226.0000 189.6000 ;
	    RECT 226.8000 191.8000 227.6000 199.8000 ;
	    RECT 230.0000 192.4000 230.8000 199.8000 ;
	    RECT 228.6000 191.8000 230.8000 192.4000 ;
	    RECT 234.2000 191.8000 236.2000 199.8000 ;
	    RECT 240.4000 193.6000 241.2000 194.4000 ;
	    RECT 240.4000 192.4000 241.0000 193.6000 ;
	    RECT 241.8000 192.4000 242.6000 199.8000 ;
	    RECT 246.8000 193.6000 247.6000 194.4000 ;
	    RECT 246.8000 192.4000 247.4000 193.6000 ;
	    RECT 248.2000 192.4000 249.0000 199.8000 ;
	    RECT 239.6000 191.8000 241.0000 192.4000 ;
	    RECT 241.6000 191.8000 242.6000 192.4000 ;
	    RECT 246.0000 191.8000 247.4000 192.4000 ;
	    RECT 248.0000 191.8000 249.0000 192.4000 ;
	    RECT 252.4000 191.8000 253.2000 199.8000 ;
	    RECT 255.6000 192.4000 256.4000 199.8000 ;
	    RECT 254.2000 191.8000 256.4000 192.4000 ;
	    RECT 226.8000 189.6000 227.4000 191.8000 ;
	    RECT 228.6000 191.2000 229.2000 191.8000 ;
	    RECT 228.0000 190.4000 229.2000 191.2000 ;
	    RECT 226.8000 182.2000 227.6000 189.6000 ;
	    RECT 228.6000 187.4000 229.2000 190.4000 ;
	    RECT 230.0000 188.8000 230.8000 190.4000 ;
	    RECT 231.6000 187.6000 232.4000 189.2000 ;
	    RECT 233.2000 188.8000 234.0000 190.4000 ;
	    RECT 235.0000 188.4000 235.6000 191.8000 ;
	    RECT 239.6000 191.6000 240.4000 191.8000 ;
	    RECT 236.4000 188.8000 237.2000 190.4000 ;
	    RECT 241.6000 188.4000 242.2000 191.8000 ;
	    RECT 246.0000 191.6000 246.8000 191.8000 ;
	    RECT 242.8000 188.8000 243.6000 190.4000 ;
	    RECT 244.4000 190.3000 245.2000 190.4000 ;
	    RECT 246.1000 190.3000 246.7000 191.6000 ;
	    RECT 244.4000 189.7000 246.7000 190.3000 ;
	    RECT 244.4000 189.6000 245.2000 189.7000 ;
	    RECT 248.0000 188.4000 248.6000 191.8000 ;
	    RECT 249.2000 188.8000 250.0000 190.4000 ;
	    RECT 252.4000 189.6000 253.0000 191.8000 ;
	    RECT 254.2000 191.2000 254.8000 191.8000 ;
	    RECT 263.6000 191.6000 264.4000 193.2000 ;
	    RECT 253.6000 190.4000 254.8000 191.2000 ;
	    RECT 234.8000 188.2000 235.6000 188.4000 ;
	    RECT 238.0000 188.3000 238.8000 188.4000 ;
	    RECT 239.6000 188.3000 242.2000 188.4000 ;
	    RECT 238.0000 188.2000 242.2000 188.3000 ;
	    RECT 244.4000 188.2000 245.2000 188.4000 ;
	    RECT 233.2000 187.6000 235.6000 188.2000 ;
	    RECT 237.2000 187.7000 242.2000 188.2000 ;
	    RECT 237.2000 187.6000 238.8000 187.7000 ;
	    RECT 239.6000 187.6000 242.2000 187.7000 ;
	    RECT 243.6000 187.6000 245.2000 188.2000 ;
	    RECT 246.0000 187.6000 248.6000 188.4000 ;
	    RECT 250.8000 188.2000 251.6000 188.4000 ;
	    RECT 250.0000 187.6000 251.6000 188.2000 ;
	    RECT 228.6000 186.8000 230.8000 187.4000 ;
	    RECT 230.0000 182.2000 230.8000 186.8000 ;
	    RECT 233.2000 186.2000 233.8000 187.6000 ;
	    RECT 237.2000 187.2000 238.0000 187.6000 ;
	    RECT 235.0000 186.2000 238.6000 186.6000 ;
	    RECT 239.8000 186.2000 240.4000 187.6000 ;
	    RECT 243.6000 187.2000 244.4000 187.6000 ;
	    RECT 241.4000 186.2000 245.0000 186.6000 ;
	    RECT 246.2000 186.2000 246.8000 187.6000 ;
	    RECT 250.0000 187.2000 250.8000 187.6000 ;
	    RECT 247.8000 186.2000 251.4000 186.6000 ;
	    RECT 231.6000 182.8000 232.4000 186.2000 ;
	    RECT 233.2000 183.4000 234.0000 186.2000 ;
	    RECT 234.8000 186.0000 238.8000 186.2000 ;
	    RECT 234.8000 182.8000 235.6000 186.0000 ;
	    RECT 231.6000 182.2000 235.6000 182.8000 ;
	    RECT 238.0000 182.2000 238.8000 186.0000 ;
	    RECT 239.6000 182.2000 240.4000 186.2000 ;
	    RECT 241.2000 186.0000 245.2000 186.2000 ;
	    RECT 241.2000 182.2000 242.0000 186.0000 ;
	    RECT 244.4000 182.2000 245.2000 186.0000 ;
	    RECT 246.0000 182.2000 246.8000 186.2000 ;
	    RECT 247.6000 186.0000 251.6000 186.2000 ;
	    RECT 247.6000 182.2000 248.4000 186.0000 ;
	    RECT 250.8000 182.2000 251.6000 186.0000 ;
	    RECT 252.4000 182.2000 253.2000 189.6000 ;
	    RECT 254.2000 187.4000 254.8000 190.4000 ;
	    RECT 255.6000 188.8000 256.4000 190.4000 ;
	    RECT 254.2000 186.8000 256.4000 187.4000 ;
	    RECT 255.6000 182.2000 256.4000 186.8000 ;
	    RECT 265.2000 186.2000 266.0000 199.8000 ;
	    RECT 266.8000 194.3000 267.6000 194.4000 ;
	    RECT 268.4000 194.3000 269.2000 199.8000 ;
	    RECT 272.6000 195.8000 273.8000 199.8000 ;
	    RECT 277.2000 195.8000 278.0000 199.8000 ;
	    RECT 281.6000 196.4000 282.4000 199.8000 ;
	    RECT 281.6000 195.8000 283.6000 196.4000 ;
	    RECT 273.2000 195.0000 274.0000 195.8000 ;
	    RECT 277.4000 195.2000 278.0000 195.8000 ;
	    RECT 276.6000 194.6000 280.2000 195.2000 ;
	    RECT 282.8000 195.0000 283.6000 195.8000 ;
	    RECT 276.6000 194.4000 277.4000 194.6000 ;
	    RECT 279.4000 194.4000 280.2000 194.6000 ;
	    RECT 266.8000 193.7000 269.2000 194.3000 ;
	    RECT 266.8000 193.6000 267.6000 193.7000 ;
	    RECT 268.4000 191.2000 269.2000 193.7000 ;
	    RECT 272.4000 193.2000 273.8000 194.0000 ;
	    RECT 273.2000 192.2000 273.8000 193.2000 ;
	    RECT 275.4000 193.0000 277.6000 193.6000 ;
	    RECT 275.4000 192.8000 276.2000 193.0000 ;
	    RECT 273.2000 191.6000 275.6000 192.2000 ;
	    RECT 268.4000 190.6000 272.6000 191.2000 ;
	    RECT 266.8000 186.8000 267.6000 188.4000 ;
	    RECT 268.4000 187.2000 269.2000 190.6000 ;
	    RECT 271.8000 190.4000 272.6000 190.6000 ;
	    RECT 270.2000 189.8000 271.0000 190.0000 ;
	    RECT 270.2000 189.2000 274.0000 189.8000 ;
	    RECT 273.2000 189.0000 274.0000 189.2000 ;
	    RECT 275.0000 188.4000 275.6000 191.6000 ;
	    RECT 277.0000 191.8000 277.6000 193.0000 ;
	    RECT 278.2000 193.0000 279.0000 193.2000 ;
	    RECT 282.8000 193.0000 283.6000 193.2000 ;
	    RECT 278.2000 192.4000 283.6000 193.0000 ;
	    RECT 277.0000 191.4000 281.8000 191.8000 ;
	    RECT 286.0000 191.4000 286.8000 199.8000 ;
	    RECT 277.0000 191.2000 286.8000 191.4000 ;
	    RECT 281.0000 191.0000 286.8000 191.2000 ;
	    RECT 281.2000 190.8000 286.8000 191.0000 ;
	    RECT 287.6000 191.8000 288.4000 199.8000 ;
	    RECT 290.8000 192.4000 291.6000 199.8000 ;
	    RECT 293.2000 193.6000 294.0000 194.4000 ;
	    RECT 293.2000 192.4000 293.8000 193.6000 ;
	    RECT 294.6000 192.4000 295.4000 199.8000 ;
	    RECT 289.4000 191.8000 291.6000 192.4000 ;
	    RECT 292.4000 191.8000 293.8000 192.4000 ;
	    RECT 294.4000 191.8000 295.4000 192.4000 ;
	    RECT 298.8000 191.8000 299.6000 199.8000 ;
	    RECT 302.0000 192.4000 302.8000 199.8000 ;
	    RECT 300.6000 191.8000 302.8000 192.4000 ;
	    RECT 303.6000 191.8000 304.4000 199.8000 ;
	    RECT 306.8000 192.4000 307.6000 199.8000 ;
	    RECT 305.4000 191.8000 307.6000 192.4000 ;
	    RECT 279.6000 190.2000 280.4000 190.4000 ;
	    RECT 279.6000 189.6000 284.6000 190.2000 ;
	    RECT 283.8000 189.4000 284.6000 189.6000 ;
	    RECT 287.6000 189.6000 288.2000 191.8000 ;
	    RECT 289.4000 191.2000 290.0000 191.8000 ;
	    RECT 292.4000 191.6000 293.2000 191.8000 ;
	    RECT 288.8000 190.4000 290.0000 191.2000 ;
	    RECT 282.2000 188.4000 283.0000 188.6000 ;
	    RECT 275.0000 187.8000 286.0000 188.4000 ;
	    RECT 275.4000 187.6000 276.2000 187.8000 ;
	    RECT 264.2000 185.6000 266.0000 186.2000 ;
	    RECT 268.4000 186.6000 272.2000 187.2000 ;
	    RECT 264.2000 184.4000 265.0000 185.6000 ;
	    RECT 263.6000 183.6000 265.0000 184.4000 ;
	    RECT 264.2000 182.2000 265.0000 183.6000 ;
	    RECT 268.4000 182.2000 269.2000 186.6000 ;
	    RECT 271.4000 186.4000 272.2000 186.6000 ;
	    RECT 281.2000 186.4000 281.8000 187.8000 ;
	    RECT 284.4000 187.6000 286.0000 187.8000 ;
	    RECT 279.4000 185.4000 280.2000 185.6000 ;
	    RECT 273.2000 184.2000 274.0000 185.0000 ;
	    RECT 277.4000 184.8000 280.2000 185.4000 ;
	    RECT 281.2000 184.8000 282.0000 186.4000 ;
	    RECT 277.4000 184.2000 278.0000 184.8000 ;
	    RECT 282.8000 184.2000 283.6000 185.0000 ;
	    RECT 272.6000 183.6000 274.0000 184.2000 ;
	    RECT 272.6000 182.2000 273.8000 183.6000 ;
	    RECT 277.2000 182.2000 278.0000 184.2000 ;
	    RECT 281.6000 183.6000 283.6000 184.2000 ;
	    RECT 281.6000 182.2000 282.4000 183.6000 ;
	    RECT 286.0000 182.2000 286.8000 187.0000 ;
	    RECT 287.6000 182.2000 288.4000 189.6000 ;
	    RECT 289.4000 187.4000 290.0000 190.4000 ;
	    RECT 290.8000 188.8000 291.6000 190.4000 ;
	    RECT 294.4000 188.4000 295.0000 191.8000 ;
	    RECT 295.6000 188.8000 296.4000 190.4000 ;
	    RECT 298.8000 189.6000 299.4000 191.8000 ;
	    RECT 300.6000 191.2000 301.2000 191.8000 ;
	    RECT 300.0000 190.4000 301.2000 191.2000 ;
	    RECT 292.4000 187.6000 295.0000 188.4000 ;
	    RECT 297.2000 188.2000 298.0000 188.4000 ;
	    RECT 296.4000 187.6000 298.0000 188.2000 ;
	    RECT 289.4000 186.8000 291.6000 187.4000 ;
	    RECT 290.8000 182.2000 291.6000 186.8000 ;
	    RECT 292.6000 186.2000 293.2000 187.6000 ;
	    RECT 296.4000 187.2000 297.2000 187.6000 ;
	    RECT 294.2000 186.2000 297.8000 186.6000 ;
	    RECT 292.4000 182.2000 293.2000 186.2000 ;
	    RECT 294.0000 186.0000 298.0000 186.2000 ;
	    RECT 294.0000 182.2000 294.8000 186.0000 ;
	    RECT 297.2000 182.2000 298.0000 186.0000 ;
	    RECT 298.8000 182.2000 299.6000 189.6000 ;
	    RECT 300.6000 187.4000 301.2000 190.4000 ;
	    RECT 302.0000 188.8000 302.8000 190.4000 ;
	    RECT 303.6000 189.6000 304.2000 191.8000 ;
	    RECT 305.4000 191.2000 306.0000 191.8000 ;
	    RECT 304.8000 190.4000 306.0000 191.2000 ;
	    RECT 300.6000 186.8000 302.8000 187.4000 ;
	    RECT 302.0000 182.2000 302.8000 186.8000 ;
	    RECT 303.6000 182.2000 304.4000 189.6000 ;
	    RECT 305.4000 187.4000 306.0000 190.4000 ;
	    RECT 306.8000 188.8000 307.6000 190.4000 ;
	    RECT 310.0000 190.3000 310.8000 199.8000 ;
	    RECT 314.0000 193.6000 314.8000 194.4000 ;
	    RECT 311.6000 191.6000 312.4000 193.2000 ;
	    RECT 314.0000 192.4000 314.6000 193.6000 ;
	    RECT 315.4000 192.4000 316.2000 199.8000 ;
	    RECT 313.2000 191.8000 314.6000 192.4000 ;
	    RECT 313.2000 191.6000 314.0000 191.8000 ;
	    RECT 315.2000 191.6000 317.2000 192.4000 ;
	    RECT 313.3000 190.3000 313.9000 191.6000 ;
	    RECT 310.0000 189.7000 313.9000 190.3000 ;
	    RECT 305.4000 186.8000 307.6000 187.4000 ;
	    RECT 308.4000 186.8000 309.2000 188.4000 ;
	    RECT 306.8000 182.2000 307.6000 186.8000 ;
	    RECT 310.0000 186.2000 310.8000 189.7000 ;
	    RECT 315.2000 188.4000 315.8000 191.6000 ;
	    RECT 319.6000 191.2000 320.4000 199.8000 ;
	    RECT 323.8000 195.8000 325.0000 199.8000 ;
	    RECT 328.4000 195.8000 329.2000 199.8000 ;
	    RECT 332.8000 196.4000 333.6000 199.8000 ;
	    RECT 332.8000 195.8000 334.8000 196.4000 ;
	    RECT 324.4000 195.0000 325.2000 195.8000 ;
	    RECT 328.6000 195.2000 329.2000 195.8000 ;
	    RECT 327.8000 194.6000 331.4000 195.2000 ;
	    RECT 334.0000 195.0000 334.8000 195.8000 ;
	    RECT 327.8000 194.4000 328.6000 194.6000 ;
	    RECT 330.6000 194.4000 331.4000 194.6000 ;
	    RECT 323.6000 193.2000 325.0000 194.0000 ;
	    RECT 324.4000 192.2000 325.0000 193.2000 ;
	    RECT 326.6000 193.0000 328.8000 193.6000 ;
	    RECT 326.6000 192.8000 327.4000 193.0000 ;
	    RECT 324.4000 191.6000 326.8000 192.2000 ;
	    RECT 319.6000 190.6000 323.8000 191.2000 ;
	    RECT 316.4000 188.8000 317.2000 190.4000 ;
	    RECT 313.2000 187.6000 315.8000 188.4000 ;
	    RECT 318.0000 188.2000 318.8000 188.4000 ;
	    RECT 317.2000 187.6000 318.8000 188.2000 ;
	    RECT 313.4000 186.2000 314.0000 187.6000 ;
	    RECT 317.2000 187.2000 318.0000 187.6000 ;
	    RECT 319.6000 187.2000 320.4000 190.6000 ;
	    RECT 323.0000 190.4000 323.8000 190.6000 ;
	    RECT 321.4000 189.8000 322.2000 190.0000 ;
	    RECT 321.4000 189.2000 325.2000 189.8000 ;
	    RECT 324.4000 189.0000 325.2000 189.2000 ;
	    RECT 326.2000 188.4000 326.8000 191.6000 ;
	    RECT 328.2000 191.8000 328.8000 193.0000 ;
	    RECT 329.4000 193.0000 330.2000 193.2000 ;
	    RECT 334.0000 193.0000 334.8000 193.2000 ;
	    RECT 329.4000 192.4000 334.8000 193.0000 ;
	    RECT 328.2000 191.4000 333.0000 191.8000 ;
	    RECT 337.2000 191.4000 338.0000 199.8000 ;
	    RECT 338.8000 192.4000 339.6000 199.8000 ;
	    RECT 338.8000 191.8000 341.0000 192.4000 ;
	    RECT 342.0000 191.8000 342.8000 199.8000 ;
	    RECT 343.6000 192.4000 344.4000 199.8000 ;
	    RECT 343.6000 191.8000 345.8000 192.4000 ;
	    RECT 346.8000 191.8000 347.6000 199.8000 ;
	    RECT 348.4000 192.4000 349.2000 199.8000 ;
	    RECT 348.4000 191.8000 350.6000 192.4000 ;
	    RECT 351.6000 191.8000 352.4000 199.8000 ;
	    RECT 328.2000 191.2000 338.0000 191.4000 ;
	    RECT 332.2000 191.0000 338.0000 191.2000 ;
	    RECT 332.4000 190.8000 338.0000 191.0000 ;
	    RECT 340.4000 191.2000 341.0000 191.8000 ;
	    RECT 340.4000 190.4000 341.6000 191.2000 ;
	    RECT 330.8000 190.2000 331.6000 190.4000 ;
	    RECT 330.8000 189.6000 335.8000 190.2000 ;
	    RECT 335.0000 189.4000 335.8000 189.6000 ;
	    RECT 338.8000 188.8000 339.6000 190.4000 ;
	    RECT 333.4000 188.4000 334.2000 188.6000 ;
	    RECT 326.2000 187.8000 337.2000 188.4000 ;
	    RECT 326.6000 187.6000 327.4000 187.8000 ;
	    RECT 319.6000 186.6000 323.4000 187.2000 ;
	    RECT 315.0000 186.2000 318.6000 186.6000 ;
	    RECT 310.0000 185.6000 311.8000 186.2000 ;
	    RECT 311.0000 182.2000 311.8000 185.6000 ;
	    RECT 313.2000 182.2000 314.0000 186.2000 ;
	    RECT 314.8000 186.0000 318.8000 186.2000 ;
	    RECT 314.8000 182.2000 315.6000 186.0000 ;
	    RECT 318.0000 182.2000 318.8000 186.0000 ;
	    RECT 319.6000 182.2000 320.4000 186.6000 ;
	    RECT 322.6000 186.4000 323.4000 186.6000 ;
	    RECT 332.4000 186.4000 333.0000 187.8000 ;
	    RECT 335.6000 187.6000 337.2000 187.8000 ;
	    RECT 340.4000 187.4000 341.0000 190.4000 ;
	    RECT 342.2000 189.6000 342.8000 191.8000 ;
	    RECT 345.2000 191.2000 345.8000 191.8000 ;
	    RECT 345.2000 190.4000 346.4000 191.2000 ;
	    RECT 330.6000 185.4000 331.4000 185.6000 ;
	    RECT 324.4000 184.2000 325.2000 185.0000 ;
	    RECT 328.6000 184.8000 331.4000 185.4000 ;
	    RECT 332.4000 184.8000 333.2000 186.4000 ;
	    RECT 328.6000 184.2000 329.2000 184.8000 ;
	    RECT 334.0000 184.2000 334.8000 185.0000 ;
	    RECT 323.8000 183.6000 325.2000 184.2000 ;
	    RECT 323.8000 182.2000 325.0000 183.6000 ;
	    RECT 328.4000 182.2000 329.2000 184.2000 ;
	    RECT 332.8000 183.6000 334.8000 184.2000 ;
	    RECT 332.8000 182.2000 333.6000 183.6000 ;
	    RECT 337.2000 182.2000 338.0000 187.0000 ;
	    RECT 338.8000 186.8000 341.0000 187.4000 ;
	    RECT 338.8000 182.2000 339.6000 186.8000 ;
	    RECT 342.0000 182.2000 342.8000 189.6000 ;
	    RECT 343.6000 188.8000 344.4000 190.4000 ;
	    RECT 345.2000 187.4000 345.8000 190.4000 ;
	    RECT 347.0000 189.6000 347.6000 191.8000 ;
	    RECT 350.0000 191.2000 350.6000 191.8000 ;
	    RECT 350.0000 190.4000 351.2000 191.2000 ;
	    RECT 343.6000 186.8000 345.8000 187.4000 ;
	    RECT 343.6000 182.2000 344.4000 186.8000 ;
	    RECT 346.8000 182.2000 347.6000 189.6000 ;
	    RECT 348.4000 188.8000 349.2000 190.4000 ;
	    RECT 350.0000 187.4000 350.6000 190.4000 ;
	    RECT 351.8000 189.6000 352.4000 191.8000 ;
	    RECT 348.4000 186.8000 350.6000 187.4000 ;
	    RECT 348.4000 182.2000 349.2000 186.8000 ;
	    RECT 351.6000 182.2000 352.4000 189.6000 ;
	    RECT 354.8000 190.3000 355.6000 199.8000 ;
	    RECT 358.8000 193.6000 359.6000 194.4000 ;
	    RECT 356.4000 191.6000 357.2000 193.2000 ;
	    RECT 358.8000 192.4000 359.4000 193.6000 ;
	    RECT 360.2000 192.4000 361.0000 199.8000 ;
	    RECT 358.0000 191.8000 359.4000 192.4000 ;
	    RECT 360.0000 191.8000 361.0000 192.4000 ;
	    RECT 358.0000 191.6000 358.8000 191.8000 ;
	    RECT 358.1000 190.3000 358.7000 191.6000 ;
	    RECT 354.8000 189.7000 358.7000 190.3000 ;
	    RECT 353.2000 186.8000 354.0000 188.4000 ;
	    RECT 354.8000 186.2000 355.6000 189.7000 ;
	    RECT 360.0000 188.4000 360.6000 191.8000 ;
	    RECT 364.4000 191.2000 365.2000 199.8000 ;
	    RECT 368.6000 195.8000 369.8000 199.8000 ;
	    RECT 373.2000 195.8000 374.0000 199.8000 ;
	    RECT 377.6000 196.4000 378.4000 199.8000 ;
	    RECT 377.6000 195.8000 379.6000 196.4000 ;
	    RECT 369.2000 195.0000 370.0000 195.8000 ;
	    RECT 373.4000 195.2000 374.0000 195.8000 ;
	    RECT 372.6000 194.6000 376.2000 195.2000 ;
	    RECT 378.8000 195.0000 379.6000 195.8000 ;
	    RECT 372.6000 194.4000 373.4000 194.6000 ;
	    RECT 375.4000 194.4000 376.2000 194.6000 ;
	    RECT 368.4000 193.2000 369.8000 194.0000 ;
	    RECT 369.2000 192.2000 369.8000 193.2000 ;
	    RECT 371.4000 193.0000 373.6000 193.6000 ;
	    RECT 371.4000 192.8000 372.2000 193.0000 ;
	    RECT 369.2000 191.6000 371.6000 192.2000 ;
	    RECT 364.4000 190.6000 368.6000 191.2000 ;
	    RECT 361.2000 190.3000 362.0000 190.4000 ;
	    RECT 362.8000 190.3000 363.6000 190.4000 ;
	    RECT 361.2000 189.7000 363.6000 190.3000 ;
	    RECT 361.2000 188.8000 362.0000 189.7000 ;
	    RECT 362.8000 189.6000 363.6000 189.7000 ;
	    RECT 358.0000 187.6000 360.6000 188.4000 ;
	    RECT 362.8000 188.2000 363.6000 188.4000 ;
	    RECT 362.0000 187.6000 363.6000 188.2000 ;
	    RECT 358.2000 186.2000 358.8000 187.6000 ;
	    RECT 362.0000 187.2000 362.8000 187.6000 ;
	    RECT 364.4000 187.2000 365.2000 190.6000 ;
	    RECT 367.8000 190.4000 368.6000 190.6000 ;
	    RECT 366.2000 189.8000 367.0000 190.0000 ;
	    RECT 366.2000 189.2000 370.0000 189.8000 ;
	    RECT 369.2000 189.0000 370.0000 189.2000 ;
	    RECT 371.0000 188.4000 371.6000 191.6000 ;
	    RECT 373.0000 191.8000 373.6000 193.0000 ;
	    RECT 374.2000 193.0000 375.0000 193.2000 ;
	    RECT 378.8000 193.0000 379.6000 193.2000 ;
	    RECT 374.2000 192.4000 379.6000 193.0000 ;
	    RECT 373.0000 191.4000 377.8000 191.8000 ;
	    RECT 382.0000 191.4000 382.8000 199.8000 ;
	    RECT 373.0000 191.2000 382.8000 191.4000 ;
	    RECT 377.0000 191.0000 382.8000 191.2000 ;
	    RECT 377.2000 190.8000 382.8000 191.0000 ;
	    RECT 375.6000 190.2000 376.4000 190.4000 ;
	    RECT 375.6000 189.6000 380.6000 190.2000 ;
	    RECT 379.8000 189.4000 380.6000 189.6000 ;
	    RECT 378.2000 188.4000 379.0000 188.6000 ;
	    RECT 371.0000 187.8000 382.0000 188.4000 ;
	    RECT 371.4000 187.6000 372.2000 187.8000 ;
	    RECT 364.4000 186.6000 368.2000 187.2000 ;
	    RECT 359.8000 186.2000 363.4000 186.6000 ;
	    RECT 354.8000 185.6000 356.6000 186.2000 ;
	    RECT 355.8000 182.2000 356.6000 185.6000 ;
	    RECT 358.0000 182.2000 358.8000 186.2000 ;
	    RECT 359.6000 186.0000 363.6000 186.2000 ;
	    RECT 359.6000 182.2000 360.4000 186.0000 ;
	    RECT 362.8000 182.2000 363.6000 186.0000 ;
	    RECT 364.4000 182.2000 365.2000 186.6000 ;
	    RECT 367.4000 186.4000 368.2000 186.6000 ;
	    RECT 377.2000 186.4000 377.8000 187.8000 ;
	    RECT 380.4000 187.6000 382.0000 187.8000 ;
	    RECT 375.4000 185.4000 376.2000 185.6000 ;
	    RECT 369.2000 184.2000 370.0000 185.0000 ;
	    RECT 373.4000 184.8000 376.2000 185.4000 ;
	    RECT 377.2000 184.8000 378.0000 186.4000 ;
	    RECT 373.4000 184.2000 374.0000 184.8000 ;
	    RECT 378.8000 184.2000 379.6000 185.0000 ;
	    RECT 368.6000 183.6000 370.0000 184.2000 ;
	    RECT 368.6000 182.2000 369.8000 183.6000 ;
	    RECT 373.2000 182.2000 374.0000 184.2000 ;
	    RECT 377.6000 183.6000 379.6000 184.2000 ;
	    RECT 377.6000 182.2000 378.4000 183.6000 ;
	    RECT 382.0000 182.2000 382.8000 187.0000 ;
	    RECT 383.6000 184.8000 384.4000 186.4000 ;
	    RECT 385.2000 182.2000 386.0000 199.8000 ;
	    RECT 386.8000 191.2000 387.6000 199.8000 ;
	    RECT 391.0000 195.8000 392.2000 199.8000 ;
	    RECT 395.6000 195.8000 396.4000 199.8000 ;
	    RECT 400.0000 196.4000 400.8000 199.8000 ;
	    RECT 400.0000 195.8000 402.0000 196.4000 ;
	    RECT 391.6000 195.0000 392.4000 195.8000 ;
	    RECT 395.8000 195.2000 396.4000 195.8000 ;
	    RECT 395.0000 194.6000 398.6000 195.2000 ;
	    RECT 401.2000 195.0000 402.0000 195.8000 ;
	    RECT 395.0000 194.4000 395.8000 194.6000 ;
	    RECT 397.8000 194.4000 398.6000 194.6000 ;
	    RECT 390.8000 193.2000 392.2000 194.0000 ;
	    RECT 391.6000 192.2000 392.2000 193.2000 ;
	    RECT 393.8000 193.0000 396.0000 193.6000 ;
	    RECT 393.8000 192.8000 394.6000 193.0000 ;
	    RECT 391.6000 191.6000 394.0000 192.2000 ;
	    RECT 386.8000 190.6000 391.0000 191.2000 ;
	    RECT 386.8000 187.2000 387.6000 190.6000 ;
	    RECT 390.2000 190.4000 391.0000 190.6000 ;
	    RECT 388.6000 189.8000 389.4000 190.0000 ;
	    RECT 388.6000 189.2000 392.4000 189.8000 ;
	    RECT 391.6000 189.0000 392.4000 189.2000 ;
	    RECT 393.4000 188.4000 394.0000 191.6000 ;
	    RECT 395.4000 191.8000 396.0000 193.0000 ;
	    RECT 396.6000 193.0000 397.4000 193.2000 ;
	    RECT 401.2000 193.0000 402.0000 193.2000 ;
	    RECT 396.6000 192.4000 402.0000 193.0000 ;
	    RECT 395.4000 191.4000 400.2000 191.8000 ;
	    RECT 404.4000 191.4000 405.2000 199.8000 ;
	    RECT 415.0000 192.4000 415.8000 199.8000 ;
	    RECT 416.4000 193.6000 417.2000 194.4000 ;
	    RECT 416.6000 192.4000 417.2000 193.6000 ;
	    RECT 418.8000 192.4000 419.6000 199.8000 ;
	    RECT 415.0000 191.8000 416.0000 192.4000 ;
	    RECT 416.6000 191.8000 418.0000 192.4000 ;
	    RECT 418.8000 191.8000 421.0000 192.4000 ;
	    RECT 422.0000 191.8000 422.8000 199.8000 ;
	    RECT 423.6000 192.4000 424.4000 199.8000 ;
	    RECT 426.8000 194.3000 427.6000 199.8000 ;
	    RECT 430.0000 195.8000 430.8000 199.8000 ;
	    RECT 430.2000 195.6000 430.8000 195.8000 ;
	    RECT 433.2000 195.8000 434.0000 199.8000 ;
	    RECT 433.2000 195.6000 433.8000 195.8000 ;
	    RECT 430.2000 195.0000 433.8000 195.6000 ;
	    RECT 430.0000 194.3000 430.8000 194.4000 ;
	    RECT 426.8000 193.7000 430.8000 194.3000 ;
	    RECT 423.6000 191.8000 425.8000 192.4000 ;
	    RECT 426.8000 191.8000 427.6000 193.7000 ;
	    RECT 430.0000 193.6000 430.8000 193.7000 ;
	    RECT 431.6000 192.8000 432.4000 194.4000 ;
	    RECT 395.4000 191.2000 405.2000 191.4000 ;
	    RECT 399.4000 191.0000 405.2000 191.2000 ;
	    RECT 399.6000 190.8000 405.2000 191.0000 ;
	    RECT 398.0000 190.2000 398.8000 190.4000 ;
	    RECT 398.0000 189.6000 403.0000 190.2000 ;
	    RECT 399.6000 189.4000 400.4000 189.6000 ;
	    RECT 402.2000 189.4000 403.0000 189.6000 ;
	    RECT 414.0000 188.8000 414.8000 190.4000 ;
	    RECT 400.6000 188.4000 401.4000 188.6000 ;
	    RECT 415.4000 188.4000 416.0000 191.8000 ;
	    RECT 417.2000 191.6000 418.0000 191.8000 ;
	    RECT 420.4000 191.2000 421.0000 191.8000 ;
	    RECT 420.4000 190.4000 421.6000 191.2000 ;
	    RECT 418.8000 188.8000 419.6000 190.4000 ;
	    RECT 393.4000 187.8000 404.4000 188.4000 ;
	    RECT 393.8000 187.6000 394.6000 187.8000 ;
	    RECT 386.8000 186.6000 390.6000 187.2000 ;
	    RECT 386.8000 182.2000 387.6000 186.6000 ;
	    RECT 389.8000 186.4000 390.6000 186.6000 ;
	    RECT 399.6000 185.6000 400.2000 187.8000 ;
	    RECT 402.8000 187.6000 404.4000 187.8000 ;
	    RECT 410.8000 188.3000 411.6000 188.4000 ;
	    RECT 412.4000 188.3000 413.2000 188.4000 ;
	    RECT 410.8000 188.2000 413.2000 188.3000 ;
	    RECT 410.8000 187.7000 414.0000 188.2000 ;
	    RECT 410.8000 187.6000 411.6000 187.7000 ;
	    RECT 412.4000 187.6000 414.0000 187.7000 ;
	    RECT 415.4000 187.6000 418.0000 188.4000 ;
	    RECT 413.2000 187.2000 414.0000 187.6000 ;
	    RECT 397.8000 185.4000 398.6000 185.6000 ;
	    RECT 391.6000 184.2000 392.4000 185.0000 ;
	    RECT 395.8000 184.8000 398.6000 185.4000 ;
	    RECT 399.6000 184.8000 400.4000 185.6000 ;
	    RECT 395.8000 184.2000 396.4000 184.8000 ;
	    RECT 401.2000 184.2000 402.0000 185.0000 ;
	    RECT 391.0000 183.6000 392.4000 184.2000 ;
	    RECT 391.0000 182.2000 392.2000 183.6000 ;
	    RECT 395.6000 182.2000 396.4000 184.2000 ;
	    RECT 400.0000 183.6000 402.0000 184.2000 ;
	    RECT 400.0000 182.2000 400.8000 183.6000 ;
	    RECT 404.4000 182.2000 405.2000 187.0000 ;
	    RECT 412.6000 186.2000 416.2000 186.6000 ;
	    RECT 417.2000 186.2000 417.8000 187.6000 ;
	    RECT 420.4000 187.4000 421.0000 190.4000 ;
	    RECT 422.2000 189.6000 422.8000 191.8000 ;
	    RECT 425.2000 191.2000 425.8000 191.8000 ;
	    RECT 425.2000 190.4000 426.4000 191.2000 ;
	    RECT 418.8000 186.8000 421.0000 187.4000 ;
	    RECT 412.4000 186.0000 416.4000 186.2000 ;
	    RECT 412.4000 182.2000 413.2000 186.0000 ;
	    RECT 415.6000 182.2000 416.4000 186.0000 ;
	    RECT 417.2000 182.2000 418.0000 186.2000 ;
	    RECT 418.8000 182.2000 419.6000 186.8000 ;
	    RECT 422.0000 182.2000 422.8000 189.6000 ;
	    RECT 423.6000 188.8000 424.4000 190.4000 ;
	    RECT 425.2000 187.4000 425.8000 190.4000 ;
	    RECT 427.0000 189.6000 427.6000 191.8000 ;
	    RECT 423.6000 186.8000 425.8000 187.4000 ;
	    RECT 423.6000 182.2000 424.4000 186.8000 ;
	    RECT 426.8000 182.2000 427.6000 189.6000 ;
	    RECT 433.2000 192.4000 433.8000 195.0000 ;
	    RECT 433.2000 191.6000 434.0000 192.4000 ;
	    RECT 433.2000 188.4000 433.8000 191.6000 ;
	    RECT 432.2000 188.2000 433.8000 188.4000 ;
	    RECT 432.0000 187.8000 433.8000 188.2000 ;
	    RECT 432.0000 182.2000 432.8000 187.8000 ;
	    RECT 436.4000 186.2000 437.2000 199.8000 ;
	    RECT 439.6000 191.6000 440.4000 194.4000 ;
	    RECT 438.0000 190.3000 438.8000 190.4000 ;
	    RECT 441.2000 190.3000 442.0000 199.8000 ;
	    RECT 438.0000 189.7000 442.0000 190.3000 ;
	    RECT 438.0000 189.6000 438.8000 189.7000 ;
	    RECT 441.2000 186.2000 442.0000 189.7000 ;
	    RECT 442.8000 186.8000 443.6000 188.4000 ;
	    RECT 435.4000 185.6000 437.2000 186.2000 ;
	    RECT 440.2000 185.6000 442.0000 186.2000 ;
	    RECT 435.4000 184.4000 436.2000 185.6000 ;
	    RECT 434.8000 183.6000 436.2000 184.4000 ;
	    RECT 435.4000 182.2000 436.2000 183.6000 ;
	    RECT 440.2000 182.2000 441.0000 185.6000 ;
	    RECT 444.4000 182.2000 445.2000 199.8000 ;
	    RECT 447.6000 192.4000 448.4000 199.8000 ;
	    RECT 447.6000 191.8000 449.8000 192.4000 ;
	    RECT 450.8000 191.8000 451.6000 199.8000 ;
	    RECT 449.2000 191.2000 449.8000 191.8000 ;
	    RECT 449.2000 190.4000 450.4000 191.2000 ;
	    RECT 447.6000 188.8000 448.4000 190.4000 ;
	    RECT 449.2000 187.4000 449.8000 190.4000 ;
	    RECT 451.0000 189.6000 451.6000 191.8000 ;
	    RECT 447.6000 186.8000 449.8000 187.4000 ;
	    RECT 447.6000 182.2000 448.4000 186.8000 ;
	    RECT 450.8000 182.2000 451.6000 189.6000 ;
	    RECT 452.4000 182.2000 453.2000 199.8000 ;
	    RECT 455.6000 195.8000 456.4000 199.8000 ;
	    RECT 455.8000 195.6000 456.4000 195.8000 ;
	    RECT 458.8000 195.6000 459.6000 199.8000 ;
	    RECT 462.0000 195.8000 462.8000 199.8000 ;
	    RECT 462.2000 195.6000 462.8000 195.8000 ;
	    RECT 465.2000 195.8000 466.0000 199.8000 ;
	    RECT 468.4000 195.8000 469.2000 199.8000 ;
	    RECT 465.2000 195.6000 465.8000 195.8000 ;
	    RECT 455.8000 195.0000 459.4000 195.6000 ;
	    RECT 462.2000 195.0000 465.8000 195.6000 ;
	    RECT 468.6000 195.6000 469.2000 195.8000 ;
	    RECT 471.6000 195.8000 472.4000 199.8000 ;
	    RECT 471.6000 195.6000 472.2000 195.8000 ;
	    RECT 468.6000 195.0000 472.2000 195.6000 ;
	    RECT 455.8000 192.4000 456.4000 195.0000 ;
	    RECT 457.2000 192.8000 458.0000 194.4000 ;
	    RECT 462.2000 192.4000 462.8000 195.0000 ;
	    RECT 463.6000 192.8000 464.4000 194.4000 ;
	    RECT 468.6000 192.4000 469.2000 195.0000 ;
	    RECT 470.0000 192.8000 470.8000 194.4000 ;
	    RECT 455.6000 191.6000 456.4000 192.4000 ;
	    RECT 462.0000 191.6000 462.8000 192.4000 ;
	    RECT 468.4000 191.6000 469.2000 192.4000 ;
	    RECT 455.8000 188.4000 456.4000 191.6000 ;
	    RECT 458.0000 189.6000 459.6000 190.4000 ;
	    RECT 462.2000 188.4000 462.8000 191.6000 ;
	    RECT 464.4000 189.6000 466.0000 190.4000 ;
	    RECT 468.6000 188.4000 469.2000 191.6000 ;
	    RECT 470.8000 189.6000 472.4000 190.4000 ;
	    RECT 455.8000 188.2000 457.4000 188.4000 ;
	    RECT 462.2000 188.2000 463.8000 188.4000 ;
	    RECT 468.6000 188.2000 470.2000 188.4000 ;
	    RECT 476.4000 188.3000 477.2000 199.8000 ;
	    RECT 480.6000 192.4000 481.4000 199.8000 ;
	    RECT 482.0000 193.6000 482.8000 194.4000 ;
	    RECT 482.2000 192.4000 482.8000 193.6000 ;
	    RECT 480.6000 191.8000 481.6000 192.4000 ;
	    RECT 482.2000 191.8000 483.6000 192.4000 ;
	    RECT 479.6000 188.8000 480.4000 190.4000 ;
	    RECT 481.0000 190.3000 481.6000 191.8000 ;
	    RECT 482.8000 191.6000 483.6000 191.8000 ;
	    RECT 484.4000 191.2000 485.2000 199.8000 ;
	    RECT 488.6000 195.8000 489.8000 199.8000 ;
	    RECT 493.2000 195.8000 494.0000 199.8000 ;
	    RECT 497.6000 196.4000 498.4000 199.8000 ;
	    RECT 497.6000 195.8000 499.6000 196.4000 ;
	    RECT 489.2000 195.0000 490.0000 195.8000 ;
	    RECT 493.4000 195.2000 494.0000 195.8000 ;
	    RECT 492.6000 194.6000 496.2000 195.2000 ;
	    RECT 498.8000 195.0000 499.6000 195.8000 ;
	    RECT 492.6000 194.4000 493.4000 194.6000 ;
	    RECT 495.4000 194.4000 496.2000 194.6000 ;
	    RECT 488.4000 193.2000 489.8000 194.0000 ;
	    RECT 489.2000 192.2000 489.8000 193.2000 ;
	    RECT 491.4000 193.0000 493.6000 193.6000 ;
	    RECT 491.4000 192.8000 492.2000 193.0000 ;
	    RECT 489.2000 191.6000 491.6000 192.2000 ;
	    RECT 484.4000 190.6000 488.6000 191.2000 ;
	    RECT 482.8000 190.3000 483.6000 190.4000 ;
	    RECT 481.0000 189.7000 483.6000 190.3000 ;
	    RECT 481.0000 188.4000 481.6000 189.7000 ;
	    RECT 482.8000 189.6000 483.6000 189.7000 ;
	    RECT 478.0000 188.3000 478.8000 188.4000 ;
	    RECT 476.4000 188.2000 478.8000 188.3000 ;
	    RECT 455.8000 187.8000 457.6000 188.2000 ;
	    RECT 462.2000 187.8000 464.0000 188.2000 ;
	    RECT 468.6000 187.8000 470.4000 188.2000 ;
	    RECT 456.8000 182.2000 457.6000 187.8000 ;
	    RECT 463.2000 182.2000 464.0000 187.8000 ;
	    RECT 469.6000 182.2000 470.4000 187.8000 ;
	    RECT 476.4000 187.7000 479.6000 188.2000 ;
	    RECT 474.8000 184.8000 475.6000 186.4000 ;
	    RECT 476.4000 182.2000 477.2000 187.7000 ;
	    RECT 478.0000 187.6000 479.6000 187.7000 ;
	    RECT 481.0000 187.6000 483.6000 188.4000 ;
	    RECT 478.8000 187.2000 479.6000 187.6000 ;
	    RECT 478.2000 186.2000 481.8000 186.6000 ;
	    RECT 482.8000 186.2000 483.4000 187.6000 ;
	    RECT 484.4000 187.2000 485.2000 190.6000 ;
	    RECT 487.8000 190.4000 488.6000 190.6000 ;
	    RECT 486.2000 189.8000 487.0000 190.0000 ;
	    RECT 486.2000 189.2000 490.0000 189.8000 ;
	    RECT 489.2000 189.0000 490.0000 189.2000 ;
	    RECT 491.0000 188.4000 491.6000 191.6000 ;
	    RECT 493.0000 191.8000 493.6000 193.0000 ;
	    RECT 494.2000 193.0000 495.0000 193.2000 ;
	    RECT 498.8000 193.0000 499.6000 193.2000 ;
	    RECT 494.2000 192.4000 499.6000 193.0000 ;
	    RECT 493.0000 191.4000 497.8000 191.8000 ;
	    RECT 502.0000 191.4000 502.8000 199.8000 ;
	    RECT 503.6000 195.8000 504.4000 199.8000 ;
	    RECT 503.8000 195.6000 504.4000 195.8000 ;
	    RECT 506.8000 195.8000 507.6000 199.8000 ;
	    RECT 506.8000 195.6000 507.4000 195.8000 ;
	    RECT 503.8000 195.0000 507.4000 195.6000 ;
	    RECT 503.8000 192.4000 504.4000 195.0000 ;
	    RECT 505.2000 192.8000 506.0000 194.4000 ;
	    RECT 503.6000 191.6000 504.4000 192.4000 ;
	    RECT 493.0000 191.2000 502.8000 191.4000 ;
	    RECT 497.0000 191.0000 502.8000 191.2000 ;
	    RECT 497.2000 190.8000 502.8000 191.0000 ;
	    RECT 492.4000 190.3000 493.2000 190.4000 ;
	    RECT 495.6000 190.3000 496.4000 190.4000 ;
	    RECT 492.4000 190.2000 496.4000 190.3000 ;
	    RECT 492.4000 189.7000 500.6000 190.2000 ;
	    RECT 492.4000 189.6000 493.2000 189.7000 ;
	    RECT 495.6000 189.6000 500.6000 189.7000 ;
	    RECT 499.8000 189.4000 500.6000 189.6000 ;
	    RECT 498.2000 188.4000 499.0000 188.6000 ;
	    RECT 503.8000 188.4000 504.4000 191.6000 ;
	    RECT 510.0000 191.8000 510.8000 199.8000 ;
	    RECT 513.2000 192.4000 514.0000 199.8000 ;
	    RECT 511.8000 191.8000 514.0000 192.4000 ;
	    RECT 506.0000 189.6000 507.6000 190.4000 ;
	    RECT 510.0000 189.6000 510.6000 191.8000 ;
	    RECT 511.8000 191.2000 512.4000 191.8000 ;
	    RECT 511.2000 190.4000 512.4000 191.2000 ;
	    RECT 491.0000 187.8000 502.0000 188.4000 ;
	    RECT 503.8000 188.2000 505.4000 188.4000 ;
	    RECT 503.8000 187.8000 505.6000 188.2000 ;
	    RECT 491.4000 187.6000 492.2000 187.8000 ;
	    RECT 484.4000 186.6000 488.2000 187.2000 ;
	    RECT 478.0000 186.0000 482.0000 186.2000 ;
	    RECT 478.0000 182.2000 478.8000 186.0000 ;
	    RECT 481.2000 182.2000 482.0000 186.0000 ;
	    RECT 482.8000 182.2000 483.6000 186.2000 ;
	    RECT 484.4000 182.2000 485.2000 186.6000 ;
	    RECT 487.4000 186.4000 488.2000 186.6000 ;
	    RECT 497.2000 186.4000 497.8000 187.8000 ;
	    RECT 500.4000 187.6000 502.0000 187.8000 ;
	    RECT 495.4000 185.4000 496.2000 185.6000 ;
	    RECT 489.2000 184.2000 490.0000 185.0000 ;
	    RECT 493.4000 184.8000 496.2000 185.4000 ;
	    RECT 497.2000 184.8000 498.0000 186.4000 ;
	    RECT 493.4000 184.2000 494.0000 184.8000 ;
	    RECT 498.8000 184.2000 499.6000 185.0000 ;
	    RECT 488.6000 183.6000 490.0000 184.2000 ;
	    RECT 488.6000 182.2000 489.8000 183.6000 ;
	    RECT 493.2000 182.2000 494.0000 184.2000 ;
	    RECT 497.6000 183.6000 499.6000 184.2000 ;
	    RECT 497.6000 182.2000 498.4000 183.6000 ;
	    RECT 502.0000 182.2000 502.8000 187.0000 ;
	    RECT 504.8000 184.3000 505.6000 187.8000 ;
	    RECT 506.8000 184.3000 507.6000 184.4000 ;
	    RECT 504.8000 183.7000 507.6000 184.3000 ;
	    RECT 504.8000 182.2000 505.6000 183.7000 ;
	    RECT 506.8000 183.6000 507.6000 183.7000 ;
	    RECT 510.0000 182.2000 510.8000 189.6000 ;
	    RECT 511.8000 187.4000 512.4000 190.4000 ;
	    RECT 513.2000 188.8000 514.0000 190.4000 ;
	    RECT 511.8000 186.8000 514.0000 187.4000 ;
	    RECT 513.2000 182.2000 514.0000 186.8000 ;
	    RECT 2.8000 175.2000 3.6000 179.8000 ;
	    RECT 6.0000 175.2000 6.8000 179.8000 ;
	    RECT 9.8000 176.4000 10.6000 179.8000 ;
	    RECT 9.8000 175.8000 11.6000 176.4000 ;
	    RECT 14.0000 175.8000 14.8000 179.8000 ;
	    RECT 18.2000 176.8000 19.0000 179.8000 ;
	    RECT 22.0000 177.6000 22.8000 179.8000 ;
	    RECT 27.8000 178.4000 28.6000 179.8000 ;
	    RECT 27.8000 177.6000 29.2000 178.4000 ;
	    RECT 18.2000 175.8000 19.6000 176.8000 ;
	    RECT 2.8000 174.4000 6.8000 175.2000 ;
	    RECT 2.8000 171.6000 3.6000 174.4000 ;
	    RECT 10.8000 172.3000 11.6000 175.8000 ;
	    RECT 14.2000 175.6000 14.8000 175.8000 ;
	    RECT 14.2000 175.2000 16.0000 175.6000 ;
	    RECT 12.4000 174.3000 13.2000 175.2000 ;
	    RECT 14.2000 175.0000 18.4000 175.2000 ;
	    RECT 15.4000 174.6000 18.4000 175.0000 ;
	    RECT 17.6000 174.4000 18.4000 174.6000 ;
	    RECT 14.0000 174.3000 14.8000 174.4000 ;
	    RECT 12.4000 173.7000 14.8000 174.3000 ;
	    RECT 12.4000 173.6000 13.2000 173.7000 ;
	    RECT 14.0000 172.8000 14.8000 173.7000 ;
	    RECT 12.4000 172.3000 13.2000 172.4000 ;
	    RECT 10.8000 171.7000 13.2000 172.3000 ;
	    RECT 2.8000 170.8000 6.8000 171.6000 ;
	    RECT 2.8000 162.2000 3.6000 170.8000 ;
	    RECT 6.0000 162.2000 6.8000 170.8000 ;
	    RECT 10.8000 162.2000 11.6000 171.7000 ;
	    RECT 12.4000 171.6000 13.2000 171.7000 ;
	    RECT 17.6000 171.0000 18.2000 174.4000 ;
	    RECT 19.0000 172.4000 19.6000 175.8000 ;
	    RECT 22.0000 174.4000 22.6000 177.6000 ;
	    RECT 27.8000 176.4000 28.6000 177.6000 ;
	    RECT 26.8000 175.8000 28.6000 176.4000 ;
	    RECT 30.0000 175.8000 30.8000 179.8000 ;
	    RECT 31.6000 176.0000 32.4000 179.8000 ;
	    RECT 34.8000 176.0000 35.6000 179.8000 ;
	    RECT 31.6000 175.8000 35.6000 176.0000 ;
	    RECT 22.0000 173.6000 22.8000 174.4000 ;
	    RECT 18.8000 171.6000 19.6000 172.4000 ;
	    RECT 15.8000 170.4000 18.2000 171.0000 ;
	    RECT 15.8000 166.2000 16.4000 170.4000 ;
	    RECT 19.0000 170.2000 19.6000 171.6000 ;
	    RECT 20.4000 170.8000 21.2000 172.4000 ;
	    RECT 22.0000 170.2000 22.6000 173.6000 ;
	    RECT 15.6000 162.2000 16.4000 166.2000 ;
	    RECT 18.8000 162.2000 19.6000 170.2000 ;
	    RECT 21.0000 169.4000 22.8000 170.2000 ;
	    RECT 21.0000 162.2000 21.8000 169.4000 ;
	    RECT 26.8000 162.2000 27.6000 175.8000 ;
	    RECT 30.2000 174.4000 30.8000 175.8000 ;
	    RECT 31.8000 175.4000 35.4000 175.8000 ;
	    RECT 36.4000 175.0000 37.2000 179.8000 ;
	    RECT 40.8000 178.4000 41.6000 179.8000 ;
	    RECT 39.6000 177.8000 41.6000 178.4000 ;
	    RECT 45.2000 177.8000 46.0000 179.8000 ;
	    RECT 49.4000 178.4000 50.6000 179.8000 ;
	    RECT 49.2000 177.8000 50.6000 178.4000 ;
	    RECT 39.6000 177.0000 40.4000 177.8000 ;
	    RECT 45.2000 177.2000 45.8000 177.8000 ;
	    RECT 41.2000 176.4000 42.0000 177.2000 ;
	    RECT 43.0000 176.6000 45.8000 177.2000 ;
	    RECT 49.2000 177.0000 50.0000 177.8000 ;
	    RECT 43.0000 176.4000 43.8000 176.6000 ;
	    RECT 34.0000 174.4000 34.8000 174.8000 ;
	    RECT 30.0000 173.6000 32.6000 174.4000 ;
	    RECT 34.0000 173.8000 35.6000 174.4000 ;
	    RECT 34.8000 173.6000 35.6000 173.8000 ;
	    RECT 37.2000 174.2000 38.8000 174.4000 ;
	    RECT 41.4000 174.2000 42.0000 176.4000 ;
	    RECT 51.0000 175.4000 51.8000 175.6000 ;
	    RECT 54.0000 175.4000 54.8000 179.8000 ;
	    RECT 51.0000 174.8000 54.8000 175.4000 ;
	    RECT 47.0000 174.2000 47.8000 174.4000 ;
	    RECT 37.2000 173.6000 48.2000 174.2000 ;
	    RECT 32.0000 172.4000 32.6000 173.6000 ;
	    RECT 40.2000 173.4000 41.0000 173.6000 ;
	    RECT 31.6000 171.6000 32.6000 172.4000 ;
	    RECT 33.2000 171.6000 34.0000 173.2000 ;
	    RECT 38.6000 172.4000 39.4000 172.6000 ;
	    RECT 38.6000 171.8000 43.6000 172.4000 ;
	    RECT 42.8000 171.6000 43.6000 171.8000 ;
	    RECT 28.4000 168.8000 29.2000 170.4000 ;
	    RECT 30.0000 170.2000 30.8000 170.4000 ;
	    RECT 32.0000 170.2000 32.6000 171.6000 ;
	    RECT 36.4000 171.0000 42.0000 171.2000 ;
	    RECT 36.4000 170.8000 42.2000 171.0000 ;
	    RECT 36.4000 170.6000 46.2000 170.8000 ;
	    RECT 30.0000 169.6000 31.4000 170.2000 ;
	    RECT 32.0000 169.6000 33.0000 170.2000 ;
	    RECT 30.8000 168.4000 31.4000 169.6000 ;
	    RECT 30.8000 167.6000 31.6000 168.4000 ;
	    RECT 32.2000 162.2000 33.0000 169.6000 ;
	    RECT 36.4000 162.2000 37.2000 170.6000 ;
	    RECT 41.4000 170.2000 46.2000 170.6000 ;
	    RECT 39.6000 169.0000 45.0000 169.6000 ;
	    RECT 39.6000 168.8000 40.4000 169.0000 ;
	    RECT 44.2000 168.8000 45.0000 169.0000 ;
	    RECT 45.6000 169.0000 46.2000 170.2000 ;
	    RECT 47.6000 170.4000 48.2000 173.6000 ;
	    RECT 49.2000 172.8000 50.0000 173.0000 ;
	    RECT 49.2000 172.2000 53.0000 172.8000 ;
	    RECT 52.2000 172.0000 53.0000 172.2000 ;
	    RECT 50.6000 171.4000 51.4000 171.6000 ;
	    RECT 54.0000 171.4000 54.8000 174.8000 ;
	    RECT 50.6000 170.8000 54.8000 171.4000 ;
	    RECT 47.6000 169.8000 50.0000 170.4000 ;
	    RECT 47.0000 169.0000 47.8000 169.2000 ;
	    RECT 45.6000 168.4000 47.8000 169.0000 ;
	    RECT 49.4000 168.8000 50.0000 169.8000 ;
	    RECT 49.4000 168.0000 50.8000 168.8000 ;
	    RECT 43.0000 167.4000 43.8000 167.6000 ;
	    RECT 45.8000 167.4000 46.6000 167.6000 ;
	    RECT 39.6000 166.2000 40.4000 167.0000 ;
	    RECT 43.0000 166.8000 46.6000 167.4000 ;
	    RECT 45.2000 166.2000 45.8000 166.8000 ;
	    RECT 49.2000 166.2000 50.0000 167.0000 ;
	    RECT 39.6000 165.6000 41.6000 166.2000 ;
	    RECT 40.8000 162.2000 41.6000 165.6000 ;
	    RECT 45.2000 162.2000 46.0000 166.2000 ;
	    RECT 49.4000 162.2000 50.6000 166.2000 ;
	    RECT 54.0000 162.2000 54.8000 170.8000 ;
	    RECT 55.6000 175.4000 56.4000 179.8000 ;
	    RECT 59.8000 178.4000 61.0000 179.8000 ;
	    RECT 59.8000 177.8000 61.2000 178.4000 ;
	    RECT 64.4000 177.8000 65.2000 179.8000 ;
	    RECT 68.8000 178.4000 69.6000 179.8000 ;
	    RECT 68.8000 177.8000 70.8000 178.4000 ;
	    RECT 60.4000 177.0000 61.2000 177.8000 ;
	    RECT 64.6000 177.2000 65.2000 177.8000 ;
	    RECT 64.6000 176.6000 67.4000 177.2000 ;
	    RECT 66.6000 176.4000 67.4000 176.6000 ;
	    RECT 68.4000 176.4000 69.2000 177.2000 ;
	    RECT 70.0000 177.0000 70.8000 177.8000 ;
	    RECT 58.6000 175.4000 59.4000 175.6000 ;
	    RECT 55.6000 174.8000 59.4000 175.4000 ;
	    RECT 55.6000 171.4000 56.4000 174.8000 ;
	    RECT 62.6000 174.2000 63.4000 174.4000 ;
	    RECT 68.4000 174.2000 69.0000 176.4000 ;
	    RECT 73.2000 175.0000 74.0000 179.8000 ;
	    RECT 77.4000 176.4000 78.2000 179.8000 ;
	    RECT 76.4000 175.8000 78.2000 176.4000 ;
	    RECT 79.6000 175.8000 80.4000 179.8000 ;
	    RECT 81.2000 176.0000 82.0000 179.8000 ;
	    RECT 84.4000 176.0000 85.2000 179.8000 ;
	    RECT 81.2000 175.8000 85.2000 176.0000 ;
	    RECT 71.6000 174.2000 73.2000 174.4000 ;
	    RECT 62.2000 173.6000 73.2000 174.2000 ;
	    RECT 74.8000 173.6000 75.6000 175.2000 ;
	    RECT 60.4000 172.8000 61.2000 173.0000 ;
	    RECT 57.4000 172.2000 61.2000 172.8000 ;
	    RECT 57.4000 172.0000 58.2000 172.2000 ;
	    RECT 59.0000 171.4000 59.8000 171.6000 ;
	    RECT 55.6000 170.8000 59.8000 171.4000 ;
	    RECT 55.6000 162.2000 56.4000 170.8000 ;
	    RECT 62.2000 170.4000 62.8000 173.6000 ;
	    RECT 69.4000 173.4000 70.2000 173.6000 ;
	    RECT 71.0000 172.4000 71.8000 172.6000 ;
	    RECT 66.8000 171.8000 71.8000 172.4000 ;
	    RECT 76.4000 172.3000 77.2000 175.8000 ;
	    RECT 79.8000 174.4000 80.4000 175.8000 ;
	    RECT 81.4000 175.4000 85.0000 175.8000 ;
	    RECT 86.0000 175.0000 86.8000 179.8000 ;
	    RECT 90.4000 178.4000 91.2000 179.8000 ;
	    RECT 89.2000 177.8000 91.2000 178.4000 ;
	    RECT 94.8000 177.8000 95.6000 179.8000 ;
	    RECT 99.0000 178.4000 100.2000 179.8000 ;
	    RECT 98.8000 177.8000 100.2000 178.4000 ;
	    RECT 89.2000 177.0000 90.0000 177.8000 ;
	    RECT 94.8000 177.2000 95.4000 177.8000 ;
	    RECT 90.8000 176.4000 91.6000 177.2000 ;
	    RECT 92.6000 176.6000 95.4000 177.2000 ;
	    RECT 98.8000 177.0000 99.6000 177.8000 ;
	    RECT 92.6000 176.4000 93.4000 176.6000 ;
	    RECT 83.6000 174.4000 84.4000 174.8000 ;
	    RECT 79.6000 173.6000 82.2000 174.4000 ;
	    RECT 83.6000 173.8000 85.2000 174.4000 ;
	    RECT 84.4000 173.6000 85.2000 173.8000 ;
	    RECT 86.8000 174.2000 88.4000 174.4000 ;
	    RECT 91.0000 174.2000 91.6000 176.4000 ;
	    RECT 100.6000 175.4000 101.4000 175.6000 ;
	    RECT 103.6000 175.4000 104.4000 179.8000 ;
	    RECT 111.6000 176.0000 112.4000 179.8000 ;
	    RECT 114.8000 176.0000 115.6000 179.8000 ;
	    RECT 111.6000 175.8000 115.6000 176.0000 ;
	    RECT 116.4000 175.8000 117.2000 179.8000 ;
	    RECT 118.6000 176.4000 119.4000 179.8000 ;
	    RECT 118.6000 175.8000 120.4000 176.4000 ;
	    RECT 111.8000 175.4000 115.4000 175.8000 ;
	    RECT 100.6000 174.8000 104.4000 175.4000 ;
	    RECT 96.6000 174.2000 97.4000 174.4000 ;
	    RECT 86.8000 173.6000 97.8000 174.2000 ;
	    RECT 66.8000 171.6000 67.6000 171.8000 ;
	    RECT 76.4000 171.7000 80.3000 172.3000 ;
	    RECT 68.4000 171.0000 74.0000 171.2000 ;
	    RECT 68.2000 170.8000 74.0000 171.0000 ;
	    RECT 60.4000 169.8000 62.8000 170.4000 ;
	    RECT 64.2000 170.6000 74.0000 170.8000 ;
	    RECT 64.2000 170.2000 69.0000 170.6000 ;
	    RECT 60.4000 168.8000 61.0000 169.8000 ;
	    RECT 59.6000 168.0000 61.0000 168.8000 ;
	    RECT 62.6000 169.0000 63.4000 169.2000 ;
	    RECT 64.2000 169.0000 64.8000 170.2000 ;
	    RECT 62.6000 168.4000 64.8000 169.0000 ;
	    RECT 65.4000 169.0000 70.8000 169.6000 ;
	    RECT 65.4000 168.8000 66.2000 169.0000 ;
	    RECT 70.0000 168.8000 70.8000 169.0000 ;
	    RECT 63.8000 167.4000 64.6000 167.6000 ;
	    RECT 66.6000 167.4000 67.4000 167.6000 ;
	    RECT 60.4000 166.2000 61.2000 167.0000 ;
	    RECT 63.8000 166.8000 67.4000 167.4000 ;
	    RECT 64.6000 166.2000 65.2000 166.8000 ;
	    RECT 70.0000 166.2000 70.8000 167.0000 ;
	    RECT 59.8000 162.2000 61.0000 166.2000 ;
	    RECT 64.4000 162.2000 65.2000 166.2000 ;
	    RECT 68.8000 165.6000 70.8000 166.2000 ;
	    RECT 68.8000 162.2000 69.6000 165.6000 ;
	    RECT 73.2000 162.2000 74.0000 170.6000 ;
	    RECT 76.4000 162.2000 77.2000 171.7000 ;
	    RECT 79.7000 170.4000 80.3000 171.7000 ;
	    RECT 78.0000 168.8000 78.8000 170.4000 ;
	    RECT 79.6000 170.2000 80.4000 170.4000 ;
	    RECT 81.6000 170.2000 82.2000 173.6000 ;
	    RECT 89.8000 173.4000 90.6000 173.6000 ;
	    RECT 82.8000 171.6000 83.6000 173.2000 ;
	    RECT 88.2000 172.4000 89.0000 172.6000 ;
	    RECT 88.2000 172.3000 93.2000 172.4000 ;
	    RECT 94.0000 172.3000 94.8000 172.4000 ;
	    RECT 88.2000 171.8000 94.8000 172.3000 ;
	    RECT 92.4000 171.7000 94.8000 171.8000 ;
	    RECT 92.4000 171.6000 93.2000 171.7000 ;
	    RECT 94.0000 171.6000 94.8000 171.7000 ;
	    RECT 86.0000 171.0000 91.6000 171.2000 ;
	    RECT 86.0000 170.8000 91.8000 171.0000 ;
	    RECT 86.0000 170.6000 95.8000 170.8000 ;
	    RECT 79.6000 169.6000 81.0000 170.2000 ;
	    RECT 81.6000 169.6000 82.6000 170.2000 ;
	    RECT 80.4000 168.4000 81.0000 169.6000 ;
	    RECT 80.4000 167.6000 81.2000 168.4000 ;
	    RECT 81.8000 162.2000 82.6000 169.6000 ;
	    RECT 86.0000 162.2000 86.8000 170.6000 ;
	    RECT 91.0000 170.2000 95.8000 170.6000 ;
	    RECT 89.2000 169.0000 94.6000 169.6000 ;
	    RECT 89.2000 168.8000 90.0000 169.0000 ;
	    RECT 93.8000 168.8000 94.6000 169.0000 ;
	    RECT 95.2000 169.0000 95.8000 170.2000 ;
	    RECT 97.2000 170.4000 97.8000 173.6000 ;
	    RECT 98.8000 172.8000 99.6000 173.0000 ;
	    RECT 98.8000 172.2000 102.6000 172.8000 ;
	    RECT 101.8000 172.0000 102.6000 172.2000 ;
	    RECT 100.2000 171.4000 101.0000 171.6000 ;
	    RECT 103.6000 171.4000 104.4000 174.8000 ;
	    RECT 112.4000 174.4000 113.2000 174.8000 ;
	    RECT 116.4000 174.4000 117.0000 175.8000 ;
	    RECT 111.6000 173.8000 113.2000 174.4000 ;
	    RECT 111.6000 173.6000 112.4000 173.8000 ;
	    RECT 114.6000 173.6000 117.2000 174.4000 ;
	    RECT 111.7000 172.4000 112.3000 173.6000 ;
	    RECT 111.6000 171.6000 112.4000 172.4000 ;
	    RECT 113.2000 171.6000 114.0000 173.2000 ;
	    RECT 114.6000 172.4000 115.2000 173.6000 ;
	    RECT 114.6000 171.6000 115.6000 172.4000 ;
	    RECT 119.6000 172.3000 120.4000 175.8000 ;
	    RECT 122.8000 175.4000 123.6000 179.8000 ;
	    RECT 127.0000 178.4000 128.2000 179.8000 ;
	    RECT 127.0000 177.8000 128.4000 178.4000 ;
	    RECT 131.6000 177.8000 132.4000 179.8000 ;
	    RECT 136.0000 178.4000 136.8000 179.8000 ;
	    RECT 136.0000 177.8000 138.0000 178.4000 ;
	    RECT 127.6000 177.0000 128.4000 177.8000 ;
	    RECT 131.8000 177.2000 132.4000 177.8000 ;
	    RECT 131.8000 176.6000 134.6000 177.2000 ;
	    RECT 133.8000 176.4000 134.6000 176.6000 ;
	    RECT 135.6000 176.4000 136.4000 177.2000 ;
	    RECT 137.2000 177.0000 138.0000 177.8000 ;
	    RECT 125.8000 175.4000 126.6000 175.6000 ;
	    RECT 121.2000 173.6000 122.0000 175.2000 ;
	    RECT 122.8000 174.8000 126.6000 175.4000 ;
	    RECT 116.5000 171.7000 120.4000 172.3000 ;
	    RECT 100.2000 170.8000 104.4000 171.4000 ;
	    RECT 97.2000 169.8000 99.6000 170.4000 ;
	    RECT 96.6000 169.0000 97.4000 169.2000 ;
	    RECT 95.2000 168.4000 97.4000 169.0000 ;
	    RECT 99.0000 168.8000 99.6000 169.8000 ;
	    RECT 99.0000 168.0000 100.4000 168.8000 ;
	    RECT 92.6000 167.4000 93.4000 167.6000 ;
	    RECT 95.4000 167.4000 96.2000 167.6000 ;
	    RECT 89.2000 166.2000 90.0000 167.0000 ;
	    RECT 92.6000 166.8000 96.2000 167.4000 ;
	    RECT 94.8000 166.2000 95.4000 166.8000 ;
	    RECT 98.8000 166.2000 99.6000 167.0000 ;
	    RECT 89.2000 165.6000 91.2000 166.2000 ;
	    RECT 90.4000 162.2000 91.2000 165.6000 ;
	    RECT 94.8000 162.2000 95.6000 166.2000 ;
	    RECT 99.0000 162.2000 100.2000 166.2000 ;
	    RECT 103.6000 162.2000 104.4000 170.8000 ;
	    RECT 114.6000 170.2000 115.2000 171.6000 ;
	    RECT 116.5000 170.4000 117.1000 171.7000 ;
	    RECT 116.4000 170.2000 117.2000 170.4000 ;
	    RECT 114.2000 169.6000 115.2000 170.2000 ;
	    RECT 115.8000 169.6000 117.2000 170.2000 ;
	    RECT 114.2000 162.2000 115.0000 169.6000 ;
	    RECT 115.8000 168.4000 116.4000 169.6000 ;
	    RECT 118.0000 168.8000 118.8000 170.4000 ;
	    RECT 115.6000 167.6000 116.4000 168.4000 ;
	    RECT 119.6000 162.2000 120.4000 171.7000 ;
	    RECT 122.8000 171.4000 123.6000 174.8000 ;
	    RECT 129.8000 174.2000 130.6000 174.4000 ;
	    RECT 132.4000 174.2000 133.2000 174.4000 ;
	    RECT 135.6000 174.2000 136.2000 176.4000 ;
	    RECT 140.4000 175.0000 141.2000 179.8000 ;
	    RECT 144.6000 176.4000 145.4000 179.8000 ;
	    RECT 143.6000 175.8000 145.4000 176.4000 ;
	    RECT 146.8000 175.8000 147.6000 179.8000 ;
	    RECT 148.4000 176.0000 149.2000 179.8000 ;
	    RECT 151.6000 176.0000 152.4000 179.8000 ;
	    RECT 148.4000 175.8000 152.4000 176.0000 ;
	    RECT 138.8000 174.2000 140.4000 174.4000 ;
	    RECT 129.4000 173.6000 140.4000 174.2000 ;
	    RECT 142.0000 173.6000 142.8000 175.2000 ;
	    RECT 127.6000 172.8000 128.4000 173.0000 ;
	    RECT 124.6000 172.2000 128.4000 172.8000 ;
	    RECT 124.6000 172.0000 125.4000 172.2000 ;
	    RECT 126.2000 171.4000 127.0000 171.6000 ;
	    RECT 122.8000 170.8000 127.0000 171.4000 ;
	    RECT 122.8000 162.2000 123.6000 170.8000 ;
	    RECT 129.4000 170.4000 130.0000 173.6000 ;
	    RECT 136.6000 173.4000 137.4000 173.6000 ;
	    RECT 135.6000 172.4000 136.4000 172.6000 ;
	    RECT 138.2000 172.4000 139.0000 172.6000 ;
	    RECT 134.0000 171.8000 139.0000 172.4000 ;
	    RECT 143.6000 172.3000 144.4000 175.8000 ;
	    RECT 147.0000 174.4000 147.6000 175.8000 ;
	    RECT 148.6000 175.4000 152.2000 175.8000 ;
	    RECT 150.8000 174.4000 151.6000 174.8000 ;
	    RECT 146.8000 173.6000 149.4000 174.4000 ;
	    RECT 150.8000 173.8000 152.4000 174.4000 ;
	    RECT 151.6000 173.6000 152.4000 173.8000 ;
	    RECT 134.0000 171.6000 134.8000 171.8000 ;
	    RECT 143.6000 171.7000 147.5000 172.3000 ;
	    RECT 135.6000 171.0000 141.2000 171.2000 ;
	    RECT 135.4000 170.8000 141.2000 171.0000 ;
	    RECT 127.6000 169.8000 130.0000 170.4000 ;
	    RECT 131.4000 170.6000 141.2000 170.8000 ;
	    RECT 131.4000 170.2000 136.2000 170.6000 ;
	    RECT 127.6000 168.8000 128.2000 169.8000 ;
	    RECT 126.8000 168.0000 128.2000 168.8000 ;
	    RECT 129.8000 169.0000 130.6000 169.2000 ;
	    RECT 131.4000 169.0000 132.0000 170.2000 ;
	    RECT 129.8000 168.4000 132.0000 169.0000 ;
	    RECT 132.6000 169.0000 138.0000 169.6000 ;
	    RECT 132.6000 168.8000 133.4000 169.0000 ;
	    RECT 137.2000 168.8000 138.0000 169.0000 ;
	    RECT 131.0000 167.4000 131.8000 167.6000 ;
	    RECT 133.8000 167.4000 134.6000 167.6000 ;
	    RECT 127.6000 166.2000 128.4000 167.0000 ;
	    RECT 131.0000 166.8000 134.6000 167.4000 ;
	    RECT 131.8000 166.2000 132.4000 166.8000 ;
	    RECT 137.2000 166.2000 138.0000 167.0000 ;
	    RECT 127.0000 162.2000 128.2000 166.2000 ;
	    RECT 131.6000 162.2000 132.4000 166.2000 ;
	    RECT 136.0000 165.6000 138.0000 166.2000 ;
	    RECT 136.0000 162.2000 136.8000 165.6000 ;
	    RECT 140.4000 162.2000 141.2000 170.6000 ;
	    RECT 143.6000 162.2000 144.4000 171.7000 ;
	    RECT 146.9000 170.4000 147.5000 171.7000 ;
	    RECT 145.2000 168.8000 146.0000 170.4000 ;
	    RECT 146.8000 170.2000 147.6000 170.4000 ;
	    RECT 148.8000 170.2000 149.4000 173.6000 ;
	    RECT 150.0000 171.6000 150.8000 173.2000 ;
	    RECT 153.2000 172.4000 154.0000 179.8000 ;
	    RECT 156.4000 175.2000 157.2000 179.8000 ;
	    RECT 155.0000 174.6000 157.2000 175.2000 ;
	    RECT 158.0000 175.4000 158.8000 179.8000 ;
	    RECT 162.2000 178.4000 163.4000 179.8000 ;
	    RECT 162.2000 177.8000 163.6000 178.4000 ;
	    RECT 166.8000 177.8000 167.6000 179.8000 ;
	    RECT 171.2000 178.4000 172.0000 179.8000 ;
	    RECT 171.2000 177.8000 173.2000 178.4000 ;
	    RECT 162.8000 177.0000 163.6000 177.8000 ;
	    RECT 167.0000 177.2000 167.6000 177.8000 ;
	    RECT 167.0000 176.6000 169.8000 177.2000 ;
	    RECT 169.0000 176.4000 169.8000 176.6000 ;
	    RECT 170.8000 176.4000 171.6000 177.2000 ;
	    RECT 172.4000 177.0000 173.2000 177.8000 ;
	    RECT 161.0000 175.4000 161.8000 175.6000 ;
	    RECT 158.0000 174.8000 161.8000 175.4000 ;
	    RECT 153.2000 170.2000 153.8000 172.4000 ;
	    RECT 155.0000 171.6000 155.6000 174.6000 ;
	    RECT 156.4000 171.6000 157.2000 173.2000 ;
	    RECT 154.4000 170.8000 155.6000 171.6000 ;
	    RECT 155.0000 170.2000 155.6000 170.8000 ;
	    RECT 158.0000 171.4000 158.8000 174.8000 ;
	    RECT 165.0000 174.2000 165.8000 174.4000 ;
	    RECT 170.8000 174.2000 171.4000 176.4000 ;
	    RECT 175.6000 175.0000 176.4000 179.8000 ;
	    RECT 174.0000 174.2000 175.6000 174.4000 ;
	    RECT 164.6000 173.6000 175.6000 174.2000 ;
	    RECT 162.8000 172.8000 163.6000 173.0000 ;
	    RECT 159.8000 172.2000 163.6000 172.8000 ;
	    RECT 164.6000 172.4000 165.2000 173.6000 ;
	    RECT 171.8000 173.4000 172.6000 173.6000 ;
	    RECT 170.8000 172.4000 171.6000 172.6000 ;
	    RECT 173.4000 172.4000 174.2000 172.6000 ;
	    RECT 159.8000 172.0000 160.6000 172.2000 ;
	    RECT 164.4000 171.6000 165.2000 172.4000 ;
	    RECT 169.2000 171.8000 174.2000 172.4000 ;
	    RECT 177.2000 172.4000 178.0000 179.8000 ;
	    RECT 180.4000 175.2000 181.2000 179.8000 ;
	    RECT 185.8000 176.0000 186.6000 179.0000 ;
	    RECT 190.0000 177.0000 190.8000 179.0000 ;
	    RECT 179.0000 174.6000 181.2000 175.2000 ;
	    RECT 185.0000 175.4000 186.6000 176.0000 ;
	    RECT 185.0000 175.0000 185.8000 175.4000 ;
	    RECT 169.2000 171.6000 170.0000 171.8000 ;
	    RECT 161.4000 171.4000 162.2000 171.6000 ;
	    RECT 158.0000 170.8000 162.2000 171.4000 ;
	    RECT 146.8000 169.6000 148.2000 170.2000 ;
	    RECT 148.8000 169.6000 149.8000 170.2000 ;
	    RECT 147.6000 168.4000 148.2000 169.6000 ;
	    RECT 147.6000 167.6000 148.4000 168.4000 ;
	    RECT 149.0000 162.2000 149.8000 169.6000 ;
	    RECT 153.2000 162.2000 154.0000 170.2000 ;
	    RECT 155.0000 169.6000 157.2000 170.2000 ;
	    RECT 156.4000 162.2000 157.2000 169.6000 ;
	    RECT 158.0000 162.2000 158.8000 170.8000 ;
	    RECT 164.6000 170.4000 165.2000 171.6000 ;
	    RECT 170.8000 171.0000 176.4000 171.2000 ;
	    RECT 170.6000 170.8000 176.4000 171.0000 ;
	    RECT 162.8000 169.8000 165.2000 170.4000 ;
	    RECT 166.6000 170.6000 176.4000 170.8000 ;
	    RECT 166.6000 170.2000 171.4000 170.6000 ;
	    RECT 162.8000 168.8000 163.4000 169.8000 ;
	    RECT 162.0000 168.0000 163.4000 168.8000 ;
	    RECT 165.0000 169.0000 165.8000 169.2000 ;
	    RECT 166.6000 169.0000 167.2000 170.2000 ;
	    RECT 165.0000 168.4000 167.2000 169.0000 ;
	    RECT 167.8000 169.0000 173.2000 169.6000 ;
	    RECT 167.8000 168.8000 168.6000 169.0000 ;
	    RECT 172.4000 168.8000 173.2000 169.0000 ;
	    RECT 166.2000 167.4000 167.0000 167.6000 ;
	    RECT 169.0000 167.4000 169.8000 167.6000 ;
	    RECT 162.8000 166.2000 163.6000 167.0000 ;
	    RECT 166.2000 166.8000 169.8000 167.4000 ;
	    RECT 167.0000 166.2000 167.6000 166.8000 ;
	    RECT 172.4000 166.2000 173.2000 167.0000 ;
	    RECT 162.2000 162.2000 163.4000 166.2000 ;
	    RECT 166.8000 162.2000 167.6000 166.2000 ;
	    RECT 171.2000 165.6000 173.2000 166.2000 ;
	    RECT 171.2000 162.2000 172.0000 165.6000 ;
	    RECT 175.6000 162.2000 176.4000 170.6000 ;
	    RECT 177.2000 170.2000 177.8000 172.4000 ;
	    RECT 179.0000 171.6000 179.6000 174.6000 ;
	    RECT 185.0000 174.4000 185.6000 175.0000 ;
	    RECT 190.2000 174.8000 190.8000 177.0000 ;
	    RECT 195.4000 176.0000 196.2000 179.0000 ;
	    RECT 199.6000 177.0000 200.4000 179.0000 ;
	    RECT 183.6000 173.6000 185.6000 174.4000 ;
	    RECT 186.6000 174.2000 190.8000 174.8000 ;
	    RECT 194.6000 175.4000 196.2000 176.0000 ;
	    RECT 194.6000 175.0000 195.4000 175.4000 ;
	    RECT 194.6000 174.4000 195.2000 175.0000 ;
	    RECT 199.8000 174.8000 200.4000 177.0000 ;
	    RECT 186.6000 173.8000 187.6000 174.2000 ;
	    RECT 180.4000 171.6000 181.2000 173.2000 ;
	    RECT 178.4000 170.8000 179.6000 171.6000 ;
	    RECT 183.6000 170.8000 184.4000 172.4000 ;
	    RECT 179.0000 170.2000 179.6000 170.8000 ;
	    RECT 177.2000 162.2000 178.0000 170.2000 ;
	    RECT 179.0000 169.6000 181.2000 170.2000 ;
	    RECT 180.4000 162.2000 181.2000 169.6000 ;
	    RECT 185.0000 169.8000 185.6000 173.6000 ;
	    RECT 186.2000 173.0000 187.6000 173.8000 ;
	    RECT 193.2000 173.6000 195.2000 174.4000 ;
	    RECT 196.2000 174.2000 200.4000 174.8000 ;
	    RECT 196.2000 173.8000 197.2000 174.2000 ;
	    RECT 187.0000 171.0000 187.6000 173.0000 ;
	    RECT 188.4000 171.6000 189.2000 173.2000 ;
	    RECT 190.0000 171.6000 190.8000 173.2000 ;
	    RECT 187.0000 170.4000 190.8000 171.0000 ;
	    RECT 193.2000 170.8000 194.0000 172.4000 ;
	    RECT 185.0000 169.2000 186.6000 169.8000 ;
	    RECT 185.8000 164.4000 186.6000 169.2000 ;
	    RECT 190.2000 167.0000 190.8000 170.4000 ;
	    RECT 194.6000 169.8000 195.2000 173.6000 ;
	    RECT 195.8000 173.0000 197.2000 173.8000 ;
	    RECT 196.6000 171.0000 197.2000 173.0000 ;
	    RECT 198.0000 171.6000 198.8000 173.2000 ;
	    RECT 199.6000 171.6000 200.4000 173.2000 ;
	    RECT 201.2000 172.4000 202.0000 179.8000 ;
	    RECT 204.4000 175.2000 205.2000 179.8000 ;
	    RECT 207.6000 175.2000 208.4000 179.8000 ;
	    RECT 210.8000 175.2000 211.6000 179.8000 ;
	    RECT 216.6000 176.4000 217.4000 179.8000 ;
	    RECT 215.6000 175.8000 217.4000 176.4000 ;
	    RECT 218.8000 175.8000 219.6000 179.8000 ;
	    RECT 220.4000 176.0000 221.2000 179.8000 ;
	    RECT 223.6000 176.0000 224.4000 179.8000 ;
	    RECT 220.4000 175.8000 224.4000 176.0000 ;
	    RECT 203.0000 174.6000 205.2000 175.2000 ;
	    RECT 196.6000 170.4000 200.4000 171.0000 ;
	    RECT 194.6000 169.2000 196.2000 169.8000 ;
	    RECT 185.2000 163.6000 186.6000 164.4000 ;
	    RECT 185.8000 162.2000 186.6000 163.6000 ;
	    RECT 190.0000 163.0000 190.8000 167.0000 ;
	    RECT 195.4000 164.4000 196.2000 169.2000 ;
	    RECT 199.8000 167.0000 200.4000 170.4000 ;
	    RECT 194.8000 163.6000 196.2000 164.4000 ;
	    RECT 195.4000 162.2000 196.2000 163.6000 ;
	    RECT 199.6000 163.0000 200.4000 167.0000 ;
	    RECT 201.2000 170.2000 201.8000 172.4000 ;
	    RECT 203.0000 171.6000 203.6000 174.6000 ;
	    RECT 206.0000 173.6000 206.8000 175.2000 ;
	    RECT 207.6000 174.4000 211.6000 175.2000 ;
	    RECT 204.4000 171.6000 205.2000 173.2000 ;
	    RECT 210.8000 171.6000 211.6000 174.4000 ;
	    RECT 214.0000 173.6000 214.8000 175.2000 ;
	    RECT 202.4000 170.8000 203.6000 171.6000 ;
	    RECT 203.0000 170.2000 203.6000 170.8000 ;
	    RECT 207.6000 170.8000 211.6000 171.6000 ;
	    RECT 201.2000 162.2000 202.0000 170.2000 ;
	    RECT 203.0000 169.6000 205.2000 170.2000 ;
	    RECT 204.4000 162.2000 205.2000 169.6000 ;
	    RECT 207.6000 162.2000 208.4000 170.8000 ;
	    RECT 210.8000 162.2000 211.6000 170.8000 ;
	    RECT 215.6000 172.3000 216.4000 175.8000 ;
	    RECT 219.0000 174.4000 219.6000 175.8000 ;
	    RECT 220.6000 175.4000 224.2000 175.8000 ;
	    RECT 225.2000 175.4000 226.0000 179.8000 ;
	    RECT 229.4000 178.4000 230.6000 179.8000 ;
	    RECT 229.4000 177.8000 230.8000 178.4000 ;
	    RECT 234.0000 177.8000 234.8000 179.8000 ;
	    RECT 238.4000 178.4000 239.2000 179.8000 ;
	    RECT 238.4000 177.8000 240.4000 178.4000 ;
	    RECT 230.0000 177.0000 230.8000 177.8000 ;
	    RECT 234.2000 177.2000 234.8000 177.8000 ;
	    RECT 234.2000 176.6000 237.0000 177.2000 ;
	    RECT 236.2000 176.4000 237.0000 176.6000 ;
	    RECT 238.0000 176.4000 238.8000 177.2000 ;
	    RECT 239.6000 177.0000 240.4000 177.8000 ;
	    RECT 228.2000 175.4000 229.0000 175.6000 ;
	    RECT 225.2000 174.8000 229.0000 175.4000 ;
	    RECT 222.8000 174.4000 223.6000 174.8000 ;
	    RECT 218.8000 173.6000 221.4000 174.4000 ;
	    RECT 222.8000 173.8000 224.4000 174.4000 ;
	    RECT 223.6000 173.6000 224.4000 173.8000 ;
	    RECT 215.6000 171.7000 219.5000 172.3000 ;
	    RECT 215.6000 162.2000 216.4000 171.7000 ;
	    RECT 218.9000 170.4000 219.5000 171.7000 ;
	    RECT 217.2000 168.8000 218.0000 170.4000 ;
	    RECT 218.8000 170.2000 219.6000 170.4000 ;
	    RECT 220.8000 170.2000 221.4000 173.6000 ;
	    RECT 222.0000 171.6000 222.8000 173.2000 ;
	    RECT 225.2000 171.4000 226.0000 174.8000 ;
	    RECT 232.2000 174.2000 233.0000 174.4000 ;
	    RECT 238.0000 174.2000 238.6000 176.4000 ;
	    RECT 242.8000 175.0000 243.6000 179.8000 ;
	    RECT 244.4000 179.2000 248.4000 179.8000 ;
	    RECT 244.4000 175.8000 245.2000 179.2000 ;
	    RECT 246.0000 175.8000 246.8000 178.6000 ;
	    RECT 247.6000 176.0000 248.4000 179.2000 ;
	    RECT 250.8000 176.0000 251.6000 179.8000 ;
	    RECT 247.6000 175.8000 251.6000 176.0000 ;
	    RECT 254.0000 177.8000 254.8000 179.8000 ;
	    RECT 265.2000 177.8000 266.0000 179.8000 ;
	    RECT 246.0000 174.4000 246.6000 175.8000 ;
	    RECT 247.8000 175.4000 251.4000 175.8000 ;
	    RECT 250.0000 174.4000 250.8000 174.8000 ;
	    RECT 254.0000 174.4000 254.6000 177.8000 ;
	    RECT 255.6000 176.3000 256.4000 177.2000 ;
	    RECT 263.6000 176.3000 264.4000 177.2000 ;
	    RECT 255.6000 175.7000 264.4000 176.3000 ;
	    RECT 255.6000 175.6000 256.4000 175.7000 ;
	    RECT 263.6000 175.6000 264.4000 175.7000 ;
	    RECT 265.4000 174.4000 266.0000 177.8000 ;
	    RECT 241.2000 174.2000 242.8000 174.4000 ;
	    RECT 231.8000 173.6000 242.8000 174.2000 ;
	    RECT 230.0000 172.8000 230.8000 173.0000 ;
	    RECT 227.0000 172.2000 230.8000 172.8000 ;
	    RECT 227.0000 172.0000 227.8000 172.2000 ;
	    RECT 228.6000 171.4000 229.4000 171.6000 ;
	    RECT 225.2000 170.8000 229.4000 171.4000 ;
	    RECT 218.8000 169.6000 220.2000 170.2000 ;
	    RECT 220.8000 169.6000 221.8000 170.2000 ;
	    RECT 219.6000 168.4000 220.2000 169.6000 ;
	    RECT 219.6000 167.6000 220.4000 168.4000 ;
	    RECT 221.0000 164.4000 221.8000 169.6000 ;
	    RECT 221.0000 163.6000 222.8000 164.4000 ;
	    RECT 221.0000 162.2000 221.8000 163.6000 ;
	    RECT 225.2000 162.2000 226.0000 170.8000 ;
	    RECT 231.8000 170.4000 232.4000 173.6000 ;
	    RECT 239.0000 173.4000 239.8000 173.6000 ;
	    RECT 244.4000 172.8000 245.2000 174.4000 ;
	    RECT 246.0000 173.8000 248.4000 174.4000 ;
	    RECT 250.0000 173.8000 251.6000 174.4000 ;
	    RECT 247.6000 173.6000 248.4000 173.8000 ;
	    RECT 250.8000 173.6000 251.6000 173.8000 ;
	    RECT 252.4000 174.3000 253.2000 174.4000 ;
	    RECT 254.0000 174.3000 254.8000 174.4000 ;
	    RECT 252.4000 173.7000 254.8000 174.3000 ;
	    RECT 252.4000 173.6000 253.2000 173.7000 ;
	    RECT 254.0000 173.6000 254.8000 173.7000 ;
	    RECT 255.6000 174.3000 256.4000 174.4000 ;
	    RECT 265.2000 174.3000 266.0000 174.4000 ;
	    RECT 255.6000 173.7000 266.0000 174.3000 ;
	    RECT 255.6000 173.6000 256.4000 173.7000 ;
	    RECT 265.2000 173.6000 266.0000 173.7000 ;
	    RECT 240.6000 172.4000 241.4000 172.6000 ;
	    RECT 234.8000 172.3000 235.6000 172.4000 ;
	    RECT 236.4000 172.3000 241.4000 172.4000 ;
	    RECT 234.8000 171.8000 241.4000 172.3000 ;
	    RECT 234.8000 171.7000 237.2000 171.8000 ;
	    RECT 234.8000 171.6000 235.6000 171.7000 ;
	    RECT 236.4000 171.6000 237.2000 171.7000 ;
	    RECT 246.0000 171.6000 246.8000 173.2000 ;
	    RECT 238.0000 171.0000 243.6000 171.2000 ;
	    RECT 237.8000 170.8000 243.6000 171.0000 ;
	    RECT 230.0000 169.8000 232.4000 170.4000 ;
	    RECT 233.8000 170.6000 243.6000 170.8000 ;
	    RECT 233.8000 170.2000 238.6000 170.6000 ;
	    RECT 230.0000 168.8000 230.6000 169.8000 ;
	    RECT 229.2000 168.0000 230.6000 168.8000 ;
	    RECT 232.2000 169.0000 233.0000 169.2000 ;
	    RECT 233.8000 169.0000 234.4000 170.2000 ;
	    RECT 232.2000 168.4000 234.4000 169.0000 ;
	    RECT 235.0000 169.0000 240.4000 169.6000 ;
	    RECT 235.0000 168.8000 235.8000 169.0000 ;
	    RECT 239.6000 168.8000 240.4000 169.0000 ;
	    RECT 233.4000 167.4000 234.2000 167.6000 ;
	    RECT 236.2000 167.4000 237.0000 167.6000 ;
	    RECT 230.0000 166.2000 230.8000 167.0000 ;
	    RECT 233.4000 166.8000 237.0000 167.4000 ;
	    RECT 234.2000 166.2000 234.8000 166.8000 ;
	    RECT 239.6000 166.2000 240.4000 167.0000 ;
	    RECT 229.4000 162.2000 230.6000 166.2000 ;
	    RECT 234.0000 162.2000 234.8000 166.2000 ;
	    RECT 238.4000 165.6000 240.4000 166.2000 ;
	    RECT 238.4000 162.2000 239.2000 165.6000 ;
	    RECT 242.8000 162.2000 243.6000 170.6000 ;
	    RECT 247.8000 170.2000 248.4000 173.6000 ;
	    RECT 249.2000 171.6000 250.0000 173.2000 ;
	    RECT 252.4000 170.8000 253.2000 172.4000 ;
	    RECT 254.0000 170.2000 254.6000 173.6000 ;
	    RECT 255.6000 172.3000 256.4000 172.4000 ;
	    RECT 263.6000 172.3000 264.4000 172.4000 ;
	    RECT 255.6000 171.7000 264.4000 172.3000 ;
	    RECT 255.6000 171.6000 256.4000 171.7000 ;
	    RECT 263.6000 171.6000 264.4000 171.7000 ;
	    RECT 265.4000 170.2000 266.0000 173.6000 ;
	    RECT 268.4000 175.4000 269.2000 179.8000 ;
	    RECT 272.6000 178.4000 273.8000 179.8000 ;
	    RECT 272.6000 177.8000 274.0000 178.4000 ;
	    RECT 277.2000 177.8000 278.0000 179.8000 ;
	    RECT 281.6000 178.4000 282.4000 179.8000 ;
	    RECT 281.6000 177.8000 283.6000 178.4000 ;
	    RECT 273.2000 177.0000 274.0000 177.8000 ;
	    RECT 277.4000 177.2000 278.0000 177.8000 ;
	    RECT 277.4000 176.6000 280.2000 177.2000 ;
	    RECT 279.4000 176.4000 280.2000 176.6000 ;
	    RECT 281.2000 176.4000 282.0000 177.2000 ;
	    RECT 282.8000 177.0000 283.6000 177.8000 ;
	    RECT 271.4000 175.4000 272.2000 175.6000 ;
	    RECT 268.4000 174.8000 272.2000 175.4000 ;
	    RECT 266.8000 170.8000 267.6000 172.4000 ;
	    RECT 268.4000 171.4000 269.2000 174.8000 ;
	    RECT 281.2000 174.4000 281.8000 176.4000 ;
	    RECT 286.0000 175.0000 286.8000 179.8000 ;
	    RECT 287.6000 176.0000 288.4000 179.8000 ;
	    RECT 290.8000 176.0000 291.6000 179.8000 ;
	    RECT 287.6000 175.8000 291.6000 176.0000 ;
	    RECT 292.4000 175.8000 293.2000 179.8000 ;
	    RECT 294.0000 175.8000 294.8000 179.8000 ;
	    RECT 295.6000 176.0000 296.4000 179.8000 ;
	    RECT 298.8000 176.0000 299.6000 179.8000 ;
	    RECT 295.6000 175.8000 299.6000 176.0000 ;
	    RECT 287.8000 175.4000 291.4000 175.8000 ;
	    RECT 288.4000 174.4000 289.2000 174.8000 ;
	    RECT 292.4000 174.4000 293.0000 175.8000 ;
	    RECT 294.2000 174.4000 294.8000 175.8000 ;
	    RECT 295.8000 175.4000 299.4000 175.8000 ;
	    RECT 300.4000 175.0000 301.2000 179.8000 ;
	    RECT 304.8000 178.4000 305.6000 179.8000 ;
	    RECT 303.6000 177.8000 305.6000 178.4000 ;
	    RECT 309.2000 177.8000 310.0000 179.8000 ;
	    RECT 313.4000 178.4000 314.6000 179.8000 ;
	    RECT 313.2000 177.8000 314.6000 178.4000 ;
	    RECT 303.6000 177.0000 304.4000 177.8000 ;
	    RECT 309.2000 177.2000 309.8000 177.8000 ;
	    RECT 305.2000 176.4000 306.0000 177.2000 ;
	    RECT 307.0000 176.6000 309.8000 177.2000 ;
	    RECT 313.2000 177.0000 314.0000 177.8000 ;
	    RECT 307.0000 176.4000 307.8000 176.6000 ;
	    RECT 298.0000 174.4000 298.8000 174.8000 ;
	    RECT 275.4000 174.2000 276.2000 174.4000 ;
	    RECT 281.2000 174.2000 282.0000 174.4000 ;
	    RECT 284.4000 174.2000 286.0000 174.4000 ;
	    RECT 275.0000 173.6000 286.0000 174.2000 ;
	    RECT 287.6000 173.8000 289.2000 174.4000 ;
	    RECT 287.6000 173.6000 288.4000 173.8000 ;
	    RECT 290.6000 173.6000 293.2000 174.4000 ;
	    RECT 294.0000 173.6000 296.6000 174.4000 ;
	    RECT 298.0000 173.8000 299.6000 174.4000 ;
	    RECT 298.8000 173.6000 299.6000 173.8000 ;
	    RECT 301.2000 174.2000 302.8000 174.4000 ;
	    RECT 305.4000 174.2000 306.0000 176.4000 ;
	    RECT 318.0000 176.3000 318.8000 179.8000 ;
	    RECT 321.2000 177.8000 322.0000 179.8000 ;
	    RECT 319.6000 176.3000 320.4000 177.2000 ;
	    RECT 318.0000 175.7000 320.4000 176.3000 ;
	    RECT 315.0000 175.4000 315.8000 175.6000 ;
	    RECT 318.0000 175.4000 318.8000 175.7000 ;
	    RECT 319.6000 175.6000 320.4000 175.7000 ;
	    RECT 315.0000 174.8000 318.8000 175.4000 ;
	    RECT 311.0000 174.2000 311.8000 174.4000 ;
	    RECT 301.2000 173.6000 312.2000 174.2000 ;
	    RECT 273.2000 172.8000 274.0000 173.0000 ;
	    RECT 270.2000 172.2000 274.0000 172.8000 ;
	    RECT 270.2000 172.0000 271.0000 172.2000 ;
	    RECT 271.8000 171.4000 272.6000 171.6000 ;
	    RECT 268.4000 170.8000 272.6000 171.4000 ;
	    RECT 247.0000 162.2000 249.0000 170.2000 ;
	    RECT 253.0000 169.4000 254.8000 170.2000 ;
	    RECT 265.2000 169.4000 267.0000 170.2000 ;
	    RECT 253.0000 162.2000 253.8000 169.4000 ;
	    RECT 266.2000 162.2000 267.0000 169.4000 ;
	    RECT 268.4000 162.2000 269.2000 170.8000 ;
	    RECT 275.0000 170.4000 275.6000 173.6000 ;
	    RECT 282.2000 173.4000 283.0000 173.6000 ;
	    RECT 283.8000 172.4000 284.6000 172.6000 ;
	    RECT 279.6000 171.8000 284.6000 172.4000 ;
	    RECT 279.6000 171.6000 280.4000 171.8000 ;
	    RECT 289.2000 171.6000 290.0000 173.2000 ;
	    RECT 290.6000 172.3000 291.2000 173.6000 ;
	    RECT 290.6000 171.7000 294.7000 172.3000 ;
	    RECT 281.2000 171.0000 286.8000 171.2000 ;
	    RECT 281.0000 170.8000 286.8000 171.0000 ;
	    RECT 273.2000 169.8000 275.6000 170.4000 ;
	    RECT 277.0000 170.6000 286.8000 170.8000 ;
	    RECT 277.0000 170.2000 281.8000 170.6000 ;
	    RECT 273.2000 168.8000 273.8000 169.8000 ;
	    RECT 272.4000 168.0000 273.8000 168.8000 ;
	    RECT 275.4000 169.0000 276.2000 169.2000 ;
	    RECT 277.0000 169.0000 277.6000 170.2000 ;
	    RECT 275.4000 168.4000 277.6000 169.0000 ;
	    RECT 278.2000 169.0000 283.6000 169.6000 ;
	    RECT 278.2000 168.8000 279.0000 169.0000 ;
	    RECT 282.8000 168.8000 283.6000 169.0000 ;
	    RECT 276.6000 167.4000 277.4000 167.6000 ;
	    RECT 279.4000 167.4000 280.2000 167.6000 ;
	    RECT 273.2000 166.2000 274.0000 167.0000 ;
	    RECT 276.6000 166.8000 280.2000 167.4000 ;
	    RECT 277.4000 166.2000 278.0000 166.8000 ;
	    RECT 282.8000 166.2000 283.6000 167.0000 ;
	    RECT 272.6000 162.2000 273.8000 166.2000 ;
	    RECT 277.2000 162.2000 278.0000 166.2000 ;
	    RECT 281.6000 165.6000 283.6000 166.2000 ;
	    RECT 281.6000 162.2000 282.4000 165.6000 ;
	    RECT 286.0000 162.2000 286.8000 170.6000 ;
	    RECT 290.6000 170.2000 291.2000 171.7000 ;
	    RECT 294.1000 170.4000 294.7000 171.7000 ;
	    RECT 292.4000 170.2000 293.2000 170.4000 ;
	    RECT 290.2000 169.6000 291.2000 170.2000 ;
	    RECT 291.8000 169.6000 293.2000 170.2000 ;
	    RECT 294.0000 170.2000 294.8000 170.4000 ;
	    RECT 296.0000 170.2000 296.6000 173.6000 ;
	    RECT 304.2000 173.4000 305.0000 173.6000 ;
	    RECT 297.2000 171.6000 298.0000 173.2000 ;
	    RECT 302.6000 172.4000 303.4000 172.6000 ;
	    RECT 305.2000 172.4000 306.0000 172.6000 ;
	    RECT 311.6000 172.4000 312.2000 173.6000 ;
	    RECT 313.2000 172.8000 314.0000 173.0000 ;
	    RECT 302.6000 171.8000 307.6000 172.4000 ;
	    RECT 306.8000 171.6000 307.6000 171.8000 ;
	    RECT 311.6000 171.6000 312.4000 172.4000 ;
	    RECT 313.2000 172.2000 317.0000 172.8000 ;
	    RECT 316.2000 172.0000 317.0000 172.2000 ;
	    RECT 300.4000 171.0000 306.0000 171.2000 ;
	    RECT 300.4000 170.8000 306.2000 171.0000 ;
	    RECT 300.4000 170.6000 310.2000 170.8000 ;
	    RECT 294.0000 169.6000 295.4000 170.2000 ;
	    RECT 296.0000 169.6000 297.0000 170.2000 ;
	    RECT 290.2000 162.2000 291.0000 169.6000 ;
	    RECT 291.8000 168.4000 292.4000 169.6000 ;
	    RECT 294.8000 168.4000 295.4000 169.6000 ;
	    RECT 291.6000 167.6000 293.2000 168.4000 ;
	    RECT 294.8000 167.6000 295.6000 168.4000 ;
	    RECT 296.2000 162.2000 297.0000 169.6000 ;
	    RECT 300.4000 162.2000 301.2000 170.6000 ;
	    RECT 305.4000 170.2000 310.2000 170.6000 ;
	    RECT 303.6000 169.0000 309.0000 169.6000 ;
	    RECT 303.6000 168.8000 304.4000 169.0000 ;
	    RECT 308.2000 168.8000 309.0000 169.0000 ;
	    RECT 309.6000 169.0000 310.2000 170.2000 ;
	    RECT 311.6000 170.4000 312.2000 171.6000 ;
	    RECT 314.6000 171.4000 315.4000 171.6000 ;
	    RECT 318.0000 171.4000 318.8000 174.8000 ;
	    RECT 321.4000 174.4000 322.0000 177.8000 ;
	    RECT 321.2000 173.6000 322.0000 174.4000 ;
	    RECT 314.6000 170.8000 318.8000 171.4000 ;
	    RECT 311.6000 169.8000 314.0000 170.4000 ;
	    RECT 311.0000 169.0000 311.8000 169.2000 ;
	    RECT 309.6000 168.4000 311.8000 169.0000 ;
	    RECT 313.4000 168.8000 314.0000 169.8000 ;
	    RECT 313.4000 168.0000 314.8000 168.8000 ;
	    RECT 307.0000 167.4000 307.8000 167.6000 ;
	    RECT 309.8000 167.4000 310.6000 167.6000 ;
	    RECT 303.6000 166.2000 304.4000 167.0000 ;
	    RECT 307.0000 166.8000 310.6000 167.4000 ;
	    RECT 309.2000 166.2000 309.8000 166.8000 ;
	    RECT 313.2000 166.2000 314.0000 167.0000 ;
	    RECT 303.6000 165.6000 305.6000 166.2000 ;
	    RECT 304.8000 162.2000 305.6000 165.6000 ;
	    RECT 309.2000 162.2000 310.0000 166.2000 ;
	    RECT 313.4000 162.2000 314.6000 166.2000 ;
	    RECT 318.0000 162.2000 318.8000 170.8000 ;
	    RECT 321.4000 170.2000 322.0000 173.6000 ;
	    RECT 324.4000 172.4000 325.2000 179.8000 ;
	    RECT 327.6000 175.2000 328.4000 179.8000 ;
	    RECT 326.2000 174.6000 328.4000 175.2000 ;
	    RECT 322.8000 170.8000 323.6000 172.4000 ;
	    RECT 324.4000 170.2000 325.0000 172.4000 ;
	    RECT 326.2000 171.6000 326.8000 174.6000 ;
	    RECT 325.6000 170.8000 326.8000 171.6000 ;
	    RECT 326.2000 170.2000 326.8000 170.8000 ;
	    RECT 321.2000 169.4000 323.0000 170.2000 ;
	    RECT 322.2000 164.4000 323.0000 169.4000 ;
	    RECT 321.2000 163.6000 323.0000 164.4000 ;
	    RECT 322.2000 162.2000 323.0000 163.6000 ;
	    RECT 324.4000 162.2000 325.2000 170.2000 ;
	    RECT 326.2000 169.6000 328.4000 170.2000 ;
	    RECT 327.6000 162.2000 328.4000 169.6000 ;
	    RECT 329.2000 162.2000 330.0000 179.8000 ;
	    RECT 336.2000 178.4000 337.0000 179.0000 ;
	    RECT 335.6000 177.6000 337.0000 178.4000 ;
	    RECT 336.2000 176.0000 337.0000 177.6000 ;
	    RECT 340.4000 177.0000 341.2000 179.0000 ;
	    RECT 335.4000 175.4000 337.0000 176.0000 ;
	    RECT 335.4000 175.0000 336.2000 175.4000 ;
	    RECT 335.4000 174.4000 336.0000 175.0000 ;
	    RECT 340.6000 174.8000 341.2000 177.0000 ;
	    RECT 345.8000 178.4000 346.6000 179.0000 ;
	    RECT 345.8000 177.6000 347.6000 178.4000 ;
	    RECT 345.8000 176.0000 346.6000 177.6000 ;
	    RECT 350.0000 177.0000 350.8000 179.0000 ;
	    RECT 334.0000 173.6000 336.0000 174.4000 ;
	    RECT 337.0000 174.2000 341.2000 174.8000 ;
	    RECT 345.0000 175.4000 346.6000 176.0000 ;
	    RECT 345.0000 175.0000 345.8000 175.4000 ;
	    RECT 345.0000 174.4000 345.6000 175.0000 ;
	    RECT 350.2000 174.8000 350.8000 177.0000 ;
	    RECT 355.4000 176.0000 356.2000 179.0000 ;
	    RECT 359.6000 177.0000 360.4000 179.0000 ;
	    RECT 337.0000 173.8000 338.0000 174.2000 ;
	    RECT 334.0000 170.8000 334.8000 172.4000 ;
	    RECT 335.4000 169.8000 336.0000 173.6000 ;
	    RECT 336.6000 173.0000 338.0000 173.8000 ;
	    RECT 343.6000 173.6000 345.6000 174.4000 ;
	    RECT 346.6000 174.2000 350.8000 174.8000 ;
	    RECT 354.6000 175.4000 356.2000 176.0000 ;
	    RECT 354.6000 175.0000 355.4000 175.4000 ;
	    RECT 354.6000 174.4000 355.2000 175.0000 ;
	    RECT 359.8000 174.8000 360.4000 177.0000 ;
	    RECT 365.0000 176.0000 365.8000 179.0000 ;
	    RECT 369.2000 177.0000 370.0000 179.0000 ;
	    RECT 346.6000 173.8000 347.6000 174.2000 ;
	    RECT 337.4000 171.0000 338.0000 173.0000 ;
	    RECT 338.8000 171.6000 339.6000 173.2000 ;
	    RECT 340.4000 171.6000 341.2000 173.2000 ;
	    RECT 337.4000 170.4000 341.2000 171.0000 ;
	    RECT 343.6000 170.8000 344.4000 172.4000 ;
	    RECT 335.4000 169.2000 337.0000 169.8000 ;
	    RECT 336.2000 162.2000 337.0000 169.2000 ;
	    RECT 340.6000 167.0000 341.2000 170.4000 ;
	    RECT 345.0000 169.8000 345.6000 173.6000 ;
	    RECT 346.2000 173.0000 347.6000 173.8000 ;
	    RECT 353.2000 173.6000 355.2000 174.4000 ;
	    RECT 356.2000 174.2000 360.4000 174.8000 ;
	    RECT 364.2000 175.4000 365.8000 176.0000 ;
	    RECT 364.2000 175.0000 365.0000 175.4000 ;
	    RECT 364.2000 174.4000 364.8000 175.0000 ;
	    RECT 369.4000 174.8000 370.0000 177.0000 ;
	    RECT 356.2000 173.8000 357.2000 174.2000 ;
	    RECT 347.0000 171.0000 347.6000 173.0000 ;
	    RECT 348.4000 171.6000 349.2000 173.2000 ;
	    RECT 350.0000 172.3000 350.8000 173.2000 ;
	    RECT 351.6000 172.3000 352.4000 172.4000 ;
	    RECT 350.0000 171.7000 352.4000 172.3000 ;
	    RECT 350.0000 171.6000 350.8000 171.7000 ;
	    RECT 351.6000 171.6000 352.4000 171.7000 ;
	    RECT 347.0000 170.4000 350.8000 171.0000 ;
	    RECT 353.2000 170.8000 354.0000 172.4000 ;
	    RECT 345.0000 169.2000 346.6000 169.8000 ;
	    RECT 340.4000 163.0000 341.2000 167.0000 ;
	    RECT 345.8000 162.2000 346.6000 169.2000 ;
	    RECT 350.2000 167.0000 350.8000 170.4000 ;
	    RECT 354.6000 170.4000 355.2000 173.6000 ;
	    RECT 355.8000 173.0000 357.2000 173.8000 ;
	    RECT 362.8000 173.6000 364.8000 174.4000 ;
	    RECT 365.8000 174.2000 370.0000 174.8000 ;
	    RECT 370.8000 175.2000 371.6000 179.8000 ;
	    RECT 370.8000 174.6000 373.0000 175.2000 ;
	    RECT 365.8000 173.8000 366.8000 174.2000 ;
	    RECT 356.6000 171.0000 357.2000 173.0000 ;
	    RECT 358.0000 171.6000 358.8000 173.2000 ;
	    RECT 359.6000 171.6000 360.4000 173.2000 ;
	    RECT 361.2000 172.3000 362.0000 172.4000 ;
	    RECT 362.8000 172.3000 363.6000 172.4000 ;
	    RECT 361.2000 171.7000 363.6000 172.3000 ;
	    RECT 361.2000 171.6000 362.0000 171.7000 ;
	    RECT 356.6000 170.4000 360.4000 171.0000 ;
	    RECT 362.8000 170.8000 363.6000 171.7000 ;
	    RECT 354.6000 169.8000 355.6000 170.4000 ;
	    RECT 354.6000 169.2000 356.2000 169.8000 ;
	    RECT 350.0000 163.0000 350.8000 167.0000 ;
	    RECT 355.4000 162.2000 356.2000 169.2000 ;
	    RECT 359.8000 167.0000 360.4000 170.4000 ;
	    RECT 364.2000 169.8000 364.8000 173.6000 ;
	    RECT 365.4000 173.0000 366.8000 173.8000 ;
	    RECT 366.2000 171.0000 366.8000 173.0000 ;
	    RECT 367.6000 171.6000 368.4000 173.2000 ;
	    RECT 369.2000 171.6000 370.0000 173.2000 ;
	    RECT 370.8000 171.6000 371.6000 173.2000 ;
	    RECT 372.4000 171.6000 373.0000 174.6000 ;
	    RECT 374.0000 172.4000 374.8000 179.8000 ;
	    RECT 377.2000 175.2000 378.0000 179.8000 ;
	    RECT 380.4000 175.2000 381.2000 179.8000 ;
	    RECT 383.6000 175.2000 384.4000 179.8000 ;
	    RECT 386.8000 175.2000 387.6000 179.8000 ;
	    RECT 390.6000 176.4000 391.4000 179.8000 ;
	    RECT 390.6000 175.8000 392.4000 176.4000 ;
	    RECT 366.2000 170.4000 370.0000 171.0000 ;
	    RECT 364.2000 169.2000 365.8000 169.8000 ;
	    RECT 359.6000 163.0000 360.4000 167.0000 ;
	    RECT 365.0000 164.4000 365.8000 169.2000 ;
	    RECT 369.4000 167.0000 370.0000 170.4000 ;
	    RECT 372.4000 170.8000 373.6000 171.6000 ;
	    RECT 372.4000 170.2000 373.0000 170.8000 ;
	    RECT 374.2000 170.2000 374.8000 172.4000 ;
	    RECT 375.6000 174.4000 378.0000 175.2000 ;
	    RECT 379.0000 174.4000 381.2000 175.2000 ;
	    RECT 382.2000 174.4000 384.4000 175.2000 ;
	    RECT 385.8000 174.4000 387.6000 175.2000 ;
	    RECT 375.6000 171.6000 376.4000 174.4000 ;
	    RECT 379.0000 173.8000 379.8000 174.4000 ;
	    RECT 382.2000 173.8000 383.0000 174.4000 ;
	    RECT 385.8000 173.8000 386.6000 174.4000 ;
	    RECT 377.2000 173.0000 379.8000 173.8000 ;
	    RECT 380.6000 173.0000 383.0000 173.8000 ;
	    RECT 384.0000 173.0000 386.6000 173.8000 ;
	    RECT 379.0000 171.6000 379.8000 173.0000 ;
	    RECT 382.2000 171.6000 383.0000 173.0000 ;
	    RECT 385.8000 171.6000 386.6000 173.0000 ;
	    RECT 375.6000 170.8000 378.0000 171.6000 ;
	    RECT 379.0000 170.8000 381.2000 171.6000 ;
	    RECT 382.2000 170.8000 384.4000 171.6000 ;
	    RECT 385.8000 170.8000 387.6000 171.6000 ;
	    RECT 364.4000 163.6000 365.8000 164.4000 ;
	    RECT 365.0000 162.2000 365.8000 163.6000 ;
	    RECT 369.2000 163.0000 370.0000 167.0000 ;
	    RECT 370.8000 169.6000 373.0000 170.2000 ;
	    RECT 370.8000 162.2000 371.6000 169.6000 ;
	    RECT 374.0000 162.2000 374.8000 170.2000 ;
	    RECT 377.2000 162.2000 378.0000 170.8000 ;
	    RECT 380.4000 162.2000 381.2000 170.8000 ;
	    RECT 383.6000 162.2000 384.4000 170.8000 ;
	    RECT 386.8000 162.2000 387.6000 170.8000 ;
	    RECT 390.0000 168.8000 390.8000 170.4000 ;
	    RECT 391.6000 162.2000 392.4000 175.8000 ;
	    RECT 394.8000 175.4000 395.6000 179.8000 ;
	    RECT 399.0000 178.4000 400.2000 179.8000 ;
	    RECT 399.0000 177.8000 400.4000 178.4000 ;
	    RECT 403.6000 177.8000 404.4000 179.8000 ;
	    RECT 408.0000 178.4000 408.8000 179.8000 ;
	    RECT 408.0000 177.8000 410.0000 178.4000 ;
	    RECT 399.6000 177.0000 400.4000 177.8000 ;
	    RECT 403.8000 177.2000 404.4000 177.8000 ;
	    RECT 403.8000 176.6000 406.6000 177.2000 ;
	    RECT 405.8000 176.4000 406.6000 176.6000 ;
	    RECT 407.6000 176.4000 408.4000 177.2000 ;
	    RECT 409.2000 177.0000 410.0000 177.8000 ;
	    RECT 397.8000 175.4000 398.6000 175.6000 ;
	    RECT 393.2000 173.6000 394.0000 175.2000 ;
	    RECT 394.8000 174.8000 398.6000 175.4000 ;
	    RECT 394.8000 171.4000 395.6000 174.8000 ;
	    RECT 401.8000 174.2000 403.6000 174.4000 ;
	    RECT 407.6000 174.2000 408.2000 176.4000 ;
	    RECT 412.4000 175.0000 413.2000 179.8000 ;
	    RECT 420.4000 175.8000 421.2000 179.8000 ;
	    RECT 422.0000 176.0000 422.8000 179.8000 ;
	    RECT 425.2000 176.0000 426.0000 179.8000 ;
	    RECT 427.4000 178.4000 428.2000 179.8000 ;
	    RECT 426.8000 177.6000 428.2000 178.4000 ;
	    RECT 422.0000 175.8000 426.0000 176.0000 ;
	    RECT 427.4000 176.4000 428.2000 177.6000 ;
	    RECT 427.4000 175.8000 429.2000 176.4000 ;
	    RECT 420.6000 174.4000 421.2000 175.8000 ;
	    RECT 422.2000 175.4000 425.8000 175.8000 ;
	    RECT 424.4000 174.4000 425.2000 174.8000 ;
	    RECT 410.8000 174.2000 412.4000 174.4000 ;
	    RECT 401.4000 173.6000 412.4000 174.2000 ;
	    RECT 414.0000 174.3000 414.8000 174.4000 ;
	    RECT 420.4000 174.3000 423.0000 174.4000 ;
	    RECT 414.0000 173.7000 423.0000 174.3000 ;
	    RECT 424.4000 173.8000 426.0000 174.4000 ;
	    RECT 414.0000 173.6000 414.8000 173.7000 ;
	    RECT 420.4000 173.6000 423.0000 173.7000 ;
	    RECT 425.2000 173.6000 426.0000 173.8000 ;
	    RECT 399.6000 172.8000 400.4000 173.0000 ;
	    RECT 396.6000 172.2000 400.4000 172.8000 ;
	    RECT 396.6000 172.0000 397.4000 172.2000 ;
	    RECT 398.2000 171.4000 399.0000 171.6000 ;
	    RECT 394.8000 170.8000 399.0000 171.4000 ;
	    RECT 393.2000 168.3000 394.0000 168.4000 ;
	    RECT 394.8000 168.3000 395.6000 170.8000 ;
	    RECT 401.4000 170.4000 402.0000 173.6000 ;
	    RECT 408.6000 173.4000 409.4000 173.6000 ;
	    RECT 407.6000 172.4000 408.4000 172.6000 ;
	    RECT 410.2000 172.4000 411.0000 172.6000 ;
	    RECT 406.0000 171.8000 411.0000 172.4000 ;
	    RECT 406.0000 171.6000 406.8000 171.8000 ;
	    RECT 407.6000 171.0000 413.2000 171.2000 ;
	    RECT 407.4000 170.8000 413.2000 171.0000 ;
	    RECT 399.6000 169.8000 402.0000 170.4000 ;
	    RECT 403.4000 170.6000 413.2000 170.8000 ;
	    RECT 403.4000 170.2000 408.2000 170.6000 ;
	    RECT 399.6000 168.8000 400.2000 169.8000 ;
	    RECT 393.2000 167.7000 395.6000 168.3000 ;
	    RECT 398.8000 168.0000 400.2000 168.8000 ;
	    RECT 401.8000 169.0000 402.6000 169.2000 ;
	    RECT 403.4000 169.0000 404.0000 170.2000 ;
	    RECT 401.8000 168.4000 404.0000 169.0000 ;
	    RECT 404.6000 169.0000 410.0000 169.6000 ;
	    RECT 404.6000 168.8000 405.4000 169.0000 ;
	    RECT 409.2000 168.8000 410.0000 169.0000 ;
	    RECT 393.2000 167.6000 394.0000 167.7000 ;
	    RECT 394.8000 162.2000 395.6000 167.7000 ;
	    RECT 403.0000 167.4000 403.8000 167.6000 ;
	    RECT 405.8000 167.4000 406.6000 167.6000 ;
	    RECT 399.6000 166.2000 400.4000 167.0000 ;
	    RECT 403.0000 166.8000 406.6000 167.4000 ;
	    RECT 403.8000 166.2000 404.4000 166.8000 ;
	    RECT 409.2000 166.2000 410.0000 167.0000 ;
	    RECT 399.0000 162.2000 400.2000 166.2000 ;
	    RECT 403.6000 162.2000 404.4000 166.2000 ;
	    RECT 408.0000 165.6000 410.0000 166.2000 ;
	    RECT 408.0000 162.2000 408.8000 165.6000 ;
	    RECT 412.4000 162.2000 413.2000 170.6000 ;
	    RECT 420.4000 170.2000 421.2000 170.4000 ;
	    RECT 422.4000 170.2000 423.0000 173.6000 ;
	    RECT 423.6000 171.6000 424.4000 173.2000 ;
	    RECT 420.4000 169.6000 421.8000 170.2000 ;
	    RECT 422.4000 169.6000 423.4000 170.2000 ;
	    RECT 421.2000 168.4000 421.8000 169.6000 ;
	    RECT 421.2000 167.6000 422.0000 168.4000 ;
	    RECT 422.6000 162.2000 423.4000 169.6000 ;
	    RECT 426.8000 168.8000 427.6000 170.4000 ;
	    RECT 428.4000 162.2000 429.2000 175.8000 ;
	    RECT 430.0000 173.6000 430.8000 175.2000 ;
	    RECT 430.0000 170.3000 430.8000 170.4000 ;
	    RECT 431.6000 170.3000 432.4000 179.8000 ;
	    RECT 436.0000 178.4000 436.8000 179.8000 ;
	    RECT 436.0000 177.6000 437.2000 178.4000 ;
	    RECT 436.0000 174.2000 436.8000 177.6000 ;
	    RECT 435.0000 173.8000 436.8000 174.2000 ;
	    RECT 435.0000 173.6000 436.6000 173.8000 ;
	    RECT 435.0000 170.4000 435.6000 173.6000 ;
	    RECT 437.2000 171.6000 438.8000 172.4000 ;
	    RECT 430.0000 169.7000 432.4000 170.3000 ;
	    RECT 430.0000 169.6000 430.8000 169.7000 ;
	    RECT 431.6000 162.2000 432.4000 169.7000 ;
	    RECT 434.8000 169.6000 435.6000 170.4000 ;
	    RECT 439.6000 170.3000 440.4000 172.4000 ;
	    RECT 441.2000 172.3000 442.0000 179.8000 ;
	    RECT 446.0000 177.8000 446.8000 179.8000 ;
	    RECT 450.8000 177.8000 451.6000 179.8000 ;
	    RECT 446.0000 174.4000 446.6000 177.8000 ;
	    RECT 450.8000 176.4000 451.4000 177.8000 ;
	    RECT 450.8000 175.6000 451.6000 176.4000 ;
	    RECT 450.8000 174.4000 451.4000 175.6000 ;
	    RECT 454.0000 175.2000 454.8000 179.8000 ;
	    RECT 454.0000 174.6000 456.2000 175.2000 ;
	    RECT 446.0000 174.3000 446.8000 174.4000 ;
	    RECT 447.6000 174.3000 448.4000 174.4000 ;
	    RECT 446.0000 173.7000 448.4000 174.3000 ;
	    RECT 446.0000 173.6000 446.8000 173.7000 ;
	    RECT 447.6000 173.6000 448.4000 173.7000 ;
	    RECT 450.8000 173.6000 451.6000 174.4000 ;
	    RECT 444.4000 172.3000 445.2000 172.4000 ;
	    RECT 441.2000 171.7000 445.2000 172.3000 ;
	    RECT 441.2000 170.3000 442.0000 171.7000 ;
	    RECT 444.4000 170.8000 445.2000 171.7000 ;
	    RECT 439.6000 169.7000 442.0000 170.3000 ;
	    RECT 446.0000 170.2000 446.6000 173.6000 ;
	    RECT 447.6000 172.3000 448.4000 172.4000 ;
	    RECT 449.2000 172.3000 450.0000 172.4000 ;
	    RECT 447.6000 171.7000 450.0000 172.3000 ;
	    RECT 447.6000 171.6000 448.4000 171.7000 ;
	    RECT 449.2000 170.8000 450.0000 171.7000 ;
	    RECT 450.8000 170.2000 451.4000 173.6000 ;
	    RECT 454.0000 171.6000 454.8000 173.2000 ;
	    RECT 455.6000 171.6000 456.2000 174.6000 ;
	    RECT 457.2000 172.4000 458.0000 179.8000 ;
	    RECT 462.4000 174.2000 463.2000 179.8000 ;
	    RECT 465.2000 175.2000 466.0000 179.8000 ;
	    RECT 465.2000 174.6000 467.4000 175.2000 ;
	    RECT 462.4000 173.8000 464.2000 174.2000 ;
	    RECT 462.6000 173.6000 464.2000 173.8000 ;
	    RECT 455.6000 170.8000 456.8000 171.6000 ;
	    RECT 455.6000 170.2000 456.2000 170.8000 ;
	    RECT 457.4000 170.2000 458.0000 172.4000 ;
	    RECT 460.4000 171.6000 462.0000 172.4000 ;
	    RECT 439.6000 169.6000 440.4000 169.7000 ;
	    RECT 435.0000 167.0000 435.6000 169.6000 ;
	    RECT 436.4000 167.6000 437.2000 169.2000 ;
	    RECT 435.0000 166.4000 438.6000 167.0000 ;
	    RECT 435.0000 166.2000 435.6000 166.4000 ;
	    RECT 434.8000 162.2000 435.6000 166.2000 ;
	    RECT 438.0000 166.2000 438.6000 166.4000 ;
	    RECT 438.0000 162.2000 438.8000 166.2000 ;
	    RECT 441.2000 162.2000 442.0000 169.7000 ;
	    RECT 445.0000 169.4000 446.8000 170.2000 ;
	    RECT 449.8000 169.4000 451.6000 170.2000 ;
	    RECT 454.0000 169.6000 456.2000 170.2000 ;
	    RECT 445.0000 162.2000 445.8000 169.4000 ;
	    RECT 449.8000 162.2000 450.6000 169.4000 ;
	    RECT 454.0000 162.2000 454.8000 169.6000 ;
	    RECT 457.2000 168.3000 458.0000 170.2000 ;
	    RECT 463.6000 170.4000 464.2000 173.6000 ;
	    RECT 465.2000 171.6000 466.0000 173.2000 ;
	    RECT 466.8000 171.6000 467.4000 174.6000 ;
	    RECT 468.4000 172.4000 469.2000 179.8000 ;
	    RECT 470.0000 175.2000 470.8000 179.8000 ;
	    RECT 470.0000 174.6000 472.2000 175.2000 ;
	    RECT 466.8000 170.8000 468.0000 171.6000 ;
	    RECT 463.6000 169.6000 464.4000 170.4000 ;
	    RECT 466.8000 170.2000 467.4000 170.8000 ;
	    RECT 468.6000 170.2000 469.2000 172.4000 ;
	    RECT 470.0000 171.6000 470.8000 173.2000 ;
	    RECT 471.6000 171.6000 472.2000 174.6000 ;
	    RECT 473.2000 172.4000 474.0000 179.8000 ;
	    RECT 476.0000 174.2000 476.8000 179.8000 ;
	    RECT 481.2000 175.2000 482.0000 179.8000 ;
	    RECT 481.2000 174.6000 483.4000 175.2000 ;
	    RECT 471.6000 170.8000 472.8000 171.6000 ;
	    RECT 471.6000 170.2000 472.2000 170.8000 ;
	    RECT 473.4000 170.2000 474.0000 172.4000 ;
	    RECT 475.0000 173.8000 476.8000 174.2000 ;
	    RECT 475.0000 173.6000 476.6000 173.8000 ;
	    RECT 475.0000 170.4000 475.6000 173.6000 ;
	    RECT 477.2000 171.6000 478.8000 172.4000 ;
	    RECT 481.2000 171.6000 482.0000 173.2000 ;
	    RECT 482.8000 171.6000 483.4000 174.6000 ;
	    RECT 484.4000 172.4000 485.2000 179.8000 ;
	    RECT 465.2000 169.6000 467.4000 170.2000 ;
	    RECT 462.0000 168.3000 462.8000 169.2000 ;
	    RECT 457.2000 167.7000 462.8000 168.3000 ;
	    RECT 457.2000 162.2000 458.0000 167.7000 ;
	    RECT 462.0000 167.6000 462.8000 167.7000 ;
	    RECT 463.6000 167.0000 464.2000 169.6000 ;
	    RECT 460.6000 166.4000 464.2000 167.0000 ;
	    RECT 460.6000 166.2000 461.2000 166.4000 ;
	    RECT 460.4000 162.2000 461.2000 166.2000 ;
	    RECT 463.6000 166.2000 464.2000 166.4000 ;
	    RECT 463.6000 162.2000 464.4000 166.2000 ;
	    RECT 465.2000 162.2000 466.0000 169.6000 ;
	    RECT 468.4000 162.2000 469.2000 170.2000 ;
	    RECT 470.0000 169.6000 472.2000 170.2000 ;
	    RECT 470.0000 162.2000 470.8000 169.6000 ;
	    RECT 473.2000 162.2000 474.0000 170.2000 ;
	    RECT 474.8000 169.6000 475.6000 170.4000 ;
	    RECT 482.8000 170.8000 484.0000 171.6000 ;
	    RECT 482.8000 170.2000 483.4000 170.8000 ;
	    RECT 484.6000 170.2000 485.2000 172.4000 ;
	    RECT 475.0000 167.0000 475.6000 169.6000 ;
	    RECT 481.2000 169.6000 483.4000 170.2000 ;
	    RECT 476.4000 167.6000 477.2000 169.2000 ;
	    RECT 475.0000 166.4000 478.6000 167.0000 ;
	    RECT 475.0000 166.2000 475.6000 166.4000 ;
	    RECT 474.8000 162.2000 475.6000 166.2000 ;
	    RECT 478.0000 166.2000 478.6000 166.4000 ;
	    RECT 478.0000 162.2000 478.8000 166.2000 ;
	    RECT 481.2000 162.2000 482.0000 169.6000 ;
	    RECT 484.4000 162.2000 485.2000 170.2000 ;
	    RECT 486.0000 175.4000 486.8000 179.8000 ;
	    RECT 490.2000 178.4000 491.4000 179.8000 ;
	    RECT 490.2000 177.8000 491.6000 178.4000 ;
	    RECT 494.8000 177.8000 495.6000 179.8000 ;
	    RECT 499.2000 178.4000 500.0000 179.8000 ;
	    RECT 499.2000 177.8000 501.2000 178.4000 ;
	    RECT 490.8000 177.0000 491.6000 177.8000 ;
	    RECT 495.0000 177.2000 495.6000 177.8000 ;
	    RECT 495.0000 176.6000 497.8000 177.2000 ;
	    RECT 497.0000 176.4000 497.8000 176.6000 ;
	    RECT 498.8000 176.4000 499.6000 177.2000 ;
	    RECT 500.4000 177.0000 501.2000 177.8000 ;
	    RECT 489.0000 175.4000 489.8000 175.6000 ;
	    RECT 486.0000 174.8000 489.8000 175.4000 ;
	    RECT 486.0000 171.4000 486.8000 174.8000 ;
	    RECT 493.0000 174.2000 493.8000 174.4000 ;
	    RECT 497.2000 174.2000 498.0000 174.4000 ;
	    RECT 498.8000 174.2000 499.4000 176.4000 ;
	    RECT 503.6000 175.0000 504.4000 179.8000 ;
	    RECT 505.2000 175.6000 506.0000 177.2000 ;
	    RECT 502.0000 174.2000 503.6000 174.4000 ;
	    RECT 492.6000 173.6000 503.6000 174.2000 ;
	    RECT 506.8000 174.3000 507.6000 179.8000 ;
	    RECT 508.4000 176.0000 509.2000 179.8000 ;
	    RECT 511.6000 176.0000 512.4000 179.8000 ;
	    RECT 508.4000 175.8000 512.4000 176.0000 ;
	    RECT 513.2000 175.8000 514.0000 179.8000 ;
	    RECT 508.6000 175.4000 512.2000 175.8000 ;
	    RECT 509.2000 174.4000 510.0000 174.8000 ;
	    RECT 513.2000 174.4000 513.8000 175.8000 ;
	    RECT 508.4000 174.3000 510.0000 174.4000 ;
	    RECT 506.8000 173.8000 510.0000 174.3000 ;
	    RECT 506.8000 173.7000 509.2000 173.8000 ;
	    RECT 490.8000 172.8000 491.6000 173.0000 ;
	    RECT 487.8000 172.2000 491.6000 172.8000 ;
	    RECT 487.8000 172.0000 488.6000 172.2000 ;
	    RECT 489.4000 171.4000 490.2000 171.6000 ;
	    RECT 486.0000 170.8000 490.2000 171.4000 ;
	    RECT 486.0000 162.2000 486.8000 170.8000 ;
	    RECT 492.6000 170.4000 493.2000 173.6000 ;
	    RECT 499.8000 173.4000 500.6000 173.6000 ;
	    RECT 498.8000 172.4000 499.6000 172.6000 ;
	    RECT 501.4000 172.4000 502.2000 172.6000 ;
	    RECT 497.2000 171.8000 502.2000 172.4000 ;
	    RECT 497.2000 171.6000 498.0000 171.8000 ;
	    RECT 498.8000 171.0000 504.4000 171.2000 ;
	    RECT 498.6000 170.8000 504.4000 171.0000 ;
	    RECT 490.8000 169.8000 493.2000 170.4000 ;
	    RECT 494.6000 170.6000 504.4000 170.8000 ;
	    RECT 494.6000 170.2000 499.4000 170.6000 ;
	    RECT 490.8000 168.8000 491.4000 169.8000 ;
	    RECT 490.0000 168.0000 491.4000 168.8000 ;
	    RECT 493.0000 169.0000 493.8000 169.2000 ;
	    RECT 494.6000 169.0000 495.2000 170.2000 ;
	    RECT 493.0000 168.4000 495.2000 169.0000 ;
	    RECT 495.8000 169.0000 501.2000 169.6000 ;
	    RECT 495.8000 168.8000 496.6000 169.0000 ;
	    RECT 500.4000 168.8000 501.2000 169.0000 ;
	    RECT 494.2000 167.4000 495.0000 167.6000 ;
	    RECT 497.0000 167.4000 497.8000 167.6000 ;
	    RECT 490.8000 166.2000 491.6000 167.0000 ;
	    RECT 494.2000 166.8000 497.8000 167.4000 ;
	    RECT 495.0000 166.2000 495.6000 166.8000 ;
	    RECT 500.4000 166.2000 501.2000 167.0000 ;
	    RECT 490.2000 162.2000 491.4000 166.2000 ;
	    RECT 494.8000 162.2000 495.6000 166.2000 ;
	    RECT 499.2000 165.6000 501.2000 166.2000 ;
	    RECT 499.2000 162.2000 500.0000 165.6000 ;
	    RECT 503.6000 162.2000 504.4000 170.6000 ;
	    RECT 506.8000 162.2000 507.6000 173.7000 ;
	    RECT 508.4000 173.6000 509.2000 173.7000 ;
	    RECT 511.4000 173.6000 514.0000 174.4000 ;
	    RECT 510.0000 171.6000 510.8000 173.2000 ;
	    RECT 511.4000 170.2000 512.0000 173.6000 ;
	    RECT 513.2000 170.2000 514.0000 170.4000 ;
	    RECT 511.0000 169.6000 512.0000 170.2000 ;
	    RECT 512.6000 169.6000 514.0000 170.2000 ;
	    RECT 511.0000 162.2000 511.8000 169.6000 ;
	    RECT 512.6000 168.4000 513.2000 169.6000 ;
	    RECT 512.4000 167.6000 513.2000 168.4000 ;
	    RECT 4.4000 152.4000 5.2000 159.8000 ;
	    RECT 3.0000 151.8000 5.2000 152.4000 ;
	    RECT 6.0000 152.4000 6.8000 159.8000 ;
	    RECT 6.0000 151.8000 8.2000 152.4000 ;
	    RECT 9.2000 151.8000 10.0000 159.8000 ;
	    RECT 10.8000 152.4000 11.6000 159.8000 ;
	    RECT 10.8000 151.8000 13.0000 152.4000 ;
	    RECT 14.0000 151.8000 14.8000 159.8000 ;
	    RECT 18.2000 158.4000 19.0000 159.8000 ;
	    RECT 17.2000 157.6000 19.0000 158.4000 ;
	    RECT 18.2000 152.4000 19.0000 157.6000 ;
	    RECT 19.6000 154.3000 20.4000 154.4000 ;
	    RECT 22.0000 154.3000 22.8000 159.8000 ;
	    RECT 26.2000 155.8000 27.4000 159.8000 ;
	    RECT 30.8000 155.8000 31.6000 159.8000 ;
	    RECT 35.2000 156.4000 36.0000 159.8000 ;
	    RECT 35.2000 155.8000 37.2000 156.4000 ;
	    RECT 26.8000 155.0000 27.6000 155.8000 ;
	    RECT 31.0000 155.2000 31.6000 155.8000 ;
	    RECT 30.2000 154.6000 33.8000 155.2000 ;
	    RECT 36.4000 155.0000 37.2000 155.8000 ;
	    RECT 30.2000 154.4000 31.0000 154.6000 ;
	    RECT 33.0000 154.4000 33.8000 154.6000 ;
	    RECT 19.6000 153.7000 22.8000 154.3000 ;
	    RECT 19.6000 153.6000 20.4000 153.7000 ;
	    RECT 19.8000 152.4000 20.4000 153.6000 ;
	    RECT 18.2000 151.8000 19.2000 152.4000 ;
	    RECT 19.8000 151.8000 21.2000 152.4000 ;
	    RECT 3.0000 151.2000 3.6000 151.8000 ;
	    RECT 2.4000 150.4000 3.6000 151.2000 ;
	    RECT 7.6000 151.2000 8.2000 151.8000 ;
	    RECT 7.6000 150.4000 8.8000 151.2000 ;
	    RECT 3.0000 147.4000 3.6000 150.4000 ;
	    RECT 4.4000 148.8000 5.2000 150.4000 ;
	    RECT 6.0000 148.8000 6.8000 150.4000 ;
	    RECT 7.6000 147.4000 8.2000 150.4000 ;
	    RECT 9.4000 149.6000 10.0000 151.8000 ;
	    RECT 3.0000 146.8000 5.2000 147.4000 ;
	    RECT 4.4000 142.2000 5.2000 146.8000 ;
	    RECT 6.0000 146.8000 8.2000 147.4000 ;
	    RECT 6.0000 142.2000 6.8000 146.8000 ;
	    RECT 9.2000 142.2000 10.0000 149.6000 ;
	    RECT 12.4000 151.2000 13.0000 151.8000 ;
	    RECT 12.4000 150.4000 13.6000 151.2000 ;
	    RECT 12.4000 147.4000 13.0000 150.4000 ;
	    RECT 14.2000 149.6000 14.8000 151.8000 ;
	    RECT 10.8000 146.8000 13.0000 147.4000 ;
	    RECT 14.0000 148.3000 14.8000 149.6000 ;
	    RECT 17.2000 148.8000 18.0000 150.4000 ;
	    RECT 18.6000 148.4000 19.2000 151.8000 ;
	    RECT 20.4000 151.6000 21.2000 151.8000 ;
	    RECT 22.0000 151.2000 22.8000 153.7000 ;
	    RECT 26.0000 153.2000 27.4000 154.0000 ;
	    RECT 26.8000 152.2000 27.4000 153.2000 ;
	    RECT 29.0000 153.0000 31.2000 153.6000 ;
	    RECT 29.0000 152.8000 29.8000 153.0000 ;
	    RECT 26.8000 151.6000 29.2000 152.2000 ;
	    RECT 22.0000 150.6000 26.2000 151.2000 ;
	    RECT 15.6000 148.3000 16.4000 148.4000 ;
	    RECT 14.0000 148.2000 16.4000 148.3000 ;
	    RECT 14.0000 147.7000 17.2000 148.2000 ;
	    RECT 10.8000 142.2000 11.6000 146.8000 ;
	    RECT 14.0000 142.2000 14.8000 147.7000 ;
	    RECT 15.6000 147.6000 17.2000 147.7000 ;
	    RECT 18.6000 147.6000 21.2000 148.4000 ;
	    RECT 16.4000 147.2000 17.2000 147.6000 ;
	    RECT 15.8000 146.2000 19.4000 146.6000 ;
	    RECT 20.4000 146.2000 21.0000 147.6000 ;
	    RECT 22.0000 147.2000 22.8000 150.6000 ;
	    RECT 25.4000 150.4000 26.2000 150.6000 ;
	    RECT 23.8000 149.8000 24.6000 150.0000 ;
	    RECT 23.8000 149.2000 27.6000 149.8000 ;
	    RECT 26.8000 149.0000 27.6000 149.2000 ;
	    RECT 28.6000 148.4000 29.2000 151.6000 ;
	    RECT 30.6000 151.8000 31.2000 153.0000 ;
	    RECT 31.8000 153.0000 32.6000 153.2000 ;
	    RECT 36.4000 153.0000 37.2000 153.2000 ;
	    RECT 31.8000 152.4000 37.2000 153.0000 ;
	    RECT 30.6000 151.4000 35.4000 151.8000 ;
	    RECT 39.6000 151.4000 40.4000 159.8000 ;
	    RECT 30.6000 151.2000 40.4000 151.4000 ;
	    RECT 34.6000 151.0000 40.4000 151.2000 ;
	    RECT 34.8000 150.8000 40.4000 151.0000 ;
	    RECT 41.2000 151.4000 42.0000 159.8000 ;
	    RECT 45.6000 156.4000 46.4000 159.8000 ;
	    RECT 44.4000 155.8000 46.4000 156.4000 ;
	    RECT 50.0000 155.8000 50.8000 159.8000 ;
	    RECT 54.2000 155.8000 55.4000 159.8000 ;
	    RECT 44.4000 155.0000 45.2000 155.8000 ;
	    RECT 50.0000 155.2000 50.6000 155.8000 ;
	    RECT 47.8000 154.6000 51.4000 155.2000 ;
	    RECT 54.0000 155.0000 54.8000 155.8000 ;
	    RECT 47.8000 154.4000 48.6000 154.6000 ;
	    RECT 50.6000 154.4000 51.4000 154.6000 ;
	    RECT 44.4000 153.0000 45.2000 153.2000 ;
	    RECT 49.0000 153.0000 49.8000 153.2000 ;
	    RECT 44.4000 152.4000 49.8000 153.0000 ;
	    RECT 50.4000 153.0000 52.6000 153.6000 ;
	    RECT 50.4000 151.8000 51.0000 153.0000 ;
	    RECT 51.8000 152.8000 52.6000 153.0000 ;
	    RECT 54.2000 153.2000 55.6000 154.0000 ;
	    RECT 54.2000 152.2000 54.8000 153.2000 ;
	    RECT 46.2000 151.4000 51.0000 151.8000 ;
	    RECT 41.2000 151.2000 51.0000 151.4000 ;
	    RECT 52.4000 151.6000 54.8000 152.2000 ;
	    RECT 41.2000 151.0000 47.0000 151.2000 ;
	    RECT 41.2000 150.8000 46.8000 151.0000 ;
	    RECT 31.6000 150.3000 32.4000 150.4000 ;
	    RECT 33.2000 150.3000 34.0000 150.4000 ;
	    RECT 31.6000 150.2000 34.0000 150.3000 ;
	    RECT 47.6000 150.2000 48.4000 150.4000 ;
	    RECT 31.6000 149.7000 38.2000 150.2000 ;
	    RECT 31.6000 149.6000 32.4000 149.7000 ;
	    RECT 33.2000 149.6000 38.2000 149.7000 ;
	    RECT 37.4000 149.4000 38.2000 149.6000 ;
	    RECT 43.4000 149.6000 48.4000 150.2000 ;
	    RECT 43.4000 149.4000 44.2000 149.6000 ;
	    RECT 35.8000 148.4000 36.6000 148.6000 ;
	    RECT 45.0000 148.4000 45.8000 148.6000 ;
	    RECT 52.4000 148.4000 53.0000 151.6000 ;
	    RECT 58.8000 151.2000 59.6000 159.8000 ;
	    RECT 55.4000 150.6000 59.6000 151.2000 ;
	    RECT 60.4000 151.4000 61.2000 159.8000 ;
	    RECT 64.8000 156.4000 65.6000 159.8000 ;
	    RECT 63.6000 155.8000 65.6000 156.4000 ;
	    RECT 69.2000 155.8000 70.0000 159.8000 ;
	    RECT 73.4000 155.8000 74.6000 159.8000 ;
	    RECT 63.6000 155.0000 64.4000 155.8000 ;
	    RECT 69.2000 155.2000 69.8000 155.8000 ;
	    RECT 67.0000 154.6000 70.6000 155.2000 ;
	    RECT 73.2000 155.0000 74.0000 155.8000 ;
	    RECT 67.0000 154.4000 67.8000 154.6000 ;
	    RECT 69.8000 154.4000 70.6000 154.6000 ;
	    RECT 63.6000 153.0000 64.4000 153.2000 ;
	    RECT 68.2000 153.0000 69.0000 153.2000 ;
	    RECT 63.6000 152.4000 69.0000 153.0000 ;
	    RECT 69.6000 153.0000 71.8000 153.6000 ;
	    RECT 69.6000 151.8000 70.2000 153.0000 ;
	    RECT 71.0000 152.8000 71.8000 153.0000 ;
	    RECT 73.4000 153.2000 74.8000 154.0000 ;
	    RECT 73.4000 152.2000 74.0000 153.2000 ;
	    RECT 65.4000 151.4000 70.2000 151.8000 ;
	    RECT 60.4000 151.2000 70.2000 151.4000 ;
	    RECT 71.6000 151.6000 74.0000 152.2000 ;
	    RECT 60.4000 151.0000 66.2000 151.2000 ;
	    RECT 60.4000 150.8000 66.0000 151.0000 ;
	    RECT 55.4000 150.4000 56.2000 150.6000 ;
	    RECT 57.0000 149.8000 57.8000 150.0000 ;
	    RECT 54.0000 149.2000 57.8000 149.8000 ;
	    RECT 54.0000 149.0000 54.8000 149.2000 ;
	    RECT 28.4000 148.3000 39.6000 148.4000 ;
	    RECT 42.0000 148.3000 53.2000 148.4000 ;
	    RECT 28.4000 147.8000 53.2000 148.3000 ;
	    RECT 28.4000 147.6000 29.8000 147.8000 ;
	    RECT 22.0000 146.6000 25.8000 147.2000 ;
	    RECT 15.6000 146.0000 19.6000 146.2000 ;
	    RECT 15.6000 142.2000 16.4000 146.0000 ;
	    RECT 18.8000 142.2000 19.6000 146.0000 ;
	    RECT 20.4000 142.2000 21.2000 146.2000 ;
	    RECT 22.0000 142.2000 22.8000 146.6000 ;
	    RECT 25.0000 146.4000 25.8000 146.6000 ;
	    RECT 34.8000 145.6000 35.4000 147.8000 ;
	    RECT 38.0000 147.7000 43.6000 147.8000 ;
	    RECT 38.0000 147.6000 39.6000 147.7000 ;
	    RECT 42.0000 147.6000 43.6000 147.7000 ;
	    RECT 33.0000 145.4000 33.8000 145.6000 ;
	    RECT 26.8000 144.2000 27.6000 145.0000 ;
	    RECT 31.0000 144.8000 33.8000 145.4000 ;
	    RECT 34.8000 144.8000 35.6000 145.6000 ;
	    RECT 31.0000 144.2000 31.6000 144.8000 ;
	    RECT 36.4000 144.2000 37.2000 145.0000 ;
	    RECT 26.2000 143.6000 27.6000 144.2000 ;
	    RECT 26.2000 142.2000 27.4000 143.6000 ;
	    RECT 30.8000 142.2000 31.6000 144.2000 ;
	    RECT 35.2000 143.6000 37.2000 144.2000 ;
	    RECT 35.2000 142.2000 36.0000 143.6000 ;
	    RECT 39.6000 142.2000 40.4000 147.0000 ;
	    RECT 41.2000 142.2000 42.0000 147.0000 ;
	    RECT 46.2000 145.6000 46.8000 147.8000 ;
	    RECT 51.8000 147.6000 53.2000 147.8000 ;
	    RECT 58.8000 147.2000 59.6000 150.6000 ;
	    RECT 66.8000 150.3000 67.6000 150.4000 ;
	    RECT 70.0000 150.3000 70.8000 150.4000 ;
	    RECT 66.8000 150.2000 70.8000 150.3000 ;
	    RECT 62.6000 149.7000 70.8000 150.2000 ;
	    RECT 62.6000 149.6000 67.6000 149.7000 ;
	    RECT 70.0000 149.6000 70.8000 149.7000 ;
	    RECT 62.6000 149.4000 63.4000 149.6000 ;
	    RECT 64.2000 148.4000 65.0000 148.6000 ;
	    RECT 71.6000 148.4000 72.2000 151.6000 ;
	    RECT 78.0000 151.2000 78.8000 159.8000 ;
	    RECT 74.6000 150.6000 78.8000 151.2000 ;
	    RECT 74.6000 150.4000 75.4000 150.6000 ;
	    RECT 76.2000 149.8000 77.0000 150.0000 ;
	    RECT 73.2000 149.2000 77.0000 149.8000 ;
	    RECT 73.2000 149.0000 74.0000 149.2000 ;
	    RECT 61.2000 147.8000 72.2000 148.4000 ;
	    RECT 61.2000 147.6000 62.8000 147.8000 ;
	    RECT 55.8000 146.6000 59.6000 147.2000 ;
	    RECT 55.8000 146.4000 56.6000 146.6000 ;
	    RECT 44.4000 144.2000 45.2000 145.0000 ;
	    RECT 46.0000 144.8000 46.8000 145.6000 ;
	    RECT 47.8000 145.4000 48.6000 145.6000 ;
	    RECT 47.8000 144.8000 50.6000 145.4000 ;
	    RECT 50.0000 144.2000 50.6000 144.8000 ;
	    RECT 54.0000 144.2000 54.8000 145.0000 ;
	    RECT 44.4000 143.6000 46.4000 144.2000 ;
	    RECT 45.6000 142.2000 46.4000 143.6000 ;
	    RECT 50.0000 142.2000 50.8000 144.2000 ;
	    RECT 54.0000 143.6000 55.4000 144.2000 ;
	    RECT 54.2000 142.2000 55.4000 143.6000 ;
	    RECT 58.8000 142.2000 59.6000 146.6000 ;
	    RECT 60.4000 142.2000 61.2000 147.0000 ;
	    RECT 65.4000 145.6000 66.0000 147.8000 ;
	    RECT 71.0000 147.6000 71.8000 147.8000 ;
	    RECT 78.0000 147.2000 78.8000 150.6000 ;
	    RECT 75.0000 146.6000 78.8000 147.2000 ;
	    RECT 75.0000 146.4000 75.8000 146.6000 ;
	    RECT 63.6000 144.2000 64.4000 145.0000 ;
	    RECT 65.2000 144.8000 66.0000 145.6000 ;
	    RECT 67.0000 145.4000 67.8000 145.6000 ;
	    RECT 67.0000 144.8000 69.8000 145.4000 ;
	    RECT 69.2000 144.2000 69.8000 144.8000 ;
	    RECT 73.2000 144.2000 74.0000 145.0000 ;
	    RECT 63.6000 143.6000 65.6000 144.2000 ;
	    RECT 64.8000 142.2000 65.6000 143.6000 ;
	    RECT 69.2000 142.2000 70.0000 144.2000 ;
	    RECT 73.2000 143.6000 74.6000 144.2000 ;
	    RECT 73.4000 142.2000 74.6000 143.6000 ;
	    RECT 78.0000 142.2000 78.8000 146.6000 ;
	    RECT 79.6000 151.8000 80.4000 159.8000 ;
	    RECT 82.8000 152.4000 83.6000 159.8000 ;
	    RECT 81.4000 151.8000 83.6000 152.4000 ;
	    RECT 79.6000 149.6000 80.2000 151.8000 ;
	    RECT 81.4000 151.2000 82.0000 151.8000 ;
	    RECT 80.8000 150.4000 82.0000 151.2000 ;
	    RECT 79.6000 142.2000 80.4000 149.6000 ;
	    RECT 81.4000 147.4000 82.0000 150.4000 ;
	    RECT 86.0000 150.3000 86.8000 159.8000 ;
	    RECT 90.0000 153.6000 90.8000 154.4000 ;
	    RECT 87.6000 151.6000 88.4000 153.2000 ;
	    RECT 90.0000 152.4000 90.6000 153.6000 ;
	    RECT 91.4000 152.4000 92.2000 159.8000 ;
	    RECT 89.2000 151.8000 90.6000 152.4000 ;
	    RECT 91.2000 151.8000 92.2000 152.4000 ;
	    RECT 98.2000 152.4000 99.0000 159.8000 ;
	    RECT 99.6000 153.6000 100.4000 154.4000 ;
	    RECT 99.8000 152.4000 100.4000 153.6000 ;
	    RECT 102.8000 153.6000 103.6000 154.4000 ;
	    RECT 102.8000 152.4000 103.4000 153.6000 ;
	    RECT 104.2000 152.4000 105.0000 159.8000 ;
	    RECT 118.6000 152.8000 119.4000 159.8000 ;
	    RECT 122.8000 155.0000 123.6000 159.0000 ;
	    RECT 98.2000 151.8000 99.2000 152.4000 ;
	    RECT 99.8000 151.8000 101.2000 152.4000 ;
	    RECT 89.2000 151.6000 90.0000 151.8000 ;
	    RECT 89.3000 150.3000 89.9000 151.6000 ;
	    RECT 91.2000 150.4000 91.8000 151.8000 ;
	    RECT 98.6000 150.4000 99.2000 151.8000 ;
	    RECT 100.4000 151.6000 101.2000 151.8000 ;
	    RECT 102.0000 151.8000 103.4000 152.4000 ;
	    RECT 104.0000 151.8000 105.0000 152.4000 ;
	    RECT 117.8000 152.2000 119.4000 152.8000 ;
	    RECT 102.0000 151.6000 102.8000 151.8000 ;
	    RECT 86.0000 149.7000 89.9000 150.3000 ;
	    RECT 81.4000 146.8000 83.6000 147.4000 ;
	    RECT 84.4000 146.8000 85.2000 148.4000 ;
	    RECT 82.8000 142.2000 83.6000 146.8000 ;
	    RECT 86.0000 146.2000 86.8000 149.7000 ;
	    RECT 90.8000 149.6000 91.8000 150.4000 ;
	    RECT 91.2000 148.4000 91.8000 149.6000 ;
	    RECT 92.4000 148.8000 93.2000 150.4000 ;
	    RECT 97.2000 148.8000 98.0000 150.4000 ;
	    RECT 98.6000 149.6000 99.6000 150.4000 ;
	    RECT 100.5000 150.3000 101.1000 151.6000 ;
	    RECT 104.0000 150.3000 104.6000 151.8000 ;
	    RECT 100.5000 149.7000 104.6000 150.3000 ;
	    RECT 98.6000 148.4000 99.2000 149.6000 ;
	    RECT 104.0000 148.4000 104.6000 149.7000 ;
	    RECT 105.2000 148.8000 106.0000 150.4000 ;
	    RECT 116.4000 149.6000 117.2000 151.2000 ;
	    RECT 117.8000 148.4000 118.4000 152.2000 ;
	    RECT 123.0000 151.6000 123.6000 155.0000 ;
	    RECT 127.0000 152.6000 127.8000 159.8000 ;
	    RECT 131.8000 152.6000 132.6000 159.8000 ;
	    RECT 136.6000 156.4000 137.4000 159.8000 ;
	    RECT 135.6000 155.6000 137.4000 156.4000 ;
	    RECT 126.0000 151.8000 127.8000 152.6000 ;
	    RECT 130.8000 151.8000 132.6000 152.6000 ;
	    RECT 136.6000 152.4000 137.4000 155.6000 ;
	    RECT 138.0000 153.6000 138.8000 154.4000 ;
	    RECT 138.2000 152.4000 138.8000 153.6000 ;
	    RECT 136.6000 151.8000 137.6000 152.4000 ;
	    RECT 138.2000 151.8000 139.6000 152.4000 ;
	    RECT 119.8000 151.0000 123.6000 151.6000 ;
	    RECT 119.8000 149.0000 120.4000 151.0000 ;
	    RECT 89.2000 147.6000 91.8000 148.4000 ;
	    RECT 94.0000 148.3000 94.8000 148.4000 ;
	    RECT 95.6000 148.3000 96.4000 148.4000 ;
	    RECT 94.0000 148.2000 96.4000 148.3000 ;
	    RECT 93.2000 147.7000 97.2000 148.2000 ;
	    RECT 93.2000 147.6000 94.8000 147.7000 ;
	    RECT 95.6000 147.6000 97.2000 147.7000 ;
	    RECT 98.6000 147.6000 101.2000 148.4000 ;
	    RECT 102.0000 147.6000 104.6000 148.4000 ;
	    RECT 106.8000 148.2000 107.6000 148.4000 ;
	    RECT 106.0000 147.6000 107.6000 148.2000 ;
	    RECT 116.4000 147.6000 118.4000 148.4000 ;
	    RECT 119.0000 148.2000 120.4000 149.0000 ;
	    RECT 121.2000 148.8000 122.0000 150.4000 ;
	    RECT 122.8000 148.8000 123.6000 150.4000 ;
	    RECT 126.2000 148.4000 126.8000 151.8000 ;
	    RECT 130.8000 151.6000 131.6000 151.8000 ;
	    RECT 127.6000 149.6000 128.4000 151.2000 ;
	    RECT 131.0000 148.4000 131.6000 151.6000 ;
	    RECT 132.4000 149.6000 133.2000 151.2000 ;
	    RECT 134.0000 150.3000 134.8000 150.4000 ;
	    RECT 135.6000 150.3000 136.4000 150.4000 ;
	    RECT 134.0000 149.7000 136.4000 150.3000 ;
	    RECT 134.0000 149.6000 134.8000 149.7000 ;
	    RECT 135.6000 148.8000 136.4000 149.7000 ;
	    RECT 137.0000 148.4000 137.6000 151.8000 ;
	    RECT 138.8000 151.6000 139.6000 151.8000 ;
	    RECT 140.4000 151.6000 141.2000 153.2000 ;
	    RECT 138.9000 150.3000 139.5000 151.6000 ;
	    RECT 142.0000 150.3000 142.8000 159.8000 ;
	    RECT 147.8000 152.4000 148.6000 159.8000 ;
	    RECT 154.2000 158.4000 156.2000 159.8000 ;
	    RECT 153.2000 157.6000 156.2000 158.4000 ;
	    RECT 149.2000 153.6000 150.0000 154.4000 ;
	    RECT 149.4000 152.4000 150.0000 153.6000 ;
	    RECT 147.8000 151.8000 148.8000 152.4000 ;
	    RECT 149.4000 151.8000 150.8000 152.4000 ;
	    RECT 154.2000 151.8000 156.2000 157.6000 ;
	    RECT 162.2000 158.4000 163.0000 159.8000 ;
	    RECT 162.2000 157.6000 163.6000 158.4000 ;
	    RECT 162.2000 152.6000 163.0000 157.6000 ;
	    RECT 161.2000 151.8000 163.0000 152.6000 ;
	    RECT 165.0000 152.6000 165.8000 159.8000 ;
	    RECT 165.0000 151.8000 166.8000 152.6000 ;
	    RECT 171.8000 152.4000 172.6000 159.8000 ;
	    RECT 173.2000 153.6000 174.0000 154.4000 ;
	    RECT 173.4000 152.4000 174.0000 153.6000 ;
	    RECT 171.8000 151.8000 172.8000 152.4000 ;
	    RECT 173.4000 151.8000 174.8000 152.4000 ;
	    RECT 178.2000 151.8000 180.2000 159.8000 ;
	    RECT 186.2000 156.4000 187.0000 159.8000 ;
	    RECT 185.2000 155.6000 187.0000 156.4000 ;
	    RECT 186.2000 152.6000 187.0000 155.6000 ;
	    RECT 185.2000 151.8000 187.0000 152.6000 ;
	    RECT 189.2000 153.6000 190.0000 154.4000 ;
	    RECT 189.2000 152.4000 189.8000 153.6000 ;
	    RECT 190.6000 152.4000 191.4000 159.8000 ;
	    RECT 197.0000 158.4000 197.8000 159.8000 ;
	    RECT 197.0000 157.6000 198.8000 158.4000 ;
	    RECT 195.6000 153.6000 196.4000 154.4000 ;
	    RECT 195.6000 152.4000 196.2000 153.6000 ;
	    RECT 197.0000 152.4000 197.8000 157.6000 ;
	    RECT 188.4000 151.8000 189.8000 152.4000 ;
	    RECT 190.4000 151.8000 191.4000 152.4000 ;
	    RECT 194.8000 151.8000 196.2000 152.4000 ;
	    RECT 196.8000 151.8000 197.8000 152.4000 ;
	    RECT 138.9000 149.7000 142.8000 150.3000 ;
	    RECT 89.4000 146.2000 90.0000 147.6000 ;
	    RECT 93.2000 147.2000 94.0000 147.6000 ;
	    RECT 96.4000 147.2000 97.2000 147.6000 ;
	    RECT 91.0000 146.2000 94.6000 146.6000 ;
	    RECT 95.8000 146.2000 99.4000 146.6000 ;
	    RECT 100.4000 146.2000 101.0000 147.6000 ;
	    RECT 102.2000 146.2000 102.8000 147.6000 ;
	    RECT 106.0000 147.2000 106.8000 147.6000 ;
	    RECT 117.8000 147.0000 118.4000 147.6000 ;
	    RECT 119.4000 147.8000 120.4000 148.2000 ;
	    RECT 119.4000 147.2000 123.6000 147.8000 ;
	    RECT 126.0000 147.6000 126.8000 148.4000 ;
	    RECT 130.8000 147.6000 131.6000 148.4000 ;
	    RECT 134.0000 148.2000 134.8000 148.4000 ;
	    RECT 134.0000 147.6000 135.6000 148.2000 ;
	    RECT 137.0000 147.6000 139.6000 148.4000 ;
	    RECT 117.8000 146.6000 118.6000 147.0000 ;
	    RECT 103.8000 146.2000 107.4000 146.6000 ;
	    RECT 86.0000 145.6000 87.8000 146.2000 ;
	    RECT 87.0000 142.2000 87.8000 145.6000 ;
	    RECT 89.2000 142.2000 90.0000 146.2000 ;
	    RECT 90.8000 146.0000 94.8000 146.2000 ;
	    RECT 90.8000 142.2000 91.6000 146.0000 ;
	    RECT 94.0000 142.2000 94.8000 146.0000 ;
	    RECT 95.6000 146.0000 99.6000 146.2000 ;
	    RECT 95.6000 142.2000 96.4000 146.0000 ;
	    RECT 98.8000 142.2000 99.6000 146.0000 ;
	    RECT 100.4000 142.2000 101.2000 146.2000 ;
	    RECT 102.0000 142.2000 102.8000 146.2000 ;
	    RECT 103.6000 146.0000 107.6000 146.2000 ;
	    RECT 117.8000 146.0000 119.4000 146.6000 ;
	    RECT 103.6000 142.2000 104.4000 146.0000 ;
	    RECT 106.8000 142.2000 107.6000 146.0000 ;
	    RECT 118.6000 144.4000 119.4000 146.0000 ;
	    RECT 123.0000 145.0000 123.6000 147.2000 ;
	    RECT 118.6000 143.6000 120.4000 144.4000 ;
	    RECT 118.6000 143.0000 119.4000 143.6000 ;
	    RECT 122.8000 143.0000 123.6000 145.0000 ;
	    RECT 124.4000 144.8000 125.2000 146.4000 ;
	    RECT 126.2000 144.4000 126.8000 147.6000 ;
	    RECT 129.2000 144.8000 130.0000 146.4000 ;
	    RECT 126.0000 142.2000 126.8000 144.4000 ;
	    RECT 131.0000 144.2000 131.6000 147.6000 ;
	    RECT 134.8000 147.2000 135.6000 147.6000 ;
	    RECT 134.2000 146.2000 137.8000 146.6000 ;
	    RECT 138.8000 146.2000 139.4000 147.6000 ;
	    RECT 142.0000 146.2000 142.8000 149.7000 ;
	    RECT 143.6000 150.3000 144.4000 150.4000 ;
	    RECT 146.8000 150.3000 147.6000 150.4000 ;
	    RECT 143.6000 149.7000 147.6000 150.3000 ;
	    RECT 143.6000 149.6000 144.4000 149.7000 ;
	    RECT 143.7000 148.4000 144.3000 149.6000 ;
	    RECT 146.8000 148.8000 147.6000 149.7000 ;
	    RECT 148.2000 148.4000 148.8000 151.8000 ;
	    RECT 150.0000 151.6000 150.8000 151.8000 ;
	    RECT 153.2000 148.8000 154.0000 150.4000 ;
	    RECT 154.8000 148.4000 155.4000 151.8000 ;
	    RECT 156.4000 148.8000 157.2000 150.4000 ;
	    RECT 143.6000 146.8000 144.4000 148.4000 ;
	    RECT 145.2000 148.2000 146.0000 148.4000 ;
	    RECT 148.2000 148.3000 150.8000 148.4000 ;
	    RECT 151.6000 148.3000 152.4000 148.4000 ;
	    RECT 148.2000 148.2000 152.4000 148.3000 ;
	    RECT 154.8000 148.2000 155.6000 148.4000 ;
	    RECT 145.2000 147.6000 146.8000 148.2000 ;
	    RECT 148.2000 147.7000 153.2000 148.2000 ;
	    RECT 148.2000 147.6000 150.8000 147.7000 ;
	    RECT 151.6000 147.6000 153.2000 147.7000 ;
	    RECT 154.8000 147.6000 157.2000 148.2000 ;
	    RECT 158.0000 147.6000 158.8000 149.2000 ;
	    RECT 161.4000 148.4000 162.0000 151.8000 ;
	    RECT 162.8000 149.6000 163.6000 151.2000 ;
	    RECT 164.4000 149.6000 165.2000 151.2000 ;
	    RECT 161.2000 147.6000 162.0000 148.4000 ;
	    RECT 146.0000 147.2000 146.8000 147.6000 ;
	    RECT 145.4000 146.2000 149.0000 146.6000 ;
	    RECT 150.0000 146.2000 150.6000 147.6000 ;
	    RECT 152.4000 147.2000 153.2000 147.6000 ;
	    RECT 151.8000 146.2000 155.4000 146.6000 ;
	    RECT 156.6000 146.2000 157.2000 147.6000 ;
	    RECT 130.8000 142.2000 131.6000 144.2000 ;
	    RECT 134.0000 146.0000 138.0000 146.2000 ;
	    RECT 134.0000 142.2000 134.8000 146.0000 ;
	    RECT 137.2000 142.2000 138.0000 146.0000 ;
	    RECT 138.8000 142.2000 139.6000 146.2000 ;
	    RECT 141.0000 145.6000 142.8000 146.2000 ;
	    RECT 145.2000 146.0000 149.2000 146.2000 ;
	    RECT 141.0000 142.2000 141.8000 145.6000 ;
	    RECT 145.2000 142.2000 146.0000 146.0000 ;
	    RECT 148.4000 142.2000 149.2000 146.0000 ;
	    RECT 150.0000 142.2000 150.8000 146.2000 ;
	    RECT 151.6000 146.0000 155.6000 146.2000 ;
	    RECT 151.6000 142.2000 152.4000 146.0000 ;
	    RECT 154.8000 142.8000 155.6000 146.0000 ;
	    RECT 156.4000 143.4000 157.2000 146.2000 ;
	    RECT 158.0000 142.8000 158.8000 146.2000 ;
	    RECT 159.6000 144.8000 160.4000 146.4000 ;
	    RECT 161.4000 144.2000 162.0000 147.6000 ;
	    RECT 166.0000 148.4000 166.6000 151.8000 ;
	    RECT 170.8000 148.8000 171.6000 150.4000 ;
	    RECT 172.2000 148.4000 172.8000 151.8000 ;
	    RECT 174.0000 151.6000 174.8000 151.8000 ;
	    RECT 175.6000 150.3000 176.4000 150.4000 ;
	    RECT 177.2000 150.3000 178.0000 150.4000 ;
	    RECT 175.6000 149.7000 178.0000 150.3000 ;
	    RECT 175.6000 149.6000 176.4000 149.7000 ;
	    RECT 177.2000 148.8000 178.0000 149.7000 ;
	    RECT 178.8000 148.4000 179.4000 151.8000 ;
	    RECT 180.4000 148.8000 181.2000 150.4000 ;
	    RECT 166.0000 147.6000 166.8000 148.4000 ;
	    RECT 169.2000 148.2000 170.0000 148.4000 ;
	    RECT 172.2000 148.3000 174.8000 148.4000 ;
	    RECT 175.6000 148.3000 176.4000 148.4000 ;
	    RECT 172.2000 148.2000 176.4000 148.3000 ;
	    RECT 178.8000 148.2000 179.6000 148.4000 ;
	    RECT 169.2000 147.6000 170.8000 148.2000 ;
	    RECT 172.2000 147.7000 177.2000 148.2000 ;
	    RECT 172.2000 147.6000 174.8000 147.7000 ;
	    RECT 175.6000 147.6000 177.2000 147.7000 ;
	    RECT 178.8000 147.6000 181.2000 148.2000 ;
	    RECT 182.0000 147.6000 182.8000 149.2000 ;
	    RECT 185.4000 148.4000 186.0000 151.8000 ;
	    RECT 188.4000 151.6000 189.2000 151.8000 ;
	    RECT 186.8000 150.3000 187.6000 151.2000 ;
	    RECT 190.4000 150.4000 191.0000 151.8000 ;
	    RECT 194.8000 151.6000 195.6000 151.8000 ;
	    RECT 188.4000 150.3000 189.2000 150.4000 ;
	    RECT 186.8000 149.7000 189.2000 150.3000 ;
	    RECT 186.8000 149.6000 187.6000 149.7000 ;
	    RECT 188.4000 149.6000 189.2000 149.7000 ;
	    RECT 190.0000 149.6000 191.0000 150.4000 ;
	    RECT 190.4000 148.4000 191.0000 149.6000 ;
	    RECT 191.6000 148.8000 192.4000 150.4000 ;
	    RECT 196.8000 148.4000 197.4000 151.8000 ;
	    RECT 201.2000 151.2000 202.0000 159.8000 ;
	    RECT 205.4000 155.8000 206.6000 159.8000 ;
	    RECT 210.0000 155.8000 210.8000 159.8000 ;
	    RECT 214.4000 156.4000 215.2000 159.8000 ;
	    RECT 214.4000 155.8000 216.4000 156.4000 ;
	    RECT 206.0000 155.0000 206.8000 155.8000 ;
	    RECT 210.2000 155.2000 210.8000 155.8000 ;
	    RECT 209.4000 154.6000 213.0000 155.2000 ;
	    RECT 215.6000 155.0000 216.4000 155.8000 ;
	    RECT 209.4000 154.4000 210.2000 154.6000 ;
	    RECT 212.2000 154.4000 213.0000 154.6000 ;
	    RECT 205.2000 153.2000 206.6000 154.0000 ;
	    RECT 206.0000 152.2000 206.6000 153.2000 ;
	    RECT 208.2000 153.0000 210.4000 153.6000 ;
	    RECT 208.2000 152.8000 209.0000 153.0000 ;
	    RECT 206.0000 151.6000 208.4000 152.2000 ;
	    RECT 201.2000 150.6000 205.4000 151.2000 ;
	    RECT 198.0000 148.8000 198.8000 150.4000 ;
	    RECT 185.2000 147.6000 186.0000 148.4000 ;
	    RECT 188.4000 147.6000 191.0000 148.4000 ;
	    RECT 193.2000 148.2000 194.0000 148.4000 ;
	    RECT 192.4000 147.6000 194.0000 148.2000 ;
	    RECT 194.8000 147.6000 197.4000 148.4000 ;
	    RECT 199.6000 148.2000 200.4000 148.4000 ;
	    RECT 198.8000 147.6000 200.4000 148.2000 ;
	    RECT 162.8000 146.3000 163.6000 146.4000 ;
	    RECT 166.0000 146.3000 166.6000 147.6000 ;
	    RECT 170.0000 147.2000 170.8000 147.6000 ;
	    RECT 162.8000 145.7000 166.7000 146.3000 ;
	    RECT 162.8000 145.6000 163.6000 145.7000 ;
	    RECT 154.8000 142.2000 158.8000 142.8000 ;
	    RECT 161.2000 142.2000 162.0000 144.2000 ;
	    RECT 166.0000 144.2000 166.6000 145.7000 ;
	    RECT 167.6000 144.8000 168.4000 146.4000 ;
	    RECT 169.4000 146.2000 173.0000 146.6000 ;
	    RECT 174.0000 146.2000 174.6000 147.6000 ;
	    RECT 176.4000 147.2000 177.2000 147.6000 ;
	    RECT 175.8000 146.2000 179.4000 146.6000 ;
	    RECT 180.6000 146.2000 181.2000 147.6000 ;
	    RECT 169.2000 146.0000 173.2000 146.2000 ;
	    RECT 166.0000 142.2000 166.8000 144.2000 ;
	    RECT 169.2000 142.2000 170.0000 146.0000 ;
	    RECT 172.4000 142.2000 173.2000 146.0000 ;
	    RECT 174.0000 142.2000 174.8000 146.2000 ;
	    RECT 175.6000 146.0000 179.6000 146.2000 ;
	    RECT 175.6000 142.2000 176.4000 146.0000 ;
	    RECT 178.8000 142.8000 179.6000 146.0000 ;
	    RECT 180.4000 143.4000 181.2000 146.2000 ;
	    RECT 182.0000 142.8000 182.8000 146.2000 ;
	    RECT 183.6000 144.8000 184.4000 146.4000 ;
	    RECT 185.4000 144.2000 186.0000 147.6000 ;
	    RECT 188.6000 146.2000 189.2000 147.6000 ;
	    RECT 192.4000 147.2000 193.2000 147.6000 ;
	    RECT 190.2000 146.2000 193.8000 146.6000 ;
	    RECT 195.0000 146.2000 195.6000 147.6000 ;
	    RECT 198.8000 147.2000 199.6000 147.6000 ;
	    RECT 201.2000 147.2000 202.0000 150.6000 ;
	    RECT 204.6000 150.4000 205.4000 150.6000 ;
	    RECT 203.0000 149.8000 203.8000 150.0000 ;
	    RECT 203.0000 149.2000 206.8000 149.8000 ;
	    RECT 206.0000 149.0000 206.8000 149.2000 ;
	    RECT 207.8000 148.4000 208.4000 151.6000 ;
	    RECT 209.8000 151.8000 210.4000 153.0000 ;
	    RECT 211.0000 153.0000 211.8000 153.2000 ;
	    RECT 215.6000 153.0000 216.4000 153.2000 ;
	    RECT 211.0000 152.4000 216.4000 153.0000 ;
	    RECT 209.8000 151.4000 214.6000 151.8000 ;
	    RECT 218.8000 151.4000 219.6000 159.8000 ;
	    RECT 220.4000 152.4000 221.2000 159.8000 ;
	    RECT 220.4000 151.8000 222.6000 152.4000 ;
	    RECT 223.6000 151.8000 224.4000 159.8000 ;
	    RECT 227.8000 152.6000 228.6000 159.8000 ;
	    RECT 226.8000 151.8000 228.6000 152.6000 ;
	    RECT 230.0000 152.4000 230.8000 159.8000 ;
	    RECT 230.0000 151.8000 232.2000 152.4000 ;
	    RECT 233.2000 151.8000 234.0000 159.8000 ;
	    RECT 209.8000 151.2000 219.6000 151.4000 ;
	    RECT 213.8000 151.0000 219.6000 151.2000 ;
	    RECT 214.0000 150.8000 219.6000 151.0000 ;
	    RECT 222.0000 151.2000 222.6000 151.8000 ;
	    RECT 222.0000 150.4000 223.2000 151.2000 ;
	    RECT 212.4000 150.2000 213.2000 150.4000 ;
	    RECT 212.4000 149.6000 217.4000 150.2000 ;
	    RECT 216.6000 149.4000 217.4000 149.6000 ;
	    RECT 215.0000 148.4000 215.8000 148.6000 ;
	    RECT 207.8000 147.8000 218.8000 148.4000 ;
	    RECT 208.2000 147.6000 209.0000 147.8000 ;
	    RECT 201.2000 146.6000 205.0000 147.2000 ;
	    RECT 196.6000 146.2000 200.2000 146.6000 ;
	    RECT 178.8000 142.2000 182.8000 142.8000 ;
	    RECT 185.2000 142.2000 186.0000 144.2000 ;
	    RECT 188.4000 142.2000 189.2000 146.2000 ;
	    RECT 190.0000 146.0000 194.0000 146.2000 ;
	    RECT 190.0000 142.2000 190.8000 146.0000 ;
	    RECT 193.2000 142.2000 194.0000 146.0000 ;
	    RECT 194.8000 142.2000 195.6000 146.2000 ;
	    RECT 196.4000 146.0000 200.4000 146.2000 ;
	    RECT 196.4000 142.2000 197.2000 146.0000 ;
	    RECT 199.6000 142.2000 200.4000 146.0000 ;
	    RECT 201.2000 142.2000 202.0000 146.6000 ;
	    RECT 204.2000 146.4000 205.0000 146.6000 ;
	    RECT 214.0000 145.6000 214.6000 147.8000 ;
	    RECT 217.2000 147.6000 218.8000 147.8000 ;
	    RECT 222.0000 147.4000 222.6000 150.4000 ;
	    RECT 223.8000 149.6000 224.4000 151.8000 ;
	    RECT 212.2000 145.4000 213.0000 145.6000 ;
	    RECT 206.0000 144.2000 206.8000 145.0000 ;
	    RECT 210.2000 144.8000 213.0000 145.4000 ;
	    RECT 214.0000 144.8000 214.8000 145.6000 ;
	    RECT 210.2000 144.2000 210.8000 144.8000 ;
	    RECT 215.6000 144.2000 216.4000 145.0000 ;
	    RECT 205.4000 143.6000 206.8000 144.2000 ;
	    RECT 205.4000 142.2000 206.6000 143.6000 ;
	    RECT 210.0000 142.2000 210.8000 144.2000 ;
	    RECT 214.4000 143.6000 216.4000 144.2000 ;
	    RECT 214.4000 142.2000 215.2000 143.6000 ;
	    RECT 218.8000 142.2000 219.6000 147.0000 ;
	    RECT 220.4000 146.8000 222.6000 147.4000 ;
	    RECT 220.4000 142.2000 221.2000 146.8000 ;
	    RECT 223.6000 142.2000 224.4000 149.6000 ;
	    RECT 227.0000 148.4000 227.6000 151.8000 ;
	    RECT 231.6000 151.2000 232.2000 151.8000 ;
	    RECT 228.4000 149.6000 229.2000 151.2000 ;
	    RECT 231.6000 150.4000 232.8000 151.2000 ;
	    RECT 226.8000 147.6000 227.6000 148.4000 ;
	    RECT 225.2000 144.8000 226.0000 146.4000 ;
	    RECT 227.0000 144.4000 227.6000 147.6000 ;
	    RECT 231.6000 147.4000 232.2000 150.4000 ;
	    RECT 233.4000 149.6000 234.0000 151.8000 ;
	    RECT 234.8000 151.4000 235.6000 159.8000 ;
	    RECT 239.2000 156.4000 240.0000 159.8000 ;
	    RECT 238.0000 155.8000 240.0000 156.4000 ;
	    RECT 243.6000 155.8000 244.4000 159.8000 ;
	    RECT 247.8000 155.8000 249.0000 159.8000 ;
	    RECT 238.0000 155.0000 238.8000 155.8000 ;
	    RECT 243.6000 155.2000 244.2000 155.8000 ;
	    RECT 241.4000 154.6000 245.0000 155.2000 ;
	    RECT 247.6000 155.0000 248.4000 155.8000 ;
	    RECT 241.4000 154.4000 242.2000 154.6000 ;
	    RECT 244.2000 154.4000 245.0000 154.6000 ;
	    RECT 238.0000 153.0000 238.8000 153.2000 ;
	    RECT 242.6000 153.0000 243.4000 153.2000 ;
	    RECT 238.0000 152.4000 243.4000 153.0000 ;
	    RECT 244.0000 153.0000 246.2000 153.6000 ;
	    RECT 244.0000 151.8000 244.6000 153.0000 ;
	    RECT 245.4000 152.8000 246.2000 153.0000 ;
	    RECT 247.8000 153.2000 249.2000 154.0000 ;
	    RECT 247.8000 152.2000 248.4000 153.2000 ;
	    RECT 239.8000 151.4000 244.6000 151.8000 ;
	    RECT 234.8000 151.2000 244.6000 151.4000 ;
	    RECT 246.0000 151.6000 248.4000 152.2000 ;
	    RECT 234.8000 151.0000 240.6000 151.2000 ;
	    RECT 234.8000 150.8000 240.4000 151.0000 ;
	    RECT 246.0000 150.4000 246.6000 151.6000 ;
	    RECT 252.4000 151.2000 253.2000 159.8000 ;
	    RECT 254.0000 158.3000 254.8000 158.4000 ;
	    RECT 260.4000 158.3000 261.2000 159.8000 ;
	    RECT 254.0000 157.7000 261.2000 158.3000 ;
	    RECT 254.0000 157.6000 254.8000 157.7000 ;
	    RECT 258.8000 154.3000 259.6000 154.4000 ;
	    RECT 260.4000 154.3000 261.2000 157.7000 ;
	    RECT 258.8000 153.7000 261.2000 154.3000 ;
	    RECT 258.8000 153.6000 259.6000 153.7000 ;
	    RECT 249.0000 150.6000 253.2000 151.2000 ;
	    RECT 249.0000 150.4000 249.8000 150.6000 ;
	    RECT 241.2000 150.3000 242.0000 150.4000 ;
	    RECT 242.8000 150.3000 243.6000 150.4000 ;
	    RECT 241.2000 150.2000 243.6000 150.3000 ;
	    RECT 226.8000 142.2000 227.6000 144.4000 ;
	    RECT 230.0000 146.8000 232.2000 147.4000 ;
	    RECT 230.0000 142.2000 230.8000 146.8000 ;
	    RECT 233.2000 142.2000 234.0000 149.6000 ;
	    RECT 237.0000 149.7000 243.6000 150.2000 ;
	    RECT 237.0000 149.6000 242.0000 149.7000 ;
	    RECT 242.8000 149.6000 243.6000 149.7000 ;
	    RECT 246.0000 149.6000 246.8000 150.4000 ;
	    RECT 250.6000 149.8000 251.4000 150.0000 ;
	    RECT 237.0000 149.4000 237.8000 149.6000 ;
	    RECT 238.6000 148.4000 239.4000 148.6000 ;
	    RECT 246.0000 148.4000 246.6000 149.6000 ;
	    RECT 247.6000 149.2000 251.4000 149.8000 ;
	    RECT 247.6000 149.0000 248.4000 149.2000 ;
	    RECT 235.6000 147.8000 246.6000 148.4000 ;
	    RECT 235.6000 147.6000 237.2000 147.8000 ;
	    RECT 234.8000 142.2000 235.6000 147.0000 ;
	    RECT 239.8000 145.6000 240.4000 147.8000 ;
	    RECT 245.4000 147.6000 246.2000 147.8000 ;
	    RECT 252.4000 147.2000 253.2000 150.6000 ;
	    RECT 249.4000 146.6000 253.2000 147.2000 ;
	    RECT 249.4000 146.4000 250.2000 146.6000 ;
	    RECT 238.0000 144.2000 238.8000 145.0000 ;
	    RECT 239.6000 144.8000 240.4000 145.6000 ;
	    RECT 241.4000 145.4000 242.2000 145.6000 ;
	    RECT 241.4000 144.8000 244.2000 145.4000 ;
	    RECT 243.6000 144.2000 244.2000 144.8000 ;
	    RECT 247.6000 144.2000 248.4000 145.0000 ;
	    RECT 238.0000 143.6000 240.0000 144.2000 ;
	    RECT 239.2000 142.2000 240.0000 143.6000 ;
	    RECT 243.6000 142.2000 244.4000 144.2000 ;
	    RECT 247.6000 143.6000 249.0000 144.2000 ;
	    RECT 247.8000 142.2000 249.0000 143.6000 ;
	    RECT 252.4000 142.2000 253.2000 146.6000 ;
	    RECT 260.4000 151.8000 261.2000 153.7000 ;
	    RECT 263.6000 152.4000 264.4000 159.8000 ;
	    RECT 262.2000 151.8000 264.4000 152.4000 ;
	    RECT 267.8000 152.4000 268.6000 159.8000 ;
	    RECT 269.2000 153.6000 270.8000 154.4000 ;
	    RECT 269.4000 152.4000 270.0000 153.6000 ;
	    RECT 267.8000 151.8000 268.8000 152.4000 ;
	    RECT 269.4000 151.8000 270.8000 152.4000 ;
	    RECT 260.4000 149.6000 261.0000 151.8000 ;
	    RECT 262.2000 151.2000 262.8000 151.8000 ;
	    RECT 261.6000 150.4000 262.8000 151.2000 ;
	    RECT 260.4000 142.2000 261.2000 149.6000 ;
	    RECT 262.2000 147.4000 262.8000 150.4000 ;
	    RECT 263.6000 150.3000 264.4000 150.4000 ;
	    RECT 265.2000 150.3000 266.0000 150.4000 ;
	    RECT 263.6000 149.7000 266.0000 150.3000 ;
	    RECT 263.6000 148.8000 264.4000 149.7000 ;
	    RECT 265.2000 149.6000 266.0000 149.7000 ;
	    RECT 266.8000 148.8000 267.6000 150.4000 ;
	    RECT 268.2000 150.3000 268.8000 151.8000 ;
	    RECT 270.0000 151.6000 270.8000 151.8000 ;
	    RECT 271.6000 151.8000 272.4000 159.8000 ;
	    RECT 274.8000 152.4000 275.6000 159.8000 ;
	    RECT 278.6000 158.4000 279.4000 159.8000 ;
	    RECT 278.6000 157.6000 280.4000 158.4000 ;
	    RECT 277.2000 153.6000 278.0000 154.4000 ;
	    RECT 277.2000 152.4000 277.8000 153.6000 ;
	    RECT 278.6000 152.4000 279.4000 157.6000 ;
	    RECT 273.4000 151.8000 275.6000 152.4000 ;
	    RECT 276.4000 151.8000 277.8000 152.4000 ;
	    RECT 278.4000 151.8000 279.4000 152.4000 ;
	    RECT 282.8000 152.4000 283.6000 159.8000 ;
	    RECT 282.8000 151.8000 285.0000 152.4000 ;
	    RECT 286.0000 151.8000 286.8000 159.8000 ;
	    RECT 288.2000 152.6000 289.0000 159.8000 ;
	    RECT 295.0000 156.4000 297.0000 159.8000 ;
	    RECT 294.0000 155.6000 297.0000 156.4000 ;
	    RECT 288.2000 151.8000 290.0000 152.6000 ;
	    RECT 295.0000 151.8000 297.0000 155.6000 ;
	    RECT 301.2000 153.6000 302.0000 154.4000 ;
	    RECT 301.2000 152.4000 301.8000 153.6000 ;
	    RECT 302.6000 152.4000 303.4000 159.8000 ;
	    RECT 309.0000 154.4000 309.8000 159.8000 ;
	    RECT 307.6000 153.6000 308.4000 154.4000 ;
	    RECT 309.0000 153.6000 310.8000 154.4000 ;
	    RECT 307.6000 152.4000 308.2000 153.6000 ;
	    RECT 309.0000 152.4000 309.8000 153.6000 ;
	    RECT 300.4000 151.8000 301.8000 152.4000 ;
	    RECT 302.4000 151.8000 303.4000 152.4000 ;
	    RECT 306.8000 151.8000 308.2000 152.4000 ;
	    RECT 308.8000 151.8000 309.8000 152.4000 ;
	    RECT 315.8000 151.8000 317.8000 159.8000 ;
	    RECT 321.8000 152.6000 322.6000 159.8000 ;
	    RECT 328.6000 156.4000 330.6000 159.8000 ;
	    RECT 327.6000 155.6000 330.6000 156.4000 ;
	    RECT 321.8000 151.8000 323.6000 152.6000 ;
	    RECT 328.6000 151.8000 330.6000 155.6000 ;
	    RECT 334.8000 153.6000 335.6000 154.4000 ;
	    RECT 334.8000 152.4000 335.4000 153.6000 ;
	    RECT 336.2000 152.4000 337.0000 159.8000 ;
	    RECT 343.0000 154.4000 343.8000 159.8000 ;
	    RECT 343.0000 153.6000 344.4000 154.4000 ;
	    RECT 343.0000 152.6000 343.8000 153.6000 ;
	    RECT 334.0000 151.8000 335.4000 152.4000 ;
	    RECT 336.0000 151.8000 337.0000 152.4000 ;
	    RECT 342.0000 151.8000 343.8000 152.6000 ;
	    RECT 347.8000 152.4000 349.8000 159.8000 ;
	    RECT 354.0000 153.6000 354.8000 154.4000 ;
	    RECT 354.0000 152.4000 354.6000 153.6000 ;
	    RECT 355.4000 152.4000 356.2000 159.8000 ;
	    RECT 346.8000 151.8000 349.8000 152.4000 ;
	    RECT 353.2000 151.8000 354.6000 152.4000 ;
	    RECT 355.2000 151.8000 356.2000 152.4000 ;
	    RECT 362.2000 152.4000 363.0000 159.8000 ;
	    RECT 363.6000 154.3000 364.4000 154.4000 ;
	    RECT 366.0000 154.3000 366.8000 154.4000 ;
	    RECT 363.6000 153.7000 366.8000 154.3000 ;
	    RECT 363.6000 153.6000 364.4000 153.7000 ;
	    RECT 366.0000 153.6000 366.8000 153.7000 ;
	    RECT 363.8000 152.4000 364.4000 153.6000 ;
	    RECT 362.2000 151.8000 363.2000 152.4000 ;
	    RECT 363.8000 151.8000 365.2000 152.4000 ;
	    RECT 270.0000 150.3000 270.8000 150.4000 ;
	    RECT 268.2000 149.7000 270.8000 150.3000 ;
	    RECT 268.2000 148.4000 268.8000 149.7000 ;
	    RECT 270.0000 149.6000 270.8000 149.7000 ;
	    RECT 271.6000 149.6000 272.2000 151.8000 ;
	    RECT 273.4000 151.2000 274.0000 151.8000 ;
	    RECT 276.4000 151.6000 277.2000 151.8000 ;
	    RECT 272.8000 150.4000 274.0000 151.2000 ;
	    RECT 265.2000 148.2000 266.0000 148.4000 ;
	    RECT 265.2000 147.6000 266.8000 148.2000 ;
	    RECT 268.2000 147.6000 270.8000 148.4000 ;
	    RECT 262.2000 146.8000 264.4000 147.4000 ;
	    RECT 266.0000 147.2000 266.8000 147.6000 ;
	    RECT 263.6000 142.2000 264.4000 146.8000 ;
	    RECT 265.4000 146.2000 269.0000 146.6000 ;
	    RECT 270.0000 146.2000 270.6000 147.6000 ;
	    RECT 265.2000 146.0000 269.2000 146.2000 ;
	    RECT 265.2000 142.2000 266.0000 146.0000 ;
	    RECT 268.4000 142.2000 269.2000 146.0000 ;
	    RECT 270.0000 142.2000 270.8000 146.2000 ;
	    RECT 271.6000 142.2000 272.4000 149.6000 ;
	    RECT 273.4000 147.4000 274.0000 150.4000 ;
	    RECT 274.8000 148.8000 275.6000 150.4000 ;
	    RECT 278.4000 148.4000 279.0000 151.8000 ;
	    RECT 284.4000 151.2000 285.0000 151.8000 ;
	    RECT 284.4000 150.4000 285.6000 151.2000 ;
	    RECT 279.6000 148.8000 280.4000 150.4000 ;
	    RECT 276.4000 147.6000 279.0000 148.4000 ;
	    RECT 281.2000 148.2000 282.0000 148.4000 ;
	    RECT 280.4000 147.6000 282.0000 148.2000 ;
	    RECT 273.4000 146.8000 275.6000 147.4000 ;
	    RECT 274.8000 142.2000 275.6000 146.8000 ;
	    RECT 276.6000 146.2000 277.2000 147.6000 ;
	    RECT 280.4000 147.2000 281.2000 147.6000 ;
	    RECT 284.4000 147.4000 285.0000 150.4000 ;
	    RECT 286.2000 149.6000 286.8000 151.8000 ;
	    RECT 287.6000 149.6000 288.4000 151.2000 ;
	    RECT 289.2000 150.3000 289.8000 151.8000 ;
	    RECT 294.0000 150.3000 294.8000 150.4000 ;
	    RECT 289.2000 149.7000 294.8000 150.3000 ;
	    RECT 282.8000 146.8000 285.0000 147.4000 ;
	    RECT 286.0000 148.3000 286.8000 149.6000 ;
	    RECT 289.2000 148.4000 289.8000 149.7000 ;
	    RECT 294.0000 148.8000 294.8000 149.7000 ;
	    RECT 295.6000 148.4000 296.2000 151.8000 ;
	    RECT 300.4000 151.6000 301.2000 151.8000 ;
	    RECT 297.2000 148.8000 298.0000 150.4000 ;
	    RECT 300.5000 150.3000 301.1000 151.6000 ;
	    RECT 298.8000 149.7000 301.1000 150.3000 ;
	    RECT 287.6000 148.3000 288.4000 148.4000 ;
	    RECT 286.0000 147.7000 288.4000 148.3000 ;
	    RECT 278.2000 146.2000 281.8000 146.6000 ;
	    RECT 276.4000 142.2000 277.2000 146.2000 ;
	    RECT 278.0000 146.0000 282.0000 146.2000 ;
	    RECT 278.0000 142.2000 278.8000 146.0000 ;
	    RECT 281.2000 142.2000 282.0000 146.0000 ;
	    RECT 282.8000 142.2000 283.6000 146.8000 ;
	    RECT 286.0000 142.2000 286.8000 147.7000 ;
	    RECT 287.6000 147.6000 288.4000 147.7000 ;
	    RECT 289.2000 147.6000 290.0000 148.4000 ;
	    RECT 292.4000 148.2000 293.2000 148.4000 ;
	    RECT 295.6000 148.2000 296.4000 148.4000 ;
	    RECT 292.4000 147.6000 294.0000 148.2000 ;
	    RECT 295.6000 147.6000 298.0000 148.2000 ;
	    RECT 298.8000 147.6000 299.6000 149.7000 ;
	    RECT 302.4000 148.4000 303.0000 151.8000 ;
	    RECT 306.8000 151.6000 307.6000 151.8000 ;
	    RECT 303.6000 150.3000 304.4000 150.4000 ;
	    RECT 305.2000 150.3000 306.0000 150.4000 ;
	    RECT 303.6000 149.7000 306.0000 150.3000 ;
	    RECT 303.6000 148.8000 304.4000 149.7000 ;
	    RECT 305.2000 149.6000 306.0000 149.7000 ;
	    RECT 308.8000 148.4000 309.4000 151.8000 ;
	    RECT 310.0000 148.8000 310.8000 150.4000 ;
	    RECT 314.8000 148.8000 315.6000 150.4000 ;
	    RECT 316.4000 148.4000 317.0000 151.8000 ;
	    RECT 318.0000 148.8000 318.8000 150.4000 ;
	    RECT 321.2000 149.6000 322.0000 151.2000 ;
	    RECT 322.8000 150.3000 323.4000 151.8000 ;
	    RECT 327.6000 150.3000 328.4000 150.4000 ;
	    RECT 322.8000 149.7000 328.4000 150.3000 ;
	    RECT 300.4000 147.6000 303.0000 148.4000 ;
	    RECT 305.2000 148.2000 306.0000 148.4000 ;
	    RECT 304.4000 147.6000 306.0000 148.2000 ;
	    RECT 306.8000 147.6000 309.4000 148.4000 ;
	    RECT 311.6000 148.2000 312.4000 148.4000 ;
	    RECT 310.8000 147.6000 312.4000 148.2000 ;
	    RECT 313.2000 148.2000 314.0000 148.4000 ;
	    RECT 316.4000 148.2000 317.2000 148.4000 ;
	    RECT 313.2000 147.6000 314.8000 148.2000 ;
	    RECT 316.4000 147.6000 318.8000 148.2000 ;
	    RECT 319.6000 147.6000 320.4000 149.2000 ;
	    RECT 322.8000 148.4000 323.4000 149.7000 ;
	    RECT 327.6000 148.8000 328.4000 149.7000 ;
	    RECT 329.2000 148.4000 329.8000 151.8000 ;
	    RECT 334.0000 151.6000 334.8000 151.8000 ;
	    RECT 330.8000 148.8000 331.6000 150.4000 ;
	    RECT 334.1000 150.3000 334.7000 151.6000 ;
	    RECT 332.4000 149.7000 334.7000 150.3000 ;
	    RECT 322.8000 147.6000 323.6000 148.4000 ;
	    RECT 326.0000 148.2000 326.8000 148.4000 ;
	    RECT 329.2000 148.2000 330.0000 148.4000 ;
	    RECT 326.0000 147.6000 327.6000 148.2000 ;
	    RECT 329.2000 147.6000 331.6000 148.2000 ;
	    RECT 332.4000 147.6000 333.2000 149.7000 ;
	    RECT 336.0000 148.4000 336.6000 151.8000 ;
	    RECT 337.2000 148.8000 338.0000 150.4000 ;
	    RECT 342.2000 148.4000 342.8000 151.8000 ;
	    RECT 346.8000 151.6000 349.0000 151.8000 ;
	    RECT 353.2000 151.6000 354.0000 151.8000 ;
	    RECT 343.6000 149.6000 344.4000 151.2000 ;
	    RECT 345.2000 150.3000 346.0000 150.4000 ;
	    RECT 346.8000 150.3000 347.6000 150.4000 ;
	    RECT 345.2000 149.7000 347.6000 150.3000 ;
	    RECT 345.2000 149.6000 346.0000 149.7000 ;
	    RECT 346.8000 148.8000 347.6000 149.7000 ;
	    RECT 348.4000 148.4000 349.0000 151.6000 ;
	    RECT 350.0000 148.8000 350.8000 150.4000 ;
	    RECT 353.3000 150.3000 353.9000 151.6000 ;
	    RECT 351.6000 149.7000 353.9000 150.3000 ;
	    RECT 334.0000 147.6000 336.6000 148.4000 ;
	    RECT 338.8000 148.2000 339.6000 148.4000 ;
	    RECT 338.0000 147.6000 339.6000 148.2000 ;
	    RECT 342.0000 147.6000 342.8000 148.4000 ;
	    RECT 345.2000 148.2000 346.0000 148.4000 ;
	    RECT 348.4000 148.2000 349.2000 148.4000 ;
	    RECT 345.2000 147.6000 346.8000 148.2000 ;
	    RECT 348.4000 147.6000 350.8000 148.2000 ;
	    RECT 351.6000 147.6000 352.4000 149.7000 ;
	    RECT 355.2000 148.4000 355.8000 151.8000 ;
	    RECT 362.6000 150.4000 363.2000 151.8000 ;
	    RECT 364.4000 151.6000 365.2000 151.8000 ;
	    RECT 356.4000 148.8000 357.2000 150.4000 ;
	    RECT 361.2000 148.8000 362.0000 150.4000 ;
	    RECT 362.6000 149.6000 363.6000 150.4000 ;
	    RECT 367.6000 150.3000 368.4000 159.8000 ;
	    RECT 371.6000 153.6000 372.4000 154.4000 ;
	    RECT 369.2000 151.6000 370.0000 153.2000 ;
	    RECT 371.6000 152.4000 372.2000 153.6000 ;
	    RECT 373.0000 152.4000 373.8000 159.8000 ;
	    RECT 370.8000 151.8000 372.2000 152.4000 ;
	    RECT 372.8000 151.8000 373.8000 152.4000 ;
	    RECT 370.8000 151.6000 371.6000 151.8000 ;
	    RECT 370.9000 150.3000 371.5000 151.6000 ;
	    RECT 372.8000 150.4000 373.4000 151.8000 ;
	    RECT 377.2000 151.2000 378.0000 159.8000 ;
	    RECT 381.4000 155.8000 382.6000 159.8000 ;
	    RECT 386.0000 155.8000 386.8000 159.8000 ;
	    RECT 390.4000 156.4000 391.2000 159.8000 ;
	    RECT 390.4000 155.8000 392.4000 156.4000 ;
	    RECT 382.0000 155.0000 382.8000 155.8000 ;
	    RECT 386.2000 155.2000 386.8000 155.8000 ;
	    RECT 385.4000 154.6000 389.0000 155.2000 ;
	    RECT 391.6000 155.0000 392.4000 155.8000 ;
	    RECT 385.4000 154.4000 386.2000 154.6000 ;
	    RECT 388.2000 154.4000 389.0000 154.6000 ;
	    RECT 381.2000 153.2000 382.6000 154.0000 ;
	    RECT 382.0000 152.2000 382.6000 153.2000 ;
	    RECT 384.2000 153.0000 386.4000 153.6000 ;
	    RECT 384.2000 152.8000 385.0000 153.0000 ;
	    RECT 382.0000 151.6000 384.4000 152.2000 ;
	    RECT 377.2000 150.6000 381.4000 151.2000 ;
	    RECT 367.6000 149.7000 371.5000 150.3000 ;
	    RECT 362.6000 148.4000 363.2000 149.6000 ;
	    RECT 353.2000 147.6000 355.8000 148.4000 ;
	    RECT 358.0000 148.2000 358.8000 148.4000 ;
	    RECT 357.2000 147.6000 358.8000 148.2000 ;
	    RECT 359.6000 148.2000 360.4000 148.4000 ;
	    RECT 359.6000 147.6000 361.2000 148.2000 ;
	    RECT 362.6000 147.6000 365.2000 148.4000 ;
	    RECT 289.2000 144.2000 289.8000 147.6000 ;
	    RECT 293.2000 147.2000 294.0000 147.6000 ;
	    RECT 290.8000 144.8000 291.6000 146.4000 ;
	    RECT 292.6000 146.2000 296.2000 146.6000 ;
	    RECT 297.4000 146.2000 298.0000 147.6000 ;
	    RECT 300.6000 146.2000 301.2000 147.6000 ;
	    RECT 304.4000 147.2000 305.2000 147.6000 ;
	    RECT 302.2000 146.2000 305.8000 146.6000 ;
	    RECT 307.0000 146.2000 307.6000 147.6000 ;
	    RECT 310.8000 147.2000 311.6000 147.6000 ;
	    RECT 314.0000 147.2000 314.8000 147.6000 ;
	    RECT 308.6000 146.2000 312.2000 146.6000 ;
	    RECT 313.4000 146.2000 317.0000 146.6000 ;
	    RECT 318.2000 146.2000 318.8000 147.6000 ;
	    RECT 292.4000 146.0000 296.4000 146.2000 ;
	    RECT 289.2000 142.2000 290.0000 144.2000 ;
	    RECT 292.4000 142.2000 293.2000 146.0000 ;
	    RECT 295.6000 142.8000 296.4000 146.0000 ;
	    RECT 297.2000 143.4000 298.0000 146.2000 ;
	    RECT 298.8000 142.8000 299.6000 146.2000 ;
	    RECT 295.6000 142.2000 299.6000 142.8000 ;
	    RECT 300.4000 142.2000 301.2000 146.2000 ;
	    RECT 302.0000 146.0000 306.0000 146.2000 ;
	    RECT 302.0000 142.2000 302.8000 146.0000 ;
	    RECT 305.2000 142.2000 306.0000 146.0000 ;
	    RECT 306.8000 142.2000 307.6000 146.2000 ;
	    RECT 308.4000 146.0000 312.4000 146.2000 ;
	    RECT 308.4000 142.2000 309.2000 146.0000 ;
	    RECT 311.6000 142.2000 312.4000 146.0000 ;
	    RECT 313.2000 146.0000 317.2000 146.2000 ;
	    RECT 313.2000 142.2000 314.0000 146.0000 ;
	    RECT 316.4000 142.8000 317.2000 146.0000 ;
	    RECT 318.0000 143.4000 318.8000 146.2000 ;
	    RECT 319.6000 142.8000 320.4000 146.2000 ;
	    RECT 316.4000 142.2000 320.4000 142.8000 ;
	    RECT 322.8000 144.2000 323.4000 147.6000 ;
	    RECT 326.8000 147.2000 327.6000 147.6000 ;
	    RECT 324.4000 144.8000 325.2000 146.4000 ;
	    RECT 326.2000 146.2000 329.8000 146.6000 ;
	    RECT 331.0000 146.2000 331.6000 147.6000 ;
	    RECT 334.2000 146.2000 334.8000 147.6000 ;
	    RECT 338.0000 147.2000 338.8000 147.6000 ;
	    RECT 335.8000 146.2000 339.4000 146.6000 ;
	    RECT 326.0000 146.0000 330.0000 146.2000 ;
	    RECT 322.8000 142.2000 323.6000 144.2000 ;
	    RECT 326.0000 142.2000 326.8000 146.0000 ;
	    RECT 329.2000 142.8000 330.0000 146.0000 ;
	    RECT 330.8000 143.4000 331.6000 146.2000 ;
	    RECT 332.4000 142.8000 333.2000 146.2000 ;
	    RECT 329.2000 142.2000 333.2000 142.8000 ;
	    RECT 334.0000 142.2000 334.8000 146.2000 ;
	    RECT 335.6000 146.0000 339.6000 146.2000 ;
	    RECT 335.6000 142.2000 336.4000 146.0000 ;
	    RECT 338.8000 142.2000 339.6000 146.0000 ;
	    RECT 340.4000 144.8000 341.2000 146.4000 ;
	    RECT 342.2000 144.2000 342.8000 147.6000 ;
	    RECT 346.0000 147.2000 346.8000 147.6000 ;
	    RECT 345.4000 146.2000 349.0000 146.6000 ;
	    RECT 350.2000 146.2000 350.8000 147.6000 ;
	    RECT 353.4000 146.2000 354.0000 147.6000 ;
	    RECT 357.2000 147.2000 358.0000 147.6000 ;
	    RECT 360.4000 147.2000 361.2000 147.6000 ;
	    RECT 355.0000 146.2000 358.6000 146.6000 ;
	    RECT 359.8000 146.2000 363.4000 146.6000 ;
	    RECT 364.4000 146.2000 365.0000 147.6000 ;
	    RECT 366.0000 146.8000 366.8000 148.4000 ;
	    RECT 367.6000 146.2000 368.4000 149.7000 ;
	    RECT 372.4000 149.6000 373.4000 150.4000 ;
	    RECT 372.8000 148.4000 373.4000 149.6000 ;
	    RECT 374.0000 150.3000 374.8000 150.4000 ;
	    RECT 375.6000 150.3000 376.4000 150.4000 ;
	    RECT 374.0000 149.7000 376.4000 150.3000 ;
	    RECT 374.0000 148.8000 374.8000 149.7000 ;
	    RECT 375.6000 149.6000 376.4000 149.7000 ;
	    RECT 370.8000 147.6000 373.4000 148.4000 ;
	    RECT 375.6000 148.2000 376.4000 148.4000 ;
	    RECT 374.8000 147.6000 376.4000 148.2000 ;
	    RECT 371.0000 146.2000 371.6000 147.6000 ;
	    RECT 374.8000 147.2000 375.6000 147.6000 ;
	    RECT 377.2000 147.2000 378.0000 150.6000 ;
	    RECT 380.6000 150.4000 381.4000 150.6000 ;
	    RECT 383.8000 150.4000 384.4000 151.6000 ;
	    RECT 385.8000 151.8000 386.4000 153.0000 ;
	    RECT 387.0000 153.0000 387.8000 153.2000 ;
	    RECT 391.6000 153.0000 392.4000 153.2000 ;
	    RECT 387.0000 152.4000 392.4000 153.0000 ;
	    RECT 385.8000 151.4000 390.6000 151.8000 ;
	    RECT 394.8000 151.4000 395.6000 159.8000 ;
	    RECT 397.2000 153.6000 398.0000 154.4000 ;
	    RECT 397.2000 152.4000 397.8000 153.6000 ;
	    RECT 398.6000 152.4000 399.4000 159.8000 ;
	    RECT 396.4000 151.8000 397.8000 152.4000 ;
	    RECT 398.4000 151.8000 399.4000 152.4000 ;
	    RECT 396.4000 151.6000 397.2000 151.8000 ;
	    RECT 385.8000 151.2000 395.6000 151.4000 ;
	    RECT 389.8000 151.0000 395.6000 151.2000 ;
	    RECT 390.0000 150.8000 395.6000 151.0000 ;
	    RECT 398.4000 150.4000 399.0000 151.8000 ;
	    RECT 409.2000 151.2000 410.0000 159.8000 ;
	    RECT 413.4000 155.8000 414.6000 159.8000 ;
	    RECT 418.0000 155.8000 418.8000 159.8000 ;
	    RECT 422.4000 156.4000 423.2000 159.8000 ;
	    RECT 422.4000 155.8000 424.4000 156.4000 ;
	    RECT 414.0000 155.0000 414.8000 155.8000 ;
	    RECT 418.2000 155.2000 418.8000 155.8000 ;
	    RECT 417.4000 154.6000 421.0000 155.2000 ;
	    RECT 423.6000 155.0000 424.4000 155.8000 ;
	    RECT 417.4000 154.4000 418.2000 154.6000 ;
	    RECT 420.2000 154.4000 421.0000 154.6000 ;
	    RECT 412.4000 154.0000 413.8000 154.4000 ;
	    RECT 412.4000 153.6000 414.6000 154.0000 ;
	    RECT 413.2000 153.2000 414.6000 153.6000 ;
	    RECT 414.0000 152.2000 414.6000 153.2000 ;
	    RECT 416.2000 153.0000 418.4000 153.6000 ;
	    RECT 416.2000 152.8000 417.0000 153.0000 ;
	    RECT 414.0000 151.6000 416.4000 152.2000 ;
	    RECT 409.2000 150.6000 413.4000 151.2000 ;
	    RECT 379.0000 149.8000 379.8000 150.0000 ;
	    RECT 379.0000 149.2000 382.8000 149.8000 ;
	    RECT 383.6000 149.6000 384.4000 150.4000 ;
	    RECT 388.4000 150.2000 389.2000 150.4000 ;
	    RECT 388.4000 149.6000 393.4000 150.2000 ;
	    RECT 398.0000 149.6000 399.0000 150.4000 ;
	    RECT 382.0000 149.0000 382.8000 149.2000 ;
	    RECT 383.8000 148.4000 384.4000 149.6000 ;
	    RECT 392.6000 149.4000 393.4000 149.6000 ;
	    RECT 391.0000 148.4000 391.8000 148.6000 ;
	    RECT 398.4000 148.4000 399.0000 149.6000 ;
	    RECT 399.6000 150.3000 400.4000 150.4000 ;
	    RECT 402.8000 150.3000 403.6000 150.4000 ;
	    RECT 399.6000 149.7000 403.6000 150.3000 ;
	    RECT 399.6000 148.8000 400.4000 149.7000 ;
	    RECT 402.8000 149.6000 403.6000 149.7000 ;
	    RECT 383.8000 147.8000 394.8000 148.4000 ;
	    RECT 384.2000 147.6000 385.0000 147.8000 ;
	    RECT 377.2000 146.6000 381.0000 147.2000 ;
	    RECT 372.6000 146.2000 376.2000 146.6000 ;
	    RECT 342.0000 142.2000 342.8000 144.2000 ;
	    RECT 345.2000 146.0000 349.2000 146.2000 ;
	    RECT 345.2000 142.2000 346.0000 146.0000 ;
	    RECT 348.4000 142.8000 349.2000 146.0000 ;
	    RECT 350.0000 143.4000 350.8000 146.2000 ;
	    RECT 351.6000 142.8000 352.4000 146.2000 ;
	    RECT 348.4000 142.2000 352.4000 142.8000 ;
	    RECT 353.2000 142.2000 354.0000 146.2000 ;
	    RECT 354.8000 146.0000 358.8000 146.2000 ;
	    RECT 354.8000 142.2000 355.6000 146.0000 ;
	    RECT 358.0000 142.2000 358.8000 146.0000 ;
	    RECT 359.6000 146.0000 363.6000 146.2000 ;
	    RECT 359.6000 142.2000 360.4000 146.0000 ;
	    RECT 362.8000 142.2000 363.6000 146.0000 ;
	    RECT 364.4000 142.2000 365.2000 146.2000 ;
	    RECT 367.6000 145.6000 369.4000 146.2000 ;
	    RECT 368.6000 142.2000 369.4000 145.6000 ;
	    RECT 370.8000 142.2000 371.6000 146.2000 ;
	    RECT 372.4000 146.0000 376.4000 146.2000 ;
	    RECT 372.4000 142.2000 373.2000 146.0000 ;
	    RECT 375.6000 142.2000 376.4000 146.0000 ;
	    RECT 377.2000 142.2000 378.0000 146.6000 ;
	    RECT 380.2000 146.4000 381.0000 146.6000 ;
	    RECT 390.0000 146.4000 390.6000 147.8000 ;
	    RECT 393.2000 147.6000 394.8000 147.8000 ;
	    RECT 396.4000 147.6000 399.0000 148.4000 ;
	    RECT 401.2000 148.2000 402.0000 148.4000 ;
	    RECT 400.4000 147.6000 402.0000 148.2000 ;
	    RECT 388.2000 145.4000 389.0000 145.6000 ;
	    RECT 382.0000 144.2000 382.8000 145.0000 ;
	    RECT 386.2000 144.8000 389.0000 145.4000 ;
	    RECT 390.0000 144.8000 390.8000 146.4000 ;
	    RECT 386.2000 144.2000 386.8000 144.8000 ;
	    RECT 391.6000 144.2000 392.4000 145.0000 ;
	    RECT 381.4000 143.6000 382.8000 144.2000 ;
	    RECT 381.4000 142.2000 382.6000 143.6000 ;
	    RECT 386.0000 142.2000 386.8000 144.2000 ;
	    RECT 390.4000 143.6000 392.4000 144.2000 ;
	    RECT 390.4000 142.2000 391.2000 143.6000 ;
	    RECT 394.8000 142.2000 395.6000 147.0000 ;
	    RECT 396.6000 146.2000 397.2000 147.6000 ;
	    RECT 400.4000 147.2000 401.2000 147.6000 ;
	    RECT 409.2000 147.2000 410.0000 150.6000 ;
	    RECT 412.6000 150.4000 413.4000 150.6000 ;
	    RECT 411.0000 149.8000 411.8000 150.0000 ;
	    RECT 411.0000 149.2000 414.8000 149.8000 ;
	    RECT 414.0000 149.0000 414.8000 149.2000 ;
	    RECT 415.8000 148.4000 416.4000 151.6000 ;
	    RECT 417.8000 151.8000 418.4000 153.0000 ;
	    RECT 419.0000 153.0000 419.8000 153.2000 ;
	    RECT 423.6000 153.0000 424.4000 153.2000 ;
	    RECT 419.0000 152.4000 424.4000 153.0000 ;
	    RECT 417.8000 151.4000 422.6000 151.8000 ;
	    RECT 426.8000 151.4000 427.6000 159.8000 ;
	    RECT 417.8000 151.2000 427.6000 151.4000 ;
	    RECT 421.8000 151.0000 427.6000 151.2000 ;
	    RECT 422.0000 150.8000 427.6000 151.0000 ;
	    RECT 428.4000 151.2000 429.2000 159.8000 ;
	    RECT 432.6000 155.8000 433.8000 159.8000 ;
	    RECT 437.2000 155.8000 438.0000 159.8000 ;
	    RECT 441.6000 156.4000 442.4000 159.8000 ;
	    RECT 441.6000 155.8000 443.6000 156.4000 ;
	    RECT 433.2000 155.0000 434.0000 155.8000 ;
	    RECT 437.4000 155.2000 438.0000 155.8000 ;
	    RECT 436.6000 154.6000 440.2000 155.2000 ;
	    RECT 442.8000 155.0000 443.6000 155.8000 ;
	    RECT 436.6000 154.4000 437.4000 154.6000 ;
	    RECT 439.4000 154.4000 440.2000 154.6000 ;
	    RECT 432.4000 153.2000 433.8000 154.0000 ;
	    RECT 433.2000 152.2000 433.8000 153.2000 ;
	    RECT 435.4000 153.0000 437.6000 153.6000 ;
	    RECT 435.4000 152.8000 436.2000 153.0000 ;
	    RECT 433.2000 151.6000 435.6000 152.2000 ;
	    RECT 428.4000 150.6000 432.6000 151.2000 ;
	    RECT 420.4000 150.2000 421.2000 150.4000 ;
	    RECT 420.4000 149.6000 425.4000 150.2000 ;
	    RECT 424.6000 149.4000 425.4000 149.6000 ;
	    RECT 423.0000 148.4000 423.8000 148.6000 ;
	    RECT 415.8000 147.8000 426.8000 148.4000 ;
	    RECT 416.2000 147.6000 417.0000 147.8000 ;
	    RECT 409.2000 146.6000 413.0000 147.2000 ;
	    RECT 398.2000 146.2000 401.8000 146.6000 ;
	    RECT 396.4000 142.2000 397.2000 146.2000 ;
	    RECT 398.0000 146.0000 402.0000 146.2000 ;
	    RECT 398.0000 142.2000 398.8000 146.0000 ;
	    RECT 401.2000 142.2000 402.0000 146.0000 ;
	    RECT 409.2000 142.2000 410.0000 146.6000 ;
	    RECT 412.2000 146.4000 413.0000 146.6000 ;
	    RECT 422.0000 145.6000 422.6000 147.8000 ;
	    RECT 425.2000 147.6000 426.8000 147.8000 ;
	    RECT 428.4000 147.2000 429.2000 150.6000 ;
	    RECT 431.8000 150.4000 432.6000 150.6000 ;
	    RECT 430.2000 149.8000 431.0000 150.0000 ;
	    RECT 430.2000 149.2000 434.0000 149.8000 ;
	    RECT 433.2000 149.0000 434.0000 149.2000 ;
	    RECT 435.0000 148.4000 435.6000 151.6000 ;
	    RECT 437.0000 151.8000 437.6000 153.0000 ;
	    RECT 438.2000 153.0000 439.0000 153.2000 ;
	    RECT 442.8000 153.0000 443.6000 153.2000 ;
	    RECT 438.2000 152.4000 443.6000 153.0000 ;
	    RECT 437.0000 151.4000 441.8000 151.8000 ;
	    RECT 446.0000 151.4000 446.8000 159.8000 ;
	    RECT 437.0000 151.2000 446.8000 151.4000 ;
	    RECT 441.0000 151.0000 446.8000 151.2000 ;
	    RECT 441.2000 150.8000 446.8000 151.0000 ;
	    RECT 439.6000 150.2000 440.4000 150.4000 ;
	    RECT 449.2000 150.3000 450.0000 159.8000 ;
	    RECT 453.2000 153.6000 454.0000 154.4000 ;
	    RECT 450.8000 151.6000 451.6000 153.2000 ;
	    RECT 453.2000 152.4000 453.8000 153.6000 ;
	    RECT 454.6000 152.4000 455.4000 159.8000 ;
	    RECT 452.4000 151.8000 453.8000 152.4000 ;
	    RECT 454.4000 151.8000 455.4000 152.4000 ;
	    RECT 452.4000 151.6000 453.2000 151.8000 ;
	    RECT 452.5000 150.3000 453.1000 151.6000 ;
	    RECT 439.6000 149.6000 444.6000 150.2000 ;
	    RECT 441.2000 149.4000 442.0000 149.6000 ;
	    RECT 443.8000 149.4000 444.6000 149.6000 ;
	    RECT 449.2000 149.7000 453.1000 150.3000 ;
	    RECT 442.2000 148.4000 443.0000 148.6000 ;
	    RECT 435.0000 147.8000 446.0000 148.4000 ;
	    RECT 435.4000 147.6000 436.2000 147.8000 ;
	    RECT 420.2000 145.4000 421.0000 145.6000 ;
	    RECT 414.0000 144.2000 414.8000 145.0000 ;
	    RECT 418.2000 144.8000 421.0000 145.4000 ;
	    RECT 422.0000 144.8000 422.8000 145.6000 ;
	    RECT 418.2000 144.2000 418.8000 144.8000 ;
	    RECT 423.6000 144.2000 424.4000 145.0000 ;
	    RECT 413.4000 143.6000 414.8000 144.2000 ;
	    RECT 413.4000 142.2000 414.6000 143.6000 ;
	    RECT 418.0000 142.2000 418.8000 144.2000 ;
	    RECT 422.4000 143.6000 424.4000 144.2000 ;
	    RECT 422.4000 142.2000 423.2000 143.6000 ;
	    RECT 426.8000 142.2000 427.6000 147.0000 ;
	    RECT 428.4000 146.6000 432.2000 147.2000 ;
	    RECT 428.4000 142.2000 429.2000 146.6000 ;
	    RECT 431.4000 146.4000 432.2000 146.6000 ;
	    RECT 441.2000 145.6000 441.8000 147.8000 ;
	    RECT 444.4000 147.6000 446.0000 147.8000 ;
	    RECT 439.4000 145.4000 440.2000 145.6000 ;
	    RECT 433.2000 144.2000 434.0000 145.0000 ;
	    RECT 437.4000 144.8000 440.2000 145.4000 ;
	    RECT 441.2000 144.8000 442.0000 145.6000 ;
	    RECT 437.4000 144.2000 438.0000 144.8000 ;
	    RECT 442.8000 144.2000 443.6000 145.0000 ;
	    RECT 432.6000 143.6000 434.0000 144.2000 ;
	    RECT 432.6000 142.2000 433.8000 143.6000 ;
	    RECT 437.2000 142.2000 438.0000 144.2000 ;
	    RECT 441.6000 143.6000 443.6000 144.2000 ;
	    RECT 441.6000 142.2000 442.4000 143.6000 ;
	    RECT 446.0000 142.2000 446.8000 147.0000 ;
	    RECT 447.6000 146.8000 448.4000 148.4000 ;
	    RECT 449.2000 146.2000 450.0000 149.7000 ;
	    RECT 454.4000 148.4000 455.0000 151.8000 ;
	    RECT 458.8000 151.2000 459.6000 159.8000 ;
	    RECT 463.0000 155.8000 464.2000 159.8000 ;
	    RECT 467.6000 155.8000 468.4000 159.8000 ;
	    RECT 472.0000 156.4000 472.8000 159.8000 ;
	    RECT 472.0000 155.8000 474.0000 156.4000 ;
	    RECT 463.6000 155.0000 464.4000 155.8000 ;
	    RECT 467.8000 155.2000 468.4000 155.8000 ;
	    RECT 467.0000 154.6000 470.6000 155.2000 ;
	    RECT 473.2000 155.0000 474.0000 155.8000 ;
	    RECT 467.0000 154.4000 467.8000 154.6000 ;
	    RECT 469.8000 154.4000 470.6000 154.6000 ;
	    RECT 462.8000 153.2000 464.2000 154.0000 ;
	    RECT 463.6000 152.2000 464.2000 153.2000 ;
	    RECT 465.8000 153.0000 468.0000 153.6000 ;
	    RECT 465.8000 152.8000 466.6000 153.0000 ;
	    RECT 463.6000 151.6000 466.0000 152.2000 ;
	    RECT 458.8000 150.6000 463.0000 151.2000 ;
	    RECT 455.6000 148.8000 456.4000 150.4000 ;
	    RECT 450.8000 148.3000 451.6000 148.4000 ;
	    RECT 452.4000 148.3000 455.0000 148.4000 ;
	    RECT 450.8000 147.7000 455.0000 148.3000 ;
	    RECT 457.2000 148.2000 458.0000 148.4000 ;
	    RECT 450.8000 147.6000 451.6000 147.7000 ;
	    RECT 452.4000 147.6000 455.0000 147.7000 ;
	    RECT 456.4000 147.6000 458.0000 148.2000 ;
	    RECT 452.6000 146.2000 453.2000 147.6000 ;
	    RECT 456.4000 147.2000 457.2000 147.6000 ;
	    RECT 458.8000 147.2000 459.6000 150.6000 ;
	    RECT 462.2000 150.4000 463.0000 150.6000 ;
	    RECT 460.6000 149.8000 461.4000 150.0000 ;
	    RECT 460.6000 149.2000 464.4000 149.8000 ;
	    RECT 463.6000 149.0000 464.4000 149.2000 ;
	    RECT 465.4000 148.4000 466.0000 151.6000 ;
	    RECT 467.4000 151.8000 468.0000 153.0000 ;
	    RECT 468.6000 153.0000 469.4000 153.2000 ;
	    RECT 473.2000 153.0000 474.0000 153.2000 ;
	    RECT 468.6000 152.4000 474.0000 153.0000 ;
	    RECT 467.4000 151.4000 472.2000 151.8000 ;
	    RECT 476.4000 151.4000 477.2000 159.8000 ;
	    RECT 478.8000 153.6000 479.6000 154.4000 ;
	    RECT 478.8000 152.4000 479.4000 153.6000 ;
	    RECT 480.2000 152.4000 481.0000 159.8000 ;
	    RECT 478.0000 151.8000 479.4000 152.4000 ;
	    RECT 480.0000 151.8000 481.0000 152.4000 ;
	    RECT 478.0000 151.6000 478.8000 151.8000 ;
	    RECT 467.4000 151.2000 477.2000 151.4000 ;
	    RECT 471.4000 151.0000 477.2000 151.2000 ;
	    RECT 471.6000 150.8000 477.2000 151.0000 ;
	    RECT 470.0000 150.2000 470.8000 150.4000 ;
	    RECT 478.0000 150.3000 478.8000 150.4000 ;
	    RECT 480.0000 150.3000 480.6000 151.8000 ;
	    RECT 470.0000 149.6000 475.0000 150.2000 ;
	    RECT 478.0000 149.7000 480.6000 150.3000 ;
	    RECT 478.0000 149.6000 478.8000 149.7000 ;
	    RECT 471.6000 149.4000 472.4000 149.6000 ;
	    RECT 474.2000 149.4000 475.0000 149.6000 ;
	    RECT 472.6000 148.4000 473.4000 148.6000 ;
	    RECT 480.0000 148.4000 480.6000 149.7000 ;
	    RECT 481.2000 148.8000 482.0000 150.4000 ;
	    RECT 465.4000 147.8000 476.4000 148.4000 ;
	    RECT 465.8000 147.6000 466.6000 147.8000 ;
	    RECT 470.0000 147.6000 470.8000 147.8000 ;
	    RECT 458.8000 146.6000 462.6000 147.2000 ;
	    RECT 454.2000 146.2000 457.8000 146.6000 ;
	    RECT 449.2000 145.6000 451.0000 146.2000 ;
	    RECT 450.2000 142.2000 451.0000 145.6000 ;
	    RECT 452.4000 142.2000 453.2000 146.2000 ;
	    RECT 454.0000 146.0000 458.0000 146.2000 ;
	    RECT 454.0000 142.2000 454.8000 146.0000 ;
	    RECT 457.2000 142.2000 458.0000 146.0000 ;
	    RECT 458.8000 142.2000 459.6000 146.6000 ;
	    RECT 461.8000 146.4000 462.6000 146.6000 ;
	    RECT 471.6000 145.6000 472.2000 147.8000 ;
	    RECT 474.8000 147.6000 476.4000 147.8000 ;
	    RECT 478.0000 147.6000 480.6000 148.4000 ;
	    RECT 482.8000 148.3000 483.6000 148.4000 ;
	    RECT 484.4000 148.3000 485.2000 159.8000 ;
	    RECT 489.2000 155.8000 490.0000 159.8000 ;
	    RECT 489.4000 151.6000 490.0000 155.8000 ;
	    RECT 492.4000 151.8000 493.2000 159.8000 ;
	    RECT 489.4000 151.0000 491.8000 151.6000 ;
	    RECT 489.2000 149.6000 490.0000 150.4000 ;
	    RECT 482.8000 148.2000 485.2000 148.3000 ;
	    RECT 482.0000 147.7000 485.2000 148.2000 ;
	    RECT 482.0000 147.6000 483.6000 147.7000 ;
	    RECT 469.8000 145.4000 470.6000 145.6000 ;
	    RECT 463.6000 144.2000 464.4000 145.0000 ;
	    RECT 467.8000 144.8000 470.6000 145.4000 ;
	    RECT 471.6000 144.8000 472.4000 145.6000 ;
	    RECT 467.8000 144.2000 468.4000 144.8000 ;
	    RECT 473.2000 144.2000 474.0000 145.0000 ;
	    RECT 463.0000 143.6000 464.4000 144.2000 ;
	    RECT 463.0000 142.2000 464.2000 143.6000 ;
	    RECT 467.6000 142.2000 468.4000 144.2000 ;
	    RECT 472.0000 143.6000 474.0000 144.2000 ;
	    RECT 472.0000 142.2000 472.8000 143.6000 ;
	    RECT 476.4000 142.2000 477.2000 147.0000 ;
	    RECT 478.2000 146.2000 478.8000 147.6000 ;
	    RECT 482.0000 147.2000 482.8000 147.6000 ;
	    RECT 479.8000 146.2000 483.4000 146.6000 ;
	    RECT 478.0000 142.2000 478.8000 146.2000 ;
	    RECT 479.6000 146.0000 483.6000 146.2000 ;
	    RECT 479.6000 142.2000 480.4000 146.0000 ;
	    RECT 482.8000 142.2000 483.6000 146.0000 ;
	    RECT 484.4000 142.2000 485.2000 147.7000 ;
	    RECT 487.6000 147.6000 488.4000 149.2000 ;
	    RECT 489.4000 148.8000 490.0000 149.6000 ;
	    RECT 489.4000 148.2000 490.4000 148.8000 ;
	    RECT 489.6000 148.0000 490.4000 148.2000 ;
	    RECT 491.2000 147.6000 491.8000 151.0000 ;
	    RECT 492.6000 150.4000 493.2000 151.8000 ;
	    RECT 492.4000 149.6000 493.2000 150.4000 ;
	    RECT 491.2000 147.4000 492.0000 147.6000 ;
	    RECT 489.0000 147.0000 492.0000 147.4000 ;
	    RECT 487.8000 146.8000 492.0000 147.0000 ;
	    RECT 487.8000 146.4000 489.6000 146.8000 ;
	    RECT 486.0000 144.8000 486.8000 146.4000 ;
	    RECT 487.8000 146.2000 488.4000 146.4000 ;
	    RECT 492.6000 146.2000 493.2000 149.6000 ;
	    RECT 487.6000 142.2000 488.4000 146.2000 ;
	    RECT 491.8000 145.2000 493.2000 146.2000 ;
	    RECT 494.0000 151.2000 494.8000 159.8000 ;
	    RECT 498.2000 155.8000 499.4000 159.8000 ;
	    RECT 502.8000 155.8000 503.6000 159.8000 ;
	    RECT 507.2000 156.4000 508.0000 159.8000 ;
	    RECT 507.2000 155.8000 509.2000 156.4000 ;
	    RECT 498.8000 155.0000 499.6000 155.8000 ;
	    RECT 503.0000 155.2000 503.6000 155.8000 ;
	    RECT 502.2000 154.6000 505.8000 155.2000 ;
	    RECT 508.4000 155.0000 509.2000 155.8000 ;
	    RECT 502.2000 154.4000 503.0000 154.6000 ;
	    RECT 505.0000 154.4000 505.8000 154.6000 ;
	    RECT 497.2000 154.0000 498.6000 154.4000 ;
	    RECT 497.2000 153.6000 499.4000 154.0000 ;
	    RECT 498.0000 153.2000 499.4000 153.6000 ;
	    RECT 498.8000 152.2000 499.4000 153.2000 ;
	    RECT 501.0000 153.0000 503.2000 153.6000 ;
	    RECT 501.0000 152.8000 501.8000 153.0000 ;
	    RECT 498.8000 151.6000 501.2000 152.2000 ;
	    RECT 494.0000 150.6000 498.2000 151.2000 ;
	    RECT 494.0000 147.2000 494.8000 150.6000 ;
	    RECT 497.4000 150.4000 498.2000 150.6000 ;
	    RECT 495.8000 149.8000 496.6000 150.0000 ;
	    RECT 495.8000 149.2000 499.6000 149.8000 ;
	    RECT 498.8000 149.0000 499.6000 149.2000 ;
	    RECT 500.6000 148.4000 501.2000 151.6000 ;
	    RECT 502.6000 151.8000 503.2000 153.0000 ;
	    RECT 503.8000 153.0000 504.6000 153.2000 ;
	    RECT 508.4000 153.0000 509.2000 153.2000 ;
	    RECT 503.8000 152.4000 509.2000 153.0000 ;
	    RECT 502.6000 151.4000 507.4000 151.8000 ;
	    RECT 511.6000 151.4000 512.4000 159.8000 ;
	    RECT 502.6000 151.2000 512.4000 151.4000 ;
	    RECT 506.6000 151.0000 512.4000 151.2000 ;
	    RECT 506.8000 150.8000 512.4000 151.0000 ;
	    RECT 505.2000 150.2000 506.0000 150.4000 ;
	    RECT 505.2000 149.6000 510.2000 150.2000 ;
	    RECT 506.8000 149.4000 507.6000 149.6000 ;
	    RECT 509.4000 149.4000 510.2000 149.6000 ;
	    RECT 507.8000 148.4000 508.6000 148.6000 ;
	    RECT 500.6000 147.8000 511.6000 148.4000 ;
	    RECT 501.0000 147.6000 501.8000 147.8000 ;
	    RECT 505.2000 147.6000 506.0000 147.8000 ;
	    RECT 494.0000 146.6000 497.8000 147.2000 ;
	    RECT 491.8000 142.2000 492.6000 145.2000 ;
	    RECT 494.0000 142.2000 494.8000 146.6000 ;
	    RECT 497.0000 146.4000 497.8000 146.6000 ;
	    RECT 506.8000 145.6000 507.4000 147.8000 ;
	    RECT 510.0000 147.6000 511.6000 147.8000 ;
	    RECT 505.0000 145.4000 505.8000 145.6000 ;
	    RECT 498.8000 144.2000 499.6000 145.0000 ;
	    RECT 503.0000 144.8000 505.8000 145.4000 ;
	    RECT 506.8000 144.8000 507.6000 145.6000 ;
	    RECT 503.0000 144.2000 503.6000 144.8000 ;
	    RECT 508.4000 144.2000 509.2000 145.0000 ;
	    RECT 498.2000 143.6000 499.6000 144.2000 ;
	    RECT 498.2000 142.2000 499.4000 143.6000 ;
	    RECT 502.8000 142.2000 503.6000 144.2000 ;
	    RECT 507.2000 143.6000 509.2000 144.2000 ;
	    RECT 507.2000 142.2000 508.0000 143.6000 ;
	    RECT 511.6000 142.2000 512.4000 147.0000 ;
	    RECT 4.4000 135.2000 5.2000 139.8000 ;
	    RECT 9.2000 135.2000 10.0000 139.8000 ;
	    RECT 3.0000 134.6000 5.2000 135.2000 ;
	    RECT 7.8000 134.6000 10.0000 135.2000 ;
	    RECT 10.8000 135.4000 11.6000 139.8000 ;
	    RECT 15.0000 138.4000 16.2000 139.8000 ;
	    RECT 15.0000 137.8000 16.4000 138.4000 ;
	    RECT 19.6000 137.8000 20.4000 139.8000 ;
	    RECT 24.0000 138.4000 24.8000 139.8000 ;
	    RECT 24.0000 137.8000 26.0000 138.4000 ;
	    RECT 15.6000 137.0000 16.4000 137.8000 ;
	    RECT 19.8000 137.2000 20.4000 137.8000 ;
	    RECT 19.8000 136.6000 22.6000 137.2000 ;
	    RECT 21.8000 136.4000 22.6000 136.6000 ;
	    RECT 23.6000 136.4000 24.4000 137.2000 ;
	    RECT 25.2000 137.0000 26.0000 137.8000 ;
	    RECT 13.8000 135.4000 14.6000 135.6000 ;
	    RECT 10.8000 134.8000 14.6000 135.4000 ;
	    RECT 3.0000 131.6000 3.6000 134.6000 ;
	    RECT 4.4000 131.6000 5.2000 133.2000 ;
	    RECT 7.8000 131.6000 8.4000 134.6000 ;
	    RECT 9.2000 131.6000 10.0000 133.2000 ;
	    RECT 2.4000 130.8000 3.6000 131.6000 ;
	    RECT 7.2000 130.8000 8.4000 131.6000 ;
	    RECT 3.0000 130.2000 3.6000 130.8000 ;
	    RECT 7.8000 130.2000 8.4000 130.8000 ;
	    RECT 10.8000 131.4000 11.6000 134.8000 ;
	    RECT 17.8000 134.2000 19.6000 134.4000 ;
	    RECT 23.6000 134.2000 24.2000 136.4000 ;
	    RECT 28.4000 135.0000 29.2000 139.8000 ;
	    RECT 30.0000 135.8000 30.8000 139.8000 ;
	    RECT 31.6000 136.0000 32.4000 139.8000 ;
	    RECT 34.8000 136.0000 35.6000 139.8000 ;
	    RECT 31.6000 135.8000 35.6000 136.0000 ;
	    RECT 36.4000 136.0000 37.2000 139.8000 ;
	    RECT 39.6000 136.0000 40.4000 139.8000 ;
	    RECT 36.4000 135.8000 40.4000 136.0000 ;
	    RECT 41.2000 135.8000 42.0000 139.8000 ;
	    RECT 30.2000 134.4000 30.8000 135.8000 ;
	    RECT 31.8000 135.4000 35.4000 135.8000 ;
	    RECT 36.6000 135.4000 40.2000 135.8000 ;
	    RECT 34.0000 134.4000 34.8000 134.8000 ;
	    RECT 37.2000 134.4000 38.0000 134.8000 ;
	    RECT 41.2000 134.4000 41.8000 135.8000 ;
	    RECT 42.8000 135.4000 43.6000 139.8000 ;
	    RECT 47.0000 138.4000 48.2000 139.8000 ;
	    RECT 47.0000 137.8000 48.4000 138.4000 ;
	    RECT 51.6000 137.8000 52.4000 139.8000 ;
	    RECT 56.0000 138.4000 56.8000 139.8000 ;
	    RECT 56.0000 137.8000 58.0000 138.4000 ;
	    RECT 47.6000 137.0000 48.4000 137.8000 ;
	    RECT 51.8000 137.2000 52.4000 137.8000 ;
	    RECT 51.8000 136.6000 54.6000 137.2000 ;
	    RECT 53.8000 136.4000 54.6000 136.6000 ;
	    RECT 55.6000 136.4000 56.4000 137.2000 ;
	    RECT 57.2000 137.0000 58.0000 137.8000 ;
	    RECT 45.8000 135.4000 46.6000 135.6000 ;
	    RECT 42.8000 134.8000 46.6000 135.4000 ;
	    RECT 26.8000 134.2000 28.4000 134.4000 ;
	    RECT 17.4000 133.6000 28.4000 134.2000 ;
	    RECT 30.0000 133.6000 32.6000 134.4000 ;
	    RECT 34.0000 134.3000 35.6000 134.4000 ;
	    RECT 36.4000 134.3000 38.0000 134.4000 ;
	    RECT 34.0000 133.8000 38.0000 134.3000 ;
	    RECT 34.8000 133.7000 37.2000 133.8000 ;
	    RECT 34.8000 133.6000 35.6000 133.7000 ;
	    RECT 36.4000 133.6000 37.2000 133.7000 ;
	    RECT 39.4000 133.6000 42.0000 134.4000 ;
	    RECT 15.6000 132.8000 16.4000 133.0000 ;
	    RECT 12.6000 132.2000 16.4000 132.8000 ;
	    RECT 12.6000 132.0000 13.4000 132.2000 ;
	    RECT 14.2000 131.4000 15.0000 131.6000 ;
	    RECT 10.8000 130.8000 15.0000 131.4000 ;
	    RECT 3.0000 129.6000 5.2000 130.2000 ;
	    RECT 7.8000 129.6000 10.0000 130.2000 ;
	    RECT 4.4000 122.2000 5.2000 129.6000 ;
	    RECT 9.2000 122.2000 10.0000 129.6000 ;
	    RECT 10.8000 122.2000 11.6000 130.8000 ;
	    RECT 17.4000 130.4000 18.0000 133.6000 ;
	    RECT 24.6000 133.4000 25.4000 133.6000 ;
	    RECT 23.6000 132.4000 24.4000 132.6000 ;
	    RECT 26.2000 132.4000 27.0000 132.6000 ;
	    RECT 22.0000 131.8000 27.0000 132.4000 ;
	    RECT 22.0000 131.6000 22.8000 131.8000 ;
	    RECT 23.6000 131.0000 29.2000 131.2000 ;
	    RECT 23.4000 130.8000 29.2000 131.0000 ;
	    RECT 15.6000 129.8000 18.0000 130.4000 ;
	    RECT 19.4000 130.6000 29.2000 130.8000 ;
	    RECT 19.4000 130.2000 24.2000 130.6000 ;
	    RECT 15.6000 128.8000 16.2000 129.8000 ;
	    RECT 14.8000 128.0000 16.2000 128.8000 ;
	    RECT 17.8000 129.0000 18.6000 129.2000 ;
	    RECT 19.4000 129.0000 20.0000 130.2000 ;
	    RECT 17.8000 128.4000 20.0000 129.0000 ;
	    RECT 20.6000 129.0000 26.0000 129.6000 ;
	    RECT 20.6000 128.8000 21.4000 129.0000 ;
	    RECT 25.2000 128.8000 26.0000 129.0000 ;
	    RECT 19.0000 127.4000 19.8000 127.6000 ;
	    RECT 21.8000 127.4000 22.6000 127.6000 ;
	    RECT 15.6000 126.2000 16.4000 127.0000 ;
	    RECT 19.0000 126.8000 22.6000 127.4000 ;
	    RECT 19.8000 126.2000 20.4000 126.8000 ;
	    RECT 25.2000 126.2000 26.0000 127.0000 ;
	    RECT 15.0000 122.2000 16.2000 126.2000 ;
	    RECT 19.6000 122.2000 20.4000 126.2000 ;
	    RECT 24.0000 125.6000 26.0000 126.2000 ;
	    RECT 24.0000 122.2000 24.8000 125.6000 ;
	    RECT 28.4000 122.2000 29.2000 130.6000 ;
	    RECT 30.0000 130.2000 30.8000 130.4000 ;
	    RECT 32.0000 130.2000 32.6000 133.6000 ;
	    RECT 33.2000 132.3000 34.0000 133.2000 ;
	    RECT 38.0000 132.3000 38.8000 133.2000 ;
	    RECT 33.2000 131.7000 38.8000 132.3000 ;
	    RECT 33.2000 131.6000 34.0000 131.7000 ;
	    RECT 38.0000 131.6000 38.8000 131.7000 ;
	    RECT 39.4000 132.3000 40.0000 133.6000 ;
	    RECT 41.2000 132.3000 42.0000 132.4000 ;
	    RECT 39.4000 131.7000 42.0000 132.3000 ;
	    RECT 39.4000 130.2000 40.0000 131.7000 ;
	    RECT 41.2000 131.6000 42.0000 131.7000 ;
	    RECT 42.8000 131.4000 43.6000 134.8000 ;
	    RECT 49.8000 134.2000 50.6000 134.4000 ;
	    RECT 52.4000 134.2000 53.2000 134.4000 ;
	    RECT 55.6000 134.2000 56.2000 136.4000 ;
	    RECT 60.4000 135.0000 61.2000 139.8000 ;
	    RECT 62.0000 135.6000 62.8000 139.8000 ;
	    RECT 63.6000 136.0000 64.4000 139.8000 ;
	    RECT 66.8000 136.0000 67.6000 139.8000 ;
	    RECT 63.6000 135.8000 67.6000 136.0000 ;
	    RECT 62.2000 134.4000 62.8000 135.6000 ;
	    RECT 63.8000 135.4000 67.4000 135.8000 ;
	    RECT 66.0000 134.4000 66.8000 134.8000 ;
	    RECT 58.8000 134.2000 60.4000 134.4000 ;
	    RECT 49.4000 133.6000 60.4000 134.2000 ;
	    RECT 62.0000 133.6000 64.6000 134.4000 ;
	    RECT 66.0000 133.8000 67.6000 134.4000 ;
	    RECT 66.8000 133.6000 67.6000 133.8000 ;
	    RECT 68.4000 133.6000 69.2000 135.2000 ;
	    RECT 47.6000 132.8000 48.4000 133.0000 ;
	    RECT 44.6000 132.2000 48.4000 132.8000 ;
	    RECT 44.6000 132.0000 45.4000 132.2000 ;
	    RECT 46.2000 131.4000 47.0000 131.6000 ;
	    RECT 42.8000 130.8000 47.0000 131.4000 ;
	    RECT 41.2000 130.2000 42.0000 130.4000 ;
	    RECT 30.0000 129.6000 31.4000 130.2000 ;
	    RECT 32.0000 129.6000 33.0000 130.2000 ;
	    RECT 30.8000 128.4000 31.4000 129.6000 ;
	    RECT 32.2000 128.4000 33.0000 129.6000 ;
	    RECT 39.0000 129.6000 40.0000 130.2000 ;
	    RECT 40.6000 129.6000 42.0000 130.2000 ;
	    RECT 30.8000 127.6000 31.6000 128.4000 ;
	    RECT 32.2000 127.6000 34.0000 128.4000 ;
	    RECT 32.2000 122.2000 33.0000 127.6000 ;
	    RECT 39.0000 122.2000 39.8000 129.6000 ;
	    RECT 40.6000 128.4000 41.2000 129.6000 ;
	    RECT 40.4000 128.3000 41.2000 128.4000 ;
	    RECT 42.8000 128.3000 43.6000 130.8000 ;
	    RECT 49.4000 130.4000 50.0000 133.6000 ;
	    RECT 56.6000 133.4000 57.4000 133.6000 ;
	    RECT 55.6000 132.4000 56.4000 132.6000 ;
	    RECT 58.2000 132.4000 59.0000 132.6000 ;
	    RECT 54.0000 131.8000 59.0000 132.4000 ;
	    RECT 54.0000 131.6000 54.8000 131.8000 ;
	    RECT 55.6000 131.0000 61.2000 131.2000 ;
	    RECT 55.4000 130.8000 61.2000 131.0000 ;
	    RECT 47.6000 129.8000 50.0000 130.4000 ;
	    RECT 51.4000 130.6000 61.2000 130.8000 ;
	    RECT 51.4000 130.2000 56.2000 130.6000 ;
	    RECT 47.6000 128.8000 48.2000 129.8000 ;
	    RECT 40.4000 127.7000 43.6000 128.3000 ;
	    RECT 46.8000 128.0000 48.2000 128.8000 ;
	    RECT 49.8000 129.0000 50.6000 129.2000 ;
	    RECT 51.4000 129.0000 52.0000 130.2000 ;
	    RECT 49.8000 128.4000 52.0000 129.0000 ;
	    RECT 52.6000 129.0000 58.0000 129.6000 ;
	    RECT 52.6000 128.8000 53.4000 129.0000 ;
	    RECT 57.2000 128.8000 58.0000 129.0000 ;
	    RECT 40.4000 127.6000 41.2000 127.7000 ;
	    RECT 42.8000 122.2000 43.6000 127.7000 ;
	    RECT 51.0000 127.4000 51.8000 127.6000 ;
	    RECT 53.8000 127.4000 54.6000 127.6000 ;
	    RECT 47.6000 126.2000 48.4000 127.0000 ;
	    RECT 51.0000 126.8000 54.6000 127.4000 ;
	    RECT 51.8000 126.2000 52.4000 126.8000 ;
	    RECT 57.2000 126.2000 58.0000 127.0000 ;
	    RECT 47.0000 122.2000 48.2000 126.2000 ;
	    RECT 51.6000 122.2000 52.4000 126.2000 ;
	    RECT 56.0000 125.6000 58.0000 126.2000 ;
	    RECT 56.0000 122.2000 56.8000 125.6000 ;
	    RECT 60.4000 122.2000 61.2000 130.6000 ;
	    RECT 62.0000 130.2000 62.8000 130.4000 ;
	    RECT 64.0000 130.2000 64.6000 133.6000 ;
	    RECT 65.2000 131.6000 66.0000 133.2000 ;
	    RECT 66.8000 132.3000 67.6000 132.4000 ;
	    RECT 70.0000 132.3000 70.8000 139.8000 ;
	    RECT 73.2000 135.8000 74.0000 139.8000 ;
	    RECT 74.8000 136.0000 75.6000 139.8000 ;
	    RECT 78.0000 136.0000 78.8000 139.8000 ;
	    RECT 81.2000 137.8000 82.0000 139.8000 ;
	    RECT 74.8000 135.8000 78.8000 136.0000 ;
	    RECT 73.4000 134.4000 74.0000 135.8000 ;
	    RECT 75.0000 135.4000 78.6000 135.8000 ;
	    RECT 79.6000 135.6000 80.4000 137.2000 ;
	    RECT 77.2000 134.4000 78.0000 134.8000 ;
	    RECT 81.4000 134.4000 82.0000 137.8000 ;
	    RECT 82.8000 136.3000 83.6000 136.4000 ;
	    RECT 84.4000 136.3000 85.2000 139.8000 ;
	    RECT 82.8000 135.7000 85.2000 136.3000 ;
	    RECT 86.0000 136.0000 86.8000 139.8000 ;
	    RECT 89.2000 136.0000 90.0000 139.8000 ;
	    RECT 86.0000 135.8000 90.0000 136.0000 ;
	    RECT 90.8000 135.8000 91.6000 139.8000 ;
	    RECT 92.4000 136.0000 93.2000 139.8000 ;
	    RECT 95.6000 136.0000 96.4000 139.8000 ;
	    RECT 92.4000 135.8000 96.4000 136.0000 ;
	    RECT 97.2000 136.0000 98.0000 139.8000 ;
	    RECT 100.4000 136.0000 101.2000 139.8000 ;
	    RECT 97.2000 135.8000 101.2000 136.0000 ;
	    RECT 102.0000 135.8000 102.8000 139.8000 ;
	    RECT 119.6000 139.2000 123.6000 139.8000 ;
	    RECT 110.0000 137.0000 110.8000 139.0000 ;
	    RECT 82.8000 135.6000 83.6000 135.7000 ;
	    RECT 84.6000 134.4000 85.2000 135.7000 ;
	    RECT 86.2000 135.4000 89.8000 135.8000 ;
	    RECT 88.4000 134.4000 89.2000 134.8000 ;
	    RECT 91.0000 134.4000 91.6000 135.8000 ;
	    RECT 92.6000 135.4000 96.2000 135.8000 ;
	    RECT 97.4000 135.4000 101.0000 135.8000 ;
	    RECT 94.8000 134.4000 95.6000 134.8000 ;
	    RECT 98.0000 134.4000 98.8000 134.8000 ;
	    RECT 102.0000 134.4000 102.6000 135.8000 ;
	    RECT 110.0000 134.8000 110.6000 137.0000 ;
	    RECT 114.2000 136.0000 115.0000 139.0000 ;
	    RECT 114.2000 135.4000 115.8000 136.0000 ;
	    RECT 119.6000 135.8000 120.4000 139.2000 ;
	    RECT 121.2000 135.8000 122.0000 138.6000 ;
	    RECT 122.8000 136.0000 123.6000 139.2000 ;
	    RECT 126.0000 136.0000 126.8000 139.8000 ;
	    RECT 122.8000 135.8000 126.8000 136.0000 ;
	    RECT 127.6000 135.8000 128.4000 139.8000 ;
	    RECT 129.2000 136.0000 130.0000 139.8000 ;
	    RECT 132.4000 136.0000 133.2000 139.8000 ;
	    RECT 129.2000 135.8000 133.2000 136.0000 ;
	    RECT 134.0000 139.2000 138.0000 139.8000 ;
	    RECT 134.0000 135.8000 134.8000 139.2000 ;
	    RECT 135.6000 135.8000 136.4000 138.6000 ;
	    RECT 137.2000 136.0000 138.0000 139.2000 ;
	    RECT 140.4000 136.0000 141.2000 139.8000 ;
	    RECT 137.2000 135.8000 141.2000 136.0000 ;
	    RECT 142.0000 139.2000 146.0000 139.8000 ;
	    RECT 142.0000 135.8000 142.8000 139.2000 ;
	    RECT 115.0000 135.0000 115.8000 135.4000 ;
	    RECT 73.2000 133.6000 75.8000 134.4000 ;
	    RECT 77.2000 133.8000 78.8000 134.4000 ;
	    RECT 78.0000 133.6000 78.8000 133.8000 ;
	    RECT 81.2000 133.6000 82.0000 134.4000 ;
	    RECT 84.4000 133.6000 87.0000 134.4000 ;
	    RECT 88.4000 133.8000 90.0000 134.4000 ;
	    RECT 89.2000 133.6000 90.0000 133.8000 ;
	    RECT 90.8000 133.6000 93.4000 134.4000 ;
	    RECT 94.8000 133.8000 96.4000 134.4000 ;
	    RECT 95.6000 133.6000 96.4000 133.8000 ;
	    RECT 97.2000 133.8000 98.8000 134.4000 ;
	    RECT 97.2000 133.6000 98.0000 133.8000 ;
	    RECT 100.2000 133.6000 102.8000 134.4000 ;
	    RECT 110.0000 134.2000 114.2000 134.8000 ;
	    RECT 113.2000 133.8000 114.2000 134.2000 ;
	    RECT 115.2000 134.4000 115.8000 135.0000 ;
	    RECT 121.2000 134.4000 121.8000 135.8000 ;
	    RECT 123.0000 135.4000 126.6000 135.8000 ;
	    RECT 125.2000 134.4000 126.0000 134.8000 ;
	    RECT 127.8000 134.4000 128.4000 135.8000 ;
	    RECT 129.4000 135.4000 133.0000 135.8000 ;
	    RECT 131.6000 134.4000 132.4000 134.8000 ;
	    RECT 135.6000 134.4000 136.2000 135.8000 ;
	    RECT 137.4000 135.4000 141.0000 135.8000 ;
	    RECT 143.6000 135.6000 144.4000 138.6000 ;
	    RECT 145.2000 136.0000 146.0000 139.2000 ;
	    RECT 148.4000 136.0000 149.2000 139.8000 ;
	    RECT 145.2000 135.8000 149.2000 136.0000 ;
	    RECT 150.0000 136.0000 150.8000 139.8000 ;
	    RECT 153.2000 136.0000 154.0000 139.8000 ;
	    RECT 150.0000 135.8000 154.0000 136.0000 ;
	    RECT 154.8000 135.8000 155.6000 139.8000 ;
	    RECT 139.6000 134.4000 140.4000 134.8000 ;
	    RECT 143.6000 134.4000 144.2000 135.6000 ;
	    RECT 145.4000 135.4000 149.0000 135.8000 ;
	    RECT 150.2000 135.4000 153.8000 135.8000 ;
	    RECT 147.6000 134.4000 148.4000 134.8000 ;
	    RECT 150.8000 134.4000 151.6000 134.8000 ;
	    RECT 154.8000 134.4000 155.4000 135.8000 ;
	    RECT 66.8000 131.7000 70.8000 132.3000 ;
	    RECT 66.8000 131.6000 67.6000 131.7000 ;
	    RECT 62.0000 129.6000 63.4000 130.2000 ;
	    RECT 64.0000 129.6000 65.0000 130.2000 ;
	    RECT 62.8000 128.4000 63.4000 129.6000 ;
	    RECT 62.8000 127.6000 63.6000 128.4000 ;
	    RECT 64.2000 122.2000 65.0000 129.6000 ;
	    RECT 70.0000 122.2000 70.8000 131.7000 ;
	    RECT 71.6000 132.3000 72.4000 132.4000 ;
	    RECT 75.2000 132.3000 75.8000 133.6000 ;
	    RECT 71.6000 131.7000 75.8000 132.3000 ;
	    RECT 71.6000 131.6000 72.4000 131.7000 ;
	    RECT 73.2000 130.2000 74.0000 130.4000 ;
	    RECT 75.2000 130.2000 75.8000 131.7000 ;
	    RECT 76.4000 132.3000 77.2000 133.2000 ;
	    RECT 79.6000 132.3000 80.4000 132.4000 ;
	    RECT 76.4000 131.7000 80.4000 132.3000 ;
	    RECT 76.4000 131.6000 77.2000 131.7000 ;
	    RECT 79.6000 131.6000 80.4000 131.7000 ;
	    RECT 81.4000 130.2000 82.0000 133.6000 ;
	    RECT 82.8000 130.8000 83.6000 132.4000 ;
	    RECT 84.4000 130.2000 85.2000 130.4000 ;
	    RECT 86.4000 130.2000 87.0000 133.6000 ;
	    RECT 87.6000 131.6000 88.4000 133.2000 ;
	    RECT 90.8000 130.2000 91.6000 130.4000 ;
	    RECT 92.8000 130.2000 93.4000 133.6000 ;
	    RECT 94.0000 131.6000 94.8000 133.2000 ;
	    RECT 98.8000 131.6000 99.6000 133.2000 ;
	    RECT 100.2000 132.4000 100.8000 133.6000 ;
	    RECT 100.2000 131.6000 101.2000 132.4000 ;
	    RECT 110.0000 131.6000 110.8000 133.2000 ;
	    RECT 111.6000 131.6000 112.4000 133.2000 ;
	    RECT 113.2000 133.0000 114.6000 133.8000 ;
	    RECT 115.2000 133.6000 117.2000 134.4000 ;
	    RECT 118.0000 134.3000 118.8000 134.4000 ;
	    RECT 119.6000 134.3000 120.4000 134.4000 ;
	    RECT 118.0000 133.7000 120.4000 134.3000 ;
	    RECT 121.2000 133.8000 123.6000 134.4000 ;
	    RECT 125.2000 134.3000 126.8000 134.4000 ;
	    RECT 127.6000 134.3000 130.2000 134.4000 ;
	    RECT 125.2000 133.8000 130.2000 134.3000 ;
	    RECT 131.6000 133.8000 133.2000 134.4000 ;
	    RECT 118.0000 133.6000 118.8000 133.7000 ;
	    RECT 100.2000 130.2000 100.8000 131.6000 ;
	    RECT 113.2000 131.0000 113.8000 133.0000 ;
	    RECT 115.2000 132.4000 115.8000 133.6000 ;
	    RECT 119.6000 132.8000 120.4000 133.7000 ;
	    RECT 122.8000 133.6000 123.6000 133.8000 ;
	    RECT 126.0000 133.7000 130.2000 133.8000 ;
	    RECT 126.0000 133.6000 126.8000 133.7000 ;
	    RECT 127.6000 133.6000 130.2000 133.7000 ;
	    RECT 132.4000 133.6000 133.2000 133.8000 ;
	    RECT 114.8000 131.6000 115.8000 132.4000 ;
	    RECT 110.0000 130.4000 113.8000 131.0000 ;
	    RECT 102.0000 130.2000 102.8000 130.4000 ;
	    RECT 73.2000 129.6000 74.6000 130.2000 ;
	    RECT 75.2000 129.6000 76.2000 130.2000 ;
	    RECT 74.0000 128.4000 74.6000 129.6000 ;
	    RECT 74.0000 127.6000 74.8000 128.4000 ;
	    RECT 75.4000 122.2000 76.2000 129.6000 ;
	    RECT 81.2000 129.4000 83.0000 130.2000 ;
	    RECT 84.4000 129.6000 85.8000 130.2000 ;
	    RECT 86.4000 129.6000 87.4000 130.2000 ;
	    RECT 90.8000 129.6000 92.2000 130.2000 ;
	    RECT 92.8000 129.6000 93.8000 130.2000 ;
	    RECT 82.2000 124.4000 83.0000 129.4000 ;
	    RECT 85.2000 128.4000 85.8000 129.6000 ;
	    RECT 85.2000 127.6000 86.0000 128.4000 ;
	    RECT 81.2000 123.6000 83.0000 124.4000 ;
	    RECT 82.2000 122.2000 83.0000 123.6000 ;
	    RECT 86.6000 122.2000 87.4000 129.6000 ;
	    RECT 91.6000 128.4000 92.2000 129.6000 ;
	    RECT 93.0000 128.4000 93.8000 129.6000 ;
	    RECT 99.8000 129.6000 100.8000 130.2000 ;
	    RECT 101.4000 129.6000 102.8000 130.2000 ;
	    RECT 91.6000 127.6000 92.4000 128.4000 ;
	    RECT 93.0000 127.6000 94.8000 128.4000 ;
	    RECT 93.0000 122.2000 93.8000 127.6000 ;
	    RECT 99.8000 122.2000 100.6000 129.6000 ;
	    RECT 101.4000 128.4000 102.0000 129.6000 ;
	    RECT 101.2000 127.6000 102.0000 128.4000 ;
	    RECT 110.0000 127.0000 110.6000 130.4000 ;
	    RECT 115.2000 129.8000 115.8000 131.6000 ;
	    RECT 116.4000 130.8000 117.2000 132.4000 ;
	    RECT 121.2000 131.6000 122.0000 133.2000 ;
	    RECT 123.0000 130.2000 123.6000 133.6000 ;
	    RECT 124.4000 132.3000 125.2000 133.2000 ;
	    RECT 127.6000 132.3000 128.4000 132.4000 ;
	    RECT 124.4000 131.7000 128.4000 132.3000 ;
	    RECT 124.4000 131.6000 125.2000 131.7000 ;
	    RECT 127.6000 131.6000 128.4000 131.7000 ;
	    RECT 127.6000 130.2000 128.4000 130.4000 ;
	    RECT 129.6000 130.2000 130.2000 133.6000 ;
	    RECT 130.8000 131.6000 131.6000 133.2000 ;
	    RECT 134.0000 132.8000 134.8000 134.4000 ;
	    RECT 135.6000 133.8000 138.0000 134.4000 ;
	    RECT 139.6000 133.8000 141.2000 134.4000 ;
	    RECT 137.2000 133.6000 138.0000 133.8000 ;
	    RECT 140.4000 133.6000 141.2000 133.8000 ;
	    RECT 135.6000 131.6000 136.4000 133.2000 ;
	    RECT 137.4000 130.2000 138.0000 133.6000 ;
	    RECT 138.8000 131.6000 139.6000 133.2000 ;
	    RECT 142.0000 132.8000 142.8000 134.4000 ;
	    RECT 143.6000 133.8000 146.0000 134.4000 ;
	    RECT 147.6000 133.8000 149.2000 134.4000 ;
	    RECT 145.2000 133.6000 146.0000 133.8000 ;
	    RECT 148.4000 133.6000 149.2000 133.8000 ;
	    RECT 150.0000 133.8000 151.6000 134.4000 ;
	    RECT 150.0000 133.6000 150.8000 133.8000 ;
	    RECT 153.0000 133.6000 155.6000 134.4000 ;
	    RECT 143.6000 131.6000 144.4000 133.2000 ;
	    RECT 145.4000 130.2000 146.0000 133.6000 ;
	    RECT 146.8000 132.3000 147.6000 133.2000 ;
	    RECT 150.0000 132.3000 150.8000 132.4000 ;
	    RECT 146.8000 131.7000 150.8000 132.3000 ;
	    RECT 146.8000 131.6000 147.6000 131.7000 ;
	    RECT 150.0000 131.6000 150.8000 131.7000 ;
	    RECT 151.6000 131.6000 152.4000 133.2000 ;
	    RECT 153.0000 130.2000 153.6000 133.6000 ;
	    RECT 156.4000 132.4000 157.2000 139.8000 ;
	    RECT 159.6000 135.2000 160.4000 139.8000 ;
	    RECT 158.2000 134.6000 160.4000 135.2000 ;
	    RECT 162.8000 137.8000 163.6000 139.8000 ;
	    RECT 167.6000 137.8000 168.4000 139.8000 ;
	    RECT 154.8000 130.2000 155.6000 130.4000 ;
	    RECT 114.2000 129.2000 115.8000 129.8000 ;
	    RECT 110.0000 123.0000 110.8000 127.0000 ;
	    RECT 114.2000 122.2000 115.0000 129.2000 ;
	    RECT 122.2000 128.4000 124.2000 130.2000 ;
	    RECT 127.6000 129.6000 129.0000 130.2000 ;
	    RECT 129.6000 129.6000 130.6000 130.2000 ;
	    RECT 121.2000 127.6000 124.2000 128.4000 ;
	    RECT 128.4000 128.4000 129.0000 129.6000 ;
	    RECT 128.4000 127.6000 129.2000 128.4000 ;
	    RECT 122.2000 122.2000 124.2000 127.6000 ;
	    RECT 129.8000 122.2000 130.6000 129.6000 ;
	    RECT 136.6000 122.2000 138.6000 130.2000 ;
	    RECT 144.6000 122.2000 146.6000 130.2000 ;
	    RECT 152.6000 129.6000 153.6000 130.2000 ;
	    RECT 154.2000 129.6000 155.6000 130.2000 ;
	    RECT 156.4000 130.2000 157.0000 132.4000 ;
	    RECT 158.2000 131.6000 158.8000 134.6000 ;
	    RECT 162.8000 134.4000 163.4000 137.8000 ;
	    RECT 164.4000 136.3000 165.2000 137.2000 ;
	    RECT 166.0000 136.3000 166.8000 137.2000 ;
	    RECT 164.4000 135.7000 166.8000 136.3000 ;
	    RECT 164.4000 135.6000 165.2000 135.7000 ;
	    RECT 166.0000 135.6000 166.8000 135.7000 ;
	    RECT 167.8000 134.4000 168.4000 137.8000 ;
	    RECT 161.2000 134.3000 162.0000 134.4000 ;
	    RECT 162.8000 134.3000 163.6000 134.4000 ;
	    RECT 161.2000 133.7000 163.6000 134.3000 ;
	    RECT 161.2000 133.6000 162.0000 133.7000 ;
	    RECT 162.8000 133.6000 163.6000 133.7000 ;
	    RECT 167.6000 133.6000 168.4000 134.4000 ;
	    RECT 157.6000 130.8000 158.8000 131.6000 ;
	    RECT 161.2000 130.8000 162.0000 132.4000 ;
	    RECT 158.2000 130.2000 158.8000 130.8000 ;
	    RECT 162.8000 130.2000 163.4000 133.6000 ;
	    RECT 167.8000 130.4000 168.4000 133.6000 ;
	    RECT 172.4000 137.6000 173.2000 139.8000 ;
	    RECT 177.2000 137.8000 178.0000 139.8000 ;
	    RECT 172.4000 134.4000 173.0000 137.6000 ;
	    RECT 174.0000 135.6000 174.8000 137.2000 ;
	    RECT 177.2000 134.4000 177.8000 137.8000 ;
	    RECT 178.8000 135.6000 179.6000 137.2000 ;
	    RECT 172.4000 133.6000 173.2000 134.4000 ;
	    RECT 174.0000 134.3000 174.8000 134.4000 ;
	    RECT 177.2000 134.3000 178.0000 134.4000 ;
	    RECT 174.0000 133.7000 178.0000 134.3000 ;
	    RECT 174.0000 133.6000 174.8000 133.7000 ;
	    RECT 177.2000 133.6000 178.0000 133.7000 ;
	    RECT 169.2000 130.8000 170.0000 132.4000 ;
	    RECT 170.8000 130.8000 171.6000 132.4000 ;
	    RECT 167.6000 130.2000 168.4000 130.4000 ;
	    RECT 172.4000 130.2000 173.0000 133.6000 ;
	    RECT 175.6000 130.8000 176.4000 132.4000 ;
	    RECT 177.2000 130.2000 177.8000 133.6000 ;
	    RECT 180.4000 132.4000 181.2000 139.8000 ;
	    RECT 183.6000 135.2000 184.4000 139.8000 ;
	    RECT 182.2000 134.6000 184.4000 135.2000 ;
	    RECT 180.4000 130.2000 181.0000 132.4000 ;
	    RECT 182.2000 131.6000 182.8000 134.6000 ;
	    RECT 181.6000 130.8000 182.8000 131.6000 ;
	    RECT 182.2000 130.2000 182.8000 130.8000 ;
	    RECT 185.2000 132.4000 186.0000 139.8000 ;
	    RECT 188.4000 135.2000 189.2000 139.8000 ;
	    RECT 187.0000 134.6000 189.2000 135.2000 ;
	    RECT 185.2000 130.2000 185.8000 132.4000 ;
	    RECT 187.0000 131.6000 187.6000 134.6000 ;
	    RECT 186.4000 130.8000 187.6000 131.6000 ;
	    RECT 187.0000 130.2000 187.6000 130.8000 ;
	    RECT 190.0000 132.4000 190.8000 139.8000 ;
	    RECT 193.2000 135.2000 194.0000 139.8000 ;
	    RECT 191.8000 134.6000 194.0000 135.2000 ;
	    RECT 190.0000 130.2000 190.6000 132.4000 ;
	    RECT 191.8000 131.6000 192.4000 134.6000 ;
	    RECT 191.2000 130.8000 192.4000 131.6000 ;
	    RECT 191.8000 130.2000 192.4000 130.8000 ;
	    RECT 194.8000 132.4000 195.6000 139.8000 ;
	    RECT 198.0000 135.2000 198.8000 139.8000 ;
	    RECT 199.6000 136.0000 200.4000 139.8000 ;
	    RECT 202.8000 136.0000 203.6000 139.8000 ;
	    RECT 199.6000 135.8000 203.6000 136.0000 ;
	    RECT 204.4000 135.8000 205.2000 139.8000 ;
	    RECT 206.0000 136.0000 206.8000 139.8000 ;
	    RECT 209.2000 136.0000 210.0000 139.8000 ;
	    RECT 206.0000 135.8000 210.0000 136.0000 ;
	    RECT 210.8000 135.8000 211.6000 139.8000 ;
	    RECT 212.4000 135.8000 213.2000 139.8000 ;
	    RECT 214.0000 136.0000 214.8000 139.8000 ;
	    RECT 217.2000 136.0000 218.0000 139.8000 ;
	    RECT 214.0000 135.8000 218.0000 136.0000 ;
	    RECT 199.8000 135.4000 203.4000 135.8000 ;
	    RECT 196.6000 134.6000 198.8000 135.2000 ;
	    RECT 194.8000 130.2000 195.4000 132.4000 ;
	    RECT 196.6000 131.6000 197.2000 134.6000 ;
	    RECT 200.4000 134.4000 201.2000 134.8000 ;
	    RECT 204.4000 134.4000 205.0000 135.8000 ;
	    RECT 206.2000 135.4000 209.8000 135.8000 ;
	    RECT 206.8000 134.4000 207.6000 134.8000 ;
	    RECT 210.8000 134.4000 211.4000 135.8000 ;
	    RECT 212.6000 134.4000 213.2000 135.8000 ;
	    RECT 214.2000 135.4000 217.8000 135.8000 ;
	    RECT 218.8000 135.4000 219.6000 139.8000 ;
	    RECT 223.0000 138.4000 224.2000 139.8000 ;
	    RECT 223.0000 137.8000 224.4000 138.4000 ;
	    RECT 227.6000 137.8000 228.4000 139.8000 ;
	    RECT 232.0000 138.4000 232.8000 139.8000 ;
	    RECT 232.0000 137.8000 234.0000 138.4000 ;
	    RECT 223.6000 137.0000 224.4000 137.8000 ;
	    RECT 227.8000 137.2000 228.4000 137.8000 ;
	    RECT 227.8000 136.6000 230.6000 137.2000 ;
	    RECT 229.8000 136.4000 230.6000 136.6000 ;
	    RECT 231.6000 135.6000 232.4000 137.2000 ;
	    RECT 233.2000 137.0000 234.0000 137.8000 ;
	    RECT 221.8000 135.4000 222.6000 135.6000 ;
	    RECT 218.8000 134.8000 222.6000 135.4000 ;
	    RECT 216.4000 134.4000 217.2000 134.8000 ;
	    RECT 199.6000 133.8000 201.2000 134.4000 ;
	    RECT 199.6000 133.6000 200.4000 133.8000 ;
	    RECT 202.6000 133.6000 205.2000 134.4000 ;
	    RECT 206.0000 133.8000 207.6000 134.4000 ;
	    RECT 206.0000 133.6000 206.8000 133.8000 ;
	    RECT 209.0000 133.6000 211.6000 134.4000 ;
	    RECT 212.4000 133.6000 215.0000 134.4000 ;
	    RECT 216.4000 133.8000 218.0000 134.4000 ;
	    RECT 217.2000 133.6000 218.0000 133.8000 ;
	    RECT 198.0000 132.3000 198.8000 133.2000 ;
	    RECT 199.6000 132.3000 200.4000 132.4000 ;
	    RECT 198.0000 131.7000 200.4000 132.3000 ;
	    RECT 198.0000 131.6000 198.8000 131.7000 ;
	    RECT 199.6000 131.6000 200.4000 131.7000 ;
	    RECT 201.2000 131.6000 202.0000 133.2000 ;
	    RECT 196.0000 130.8000 197.2000 131.6000 ;
	    RECT 196.6000 130.2000 197.2000 130.8000 ;
	    RECT 202.6000 130.2000 203.2000 133.6000 ;
	    RECT 207.6000 131.6000 208.4000 133.2000 ;
	    RECT 209.0000 132.3000 209.6000 133.6000 ;
	    RECT 209.0000 131.7000 213.1000 132.3000 ;
	    RECT 204.4000 130.2000 205.2000 130.4000 ;
	    RECT 209.0000 130.2000 209.6000 131.7000 ;
	    RECT 212.5000 130.4000 213.1000 131.7000 ;
	    RECT 210.8000 130.2000 211.6000 130.4000 ;
	    RECT 152.6000 128.4000 153.4000 129.6000 ;
	    RECT 154.2000 128.4000 154.8000 129.6000 ;
	    RECT 151.6000 127.6000 153.4000 128.4000 ;
	    RECT 154.0000 127.6000 154.8000 128.4000 ;
	    RECT 152.6000 122.2000 153.4000 127.6000 ;
	    RECT 156.4000 122.2000 157.2000 130.2000 ;
	    RECT 158.2000 129.6000 160.4000 130.2000 ;
	    RECT 159.6000 122.2000 160.4000 129.6000 ;
	    RECT 161.8000 129.4000 163.6000 130.2000 ;
	    RECT 167.6000 129.4000 169.4000 130.2000 ;
	    RECT 161.8000 122.2000 162.6000 129.4000 ;
	    RECT 168.6000 122.2000 169.4000 129.4000 ;
	    RECT 171.4000 129.4000 173.2000 130.2000 ;
	    RECT 176.2000 129.4000 178.0000 130.2000 ;
	    RECT 171.4000 122.2000 172.2000 129.4000 ;
	    RECT 176.2000 122.2000 177.0000 129.4000 ;
	    RECT 180.4000 122.2000 181.2000 130.2000 ;
	    RECT 182.2000 129.6000 184.4000 130.2000 ;
	    RECT 183.6000 122.2000 184.4000 129.6000 ;
	    RECT 185.2000 122.2000 186.0000 130.2000 ;
	    RECT 187.0000 129.6000 189.2000 130.2000 ;
	    RECT 188.4000 122.2000 189.2000 129.6000 ;
	    RECT 190.0000 122.2000 190.8000 130.2000 ;
	    RECT 191.8000 129.6000 194.0000 130.2000 ;
	    RECT 193.2000 122.2000 194.0000 129.6000 ;
	    RECT 194.8000 122.2000 195.6000 130.2000 ;
	    RECT 196.6000 129.6000 198.8000 130.2000 ;
	    RECT 198.0000 122.2000 198.8000 129.6000 ;
	    RECT 202.2000 129.6000 203.2000 130.2000 ;
	    RECT 203.8000 129.6000 205.2000 130.2000 ;
	    RECT 208.6000 129.6000 209.6000 130.2000 ;
	    RECT 210.2000 129.6000 211.6000 130.2000 ;
	    RECT 212.4000 130.2000 213.2000 130.4000 ;
	    RECT 214.4000 130.2000 215.0000 133.6000 ;
	    RECT 215.6000 131.6000 216.4000 133.2000 ;
	    RECT 218.8000 131.4000 219.6000 134.8000 ;
	    RECT 225.8000 134.2000 226.6000 134.4000 ;
	    RECT 231.6000 134.2000 232.2000 135.6000 ;
	    RECT 236.4000 135.0000 237.2000 139.8000 ;
	    RECT 238.0000 135.2000 238.8000 139.8000 ;
	    RECT 238.0000 134.6000 240.2000 135.2000 ;
	    RECT 234.8000 134.2000 236.4000 134.4000 ;
	    RECT 225.4000 133.6000 236.4000 134.2000 ;
	    RECT 223.6000 132.8000 224.4000 133.0000 ;
	    RECT 220.6000 132.2000 224.4000 132.8000 ;
	    RECT 220.6000 132.0000 221.4000 132.2000 ;
	    RECT 222.2000 131.4000 223.0000 131.6000 ;
	    RECT 218.8000 130.8000 223.0000 131.4000 ;
	    RECT 212.4000 129.6000 213.8000 130.2000 ;
	    RECT 214.4000 129.6000 215.4000 130.2000 ;
	    RECT 202.2000 124.4000 203.0000 129.6000 ;
	    RECT 203.8000 128.4000 204.4000 129.6000 ;
	    RECT 203.6000 127.6000 205.2000 128.4000 ;
	    RECT 201.2000 123.6000 203.0000 124.4000 ;
	    RECT 202.2000 122.2000 203.0000 123.6000 ;
	    RECT 208.6000 122.2000 209.4000 129.6000 ;
	    RECT 210.2000 128.4000 210.8000 129.6000 ;
	    RECT 213.2000 128.4000 213.8000 129.6000 ;
	    RECT 210.0000 127.6000 211.6000 128.4000 ;
	    RECT 213.2000 127.6000 214.0000 128.4000 ;
	    RECT 214.6000 126.4000 215.4000 129.6000 ;
	    RECT 214.6000 125.6000 216.4000 126.4000 ;
	    RECT 214.6000 122.2000 215.4000 125.6000 ;
	    RECT 218.8000 122.2000 219.6000 130.8000 ;
	    RECT 225.4000 130.4000 226.0000 133.6000 ;
	    RECT 232.6000 133.4000 233.4000 133.6000 ;
	    RECT 234.2000 132.4000 235.0000 132.6000 ;
	    RECT 228.4000 132.3000 229.2000 132.4000 ;
	    RECT 230.0000 132.3000 235.0000 132.4000 ;
	    RECT 228.4000 131.8000 235.0000 132.3000 ;
	    RECT 228.4000 131.7000 230.8000 131.8000 ;
	    RECT 228.4000 131.6000 229.2000 131.7000 ;
	    RECT 230.0000 131.6000 230.8000 131.7000 ;
	    RECT 238.0000 131.6000 238.8000 133.2000 ;
	    RECT 239.6000 131.6000 240.2000 134.6000 ;
	    RECT 241.2000 132.4000 242.0000 139.8000 ;
	    RECT 231.6000 131.0000 237.2000 131.2000 ;
	    RECT 231.4000 130.8000 237.2000 131.0000 ;
	    RECT 223.6000 129.8000 226.0000 130.4000 ;
	    RECT 227.4000 130.6000 237.2000 130.8000 ;
	    RECT 227.4000 130.2000 232.2000 130.6000 ;
	    RECT 223.6000 128.8000 224.2000 129.8000 ;
	    RECT 222.8000 128.0000 224.2000 128.8000 ;
	    RECT 225.8000 129.0000 226.6000 129.2000 ;
	    RECT 227.4000 129.0000 228.0000 130.2000 ;
	    RECT 225.8000 128.4000 228.0000 129.0000 ;
	    RECT 228.6000 129.0000 234.0000 129.6000 ;
	    RECT 228.6000 128.8000 229.4000 129.0000 ;
	    RECT 233.2000 128.8000 234.0000 129.0000 ;
	    RECT 227.0000 127.4000 227.8000 127.6000 ;
	    RECT 229.8000 127.4000 230.6000 127.6000 ;
	    RECT 223.6000 126.2000 224.4000 127.0000 ;
	    RECT 227.0000 126.8000 230.6000 127.4000 ;
	    RECT 227.8000 126.2000 228.4000 126.8000 ;
	    RECT 233.2000 126.2000 234.0000 127.0000 ;
	    RECT 223.0000 122.2000 224.2000 126.2000 ;
	    RECT 227.6000 122.2000 228.4000 126.2000 ;
	    RECT 232.0000 125.6000 234.0000 126.2000 ;
	    RECT 232.0000 122.2000 232.8000 125.6000 ;
	    RECT 236.4000 122.2000 237.2000 130.6000 ;
	    RECT 239.6000 130.8000 240.8000 131.6000 ;
	    RECT 239.6000 130.2000 240.2000 130.8000 ;
	    RECT 241.4000 130.2000 242.0000 132.4000 ;
	    RECT 238.0000 129.6000 240.2000 130.2000 ;
	    RECT 238.0000 122.2000 238.8000 129.6000 ;
	    RECT 241.2000 122.2000 242.0000 130.2000 ;
	    RECT 242.8000 132.4000 243.6000 139.8000 ;
	    RECT 246.0000 135.2000 246.8000 139.8000 ;
	    RECT 247.6000 136.0000 248.4000 139.8000 ;
	    RECT 250.8000 136.0000 251.6000 139.8000 ;
	    RECT 247.6000 135.8000 251.6000 136.0000 ;
	    RECT 252.4000 135.8000 253.2000 139.8000 ;
	    RECT 260.4000 135.8000 261.2000 139.8000 ;
	    RECT 262.0000 136.0000 262.8000 139.8000 ;
	    RECT 265.2000 136.0000 266.0000 139.8000 ;
	    RECT 262.0000 135.8000 266.0000 136.0000 ;
	    RECT 247.8000 135.4000 251.4000 135.8000 ;
	    RECT 244.6000 134.6000 246.8000 135.2000 ;
	    RECT 242.8000 130.2000 243.4000 132.4000 ;
	    RECT 244.6000 131.6000 245.2000 134.6000 ;
	    RECT 248.4000 134.4000 249.2000 134.8000 ;
	    RECT 252.4000 134.4000 253.0000 135.8000 ;
	    RECT 260.6000 134.4000 261.2000 135.8000 ;
	    RECT 262.2000 135.4000 265.8000 135.8000 ;
	    RECT 266.8000 135.2000 267.6000 139.8000 ;
	    RECT 264.4000 134.4000 265.2000 134.8000 ;
	    RECT 266.8000 134.6000 269.0000 135.2000 ;
	    RECT 247.6000 133.8000 249.2000 134.4000 ;
	    RECT 247.6000 133.6000 248.4000 133.8000 ;
	    RECT 250.6000 133.6000 253.2000 134.4000 ;
	    RECT 258.8000 134.3000 259.6000 134.4000 ;
	    RECT 260.4000 134.3000 263.0000 134.4000 ;
	    RECT 258.8000 133.7000 263.0000 134.3000 ;
	    RECT 264.4000 133.8000 266.0000 134.4000 ;
	    RECT 258.8000 133.6000 259.6000 133.7000 ;
	    RECT 260.4000 133.6000 263.0000 133.7000 ;
	    RECT 265.2000 133.6000 266.0000 133.8000 ;
	    RECT 246.0000 131.6000 246.8000 133.2000 ;
	    RECT 249.2000 131.6000 250.0000 133.2000 ;
	    RECT 250.6000 132.3000 251.2000 133.6000 ;
	    RECT 250.6000 131.7000 261.1000 132.3000 ;
	    RECT 244.0000 130.8000 245.2000 131.6000 ;
	    RECT 244.6000 130.2000 245.2000 130.8000 ;
	    RECT 250.6000 130.2000 251.2000 131.7000 ;
	    RECT 260.5000 130.4000 261.1000 131.7000 ;
	    RECT 252.4000 130.2000 253.2000 130.4000 ;
	    RECT 242.8000 122.2000 243.6000 130.2000 ;
	    RECT 244.6000 129.6000 246.8000 130.2000 ;
	    RECT 246.0000 122.2000 246.8000 129.6000 ;
	    RECT 250.2000 129.6000 251.2000 130.2000 ;
	    RECT 251.8000 129.6000 253.2000 130.2000 ;
	    RECT 260.4000 130.2000 261.2000 130.4000 ;
	    RECT 262.4000 130.2000 263.0000 133.6000 ;
	    RECT 263.6000 131.6000 264.4000 133.2000 ;
	    RECT 266.8000 131.6000 267.6000 133.2000 ;
	    RECT 268.4000 131.6000 269.0000 134.6000 ;
	    RECT 270.0000 132.4000 270.8000 139.8000 ;
	    RECT 273.2000 135.2000 274.0000 139.8000 ;
	    RECT 276.4000 135.2000 277.2000 139.8000 ;
	    RECT 271.6000 133.6000 272.4000 135.2000 ;
	    RECT 273.2000 134.4000 277.2000 135.2000 ;
	    RECT 279.6000 135.2000 280.4000 139.8000 ;
	    RECT 279.6000 134.6000 281.8000 135.2000 ;
	    RECT 268.4000 130.8000 269.6000 131.6000 ;
	    RECT 268.4000 130.2000 269.0000 130.8000 ;
	    RECT 270.2000 130.2000 270.8000 132.4000 ;
	    RECT 276.4000 131.6000 277.2000 134.4000 ;
	    RECT 260.4000 129.6000 261.8000 130.2000 ;
	    RECT 262.4000 129.6000 263.4000 130.2000 ;
	    RECT 250.2000 122.2000 251.0000 129.6000 ;
	    RECT 251.8000 128.4000 252.4000 129.6000 ;
	    RECT 251.6000 127.6000 252.4000 128.4000 ;
	    RECT 261.2000 128.4000 261.8000 129.6000 ;
	    RECT 261.2000 127.6000 262.0000 128.4000 ;
	    RECT 262.6000 122.2000 263.4000 129.6000 ;
	    RECT 266.8000 129.6000 269.0000 130.2000 ;
	    RECT 266.8000 122.2000 267.6000 129.6000 ;
	    RECT 270.0000 122.2000 270.8000 130.2000 ;
	    RECT 273.2000 130.8000 277.2000 131.6000 ;
	    RECT 273.2000 122.2000 274.0000 130.8000 ;
	    RECT 276.4000 122.2000 277.2000 130.8000 ;
	    RECT 281.2000 131.6000 281.8000 134.6000 ;
	    RECT 282.8000 132.4000 283.6000 139.8000 ;
	    RECT 286.0000 137.8000 286.8000 139.8000 ;
	    RECT 290.8000 137.8000 291.6000 139.8000 ;
	    RECT 294.0000 139.2000 298.0000 139.8000 ;
	    RECT 286.0000 134.4000 286.6000 137.8000 ;
	    RECT 287.6000 135.6000 288.4000 137.2000 ;
	    RECT 290.8000 134.4000 291.4000 137.8000 ;
	    RECT 292.4000 135.6000 293.2000 137.2000 ;
	    RECT 294.0000 135.8000 294.8000 139.2000 ;
	    RECT 295.6000 135.8000 296.4000 138.6000 ;
	    RECT 297.2000 136.0000 298.0000 139.2000 ;
	    RECT 300.4000 136.0000 301.2000 139.8000 ;
	    RECT 297.2000 135.8000 301.2000 136.0000 ;
	    RECT 303.6000 137.8000 304.4000 139.8000 ;
	    RECT 295.6000 134.4000 296.2000 135.8000 ;
	    RECT 297.4000 135.4000 301.0000 135.8000 ;
	    RECT 299.6000 134.4000 300.4000 134.8000 ;
	    RECT 303.6000 134.4000 304.2000 137.8000 ;
	    RECT 305.2000 135.6000 306.0000 137.2000 ;
	    RECT 306.8000 135.8000 307.6000 139.8000 ;
	    RECT 308.4000 136.0000 309.2000 139.8000 ;
	    RECT 311.6000 136.0000 312.4000 139.8000 ;
	    RECT 314.8000 137.8000 315.6000 139.8000 ;
	    RECT 308.4000 135.8000 312.4000 136.0000 ;
	    RECT 307.0000 134.4000 307.6000 135.8000 ;
	    RECT 308.6000 135.4000 312.2000 135.8000 ;
	    RECT 313.2000 135.6000 314.0000 137.2000 ;
	    RECT 310.8000 134.4000 311.6000 134.8000 ;
	    RECT 315.0000 134.4000 315.6000 137.8000 ;
	    RECT 318.0000 136.0000 318.8000 139.8000 ;
	    RECT 321.2000 139.2000 325.2000 139.8000 ;
	    RECT 321.2000 136.0000 322.0000 139.2000 ;
	    RECT 318.0000 135.8000 322.0000 136.0000 ;
	    RECT 322.8000 135.8000 323.6000 138.6000 ;
	    RECT 324.4000 135.8000 325.2000 139.2000 ;
	    RECT 326.0000 135.8000 326.8000 139.8000 ;
	    RECT 327.6000 136.0000 328.4000 139.8000 ;
	    RECT 330.8000 136.0000 331.6000 139.8000 ;
	    RECT 327.6000 135.8000 331.6000 136.0000 ;
	    RECT 318.2000 135.4000 321.8000 135.8000 ;
	    RECT 318.8000 134.4000 319.6000 134.8000 ;
	    RECT 323.0000 134.4000 323.6000 135.8000 ;
	    RECT 326.2000 134.4000 326.8000 135.8000 ;
	    RECT 327.8000 135.4000 331.4000 135.8000 ;
	    RECT 332.4000 135.2000 333.2000 139.8000 ;
	    RECT 330.0000 134.4000 330.8000 134.8000 ;
	    RECT 332.4000 134.6000 334.6000 135.2000 ;
	    RECT 286.0000 133.6000 286.8000 134.4000 ;
	    RECT 290.8000 133.6000 291.6000 134.4000 ;
	    RECT 281.2000 130.8000 282.4000 131.6000 ;
	    RECT 281.2000 130.2000 281.8000 130.8000 ;
	    RECT 283.0000 130.2000 283.6000 132.4000 ;
	    RECT 284.4000 130.8000 285.2000 132.4000 ;
	    RECT 286.0000 130.2000 286.6000 133.6000 ;
	    RECT 289.2000 130.8000 290.0000 132.4000 ;
	    RECT 290.8000 130.4000 291.4000 133.6000 ;
	    RECT 294.0000 132.8000 294.8000 134.4000 ;
	    RECT 295.6000 133.8000 298.0000 134.4000 ;
	    RECT 299.6000 133.8000 301.2000 134.4000 ;
	    RECT 297.2000 133.6000 298.0000 133.8000 ;
	    RECT 300.4000 133.6000 301.2000 133.8000 ;
	    RECT 303.6000 133.6000 304.4000 134.4000 ;
	    RECT 305.2000 134.3000 306.0000 134.4000 ;
	    RECT 306.8000 134.3000 309.4000 134.4000 ;
	    RECT 305.2000 133.7000 309.4000 134.3000 ;
	    RECT 310.8000 133.8000 312.4000 134.4000 ;
	    RECT 305.2000 133.6000 306.0000 133.7000 ;
	    RECT 306.8000 133.6000 309.4000 133.7000 ;
	    RECT 311.6000 133.6000 312.4000 133.8000 ;
	    RECT 314.8000 133.6000 315.6000 134.4000 ;
	    RECT 318.0000 133.8000 319.6000 134.4000 ;
	    RECT 321.2000 133.8000 323.6000 134.4000 ;
	    RECT 318.0000 133.6000 318.8000 133.8000 ;
	    RECT 321.2000 133.6000 322.0000 133.8000 ;
	    RECT 295.6000 131.6000 296.4000 133.2000 ;
	    RECT 297.4000 132.4000 298.0000 133.6000 ;
	    RECT 297.2000 131.6000 298.0000 132.4000 ;
	    RECT 298.8000 132.3000 299.6000 133.2000 ;
	    RECT 300.4000 132.3000 301.2000 132.4000 ;
	    RECT 298.8000 131.7000 301.2000 132.3000 ;
	    RECT 298.8000 131.6000 299.6000 131.7000 ;
	    RECT 300.4000 131.6000 301.2000 131.7000 ;
	    RECT 290.8000 130.2000 291.6000 130.4000 ;
	    RECT 297.4000 130.2000 298.0000 131.6000 ;
	    RECT 302.0000 130.8000 302.8000 132.4000 ;
	    RECT 303.6000 130.2000 304.2000 133.6000 ;
	    RECT 306.8000 130.2000 307.6000 130.4000 ;
	    RECT 308.8000 130.2000 309.4000 133.6000 ;
	    RECT 310.0000 131.6000 310.8000 133.2000 ;
	    RECT 315.0000 130.2000 315.6000 133.6000 ;
	    RECT 316.4000 130.8000 317.2000 132.4000 ;
	    RECT 319.6000 131.6000 320.4000 133.2000 ;
	    RECT 321.2000 130.2000 321.8000 133.6000 ;
	    RECT 322.8000 131.6000 323.6000 133.2000 ;
	    RECT 324.4000 132.8000 325.2000 134.4000 ;
	    RECT 326.0000 133.6000 328.6000 134.4000 ;
	    RECT 330.0000 133.8000 331.6000 134.4000 ;
	    RECT 330.8000 133.6000 331.6000 133.8000 ;
	    RECT 326.0000 130.2000 326.8000 130.4000 ;
	    RECT 328.0000 130.2000 328.6000 133.6000 ;
	    RECT 329.2000 131.6000 330.0000 133.2000 ;
	    RECT 332.4000 131.6000 333.2000 133.2000 ;
	    RECT 334.0000 131.6000 334.6000 134.6000 ;
	    RECT 335.6000 132.4000 336.4000 139.8000 ;
	    RECT 337.2000 139.2000 341.2000 139.8000 ;
	    RECT 337.2000 135.8000 338.0000 139.2000 ;
	    RECT 338.8000 135.8000 339.6000 138.6000 ;
	    RECT 340.4000 136.0000 341.2000 139.2000 ;
	    RECT 343.6000 136.0000 344.4000 139.8000 ;
	    RECT 340.4000 135.8000 344.4000 136.0000 ;
	    RECT 346.8000 137.8000 347.6000 139.8000 ;
	    RECT 338.8000 134.4000 339.4000 135.8000 ;
	    RECT 340.6000 135.4000 344.2000 135.8000 ;
	    RECT 342.8000 134.4000 343.6000 134.8000 ;
	    RECT 346.8000 134.4000 347.4000 137.8000 ;
	    RECT 348.4000 135.6000 349.2000 137.2000 ;
	    RECT 350.0000 135.6000 350.8000 139.8000 ;
	    RECT 351.6000 136.0000 352.4000 139.8000 ;
	    RECT 354.8000 136.0000 355.6000 139.8000 ;
	    RECT 351.6000 135.8000 355.6000 136.0000 ;
	    RECT 356.4000 135.8000 357.2000 139.8000 ;
	    RECT 358.0000 136.0000 358.8000 139.8000 ;
	    RECT 361.2000 136.0000 362.0000 139.8000 ;
	    RECT 358.0000 135.8000 362.0000 136.0000 ;
	    RECT 362.8000 137.0000 363.6000 139.0000 ;
	    RECT 350.2000 134.4000 350.8000 135.6000 ;
	    RECT 351.8000 135.4000 355.4000 135.8000 ;
	    RECT 354.0000 134.4000 354.8000 134.8000 ;
	    RECT 356.6000 134.4000 357.2000 135.8000 ;
	    RECT 358.2000 135.4000 361.8000 135.8000 ;
	    RECT 362.8000 134.8000 363.4000 137.0000 ;
	    RECT 367.0000 136.0000 367.8000 139.0000 ;
	    RECT 372.4000 137.0000 373.2000 139.0000 ;
	    RECT 376.6000 138.4000 377.4000 139.0000 ;
	    RECT 376.6000 137.6000 378.0000 138.4000 ;
	    RECT 367.0000 135.4000 368.6000 136.0000 ;
	    RECT 367.8000 135.0000 368.6000 135.4000 ;
	    RECT 360.4000 134.4000 361.2000 134.8000 ;
	    RECT 337.2000 132.8000 338.0000 134.4000 ;
	    RECT 338.8000 133.8000 341.2000 134.4000 ;
	    RECT 342.8000 133.8000 344.4000 134.4000 ;
	    RECT 340.4000 133.6000 341.2000 133.8000 ;
	    RECT 343.6000 133.6000 344.4000 133.8000 ;
	    RECT 346.8000 133.6000 347.6000 134.4000 ;
	    RECT 350.0000 133.6000 352.6000 134.4000 ;
	    RECT 354.0000 133.8000 355.6000 134.4000 ;
	    RECT 354.8000 133.6000 355.6000 133.8000 ;
	    RECT 356.4000 133.6000 359.0000 134.4000 ;
	    RECT 360.4000 133.8000 362.0000 134.4000 ;
	    RECT 362.8000 134.2000 367.0000 134.8000 ;
	    RECT 361.2000 133.6000 362.0000 133.8000 ;
	    RECT 366.0000 133.8000 367.0000 134.2000 ;
	    RECT 368.0000 134.4000 368.6000 135.0000 ;
	    RECT 372.4000 134.8000 373.0000 137.0000 ;
	    RECT 376.6000 136.0000 377.4000 137.6000 ;
	    RECT 376.6000 135.4000 378.2000 136.0000 ;
	    RECT 377.4000 135.0000 378.2000 135.4000 ;
	    RECT 334.0000 130.8000 335.2000 131.6000 ;
	    RECT 334.0000 130.2000 334.6000 130.8000 ;
	    RECT 335.8000 130.2000 336.4000 132.4000 ;
	    RECT 338.8000 131.6000 339.6000 133.2000 ;
	    RECT 340.6000 130.2000 341.2000 133.6000 ;
	    RECT 342.0000 132.3000 342.8000 133.2000 ;
	    RECT 343.6000 132.3000 344.4000 132.4000 ;
	    RECT 342.0000 131.7000 344.4000 132.3000 ;
	    RECT 342.0000 131.6000 342.8000 131.7000 ;
	    RECT 343.6000 131.6000 344.4000 131.7000 ;
	    RECT 345.2000 130.8000 346.0000 132.4000 ;
	    RECT 346.8000 130.2000 347.4000 133.6000 ;
	    RECT 350.0000 130.2000 350.8000 130.4000 ;
	    RECT 352.0000 130.2000 352.6000 133.6000 ;
	    RECT 353.2000 132.3000 354.0000 133.2000 ;
	    RECT 358.4000 132.4000 359.0000 133.6000 ;
	    RECT 356.4000 132.3000 357.2000 132.4000 ;
	    RECT 353.2000 131.7000 357.2000 132.3000 ;
	    RECT 353.2000 131.6000 354.0000 131.7000 ;
	    RECT 356.4000 131.6000 357.2000 131.7000 ;
	    RECT 358.0000 131.6000 359.0000 132.4000 ;
	    RECT 359.6000 131.6000 360.4000 133.2000 ;
	    RECT 362.8000 131.6000 363.6000 133.2000 ;
	    RECT 364.4000 131.6000 365.2000 133.2000 ;
	    RECT 366.0000 133.0000 367.4000 133.8000 ;
	    RECT 368.0000 133.6000 370.0000 134.4000 ;
	    RECT 372.4000 134.2000 376.6000 134.8000 ;
	    RECT 375.6000 133.8000 376.6000 134.2000 ;
	    RECT 377.6000 134.4000 378.2000 135.0000 ;
	    RECT 356.4000 130.2000 357.2000 130.4000 ;
	    RECT 358.4000 130.2000 359.0000 131.6000 ;
	    RECT 366.0000 131.0000 366.6000 133.0000 ;
	    RECT 362.8000 130.4000 366.6000 131.0000 ;
	    RECT 279.6000 129.6000 281.8000 130.2000 ;
	    RECT 279.6000 122.2000 280.4000 129.6000 ;
	    RECT 282.8000 122.2000 283.6000 130.2000 ;
	    RECT 285.0000 129.4000 286.8000 130.2000 ;
	    RECT 289.8000 129.4000 291.6000 130.2000 ;
	    RECT 285.0000 124.4000 285.8000 129.4000 ;
	    RECT 284.4000 123.6000 285.8000 124.4000 ;
	    RECT 285.0000 122.2000 285.8000 123.6000 ;
	    RECT 289.8000 122.2000 290.6000 129.4000 ;
	    RECT 296.6000 122.2000 298.6000 130.2000 ;
	    RECT 302.6000 129.4000 304.4000 130.2000 ;
	    RECT 306.8000 129.6000 308.2000 130.2000 ;
	    RECT 308.8000 129.6000 309.8000 130.2000 ;
	    RECT 302.6000 128.4000 303.4000 129.4000 ;
	    RECT 302.0000 127.6000 303.4000 128.4000 ;
	    RECT 307.6000 128.4000 308.2000 129.6000 ;
	    RECT 307.6000 127.6000 308.4000 128.4000 ;
	    RECT 302.6000 122.2000 303.4000 127.6000 ;
	    RECT 309.0000 122.2000 309.8000 129.6000 ;
	    RECT 314.8000 129.4000 316.6000 130.2000 ;
	    RECT 315.8000 128.4000 316.6000 129.4000 ;
	    RECT 315.8000 127.6000 317.2000 128.4000 ;
	    RECT 315.8000 122.2000 316.6000 127.6000 ;
	    RECT 320.6000 124.4000 322.6000 130.2000 ;
	    RECT 326.0000 129.6000 327.4000 130.2000 ;
	    RECT 328.0000 129.6000 329.0000 130.2000 ;
	    RECT 326.8000 128.4000 327.4000 129.6000 ;
	    RECT 326.8000 127.6000 327.6000 128.4000 ;
	    RECT 319.6000 123.6000 322.6000 124.4000 ;
	    RECT 320.6000 122.2000 322.6000 123.6000 ;
	    RECT 328.2000 122.2000 329.0000 129.6000 ;
	    RECT 332.4000 129.6000 334.6000 130.2000 ;
	    RECT 332.4000 122.2000 333.2000 129.6000 ;
	    RECT 335.6000 122.2000 336.4000 130.2000 ;
	    RECT 339.8000 122.2000 341.8000 130.2000 ;
	    RECT 345.8000 129.4000 347.6000 130.2000 ;
	    RECT 350.0000 129.6000 351.4000 130.2000 ;
	    RECT 352.0000 129.6000 353.0000 130.2000 ;
	    RECT 356.4000 129.6000 357.8000 130.2000 ;
	    RECT 358.4000 129.6000 359.4000 130.2000 ;
	    RECT 345.8000 128.4000 346.6000 129.4000 ;
	    RECT 345.2000 127.6000 346.6000 128.4000 ;
	    RECT 350.8000 128.4000 351.4000 129.6000 ;
	    RECT 350.8000 127.6000 351.6000 128.4000 ;
	    RECT 345.8000 122.2000 346.6000 127.6000 ;
	    RECT 352.2000 122.2000 353.0000 129.6000 ;
	    RECT 357.2000 128.4000 357.8000 129.6000 ;
	    RECT 356.4000 127.6000 358.0000 128.4000 ;
	    RECT 358.6000 122.2000 359.4000 129.6000 ;
	    RECT 362.8000 127.0000 363.4000 130.4000 ;
	    RECT 368.0000 129.8000 368.6000 133.6000 ;
	    RECT 369.2000 132.3000 370.0000 132.4000 ;
	    RECT 370.8000 132.3000 371.6000 132.4000 ;
	    RECT 369.2000 131.7000 371.6000 132.3000 ;
	    RECT 369.2000 130.8000 370.0000 131.7000 ;
	    RECT 370.8000 131.6000 371.6000 131.7000 ;
	    RECT 372.4000 131.6000 373.2000 133.2000 ;
	    RECT 374.0000 131.6000 374.8000 133.2000 ;
	    RECT 375.6000 133.0000 377.0000 133.8000 ;
	    RECT 377.6000 133.6000 379.6000 134.4000 ;
	    RECT 375.6000 131.0000 376.2000 133.0000 ;
	    RECT 367.0000 129.2000 368.6000 129.8000 ;
	    RECT 372.4000 130.4000 376.2000 131.0000 ;
	    RECT 362.8000 123.0000 363.6000 127.0000 ;
	    RECT 367.0000 124.4000 367.8000 129.2000 ;
	    RECT 366.0000 123.6000 367.8000 124.4000 ;
	    RECT 367.0000 122.2000 367.8000 123.6000 ;
	    RECT 372.4000 127.0000 373.0000 130.4000 ;
	    RECT 377.6000 129.8000 378.2000 133.6000 ;
	    RECT 382.0000 132.4000 382.8000 139.8000 ;
	    RECT 385.2000 135.2000 386.0000 139.8000 ;
	    RECT 386.8000 135.8000 387.6000 139.8000 ;
	    RECT 388.4000 136.0000 389.2000 139.8000 ;
	    RECT 391.6000 136.0000 392.4000 139.8000 ;
	    RECT 388.4000 135.8000 392.4000 136.0000 ;
	    RECT 393.2000 136.0000 394.0000 139.8000 ;
	    RECT 396.4000 136.0000 397.2000 139.8000 ;
	    RECT 393.2000 135.8000 397.2000 136.0000 ;
	    RECT 398.0000 135.8000 398.8000 139.8000 ;
	    RECT 399.6000 135.8000 400.4000 139.8000 ;
	    RECT 401.2000 136.0000 402.0000 139.8000 ;
	    RECT 404.4000 136.0000 405.2000 139.8000 ;
	    RECT 401.2000 135.8000 405.2000 136.0000 ;
	    RECT 383.8000 134.6000 386.0000 135.2000 ;
	    RECT 378.8000 130.8000 379.6000 132.4000 ;
	    RECT 376.6000 129.2000 378.2000 129.8000 ;
	    RECT 382.0000 130.2000 382.6000 132.4000 ;
	    RECT 383.8000 131.6000 384.4000 134.6000 ;
	    RECT 387.0000 134.4000 387.6000 135.8000 ;
	    RECT 388.6000 135.4000 392.2000 135.8000 ;
	    RECT 393.4000 135.4000 397.0000 135.8000 ;
	    RECT 390.8000 134.4000 391.6000 134.8000 ;
	    RECT 394.0000 134.4000 394.8000 134.8000 ;
	    RECT 398.0000 134.4000 398.6000 135.8000 ;
	    RECT 399.8000 134.4000 400.4000 135.8000 ;
	    RECT 401.4000 135.4000 405.0000 135.8000 ;
	    RECT 412.4000 135.4000 413.2000 139.8000 ;
	    RECT 416.6000 138.4000 417.8000 139.8000 ;
	    RECT 416.6000 137.8000 418.0000 138.4000 ;
	    RECT 421.2000 137.8000 422.0000 139.8000 ;
	    RECT 425.6000 138.4000 426.4000 139.8000 ;
	    RECT 425.6000 137.8000 427.6000 138.4000 ;
	    RECT 417.2000 137.0000 418.0000 137.8000 ;
	    RECT 421.4000 137.2000 422.0000 137.8000 ;
	    RECT 421.4000 136.6000 424.2000 137.2000 ;
	    RECT 423.4000 136.4000 424.2000 136.6000 ;
	    RECT 425.2000 135.6000 426.0000 137.2000 ;
	    RECT 426.8000 137.0000 427.6000 137.8000 ;
	    RECT 415.4000 135.4000 416.2000 135.6000 ;
	    RECT 412.4000 134.8000 416.2000 135.4000 ;
	    RECT 403.6000 134.4000 404.4000 134.8000 ;
	    RECT 386.8000 133.6000 389.4000 134.4000 ;
	    RECT 390.8000 134.3000 392.4000 134.4000 ;
	    RECT 393.2000 134.3000 394.8000 134.4000 ;
	    RECT 390.8000 133.8000 394.8000 134.3000 ;
	    RECT 391.6000 133.7000 394.0000 133.8000 ;
	    RECT 391.6000 133.6000 392.4000 133.7000 ;
	    RECT 393.2000 133.6000 394.0000 133.7000 ;
	    RECT 396.2000 133.6000 398.8000 134.4000 ;
	    RECT 399.6000 133.6000 402.2000 134.4000 ;
	    RECT 403.6000 133.8000 405.2000 134.4000 ;
	    RECT 404.4000 133.6000 405.2000 133.8000 ;
	    RECT 385.2000 131.6000 386.0000 133.2000 ;
	    RECT 383.2000 130.8000 384.4000 131.6000 ;
	    RECT 383.8000 130.2000 384.4000 130.8000 ;
	    RECT 386.8000 130.2000 387.6000 130.4000 ;
	    RECT 388.8000 130.2000 389.4000 133.6000 ;
	    RECT 390.0000 132.3000 390.8000 133.2000 ;
	    RECT 391.6000 132.3000 392.4000 132.4000 ;
	    RECT 394.8000 132.3000 395.6000 133.2000 ;
	    RECT 390.0000 131.7000 395.6000 132.3000 ;
	    RECT 390.0000 131.6000 390.8000 131.7000 ;
	    RECT 391.6000 131.6000 392.4000 131.7000 ;
	    RECT 394.8000 131.6000 395.6000 131.7000 ;
	    RECT 396.2000 132.3000 396.8000 133.6000 ;
	    RECT 401.6000 132.4000 402.2000 133.6000 ;
	    RECT 396.2000 131.7000 400.3000 132.3000 ;
	    RECT 396.2000 130.2000 396.8000 131.7000 ;
	    RECT 399.7000 130.4000 400.3000 131.7000 ;
	    RECT 401.2000 131.6000 402.2000 132.4000 ;
	    RECT 402.8000 131.6000 403.6000 133.2000 ;
	    RECT 398.0000 130.2000 398.8000 130.4000 ;
	    RECT 372.4000 123.0000 373.2000 127.0000 ;
	    RECT 376.6000 122.2000 377.4000 129.2000 ;
	    RECT 382.0000 122.2000 382.8000 130.2000 ;
	    RECT 383.8000 129.6000 386.0000 130.2000 ;
	    RECT 386.8000 129.6000 388.2000 130.2000 ;
	    RECT 388.8000 129.6000 389.8000 130.2000 ;
	    RECT 385.2000 122.2000 386.0000 129.6000 ;
	    RECT 387.6000 128.4000 388.2000 129.6000 ;
	    RECT 386.8000 127.6000 388.4000 128.4000 ;
	    RECT 389.0000 124.4000 389.8000 129.6000 ;
	    RECT 395.8000 129.6000 396.8000 130.2000 ;
	    RECT 397.4000 129.6000 398.8000 130.2000 ;
	    RECT 399.6000 130.2000 400.4000 130.4000 ;
	    RECT 401.6000 130.2000 402.2000 131.6000 ;
	    RECT 412.4000 131.4000 413.2000 134.8000 ;
	    RECT 419.4000 134.2000 420.2000 134.4000 ;
	    RECT 425.2000 134.2000 425.8000 135.6000 ;
	    RECT 430.0000 135.0000 430.8000 139.8000 ;
	    RECT 432.2000 136.4000 433.0000 139.8000 ;
	    RECT 432.2000 135.8000 434.0000 136.4000 ;
	    RECT 436.4000 135.8000 437.2000 139.8000 ;
	    RECT 438.0000 136.0000 438.8000 139.8000 ;
	    RECT 441.2000 136.0000 442.0000 139.8000 ;
	    RECT 438.0000 135.8000 442.0000 136.0000 ;
	    RECT 442.8000 136.0000 443.6000 139.8000 ;
	    RECT 446.0000 136.0000 446.8000 139.8000 ;
	    RECT 442.8000 135.8000 446.8000 136.0000 ;
	    RECT 447.6000 135.8000 448.4000 139.8000 ;
	    RECT 449.8000 136.4000 450.6000 139.8000 ;
	    RECT 449.8000 135.8000 451.6000 136.4000 ;
	    RECT 428.4000 134.2000 430.0000 134.4000 ;
	    RECT 419.0000 133.6000 430.0000 134.2000 ;
	    RECT 417.2000 132.8000 418.0000 133.0000 ;
	    RECT 414.2000 132.2000 418.0000 132.8000 ;
	    RECT 414.2000 132.0000 415.0000 132.2000 ;
	    RECT 415.8000 131.4000 416.6000 131.6000 ;
	    RECT 412.4000 130.8000 416.6000 131.4000 ;
	    RECT 399.6000 129.6000 401.0000 130.2000 ;
	    RECT 401.6000 129.6000 402.6000 130.2000 ;
	    RECT 389.0000 123.6000 390.8000 124.4000 ;
	    RECT 389.0000 122.2000 389.8000 123.6000 ;
	    RECT 395.8000 122.2000 396.6000 129.6000 ;
	    RECT 397.4000 128.4000 398.0000 129.6000 ;
	    RECT 400.4000 128.4000 401.0000 129.6000 ;
	    RECT 397.2000 127.6000 398.8000 128.4000 ;
	    RECT 400.4000 127.6000 401.2000 128.4000 ;
	    RECT 401.8000 122.2000 402.6000 129.6000 ;
	    RECT 412.4000 122.2000 413.2000 130.8000 ;
	    RECT 419.0000 130.4000 419.6000 133.6000 ;
	    RECT 426.2000 133.4000 427.0000 133.6000 ;
	    RECT 425.2000 132.4000 426.0000 132.6000 ;
	    RECT 427.8000 132.4000 428.6000 132.6000 ;
	    RECT 423.6000 131.8000 428.6000 132.4000 ;
	    RECT 423.6000 131.6000 424.4000 131.8000 ;
	    RECT 425.2000 131.0000 430.8000 131.2000 ;
	    RECT 425.0000 130.8000 430.8000 131.0000 ;
	    RECT 417.2000 129.8000 419.6000 130.4000 ;
	    RECT 421.0000 130.6000 430.8000 130.8000 ;
	    RECT 421.0000 130.2000 425.8000 130.6000 ;
	    RECT 417.2000 128.8000 417.8000 129.8000 ;
	    RECT 416.4000 128.0000 417.8000 128.8000 ;
	    RECT 419.4000 129.0000 420.2000 129.2000 ;
	    RECT 421.0000 129.0000 421.6000 130.2000 ;
	    RECT 419.4000 128.4000 421.6000 129.0000 ;
	    RECT 422.2000 129.0000 427.6000 129.6000 ;
	    RECT 422.2000 128.8000 423.0000 129.0000 ;
	    RECT 426.8000 128.8000 427.6000 129.0000 ;
	    RECT 420.6000 127.4000 421.4000 127.6000 ;
	    RECT 423.4000 127.4000 424.2000 127.6000 ;
	    RECT 417.2000 126.2000 418.0000 127.0000 ;
	    RECT 420.6000 126.8000 424.2000 127.4000 ;
	    RECT 421.4000 126.2000 422.0000 126.8000 ;
	    RECT 426.8000 126.2000 427.6000 127.0000 ;
	    RECT 416.6000 122.2000 417.8000 126.2000 ;
	    RECT 421.2000 122.2000 422.0000 126.2000 ;
	    RECT 425.6000 125.6000 427.6000 126.2000 ;
	    RECT 425.6000 122.2000 426.4000 125.6000 ;
	    RECT 430.0000 122.2000 430.8000 130.6000 ;
	    RECT 431.6000 128.8000 432.4000 130.4000 ;
	    RECT 433.2000 130.3000 434.0000 135.8000 ;
	    RECT 434.8000 133.6000 435.6000 135.2000 ;
	    RECT 436.6000 134.4000 437.2000 135.8000 ;
	    RECT 438.2000 135.4000 441.8000 135.8000 ;
	    RECT 443.0000 135.4000 446.6000 135.8000 ;
	    RECT 440.4000 134.4000 441.2000 134.8000 ;
	    RECT 443.6000 134.4000 444.4000 134.8000 ;
	    RECT 447.6000 134.4000 448.2000 135.8000 ;
	    RECT 436.4000 133.6000 439.0000 134.4000 ;
	    RECT 440.4000 134.3000 442.0000 134.4000 ;
	    RECT 442.8000 134.3000 444.4000 134.4000 ;
	    RECT 440.4000 133.8000 444.4000 134.3000 ;
	    RECT 445.8000 134.3000 448.4000 134.4000 ;
	    RECT 449.2000 134.3000 450.0000 134.4000 ;
	    RECT 441.2000 133.7000 443.6000 133.8000 ;
	    RECT 441.2000 133.6000 442.0000 133.7000 ;
	    RECT 442.8000 133.6000 443.6000 133.7000 ;
	    RECT 445.8000 133.7000 450.0000 134.3000 ;
	    RECT 445.8000 133.6000 448.4000 133.7000 ;
	    RECT 449.2000 133.6000 450.0000 133.7000 ;
	    RECT 434.8000 132.3000 435.6000 132.4000 ;
	    RECT 438.4000 132.3000 439.0000 133.6000 ;
	    RECT 434.8000 131.7000 439.0000 132.3000 ;
	    RECT 434.8000 131.6000 435.6000 131.7000 ;
	    RECT 436.4000 130.3000 437.2000 130.4000 ;
	    RECT 433.2000 130.2000 437.2000 130.3000 ;
	    RECT 438.4000 130.2000 439.0000 131.7000 ;
	    RECT 439.6000 131.6000 440.4000 133.2000 ;
	    RECT 444.4000 131.6000 445.2000 133.2000 ;
	    RECT 445.8000 130.2000 446.4000 133.6000 ;
	    RECT 450.8000 132.3000 451.6000 135.8000 ;
	    RECT 454.0000 135.4000 454.8000 139.8000 ;
	    RECT 458.2000 138.4000 459.4000 139.8000 ;
	    RECT 458.2000 137.8000 459.6000 138.4000 ;
	    RECT 462.8000 137.8000 463.6000 139.8000 ;
	    RECT 467.2000 138.4000 468.0000 139.8000 ;
	    RECT 467.2000 137.8000 469.2000 138.4000 ;
	    RECT 458.8000 137.0000 459.6000 137.8000 ;
	    RECT 463.0000 137.2000 463.6000 137.8000 ;
	    RECT 463.0000 136.6000 465.8000 137.2000 ;
	    RECT 465.0000 136.4000 465.8000 136.6000 ;
	    RECT 466.8000 136.4000 467.6000 137.2000 ;
	    RECT 468.4000 137.0000 469.2000 137.8000 ;
	    RECT 457.0000 135.4000 457.8000 135.6000 ;
	    RECT 452.4000 133.6000 453.2000 135.2000 ;
	    RECT 454.0000 134.8000 457.8000 135.4000 ;
	    RECT 447.7000 131.7000 451.6000 132.3000 ;
	    RECT 447.7000 130.4000 448.3000 131.7000 ;
	    RECT 447.6000 130.2000 448.4000 130.4000 ;
	    RECT 433.2000 129.7000 437.8000 130.2000 ;
	    RECT 433.2000 122.2000 434.0000 129.7000 ;
	    RECT 436.4000 129.6000 437.8000 129.7000 ;
	    RECT 438.4000 129.6000 439.4000 130.2000 ;
	    RECT 437.2000 128.4000 437.8000 129.6000 ;
	    RECT 437.2000 127.6000 438.0000 128.4000 ;
	    RECT 438.6000 122.2000 439.4000 129.6000 ;
	    RECT 445.4000 129.6000 446.4000 130.2000 ;
	    RECT 447.0000 129.6000 448.4000 130.2000 ;
	    RECT 445.4000 122.2000 446.2000 129.6000 ;
	    RECT 447.0000 128.4000 447.6000 129.6000 ;
	    RECT 449.2000 128.8000 450.0000 130.4000 ;
	    RECT 446.8000 127.6000 447.6000 128.4000 ;
	    RECT 450.8000 122.2000 451.6000 131.7000 ;
	    RECT 454.0000 131.4000 454.8000 134.8000 ;
	    RECT 461.0000 134.2000 461.8000 134.4000 ;
	    RECT 466.8000 134.2000 467.4000 136.4000 ;
	    RECT 471.6000 135.0000 472.4000 139.8000 ;
	    RECT 473.2000 135.4000 474.0000 139.8000 ;
	    RECT 477.4000 138.4000 478.6000 139.8000 ;
	    RECT 477.4000 137.8000 478.8000 138.4000 ;
	    RECT 482.0000 137.8000 482.8000 139.8000 ;
	    RECT 486.4000 138.4000 487.2000 139.8000 ;
	    RECT 486.4000 137.8000 488.4000 138.4000 ;
	    RECT 478.0000 137.0000 478.8000 137.8000 ;
	    RECT 482.2000 137.2000 482.8000 137.8000 ;
	    RECT 482.2000 136.6000 485.0000 137.2000 ;
	    RECT 484.2000 136.4000 485.0000 136.6000 ;
	    RECT 486.0000 136.4000 486.8000 137.2000 ;
	    RECT 487.6000 137.0000 488.4000 137.8000 ;
	    RECT 476.2000 135.4000 477.0000 135.6000 ;
	    RECT 473.2000 134.8000 477.0000 135.4000 ;
	    RECT 470.0000 134.2000 471.6000 134.4000 ;
	    RECT 460.6000 133.6000 471.6000 134.2000 ;
	    RECT 458.8000 132.8000 459.6000 133.0000 ;
	    RECT 455.8000 132.2000 459.6000 132.8000 ;
	    RECT 455.8000 132.0000 456.6000 132.2000 ;
	    RECT 457.4000 131.4000 458.2000 131.6000 ;
	    RECT 454.0000 130.8000 458.2000 131.4000 ;
	    RECT 452.4000 128.3000 453.2000 128.4000 ;
	    RECT 454.0000 128.3000 454.8000 130.8000 ;
	    RECT 460.6000 130.4000 461.2000 133.6000 ;
	    RECT 467.8000 133.4000 468.6000 133.6000 ;
	    RECT 469.4000 132.4000 470.2000 132.6000 ;
	    RECT 463.6000 132.3000 464.4000 132.4000 ;
	    RECT 465.2000 132.3000 470.2000 132.4000 ;
	    RECT 463.6000 131.8000 470.2000 132.3000 ;
	    RECT 463.6000 131.7000 466.0000 131.8000 ;
	    RECT 463.6000 131.6000 464.4000 131.7000 ;
	    RECT 465.2000 131.6000 466.0000 131.7000 ;
	    RECT 473.2000 131.4000 474.0000 134.8000 ;
	    RECT 480.2000 134.2000 481.0000 134.4000 ;
	    RECT 486.0000 134.2000 486.6000 136.4000 ;
	    RECT 490.8000 135.0000 491.6000 139.8000 ;
	    RECT 492.4000 135.6000 493.2000 137.2000 ;
	    RECT 489.2000 134.2000 490.8000 134.4000 ;
	    RECT 479.8000 133.6000 490.8000 134.2000 ;
	    RECT 494.0000 134.3000 494.8000 139.8000 ;
	    RECT 495.6000 136.0000 496.4000 139.8000 ;
	    RECT 498.8000 136.0000 499.6000 139.8000 ;
	    RECT 495.6000 135.8000 499.6000 136.0000 ;
	    RECT 500.4000 135.8000 501.2000 139.8000 ;
	    RECT 502.0000 136.0000 502.8000 139.8000 ;
	    RECT 505.2000 136.0000 506.0000 139.8000 ;
	    RECT 502.0000 135.8000 506.0000 136.0000 ;
	    RECT 506.8000 135.8000 507.6000 139.8000 ;
	    RECT 495.8000 135.4000 499.4000 135.8000 ;
	    RECT 496.4000 134.4000 497.2000 134.8000 ;
	    RECT 500.4000 134.4000 501.0000 135.8000 ;
	    RECT 502.2000 135.4000 505.8000 135.8000 ;
	    RECT 502.8000 134.4000 503.6000 134.8000 ;
	    RECT 506.8000 134.4000 507.4000 135.8000 ;
	    RECT 495.6000 134.3000 497.2000 134.4000 ;
	    RECT 494.0000 133.8000 497.2000 134.3000 ;
	    RECT 494.0000 133.7000 496.4000 133.8000 ;
	    RECT 478.0000 132.8000 478.8000 133.0000 ;
	    RECT 475.0000 132.2000 478.8000 132.8000 ;
	    RECT 475.0000 132.0000 475.8000 132.2000 ;
	    RECT 476.6000 131.4000 477.4000 131.6000 ;
	    RECT 466.8000 131.0000 472.4000 131.2000 ;
	    RECT 466.6000 130.8000 472.4000 131.0000 ;
	    RECT 458.8000 129.8000 461.2000 130.4000 ;
	    RECT 462.6000 130.6000 472.4000 130.8000 ;
	    RECT 462.6000 130.2000 467.4000 130.6000 ;
	    RECT 458.8000 128.8000 459.4000 129.8000 ;
	    RECT 452.4000 127.7000 454.8000 128.3000 ;
	    RECT 458.0000 128.0000 459.4000 128.8000 ;
	    RECT 461.0000 129.0000 461.8000 129.2000 ;
	    RECT 462.6000 129.0000 463.2000 130.2000 ;
	    RECT 461.0000 128.4000 463.2000 129.0000 ;
	    RECT 463.8000 129.0000 469.2000 129.6000 ;
	    RECT 463.8000 128.8000 464.6000 129.0000 ;
	    RECT 468.4000 128.8000 469.2000 129.0000 ;
	    RECT 452.4000 127.6000 453.2000 127.7000 ;
	    RECT 454.0000 122.2000 454.8000 127.7000 ;
	    RECT 462.2000 127.4000 463.0000 127.6000 ;
	    RECT 465.0000 127.4000 465.8000 127.6000 ;
	    RECT 458.8000 126.2000 459.6000 127.0000 ;
	    RECT 462.2000 126.8000 465.8000 127.4000 ;
	    RECT 463.0000 126.2000 463.6000 126.8000 ;
	    RECT 468.4000 126.2000 469.2000 127.0000 ;
	    RECT 458.2000 122.2000 459.4000 126.2000 ;
	    RECT 462.8000 122.2000 463.6000 126.2000 ;
	    RECT 467.2000 125.6000 469.2000 126.2000 ;
	    RECT 467.2000 122.2000 468.0000 125.6000 ;
	    RECT 471.6000 122.2000 472.4000 130.6000 ;
	    RECT 473.2000 130.8000 477.4000 131.4000 ;
	    RECT 473.2000 122.2000 474.0000 130.8000 ;
	    RECT 479.8000 130.4000 480.4000 133.6000 ;
	    RECT 487.0000 133.4000 487.8000 133.6000 ;
	    RECT 486.0000 132.4000 486.8000 132.6000 ;
	    RECT 488.6000 132.4000 489.4000 132.6000 ;
	    RECT 484.4000 131.8000 489.4000 132.4000 ;
	    RECT 484.4000 131.6000 485.2000 131.8000 ;
	    RECT 486.0000 131.0000 491.6000 131.2000 ;
	    RECT 485.8000 130.8000 491.6000 131.0000 ;
	    RECT 478.0000 129.8000 480.4000 130.4000 ;
	    RECT 481.8000 130.6000 491.6000 130.8000 ;
	    RECT 481.8000 130.2000 486.6000 130.6000 ;
	    RECT 478.0000 128.8000 478.6000 129.8000 ;
	    RECT 477.2000 128.0000 478.6000 128.8000 ;
	    RECT 480.2000 129.0000 481.0000 129.2000 ;
	    RECT 481.8000 129.0000 482.4000 130.2000 ;
	    RECT 480.2000 128.4000 482.4000 129.0000 ;
	    RECT 483.0000 129.0000 488.4000 129.6000 ;
	    RECT 483.0000 128.8000 483.8000 129.0000 ;
	    RECT 487.6000 128.8000 488.4000 129.0000 ;
	    RECT 481.4000 127.4000 482.2000 127.6000 ;
	    RECT 484.2000 127.4000 485.0000 127.6000 ;
	    RECT 478.0000 126.2000 478.8000 127.0000 ;
	    RECT 481.4000 126.8000 485.0000 127.4000 ;
	    RECT 482.2000 126.2000 482.8000 126.8000 ;
	    RECT 487.6000 126.2000 488.4000 127.0000 ;
	    RECT 477.4000 122.2000 478.6000 126.2000 ;
	    RECT 482.0000 122.2000 482.8000 126.2000 ;
	    RECT 486.4000 125.6000 488.4000 126.2000 ;
	    RECT 486.4000 122.2000 487.2000 125.6000 ;
	    RECT 490.8000 122.2000 491.6000 130.6000 ;
	    RECT 494.0000 122.2000 494.8000 133.7000 ;
	    RECT 495.6000 133.6000 496.4000 133.7000 ;
	    RECT 498.6000 133.6000 501.2000 134.4000 ;
	    RECT 502.0000 133.8000 503.6000 134.4000 ;
	    RECT 502.0000 133.6000 502.8000 133.8000 ;
	    RECT 505.0000 133.6000 507.6000 134.4000 ;
	    RECT 512.0000 134.2000 512.8000 139.8000 ;
	    RECT 512.0000 133.8000 513.8000 134.2000 ;
	    RECT 512.2000 133.6000 513.8000 133.8000 ;
	    RECT 495.6000 132.3000 496.4000 132.4000 ;
	    RECT 497.2000 132.3000 498.0000 133.2000 ;
	    RECT 495.6000 131.7000 498.0000 132.3000 ;
	    RECT 495.6000 131.6000 496.4000 131.7000 ;
	    RECT 497.2000 131.6000 498.0000 131.7000 ;
	    RECT 498.6000 130.2000 499.2000 133.6000 ;
	    RECT 503.6000 131.6000 504.4000 133.2000 ;
	    RECT 500.4000 130.2000 501.2000 130.4000 ;
	    RECT 505.0000 130.2000 505.6000 133.6000 ;
	    RECT 510.0000 131.6000 511.6000 132.4000 ;
	    RECT 513.2000 130.4000 513.8000 133.6000 ;
	    RECT 506.8000 130.2000 507.6000 130.4000 ;
	    RECT 498.2000 129.6000 499.2000 130.2000 ;
	    RECT 499.8000 129.6000 501.2000 130.2000 ;
	    RECT 504.6000 129.6000 505.6000 130.2000 ;
	    RECT 506.2000 129.6000 507.6000 130.2000 ;
	    RECT 513.2000 129.6000 514.0000 130.4000 ;
	    RECT 498.2000 122.2000 499.0000 129.6000 ;
	    RECT 499.8000 128.4000 500.4000 129.6000 ;
	    RECT 499.6000 127.6000 500.4000 128.4000 ;
	    RECT 504.6000 122.2000 505.4000 129.6000 ;
	    RECT 506.2000 128.4000 506.8000 129.6000 ;
	    RECT 506.0000 127.6000 506.8000 128.4000 ;
	    RECT 511.6000 127.6000 512.4000 129.2000 ;
	    RECT 513.2000 127.0000 513.8000 129.6000 ;
	    RECT 510.2000 126.4000 513.8000 127.0000 ;
	    RECT 510.0000 122.2000 510.8000 126.4000 ;
	    RECT 513.2000 126.2000 513.8000 126.4000 ;
	    RECT 513.2000 122.2000 514.0000 126.2000 ;
	    RECT 4.4000 112.4000 5.2000 119.8000 ;
	    RECT 3.0000 111.8000 5.2000 112.4000 ;
	    RECT 3.0000 111.2000 3.6000 111.8000 ;
	    RECT 2.4000 110.4000 3.6000 111.2000 ;
	    RECT 6.0000 111.2000 6.8000 119.8000 ;
	    RECT 10.2000 115.8000 11.4000 119.8000 ;
	    RECT 14.8000 115.8000 15.6000 119.8000 ;
	    RECT 19.2000 116.4000 20.0000 119.8000 ;
	    RECT 19.2000 115.8000 21.2000 116.4000 ;
	    RECT 10.8000 115.0000 11.6000 115.8000 ;
	    RECT 15.0000 115.2000 15.6000 115.8000 ;
	    RECT 14.2000 114.6000 17.8000 115.2000 ;
	    RECT 20.4000 115.0000 21.2000 115.8000 ;
	    RECT 14.2000 114.4000 15.0000 114.6000 ;
	    RECT 17.0000 114.4000 17.8000 114.6000 ;
	    RECT 10.0000 113.2000 11.4000 114.0000 ;
	    RECT 10.8000 112.2000 11.4000 113.2000 ;
	    RECT 13.0000 113.0000 15.2000 113.6000 ;
	    RECT 13.0000 112.8000 13.8000 113.0000 ;
	    RECT 10.8000 111.6000 13.2000 112.2000 ;
	    RECT 6.0000 110.6000 10.2000 111.2000 ;
	    RECT 3.0000 107.4000 3.6000 110.4000 ;
	    RECT 4.4000 108.8000 5.2000 110.4000 ;
	    RECT 3.0000 106.8000 5.2000 107.4000 ;
	    RECT 4.4000 102.2000 5.2000 106.8000 ;
	    RECT 6.0000 107.2000 6.8000 110.6000 ;
	    RECT 9.4000 110.4000 10.2000 110.6000 ;
	    RECT 7.8000 109.8000 8.6000 110.0000 ;
	    RECT 7.8000 109.2000 11.6000 109.8000 ;
	    RECT 10.8000 109.0000 11.6000 109.2000 ;
	    RECT 12.6000 108.4000 13.2000 111.6000 ;
	    RECT 14.6000 111.8000 15.2000 113.0000 ;
	    RECT 15.8000 113.0000 16.6000 113.2000 ;
	    RECT 20.4000 113.0000 21.2000 113.2000 ;
	    RECT 15.8000 112.4000 21.2000 113.0000 ;
	    RECT 14.6000 111.4000 19.4000 111.8000 ;
	    RECT 23.6000 111.4000 24.4000 119.8000 ;
	    RECT 27.8000 114.4000 28.6000 119.8000 ;
	    RECT 32.2000 118.4000 33.0000 119.8000 ;
	    RECT 32.2000 117.6000 34.0000 118.4000 ;
	    RECT 26.8000 113.6000 28.6000 114.4000 ;
	    RECT 29.2000 113.6000 30.0000 114.4000 ;
	    RECT 27.8000 112.4000 28.6000 113.6000 ;
	    RECT 29.4000 112.4000 30.0000 113.6000 ;
	    RECT 32.2000 112.6000 33.0000 117.6000 ;
	    RECT 27.8000 111.8000 28.8000 112.4000 ;
	    RECT 29.4000 111.8000 30.8000 112.4000 ;
	    RECT 32.2000 111.8000 34.0000 112.6000 ;
	    RECT 14.6000 111.2000 24.4000 111.4000 ;
	    RECT 18.6000 111.0000 24.4000 111.2000 ;
	    RECT 18.8000 110.8000 24.4000 111.0000 ;
	    RECT 17.2000 110.2000 18.0000 110.4000 ;
	    RECT 17.2000 109.6000 22.2000 110.2000 ;
	    RECT 21.4000 109.4000 22.2000 109.6000 ;
	    RECT 26.8000 108.8000 27.6000 110.4000 ;
	    RECT 19.8000 108.4000 20.6000 108.6000 ;
	    RECT 28.2000 108.4000 28.8000 111.8000 ;
	    RECT 30.0000 111.6000 30.8000 111.8000 ;
	    RECT 31.6000 109.6000 32.4000 111.2000 ;
	    RECT 33.2000 108.4000 33.8000 111.8000 ;
	    RECT 36.4000 111.2000 37.2000 119.8000 ;
	    RECT 40.6000 115.8000 41.8000 119.8000 ;
	    RECT 45.2000 115.8000 46.0000 119.8000 ;
	    RECT 49.6000 116.4000 50.4000 119.8000 ;
	    RECT 49.6000 115.8000 51.6000 116.4000 ;
	    RECT 41.2000 115.0000 42.0000 115.8000 ;
	    RECT 45.4000 115.2000 46.0000 115.8000 ;
	    RECT 44.6000 114.6000 48.2000 115.2000 ;
	    RECT 50.8000 115.0000 51.6000 115.8000 ;
	    RECT 44.6000 114.4000 45.4000 114.6000 ;
	    RECT 47.4000 114.4000 48.2000 114.6000 ;
	    RECT 40.4000 113.2000 41.8000 114.0000 ;
	    RECT 41.2000 112.2000 41.8000 113.2000 ;
	    RECT 43.4000 113.0000 45.6000 113.6000 ;
	    RECT 43.4000 112.8000 44.2000 113.0000 ;
	    RECT 41.2000 111.6000 43.6000 112.2000 ;
	    RECT 36.4000 110.6000 40.6000 111.2000 ;
	    RECT 12.6000 107.8000 23.6000 108.4000 ;
	    RECT 13.0000 107.6000 13.8000 107.8000 ;
	    RECT 18.8000 107.6000 19.6000 107.8000 ;
	    RECT 22.0000 107.6000 23.6000 107.8000 ;
	    RECT 25.2000 108.2000 26.0000 108.4000 ;
	    RECT 25.2000 107.6000 26.8000 108.2000 ;
	    RECT 28.2000 107.6000 30.8000 108.4000 ;
	    RECT 33.2000 107.6000 34.0000 108.4000 ;
	    RECT 6.0000 106.6000 9.8000 107.2000 ;
	    RECT 6.0000 102.2000 6.8000 106.6000 ;
	    RECT 9.0000 106.4000 9.8000 106.6000 ;
	    RECT 18.8000 105.6000 19.4000 107.6000 ;
	    RECT 26.0000 107.2000 26.8000 107.6000 ;
	    RECT 17.0000 105.4000 17.8000 105.6000 ;
	    RECT 10.8000 104.2000 11.6000 105.0000 ;
	    RECT 15.0000 104.8000 17.8000 105.4000 ;
	    RECT 18.8000 104.8000 19.6000 105.6000 ;
	    RECT 15.0000 104.2000 15.6000 104.8000 ;
	    RECT 20.4000 104.2000 21.2000 105.0000 ;
	    RECT 10.2000 103.6000 11.6000 104.2000 ;
	    RECT 10.2000 102.2000 11.4000 103.6000 ;
	    RECT 14.8000 102.2000 15.6000 104.2000 ;
	    RECT 19.2000 103.6000 21.2000 104.2000 ;
	    RECT 19.2000 102.2000 20.0000 103.6000 ;
	    RECT 23.6000 102.2000 24.4000 107.0000 ;
	    RECT 25.4000 106.2000 29.0000 106.6000 ;
	    RECT 30.0000 106.2000 30.6000 107.6000 ;
	    RECT 25.2000 106.0000 29.2000 106.2000 ;
	    RECT 25.2000 102.2000 26.0000 106.0000 ;
	    RECT 28.4000 102.2000 29.2000 106.0000 ;
	    RECT 30.0000 102.2000 30.8000 106.2000 ;
	    RECT 33.2000 104.4000 33.8000 107.6000 ;
	    RECT 36.4000 107.2000 37.2000 110.6000 ;
	    RECT 39.8000 110.4000 40.6000 110.6000 ;
	    RECT 38.2000 109.8000 39.0000 110.0000 ;
	    RECT 38.2000 109.2000 42.0000 109.8000 ;
	    RECT 41.2000 109.0000 42.0000 109.2000 ;
	    RECT 43.0000 108.4000 43.6000 111.6000 ;
	    RECT 45.0000 111.8000 45.6000 113.0000 ;
	    RECT 46.2000 113.0000 47.0000 113.2000 ;
	    RECT 50.8000 113.0000 51.6000 113.2000 ;
	    RECT 46.2000 112.4000 51.6000 113.0000 ;
	    RECT 45.0000 111.4000 49.8000 111.8000 ;
	    RECT 54.0000 111.4000 54.8000 119.8000 ;
	    RECT 56.4000 113.6000 57.2000 114.4000 ;
	    RECT 56.4000 112.4000 57.0000 113.6000 ;
	    RECT 57.8000 112.4000 58.6000 119.8000 ;
	    RECT 55.6000 111.8000 57.0000 112.4000 ;
	    RECT 57.6000 111.8000 58.6000 112.4000 ;
	    RECT 55.6000 111.6000 56.4000 111.8000 ;
	    RECT 45.0000 111.2000 54.8000 111.4000 ;
	    RECT 49.0000 111.0000 54.8000 111.2000 ;
	    RECT 49.2000 110.8000 54.8000 111.0000 ;
	    RECT 47.6000 110.2000 48.4000 110.4000 ;
	    RECT 47.6000 109.6000 52.6000 110.2000 ;
	    RECT 49.2000 109.4000 50.0000 109.6000 ;
	    RECT 51.8000 109.4000 52.6000 109.6000 ;
	    RECT 50.2000 108.4000 51.0000 108.6000 ;
	    RECT 57.6000 108.4000 58.2000 111.8000 ;
	    RECT 62.0000 111.4000 62.8000 119.8000 ;
	    RECT 66.4000 116.4000 67.2000 119.8000 ;
	    RECT 65.2000 115.8000 67.2000 116.4000 ;
	    RECT 70.8000 115.8000 71.6000 119.8000 ;
	    RECT 75.0000 115.8000 76.2000 119.8000 ;
	    RECT 65.2000 115.0000 66.0000 115.8000 ;
	    RECT 70.8000 115.2000 71.4000 115.8000 ;
	    RECT 68.6000 114.6000 72.2000 115.2000 ;
	    RECT 74.8000 115.0000 75.6000 115.8000 ;
	    RECT 68.6000 114.4000 69.4000 114.6000 ;
	    RECT 71.4000 114.4000 72.2000 114.6000 ;
	    RECT 65.2000 113.0000 66.0000 113.2000 ;
	    RECT 69.8000 113.0000 70.6000 113.2000 ;
	    RECT 65.2000 112.4000 70.6000 113.0000 ;
	    RECT 71.2000 113.0000 73.4000 113.6000 ;
	    RECT 71.2000 111.8000 71.8000 113.0000 ;
	    RECT 72.6000 112.8000 73.4000 113.0000 ;
	    RECT 75.0000 113.2000 76.4000 114.0000 ;
	    RECT 75.0000 112.2000 75.6000 113.2000 ;
	    RECT 67.0000 111.4000 71.8000 111.8000 ;
	    RECT 62.0000 111.2000 71.8000 111.4000 ;
	    RECT 73.2000 111.6000 75.6000 112.2000 ;
	    RECT 62.0000 111.0000 67.8000 111.2000 ;
	    RECT 62.0000 110.8000 67.6000 111.0000 ;
	    RECT 58.8000 108.8000 59.6000 110.4000 ;
	    RECT 68.4000 110.3000 69.2000 110.4000 ;
	    RECT 71.6000 110.3000 72.4000 110.4000 ;
	    RECT 68.4000 110.2000 72.4000 110.3000 ;
	    RECT 64.2000 109.7000 72.4000 110.2000 ;
	    RECT 64.2000 109.6000 69.2000 109.7000 ;
	    RECT 71.6000 109.6000 72.4000 109.7000 ;
	    RECT 64.2000 109.4000 65.0000 109.6000 ;
	    RECT 65.8000 108.4000 66.6000 108.6000 ;
	    RECT 73.2000 108.4000 73.8000 111.6000 ;
	    RECT 79.6000 111.2000 80.4000 119.8000 ;
	    RECT 76.2000 110.6000 80.4000 111.2000 ;
	    RECT 76.2000 110.4000 77.0000 110.6000 ;
	    RECT 77.8000 109.8000 78.6000 110.0000 ;
	    RECT 74.8000 109.2000 78.6000 109.8000 ;
	    RECT 74.8000 109.0000 75.6000 109.2000 ;
	    RECT 43.0000 107.8000 54.0000 108.4000 ;
	    RECT 43.4000 107.6000 44.2000 107.8000 ;
	    RECT 36.4000 106.6000 40.2000 107.2000 ;
	    RECT 34.8000 104.8000 35.6000 106.4000 ;
	    RECT 33.2000 102.2000 34.0000 104.4000 ;
	    RECT 36.4000 102.2000 37.2000 106.6000 ;
	    RECT 39.4000 106.4000 40.2000 106.6000 ;
	    RECT 49.2000 105.6000 49.8000 107.8000 ;
	    RECT 52.4000 107.6000 54.0000 107.8000 ;
	    RECT 55.6000 107.6000 58.2000 108.4000 ;
	    RECT 60.4000 108.2000 61.2000 108.4000 ;
	    RECT 59.6000 107.6000 61.2000 108.2000 ;
	    RECT 62.8000 107.8000 73.8000 108.4000 ;
	    RECT 79.6000 108.3000 80.4000 110.6000 ;
	    RECT 82.8000 110.3000 83.6000 119.8000 ;
	    RECT 86.8000 113.6000 87.6000 114.4000 ;
	    RECT 84.4000 111.6000 85.2000 113.2000 ;
	    RECT 86.8000 112.4000 87.4000 113.6000 ;
	    RECT 88.2000 112.4000 89.0000 119.8000 ;
	    RECT 96.2000 112.8000 97.0000 119.8000 ;
	    RECT 100.4000 115.0000 101.2000 119.0000 ;
	    RECT 86.0000 111.8000 87.4000 112.4000 ;
	    RECT 88.0000 111.8000 89.0000 112.4000 ;
	    RECT 95.4000 112.2000 97.0000 112.8000 ;
	    RECT 86.0000 111.6000 86.8000 111.8000 ;
	    RECT 86.1000 110.3000 86.7000 111.6000 ;
	    RECT 82.8000 109.7000 86.7000 110.3000 ;
	    RECT 81.2000 108.3000 82.0000 108.4000 ;
	    RECT 62.8000 107.6000 64.4000 107.8000 ;
	    RECT 47.4000 105.4000 48.2000 105.6000 ;
	    RECT 41.2000 104.2000 42.0000 105.0000 ;
	    RECT 45.4000 104.8000 48.2000 105.4000 ;
	    RECT 49.2000 104.8000 50.0000 105.6000 ;
	    RECT 45.4000 104.2000 46.0000 104.8000 ;
	    RECT 50.8000 104.2000 51.6000 105.0000 ;
	    RECT 40.6000 103.6000 42.0000 104.2000 ;
	    RECT 40.6000 102.2000 41.8000 103.6000 ;
	    RECT 45.2000 102.2000 46.0000 104.2000 ;
	    RECT 49.6000 103.6000 51.6000 104.2000 ;
	    RECT 49.6000 102.2000 50.4000 103.6000 ;
	    RECT 54.0000 102.2000 54.8000 107.0000 ;
	    RECT 55.8000 106.2000 56.4000 107.6000 ;
	    RECT 59.6000 107.2000 60.4000 107.6000 ;
	    RECT 57.4000 106.2000 61.0000 106.6000 ;
	    RECT 55.6000 102.2000 56.4000 106.2000 ;
	    RECT 57.2000 106.0000 61.2000 106.2000 ;
	    RECT 57.2000 102.2000 58.0000 106.0000 ;
	    RECT 60.4000 102.2000 61.2000 106.0000 ;
	    RECT 62.0000 102.2000 62.8000 107.0000 ;
	    RECT 67.0000 105.6000 67.6000 107.8000 ;
	    RECT 68.4000 107.6000 69.2000 107.8000 ;
	    RECT 72.6000 107.6000 73.4000 107.8000 ;
	    RECT 79.6000 107.7000 82.0000 108.3000 ;
	    RECT 79.6000 107.2000 80.4000 107.7000 ;
	    RECT 76.6000 106.6000 80.4000 107.2000 ;
	    RECT 81.2000 106.8000 82.0000 107.7000 ;
	    RECT 76.6000 106.4000 77.4000 106.6000 ;
	    RECT 65.2000 104.2000 66.0000 105.0000 ;
	    RECT 66.8000 104.8000 67.6000 105.6000 ;
	    RECT 68.6000 105.4000 69.4000 105.6000 ;
	    RECT 68.6000 104.8000 71.4000 105.4000 ;
	    RECT 70.8000 104.2000 71.4000 104.8000 ;
	    RECT 74.8000 104.2000 75.6000 105.0000 ;
	    RECT 65.2000 103.6000 67.2000 104.2000 ;
	    RECT 66.4000 102.2000 67.2000 103.6000 ;
	    RECT 70.8000 102.2000 71.6000 104.2000 ;
	    RECT 74.8000 103.6000 76.2000 104.2000 ;
	    RECT 75.0000 102.2000 76.2000 103.6000 ;
	    RECT 79.6000 102.2000 80.4000 106.6000 ;
	    RECT 82.8000 106.2000 83.6000 109.7000 ;
	    RECT 88.0000 108.4000 88.6000 111.8000 ;
	    RECT 89.2000 108.8000 90.0000 110.4000 ;
	    RECT 94.0000 109.6000 94.8000 111.2000 ;
	    RECT 95.4000 110.4000 96.0000 112.2000 ;
	    RECT 100.6000 111.6000 101.2000 115.0000 ;
	    RECT 111.0000 111.8000 113.0000 119.8000 ;
	    RECT 117.2000 113.6000 118.0000 114.4000 ;
	    RECT 117.2000 112.4000 117.8000 113.6000 ;
	    RECT 118.6000 112.4000 119.4000 119.8000 ;
	    RECT 116.4000 111.8000 117.8000 112.4000 ;
	    RECT 118.4000 111.8000 119.4000 112.4000 ;
	    RECT 122.8000 115.0000 123.6000 119.0000 ;
	    RECT 127.0000 118.4000 127.8000 119.8000 ;
	    RECT 135.0000 118.4000 135.8000 119.8000 ;
	    RECT 127.0000 117.6000 128.4000 118.4000 ;
	    RECT 134.0000 117.6000 135.8000 118.4000 ;
	    RECT 97.4000 111.0000 101.2000 111.6000 ;
	    RECT 95.4000 109.6000 96.4000 110.4000 ;
	    RECT 95.4000 108.4000 96.0000 109.6000 ;
	    RECT 97.4000 109.0000 98.0000 111.0000 ;
	    RECT 86.0000 107.6000 88.6000 108.4000 ;
	    RECT 90.8000 108.2000 91.6000 108.4000 ;
	    RECT 90.0000 107.6000 91.6000 108.2000 ;
	    RECT 94.0000 107.6000 96.0000 108.4000 ;
	    RECT 96.6000 108.2000 98.0000 109.0000 ;
	    RECT 98.8000 108.8000 99.6000 110.4000 ;
	    RECT 100.4000 108.8000 101.2000 110.4000 ;
	    RECT 86.2000 106.2000 86.8000 107.6000 ;
	    RECT 90.0000 107.2000 90.8000 107.6000 ;
	    RECT 95.4000 107.0000 96.0000 107.6000 ;
	    RECT 97.0000 107.8000 98.0000 108.2000 ;
	    RECT 97.0000 107.2000 101.2000 107.8000 ;
	    RECT 108.4000 107.6000 109.2000 109.2000 ;
	    RECT 110.0000 108.8000 110.8000 110.4000 ;
	    RECT 111.8000 108.4000 112.4000 111.8000 ;
	    RECT 116.4000 111.6000 117.2000 111.8000 ;
	    RECT 113.2000 110.3000 114.0000 110.4000 ;
	    RECT 114.8000 110.3000 115.6000 110.4000 ;
	    RECT 113.2000 109.7000 115.6000 110.3000 ;
	    RECT 113.2000 108.8000 114.0000 109.7000 ;
	    RECT 114.8000 109.6000 115.6000 109.7000 ;
	    RECT 118.4000 108.4000 119.0000 111.8000 ;
	    RECT 122.8000 111.6000 123.4000 115.0000 ;
	    RECT 127.0000 112.8000 127.8000 117.6000 ;
	    RECT 127.0000 112.2000 128.6000 112.8000 ;
	    RECT 122.8000 111.0000 126.6000 111.6000 ;
	    RECT 119.6000 108.8000 120.4000 110.4000 ;
	    RECT 122.8000 108.8000 123.6000 110.4000 ;
	    RECT 124.4000 108.8000 125.2000 110.4000 ;
	    RECT 126.0000 109.0000 126.6000 111.0000 ;
	    RECT 111.6000 108.2000 112.4000 108.4000 ;
	    RECT 114.8000 108.3000 115.6000 108.4000 ;
	    RECT 116.4000 108.3000 119.0000 108.4000 ;
	    RECT 114.8000 108.2000 119.0000 108.3000 ;
	    RECT 121.2000 108.2000 122.0000 108.4000 ;
	    RECT 110.0000 107.6000 112.4000 108.2000 ;
	    RECT 114.0000 107.7000 119.0000 108.2000 ;
	    RECT 114.0000 107.6000 115.6000 107.7000 ;
	    RECT 116.4000 107.6000 119.0000 107.7000 ;
	    RECT 120.4000 107.6000 122.0000 108.2000 ;
	    RECT 126.0000 108.2000 127.4000 109.0000 ;
	    RECT 128.0000 108.4000 128.6000 112.2000 ;
	    RECT 135.0000 112.4000 135.8000 117.6000 ;
	    RECT 136.4000 113.6000 137.2000 114.4000 ;
	    RECT 136.6000 112.4000 137.2000 113.6000 ;
	    RECT 135.0000 111.8000 136.0000 112.4000 ;
	    RECT 136.6000 111.8000 138.0000 112.4000 ;
	    RECT 129.2000 109.6000 130.0000 111.2000 ;
	    RECT 134.0000 108.8000 134.8000 110.4000 ;
	    RECT 135.4000 108.4000 136.0000 111.8000 ;
	    RECT 137.2000 111.6000 138.0000 111.8000 ;
	    RECT 138.8000 111.2000 139.6000 119.8000 ;
	    RECT 143.0000 115.8000 144.2000 119.8000 ;
	    RECT 147.6000 115.8000 148.4000 119.8000 ;
	    RECT 152.0000 116.4000 152.8000 119.8000 ;
	    RECT 152.0000 115.8000 154.0000 116.4000 ;
	    RECT 143.6000 115.0000 144.4000 115.8000 ;
	    RECT 147.8000 115.2000 148.4000 115.8000 ;
	    RECT 147.0000 114.6000 150.6000 115.2000 ;
	    RECT 153.2000 115.0000 154.0000 115.8000 ;
	    RECT 147.0000 114.4000 147.8000 114.6000 ;
	    RECT 149.8000 114.4000 150.6000 114.6000 ;
	    RECT 142.8000 113.2000 144.2000 114.0000 ;
	    RECT 143.6000 112.2000 144.2000 113.2000 ;
	    RECT 145.8000 113.0000 148.0000 113.6000 ;
	    RECT 145.8000 112.8000 146.6000 113.0000 ;
	    RECT 143.6000 111.6000 146.0000 112.2000 ;
	    RECT 138.8000 110.6000 143.0000 111.2000 ;
	    RECT 126.0000 107.8000 127.0000 108.2000 ;
	    RECT 95.4000 106.6000 96.2000 107.0000 ;
	    RECT 87.8000 106.2000 91.4000 106.6000 ;
	    RECT 82.8000 105.6000 84.6000 106.2000 ;
	    RECT 83.8000 102.2000 84.6000 105.6000 ;
	    RECT 86.0000 102.2000 86.8000 106.2000 ;
	    RECT 87.6000 106.0000 91.6000 106.2000 ;
	    RECT 95.4000 106.0000 97.0000 106.6000 ;
	    RECT 87.6000 102.2000 88.4000 106.0000 ;
	    RECT 90.8000 102.2000 91.6000 106.0000 ;
	    RECT 96.2000 103.0000 97.0000 106.0000 ;
	    RECT 100.6000 105.0000 101.2000 107.2000 ;
	    RECT 110.0000 106.4000 110.6000 107.6000 ;
	    RECT 114.0000 107.2000 114.8000 107.6000 ;
	    RECT 100.4000 103.0000 101.2000 105.0000 ;
	    RECT 108.4000 102.8000 109.2000 106.2000 ;
	    RECT 110.0000 103.4000 110.8000 106.4000 ;
	    RECT 111.8000 106.2000 115.4000 106.6000 ;
	    RECT 116.6000 106.2000 117.2000 107.6000 ;
	    RECT 120.4000 107.2000 121.2000 107.6000 ;
	    RECT 122.8000 107.2000 127.0000 107.8000 ;
	    RECT 128.0000 107.6000 130.0000 108.4000 ;
	    RECT 132.4000 108.2000 133.2000 108.4000 ;
	    RECT 132.4000 107.6000 134.0000 108.2000 ;
	    RECT 135.4000 107.6000 138.0000 108.4000 ;
	    RECT 118.2000 106.2000 121.8000 106.6000 ;
	    RECT 111.6000 106.0000 115.6000 106.2000 ;
	    RECT 111.6000 102.8000 112.4000 106.0000 ;
	    RECT 108.4000 102.2000 112.4000 102.8000 ;
	    RECT 114.8000 102.2000 115.6000 106.0000 ;
	    RECT 116.4000 102.2000 117.2000 106.2000 ;
	    RECT 118.0000 106.0000 122.0000 106.2000 ;
	    RECT 118.0000 102.2000 118.8000 106.0000 ;
	    RECT 121.2000 102.2000 122.0000 106.0000 ;
	    RECT 122.8000 105.0000 123.4000 107.2000 ;
	    RECT 128.0000 107.0000 128.6000 107.6000 ;
	    RECT 133.2000 107.2000 134.0000 107.6000 ;
	    RECT 127.8000 106.6000 128.6000 107.0000 ;
	    RECT 127.0000 106.0000 128.6000 106.6000 ;
	    RECT 132.6000 106.2000 136.2000 106.6000 ;
	    RECT 137.2000 106.2000 137.8000 107.6000 ;
	    RECT 138.8000 107.2000 139.6000 110.6000 ;
	    RECT 142.2000 110.4000 143.0000 110.6000 ;
	    RECT 145.4000 110.4000 146.0000 111.6000 ;
	    RECT 147.4000 111.8000 148.0000 113.0000 ;
	    RECT 148.6000 113.0000 149.4000 113.2000 ;
	    RECT 153.2000 113.0000 154.0000 113.2000 ;
	    RECT 148.6000 112.4000 154.0000 113.0000 ;
	    RECT 147.4000 111.4000 152.2000 111.8000 ;
	    RECT 156.4000 111.4000 157.2000 119.8000 ;
	    RECT 147.4000 111.2000 157.2000 111.4000 ;
	    RECT 151.4000 111.0000 157.2000 111.2000 ;
	    RECT 151.6000 110.8000 157.2000 111.0000 ;
	    RECT 140.6000 109.8000 141.4000 110.0000 ;
	    RECT 140.6000 109.2000 144.4000 109.8000 ;
	    RECT 145.2000 109.6000 146.0000 110.4000 ;
	    RECT 150.0000 110.2000 150.8000 110.4000 ;
	    RECT 159.6000 110.3000 160.4000 119.8000 ;
	    RECT 163.6000 113.6000 164.4000 114.4000 ;
	    RECT 161.2000 111.6000 162.0000 113.2000 ;
	    RECT 163.6000 112.4000 164.2000 113.6000 ;
	    RECT 165.0000 112.4000 165.8000 119.8000 ;
	    RECT 162.8000 111.8000 164.2000 112.4000 ;
	    RECT 164.8000 111.8000 165.8000 112.4000 ;
	    RECT 169.8000 112.6000 170.6000 119.8000 ;
	    RECT 174.6000 112.6000 175.4000 119.8000 ;
	    RECT 179.4000 112.6000 180.2000 119.8000 ;
	    RECT 186.2000 112.6000 187.0000 119.8000 ;
	    RECT 191.0000 112.6000 191.8000 119.8000 ;
	    RECT 169.8000 111.8000 171.6000 112.6000 ;
	    RECT 174.6000 111.8000 176.4000 112.6000 ;
	    RECT 179.4000 111.8000 181.2000 112.6000 ;
	    RECT 185.2000 111.8000 187.0000 112.6000 ;
	    RECT 190.0000 111.8000 191.8000 112.6000 ;
	    RECT 162.8000 111.6000 163.6000 111.8000 ;
	    RECT 162.9000 110.3000 163.5000 111.6000 ;
	    RECT 150.0000 109.6000 155.0000 110.2000 ;
	    RECT 143.6000 109.0000 144.4000 109.2000 ;
	    RECT 145.4000 108.4000 146.0000 109.6000 ;
	    RECT 151.6000 109.4000 152.4000 109.6000 ;
	    RECT 154.2000 109.4000 155.0000 109.6000 ;
	    RECT 159.6000 109.7000 163.5000 110.3000 ;
	    RECT 152.6000 108.4000 153.4000 108.6000 ;
	    RECT 145.4000 107.8000 156.4000 108.4000 ;
	    RECT 145.8000 107.6000 146.6000 107.8000 ;
	    RECT 138.8000 106.6000 142.6000 107.2000 ;
	    RECT 132.4000 106.0000 136.4000 106.2000 ;
	    RECT 122.8000 103.0000 123.6000 105.0000 ;
	    RECT 127.0000 103.0000 127.8000 106.0000 ;
	    RECT 132.4000 102.2000 133.2000 106.0000 ;
	    RECT 135.6000 102.2000 136.4000 106.0000 ;
	    RECT 137.2000 102.2000 138.0000 106.2000 ;
	    RECT 138.8000 102.2000 139.6000 106.6000 ;
	    RECT 141.8000 106.4000 142.6000 106.6000 ;
	    RECT 151.6000 105.6000 152.2000 107.8000 ;
	    RECT 154.8000 107.6000 156.4000 107.8000 ;
	    RECT 149.8000 105.4000 150.6000 105.6000 ;
	    RECT 143.6000 104.2000 144.4000 105.0000 ;
	    RECT 147.8000 104.8000 150.6000 105.4000 ;
	    RECT 151.6000 104.8000 152.4000 105.6000 ;
	    RECT 147.8000 104.2000 148.4000 104.8000 ;
	    RECT 153.2000 104.2000 154.0000 105.0000 ;
	    RECT 143.0000 103.6000 144.4000 104.2000 ;
	    RECT 143.0000 102.2000 144.2000 103.6000 ;
	    RECT 147.6000 102.2000 148.4000 104.2000 ;
	    RECT 152.0000 103.6000 154.0000 104.2000 ;
	    RECT 152.0000 102.2000 152.8000 103.6000 ;
	    RECT 156.4000 102.2000 157.2000 107.0000 ;
	    RECT 158.0000 106.8000 158.8000 108.4000 ;
	    RECT 159.6000 106.2000 160.4000 109.7000 ;
	    RECT 164.8000 108.4000 165.4000 111.8000 ;
	    RECT 166.0000 108.8000 166.8000 110.4000 ;
	    RECT 169.2000 109.6000 170.0000 111.2000 ;
	    RECT 170.8000 108.4000 171.4000 111.8000 ;
	    RECT 174.0000 109.6000 174.8000 111.2000 ;
	    RECT 175.6000 108.4000 176.2000 111.8000 ;
	    RECT 178.8000 109.6000 179.6000 111.2000 ;
	    RECT 180.4000 108.4000 181.0000 111.8000 ;
	    RECT 185.4000 108.4000 186.0000 111.8000 ;
	    RECT 186.8000 109.6000 187.6000 111.2000 ;
	    RECT 190.2000 108.4000 190.8000 111.8000 ;
	    RECT 193.2000 111.2000 194.0000 119.8000 ;
	    RECT 197.4000 115.8000 198.6000 119.8000 ;
	    RECT 202.0000 115.8000 202.8000 119.8000 ;
	    RECT 206.4000 116.4000 207.2000 119.8000 ;
	    RECT 206.4000 115.8000 208.4000 116.4000 ;
	    RECT 198.0000 115.0000 198.8000 115.8000 ;
	    RECT 202.2000 115.2000 202.8000 115.8000 ;
	    RECT 201.4000 114.6000 205.0000 115.2000 ;
	    RECT 207.6000 115.0000 208.4000 115.8000 ;
	    RECT 201.4000 114.4000 202.2000 114.6000 ;
	    RECT 204.2000 114.4000 205.0000 114.6000 ;
	    RECT 197.2000 113.2000 198.6000 114.0000 ;
	    RECT 198.0000 112.2000 198.6000 113.2000 ;
	    RECT 200.2000 113.0000 202.4000 113.6000 ;
	    RECT 200.2000 112.8000 201.0000 113.0000 ;
	    RECT 198.0000 111.6000 200.4000 112.2000 ;
	    RECT 191.6000 109.6000 192.4000 111.2000 ;
	    RECT 193.2000 110.6000 197.4000 111.2000 ;
	    RECT 161.2000 108.3000 162.0000 108.4000 ;
	    RECT 162.8000 108.3000 165.4000 108.4000 ;
	    RECT 161.2000 107.7000 165.4000 108.3000 ;
	    RECT 167.6000 108.3000 168.4000 108.4000 ;
	    RECT 169.2000 108.3000 170.0000 108.4000 ;
	    RECT 167.6000 108.2000 170.0000 108.3000 ;
	    RECT 161.2000 107.6000 162.0000 107.7000 ;
	    RECT 162.8000 107.6000 165.4000 107.7000 ;
	    RECT 166.8000 107.7000 170.0000 108.2000 ;
	    RECT 166.8000 107.6000 168.4000 107.7000 ;
	    RECT 169.2000 107.6000 170.0000 107.7000 ;
	    RECT 170.8000 107.6000 171.6000 108.4000 ;
	    RECT 175.6000 107.6000 176.4000 108.4000 ;
	    RECT 180.4000 107.6000 181.2000 108.4000 ;
	    RECT 183.6000 108.3000 184.4000 108.4000 ;
	    RECT 182.1000 107.7000 184.4000 108.3000 ;
	    RECT 163.0000 106.2000 163.6000 107.6000 ;
	    RECT 166.8000 107.2000 167.6000 107.6000 ;
	    RECT 164.6000 106.2000 168.2000 106.6000 ;
	    RECT 159.6000 105.6000 161.4000 106.2000 ;
	    RECT 160.6000 102.2000 161.4000 105.6000 ;
	    RECT 162.8000 102.2000 163.6000 106.2000 ;
	    RECT 164.4000 106.0000 168.4000 106.2000 ;
	    RECT 164.4000 102.2000 165.2000 106.0000 ;
	    RECT 167.6000 102.2000 168.4000 106.0000 ;
	    RECT 170.8000 104.4000 171.4000 107.6000 ;
	    RECT 172.4000 104.8000 173.2000 106.4000 ;
	    RECT 175.6000 104.4000 176.2000 107.6000 ;
	    RECT 177.2000 104.8000 178.0000 106.4000 ;
	    RECT 178.8000 106.3000 179.6000 106.4000 ;
	    RECT 180.4000 106.3000 181.0000 107.6000 ;
	    RECT 182.1000 106.4000 182.7000 107.7000 ;
	    RECT 183.6000 107.6000 184.4000 107.7000 ;
	    RECT 185.2000 107.6000 186.0000 108.4000 ;
	    RECT 190.0000 107.6000 190.8000 108.4000 ;
	    RECT 178.8000 105.7000 181.1000 106.3000 ;
	    RECT 178.8000 105.6000 179.6000 105.7000 ;
	    RECT 170.8000 102.2000 171.6000 104.4000 ;
	    RECT 175.6000 102.2000 176.4000 104.4000 ;
	    RECT 180.4000 104.2000 181.0000 105.7000 ;
	    RECT 182.0000 104.8000 182.8000 106.4000 ;
	    RECT 183.6000 104.8000 184.4000 106.4000 ;
	    RECT 185.4000 104.4000 186.0000 107.6000 ;
	    RECT 188.4000 104.8000 189.2000 106.4000 ;
	    RECT 190.2000 104.4000 190.8000 107.6000 ;
	    RECT 180.4000 102.2000 181.2000 104.2000 ;
	    RECT 185.2000 102.2000 186.0000 104.4000 ;
	    RECT 190.0000 102.2000 190.8000 104.4000 ;
	    RECT 193.2000 107.2000 194.0000 110.6000 ;
	    RECT 196.6000 110.4000 197.4000 110.6000 ;
	    RECT 195.0000 109.8000 195.8000 110.0000 ;
	    RECT 195.0000 109.2000 198.8000 109.8000 ;
	    RECT 198.0000 109.0000 198.8000 109.2000 ;
	    RECT 199.8000 108.4000 200.4000 111.6000 ;
	    RECT 201.8000 111.8000 202.4000 113.0000 ;
	    RECT 203.0000 113.0000 203.8000 113.2000 ;
	    RECT 207.6000 113.0000 208.4000 113.2000 ;
	    RECT 203.0000 112.4000 208.4000 113.0000 ;
	    RECT 201.8000 111.4000 206.6000 111.8000 ;
	    RECT 210.8000 111.4000 211.6000 119.8000 ;
	    RECT 213.2000 113.6000 214.0000 114.4000 ;
	    RECT 213.2000 112.4000 213.8000 113.6000 ;
	    RECT 214.6000 112.4000 215.4000 119.8000 ;
	    RECT 221.4000 112.6000 222.2000 119.8000 ;
	    RECT 226.2000 112.6000 227.0000 119.8000 ;
	    RECT 231.0000 112.6000 231.8000 119.8000 ;
	    RECT 212.4000 111.8000 213.8000 112.4000 ;
	    RECT 214.4000 111.8000 215.4000 112.4000 ;
	    RECT 220.4000 111.8000 222.2000 112.6000 ;
	    RECT 225.2000 111.8000 227.0000 112.6000 ;
	    RECT 230.0000 111.8000 231.8000 112.6000 ;
	    RECT 233.8000 112.6000 234.6000 119.8000 ;
	    RECT 240.6000 112.6000 241.4000 119.8000 ;
	    RECT 233.8000 111.8000 235.6000 112.6000 ;
	    RECT 239.6000 111.8000 241.4000 112.6000 ;
	    RECT 245.4000 112.4000 246.2000 119.8000 ;
	    RECT 246.8000 113.6000 247.6000 114.4000 ;
	    RECT 247.0000 112.4000 247.6000 113.6000 ;
	    RECT 245.4000 111.8000 246.4000 112.4000 ;
	    RECT 247.0000 111.8000 248.4000 112.4000 ;
	    RECT 212.4000 111.6000 213.2000 111.8000 ;
	    RECT 201.8000 111.2000 211.6000 111.4000 ;
	    RECT 205.8000 111.0000 211.6000 111.2000 ;
	    RECT 206.0000 110.8000 211.6000 111.0000 ;
	    RECT 204.4000 110.2000 205.2000 110.4000 ;
	    RECT 212.4000 110.3000 213.2000 110.4000 ;
	    RECT 214.4000 110.3000 215.0000 111.8000 ;
	    RECT 204.4000 109.6000 209.4000 110.2000 ;
	    RECT 212.4000 109.7000 215.0000 110.3000 ;
	    RECT 212.4000 109.6000 213.2000 109.7000 ;
	    RECT 206.0000 109.4000 206.8000 109.6000 ;
	    RECT 208.6000 109.4000 209.4000 109.6000 ;
	    RECT 207.0000 108.4000 207.8000 108.6000 ;
	    RECT 214.4000 108.4000 215.0000 109.7000 ;
	    RECT 215.6000 110.3000 216.4000 110.4000 ;
	    RECT 217.2000 110.3000 218.0000 110.4000 ;
	    RECT 215.6000 109.7000 218.0000 110.3000 ;
	    RECT 215.6000 108.8000 216.4000 109.7000 ;
	    RECT 217.2000 109.6000 218.0000 109.7000 ;
	    RECT 220.6000 108.4000 221.2000 111.8000 ;
	    RECT 222.0000 109.6000 222.8000 111.2000 ;
	    RECT 225.4000 108.4000 226.0000 111.8000 ;
	    RECT 226.8000 110.3000 227.6000 111.2000 ;
	    RECT 228.4000 110.3000 229.2000 110.4000 ;
	    RECT 226.8000 109.7000 229.2000 110.3000 ;
	    RECT 226.8000 109.6000 227.6000 109.7000 ;
	    RECT 228.4000 109.6000 229.2000 109.7000 ;
	    RECT 230.2000 108.4000 230.8000 111.8000 ;
	    RECT 231.6000 109.6000 232.4000 111.2000 ;
	    RECT 233.2000 109.6000 234.0000 111.2000 ;
	    RECT 199.8000 107.8000 210.8000 108.4000 ;
	    RECT 200.2000 107.6000 201.0000 107.8000 ;
	    RECT 202.8000 107.6000 203.6000 107.8000 ;
	    RECT 193.2000 106.6000 197.0000 107.2000 ;
	    RECT 193.2000 102.2000 194.0000 106.6000 ;
	    RECT 196.2000 106.4000 197.0000 106.6000 ;
	    RECT 206.0000 105.6000 206.6000 107.8000 ;
	    RECT 209.2000 107.6000 210.8000 107.8000 ;
	    RECT 212.4000 107.6000 215.0000 108.4000 ;
	    RECT 217.2000 108.2000 218.0000 108.4000 ;
	    RECT 216.4000 107.6000 218.0000 108.2000 ;
	    RECT 220.4000 107.6000 221.2000 108.4000 ;
	    RECT 225.2000 107.6000 226.0000 108.4000 ;
	    RECT 230.0000 107.6000 230.8000 108.4000 ;
	    RECT 204.2000 105.4000 205.0000 105.6000 ;
	    RECT 198.0000 104.2000 198.8000 105.0000 ;
	    RECT 202.2000 104.8000 205.0000 105.4000 ;
	    RECT 206.0000 104.8000 206.8000 105.6000 ;
	    RECT 202.2000 104.2000 202.8000 104.8000 ;
	    RECT 207.6000 104.2000 208.4000 105.0000 ;
	    RECT 197.4000 103.6000 198.8000 104.2000 ;
	    RECT 197.4000 102.2000 198.6000 103.6000 ;
	    RECT 202.0000 102.2000 202.8000 104.2000 ;
	    RECT 206.4000 103.6000 208.4000 104.2000 ;
	    RECT 206.4000 102.2000 207.2000 103.6000 ;
	    RECT 210.8000 102.2000 211.6000 107.0000 ;
	    RECT 212.6000 106.2000 213.2000 107.6000 ;
	    RECT 216.4000 107.2000 217.2000 107.6000 ;
	    RECT 214.2000 106.2000 217.8000 106.6000 ;
	    RECT 212.4000 102.2000 213.2000 106.2000 ;
	    RECT 214.0000 106.0000 218.0000 106.2000 ;
	    RECT 214.0000 102.2000 214.8000 106.0000 ;
	    RECT 217.2000 102.2000 218.0000 106.0000 ;
	    RECT 218.8000 104.8000 219.6000 106.4000 ;
	    RECT 220.6000 104.4000 221.2000 107.6000 ;
	    RECT 223.6000 104.8000 224.4000 106.4000 ;
	    RECT 225.4000 104.4000 226.0000 107.6000 ;
	    RECT 228.4000 104.8000 229.2000 106.4000 ;
	    RECT 230.2000 106.3000 230.8000 107.6000 ;
	    RECT 234.8000 108.4000 235.4000 111.8000 ;
	    RECT 236.4000 110.3000 237.2000 110.4000 ;
	    RECT 239.8000 110.3000 240.4000 111.8000 ;
	    RECT 236.4000 109.7000 240.4000 110.3000 ;
	    RECT 236.4000 109.6000 237.2000 109.7000 ;
	    RECT 239.8000 108.4000 240.4000 109.7000 ;
	    RECT 241.2000 109.6000 242.0000 111.2000 ;
	    RECT 245.8000 110.4000 246.4000 111.8000 ;
	    RECT 247.6000 111.6000 248.4000 111.8000 ;
	    RECT 255.6000 111.4000 256.4000 119.8000 ;
	    RECT 260.0000 116.4000 260.8000 119.8000 ;
	    RECT 258.8000 115.8000 260.8000 116.4000 ;
	    RECT 264.4000 115.8000 265.2000 119.8000 ;
	    RECT 268.6000 115.8000 269.8000 119.8000 ;
	    RECT 258.8000 115.0000 259.6000 115.8000 ;
	    RECT 264.4000 115.2000 265.0000 115.8000 ;
	    RECT 262.2000 114.6000 265.8000 115.2000 ;
	    RECT 268.4000 115.0000 269.2000 115.8000 ;
	    RECT 262.2000 114.4000 263.0000 114.6000 ;
	    RECT 265.0000 114.4000 265.8000 114.6000 ;
	    RECT 258.8000 113.0000 259.6000 113.2000 ;
	    RECT 263.4000 113.0000 264.2000 113.2000 ;
	    RECT 258.8000 112.4000 264.2000 113.0000 ;
	    RECT 264.8000 113.0000 267.0000 113.6000 ;
	    RECT 264.8000 111.8000 265.4000 113.0000 ;
	    RECT 266.2000 112.8000 267.0000 113.0000 ;
	    RECT 268.6000 113.2000 270.0000 114.0000 ;
	    RECT 268.6000 112.2000 269.2000 113.2000 ;
	    RECT 260.6000 111.4000 265.4000 111.8000 ;
	    RECT 255.6000 111.2000 265.4000 111.4000 ;
	    RECT 266.8000 111.6000 269.2000 112.2000 ;
	    RECT 255.6000 111.0000 261.4000 111.2000 ;
	    RECT 255.6000 110.8000 261.2000 111.0000 ;
	    RECT 242.8000 110.3000 243.6000 110.4000 ;
	    RECT 244.4000 110.3000 245.2000 110.4000 ;
	    RECT 242.8000 109.7000 245.2000 110.3000 ;
	    RECT 242.8000 109.6000 243.6000 109.7000 ;
	    RECT 244.4000 108.8000 245.2000 109.7000 ;
	    RECT 245.8000 109.6000 246.8000 110.4000 ;
	    RECT 262.0000 110.2000 262.8000 110.4000 ;
	    RECT 257.8000 109.6000 262.8000 110.2000 ;
	    RECT 245.8000 108.4000 246.4000 109.6000 ;
	    RECT 257.8000 109.4000 258.6000 109.6000 ;
	    RECT 260.4000 109.4000 261.2000 109.6000 ;
	    RECT 259.4000 108.4000 260.2000 108.6000 ;
	    RECT 266.8000 108.4000 267.4000 111.6000 ;
	    RECT 273.2000 111.2000 274.0000 119.8000 ;
	    RECT 274.8000 112.4000 275.6000 119.8000 ;
	    RECT 274.8000 111.8000 277.0000 112.4000 ;
	    RECT 278.0000 111.8000 278.8000 119.8000 ;
	    RECT 283.4000 112.8000 284.2000 119.8000 ;
	    RECT 287.6000 115.0000 288.4000 119.0000 ;
	    RECT 269.8000 110.6000 274.0000 111.2000 ;
	    RECT 269.8000 110.4000 270.6000 110.6000 ;
	    RECT 271.4000 109.8000 272.2000 110.0000 ;
	    RECT 268.4000 109.2000 272.2000 109.8000 ;
	    RECT 268.4000 109.0000 269.2000 109.2000 ;
	    RECT 234.8000 107.6000 235.6000 108.4000 ;
	    RECT 239.6000 107.6000 240.4000 108.4000 ;
	    RECT 242.8000 108.2000 243.6000 108.4000 ;
	    RECT 242.8000 107.6000 244.4000 108.2000 ;
	    RECT 245.8000 107.6000 248.4000 108.4000 ;
	    RECT 256.4000 107.8000 267.4000 108.4000 ;
	    RECT 256.4000 107.6000 258.0000 107.8000 ;
	    RECT 231.6000 106.3000 232.4000 106.4000 ;
	    RECT 230.1000 105.7000 232.4000 106.3000 ;
	    RECT 220.4000 102.2000 221.2000 104.4000 ;
	    RECT 225.2000 102.2000 226.0000 104.4000 ;
	    RECT 230.2000 104.2000 230.8000 105.7000 ;
	    RECT 231.6000 105.6000 232.4000 105.7000 ;
	    RECT 233.2000 106.3000 234.0000 106.4000 ;
	    RECT 234.8000 106.3000 235.4000 107.6000 ;
	    RECT 236.4000 106.3000 237.2000 106.4000 ;
	    RECT 238.0000 106.3000 238.8000 106.4000 ;
	    RECT 233.2000 105.7000 235.5000 106.3000 ;
	    RECT 236.4000 105.7000 238.8000 106.3000 ;
	    RECT 233.2000 105.6000 234.0000 105.7000 ;
	    RECT 230.0000 102.2000 230.8000 104.2000 ;
	    RECT 234.8000 104.2000 235.4000 105.7000 ;
	    RECT 236.4000 104.8000 237.2000 105.7000 ;
	    RECT 238.0000 104.8000 238.8000 105.7000 ;
	    RECT 239.8000 104.2000 240.4000 107.6000 ;
	    RECT 243.6000 107.2000 244.4000 107.6000 ;
	    RECT 243.0000 106.2000 246.6000 106.6000 ;
	    RECT 247.6000 106.2000 248.2000 107.6000 ;
	    RECT 234.8000 102.2000 235.6000 104.2000 ;
	    RECT 239.6000 102.2000 240.4000 104.2000 ;
	    RECT 242.8000 106.0000 246.8000 106.2000 ;
	    RECT 242.8000 102.2000 243.6000 106.0000 ;
	    RECT 246.0000 102.2000 246.8000 106.0000 ;
	    RECT 247.6000 102.2000 248.4000 106.2000 ;
	    RECT 255.6000 102.2000 256.4000 107.0000 ;
	    RECT 260.6000 105.6000 261.2000 107.8000 ;
	    RECT 262.0000 107.6000 262.8000 107.8000 ;
	    RECT 266.2000 107.6000 267.0000 107.8000 ;
	    RECT 273.2000 107.2000 274.0000 110.6000 ;
	    RECT 276.4000 111.2000 277.0000 111.8000 ;
	    RECT 276.4000 110.4000 277.6000 111.2000 ;
	    RECT 274.8000 108.8000 275.6000 110.4000 ;
	    RECT 276.4000 107.4000 277.0000 110.4000 ;
	    RECT 278.2000 109.6000 278.8000 111.8000 ;
	    RECT 282.6000 112.2000 284.2000 112.8000 ;
	    RECT 281.2000 109.6000 282.0000 111.2000 ;
	    RECT 270.0000 106.6000 274.0000 107.2000 ;
	    RECT 270.0000 106.4000 271.0000 106.6000 ;
	    RECT 270.0000 105.6000 270.8000 106.4000 ;
	    RECT 258.8000 104.2000 259.6000 105.0000 ;
	    RECT 260.4000 104.8000 261.2000 105.6000 ;
	    RECT 262.2000 105.4000 263.0000 105.6000 ;
	    RECT 262.2000 104.8000 265.0000 105.4000 ;
	    RECT 264.4000 104.2000 265.0000 104.8000 ;
	    RECT 268.4000 104.2000 269.2000 105.0000 ;
	    RECT 258.8000 103.6000 260.8000 104.2000 ;
	    RECT 260.0000 102.2000 260.8000 103.6000 ;
	    RECT 264.4000 102.2000 265.2000 104.2000 ;
	    RECT 268.4000 103.6000 269.8000 104.2000 ;
	    RECT 268.6000 102.2000 269.8000 103.6000 ;
	    RECT 273.2000 102.2000 274.0000 106.6000 ;
	    RECT 274.8000 106.8000 277.0000 107.4000 ;
	    RECT 274.8000 102.2000 275.6000 106.8000 ;
	    RECT 278.0000 102.2000 278.8000 109.6000 ;
	    RECT 282.6000 108.4000 283.2000 112.2000 ;
	    RECT 287.8000 111.6000 288.4000 115.0000 ;
	    RECT 284.6000 111.0000 288.4000 111.6000 ;
	    RECT 289.2000 115.0000 290.0000 119.0000 ;
	    RECT 289.2000 111.6000 289.8000 115.0000 ;
	    RECT 293.4000 114.4000 294.2000 119.8000 ;
	    RECT 301.4000 116.4000 303.4000 119.8000 ;
	    RECT 300.4000 115.6000 303.4000 116.4000 ;
	    RECT 293.4000 113.6000 294.8000 114.4000 ;
	    RECT 293.4000 112.8000 294.2000 113.6000 ;
	    RECT 293.4000 112.2000 295.0000 112.8000 ;
	    RECT 289.2000 111.0000 293.0000 111.6000 ;
	    RECT 284.6000 109.0000 285.2000 111.0000 ;
	    RECT 281.2000 107.6000 283.2000 108.4000 ;
	    RECT 283.8000 108.2000 285.2000 109.0000 ;
	    RECT 286.0000 108.8000 286.8000 110.4000 ;
	    RECT 287.6000 108.8000 288.4000 110.4000 ;
	    RECT 289.2000 108.8000 290.0000 110.4000 ;
	    RECT 290.8000 108.8000 291.6000 110.4000 ;
	    RECT 292.4000 109.0000 293.0000 111.0000 ;
	    RECT 282.6000 107.0000 283.2000 107.6000 ;
	    RECT 284.2000 107.8000 285.2000 108.2000 ;
	    RECT 292.4000 108.2000 293.8000 109.0000 ;
	    RECT 294.4000 108.4000 295.0000 112.2000 ;
	    RECT 301.4000 111.8000 303.4000 115.6000 ;
	    RECT 309.4000 112.4000 310.2000 119.8000 ;
	    RECT 310.8000 113.6000 311.6000 114.4000 ;
	    RECT 311.0000 112.4000 311.6000 113.6000 ;
	    RECT 313.8000 112.6000 314.6000 119.8000 ;
	    RECT 309.4000 111.8000 310.4000 112.4000 ;
	    RECT 311.0000 111.8000 312.4000 112.4000 ;
	    RECT 313.8000 111.8000 315.6000 112.6000 ;
	    RECT 320.6000 112.4000 321.4000 119.8000 ;
	    RECT 322.0000 113.6000 322.8000 114.4000 ;
	    RECT 322.2000 112.4000 322.8000 113.6000 ;
	    RECT 320.6000 111.8000 321.6000 112.4000 ;
	    RECT 322.2000 111.8000 323.6000 112.4000 ;
	    RECT 295.6000 109.6000 296.4000 111.2000 ;
	    RECT 292.4000 107.8000 293.4000 108.2000 ;
	    RECT 284.2000 107.2000 288.4000 107.8000 ;
	    RECT 282.6000 106.6000 283.4000 107.0000 ;
	    RECT 282.6000 106.0000 284.2000 106.6000 ;
	    RECT 283.4000 104.4000 284.2000 106.0000 ;
	    RECT 287.8000 105.0000 288.4000 107.2000 ;
	    RECT 282.8000 103.6000 284.2000 104.4000 ;
	    RECT 283.4000 103.0000 284.2000 103.6000 ;
	    RECT 287.6000 103.0000 288.4000 105.0000 ;
	    RECT 289.2000 107.2000 293.4000 107.8000 ;
	    RECT 294.4000 107.6000 296.4000 108.4000 ;
	    RECT 297.2000 108.3000 298.0000 108.4000 ;
	    RECT 298.8000 108.3000 299.6000 109.2000 ;
	    RECT 300.4000 108.8000 301.2000 110.4000 ;
	    RECT 302.2000 108.4000 302.8000 111.8000 ;
	    RECT 303.6000 108.8000 304.4000 110.4000 ;
	    RECT 306.8000 110.3000 307.6000 110.4000 ;
	    RECT 308.4000 110.3000 309.2000 110.4000 ;
	    RECT 306.8000 109.7000 309.2000 110.3000 ;
	    RECT 306.8000 109.6000 307.6000 109.7000 ;
	    RECT 308.4000 108.8000 309.2000 109.7000 ;
	    RECT 309.8000 108.4000 310.4000 111.8000 ;
	    RECT 311.6000 111.6000 312.4000 111.8000 ;
	    RECT 313.2000 109.6000 314.0000 111.2000 ;
	    RECT 314.8000 108.4000 315.4000 111.8000 ;
	    RECT 319.6000 108.8000 320.4000 110.4000 ;
	    RECT 321.0000 108.4000 321.6000 111.8000 ;
	    RECT 322.8000 111.6000 323.6000 111.8000 ;
	    RECT 324.4000 111.8000 325.2000 119.8000 ;
	    RECT 327.6000 112.4000 328.4000 119.8000 ;
	    RECT 326.2000 111.8000 328.4000 112.4000 ;
	    RECT 329.2000 112.4000 330.0000 119.8000 ;
	    RECT 329.2000 111.8000 331.4000 112.4000 ;
	    RECT 332.4000 111.8000 333.2000 119.8000 ;
	    RECT 324.4000 109.6000 325.0000 111.8000 ;
	    RECT 326.2000 111.2000 326.8000 111.8000 ;
	    RECT 325.6000 110.4000 326.8000 111.2000 ;
	    RECT 297.2000 107.7000 299.6000 108.3000 ;
	    RECT 302.0000 108.2000 302.8000 108.4000 ;
	    RECT 305.2000 108.2000 306.0000 108.4000 ;
	    RECT 297.2000 107.6000 298.0000 107.7000 ;
	    RECT 298.8000 107.6000 299.6000 107.7000 ;
	    RECT 300.4000 107.6000 302.8000 108.2000 ;
	    RECT 304.4000 107.6000 306.0000 108.2000 ;
	    RECT 306.8000 108.2000 307.6000 108.4000 ;
	    RECT 306.8000 107.6000 308.4000 108.2000 ;
	    RECT 309.8000 107.6000 312.4000 108.4000 ;
	    RECT 314.8000 107.6000 315.6000 108.4000 ;
	    RECT 318.0000 108.2000 318.8000 108.4000 ;
	    RECT 318.0000 107.6000 319.6000 108.2000 ;
	    RECT 321.0000 107.6000 323.6000 108.4000 ;
	    RECT 289.2000 105.0000 289.8000 107.2000 ;
	    RECT 294.4000 107.0000 295.0000 107.6000 ;
	    RECT 294.2000 106.6000 295.0000 107.0000 ;
	    RECT 293.4000 106.0000 295.0000 106.6000 ;
	    RECT 300.4000 106.2000 301.0000 107.6000 ;
	    RECT 304.4000 107.2000 305.2000 107.6000 ;
	    RECT 307.6000 107.2000 308.4000 107.6000 ;
	    RECT 302.2000 106.2000 305.8000 106.6000 ;
	    RECT 307.0000 106.2000 310.6000 106.6000 ;
	    RECT 311.6000 106.2000 312.2000 107.6000 ;
	    RECT 313.2000 106.3000 314.0000 106.4000 ;
	    RECT 314.8000 106.3000 315.4000 107.6000 ;
	    RECT 318.8000 107.2000 319.6000 107.6000 ;
	    RECT 289.2000 103.0000 290.0000 105.0000 ;
	    RECT 293.4000 103.0000 294.2000 106.0000 ;
	    RECT 298.8000 102.8000 299.6000 106.2000 ;
	    RECT 300.4000 103.4000 301.2000 106.2000 ;
	    RECT 302.0000 106.0000 306.0000 106.2000 ;
	    RECT 302.0000 102.8000 302.8000 106.0000 ;
	    RECT 298.8000 102.2000 302.8000 102.8000 ;
	    RECT 305.2000 102.2000 306.0000 106.0000 ;
	    RECT 306.8000 106.0000 310.8000 106.2000 ;
	    RECT 306.8000 102.2000 307.6000 106.0000 ;
	    RECT 310.0000 102.2000 310.8000 106.0000 ;
	    RECT 311.6000 102.2000 312.4000 106.2000 ;
	    RECT 313.2000 105.7000 315.5000 106.3000 ;
	    RECT 313.2000 105.6000 314.0000 105.7000 ;
	    RECT 314.8000 104.2000 315.4000 105.7000 ;
	    RECT 316.4000 104.8000 317.2000 106.4000 ;
	    RECT 318.2000 106.2000 321.8000 106.6000 ;
	    RECT 322.8000 106.2000 323.4000 107.6000 ;
	    RECT 318.0000 106.0000 322.0000 106.2000 ;
	    RECT 314.8000 102.2000 315.6000 104.2000 ;
	    RECT 318.0000 102.2000 318.8000 106.0000 ;
	    RECT 321.2000 102.2000 322.0000 106.0000 ;
	    RECT 322.8000 102.2000 323.6000 106.2000 ;
	    RECT 324.4000 102.2000 325.2000 109.6000 ;
	    RECT 326.2000 107.4000 326.8000 110.4000 ;
	    RECT 330.8000 111.2000 331.4000 111.8000 ;
	    RECT 330.8000 110.4000 332.0000 111.2000 ;
	    RECT 330.8000 107.4000 331.4000 110.4000 ;
	    RECT 332.6000 109.6000 333.2000 111.8000 ;
	    RECT 326.2000 106.8000 328.4000 107.4000 ;
	    RECT 327.6000 102.2000 328.4000 106.8000 ;
	    RECT 329.2000 106.8000 331.4000 107.4000 ;
	    RECT 329.2000 102.2000 330.0000 106.8000 ;
	    RECT 332.4000 102.2000 333.2000 109.6000 ;
	    RECT 334.0000 111.2000 334.8000 119.8000 ;
	    RECT 338.2000 115.8000 339.4000 119.8000 ;
	    RECT 342.8000 115.8000 343.6000 119.8000 ;
	    RECT 347.2000 116.4000 348.0000 119.8000 ;
	    RECT 347.2000 115.8000 349.2000 116.4000 ;
	    RECT 338.8000 115.0000 339.6000 115.8000 ;
	    RECT 343.0000 115.2000 343.6000 115.8000 ;
	    RECT 342.2000 114.6000 345.8000 115.2000 ;
	    RECT 348.4000 115.0000 349.2000 115.8000 ;
	    RECT 342.2000 114.4000 343.0000 114.6000 ;
	    RECT 345.0000 114.4000 345.8000 114.6000 ;
	    RECT 338.0000 113.2000 339.4000 114.0000 ;
	    RECT 338.8000 112.2000 339.4000 113.2000 ;
	    RECT 341.0000 113.0000 343.2000 113.6000 ;
	    RECT 341.0000 112.8000 341.8000 113.0000 ;
	    RECT 338.8000 111.6000 341.2000 112.2000 ;
	    RECT 334.0000 110.6000 338.2000 111.2000 ;
	    RECT 334.0000 107.2000 334.8000 110.6000 ;
	    RECT 337.4000 110.4000 338.2000 110.6000 ;
	    RECT 335.8000 109.8000 336.6000 110.0000 ;
	    RECT 335.8000 109.2000 339.6000 109.8000 ;
	    RECT 338.8000 109.0000 339.6000 109.2000 ;
	    RECT 340.6000 108.4000 341.2000 111.6000 ;
	    RECT 342.6000 111.8000 343.2000 113.0000 ;
	    RECT 343.8000 113.0000 344.6000 113.2000 ;
	    RECT 348.4000 113.0000 349.2000 113.2000 ;
	    RECT 343.8000 112.4000 349.2000 113.0000 ;
	    RECT 342.6000 111.4000 347.4000 111.8000 ;
	    RECT 351.6000 111.4000 352.4000 119.8000 ;
	    RECT 355.8000 112.4000 356.6000 119.8000 ;
	    RECT 359.6000 115.0000 360.4000 119.0000 ;
	    RECT 357.2000 113.6000 358.0000 114.4000 ;
	    RECT 357.4000 112.4000 358.0000 113.6000 ;
	    RECT 354.8000 111.6000 356.8000 112.4000 ;
	    RECT 357.4000 111.8000 358.8000 112.4000 ;
	    RECT 358.0000 111.6000 358.8000 111.8000 ;
	    RECT 359.6000 111.6000 360.2000 115.0000 ;
	    RECT 363.8000 112.8000 364.6000 119.8000 ;
	    RECT 369.2000 115.0000 370.0000 119.0000 ;
	    RECT 363.8000 112.2000 365.4000 112.8000 ;
	    RECT 342.6000 111.2000 352.4000 111.4000 ;
	    RECT 346.6000 111.0000 352.4000 111.2000 ;
	    RECT 346.8000 110.8000 352.4000 111.0000 ;
	    RECT 345.2000 110.2000 346.0000 110.4000 ;
	    RECT 345.2000 109.6000 350.2000 110.2000 ;
	    RECT 346.8000 109.4000 347.6000 109.6000 ;
	    RECT 349.4000 109.4000 350.2000 109.6000 ;
	    RECT 354.8000 108.8000 355.6000 110.4000 ;
	    RECT 347.8000 108.4000 348.6000 108.6000 ;
	    RECT 356.2000 108.4000 356.8000 111.6000 ;
	    RECT 359.6000 111.0000 363.4000 111.6000 ;
	    RECT 359.6000 108.8000 360.4000 110.4000 ;
	    RECT 361.2000 108.8000 362.0000 110.4000 ;
	    RECT 362.8000 109.0000 363.4000 111.0000 ;
	    RECT 340.6000 107.8000 351.6000 108.4000 ;
	    RECT 341.0000 107.6000 341.8000 107.8000 ;
	    RECT 346.8000 107.6000 347.6000 107.8000 ;
	    RECT 350.0000 107.6000 351.6000 107.8000 ;
	    RECT 353.2000 108.2000 354.0000 108.4000 ;
	    RECT 353.2000 107.6000 354.8000 108.2000 ;
	    RECT 356.2000 107.6000 358.8000 108.4000 ;
	    RECT 362.8000 108.2000 364.2000 109.0000 ;
	    RECT 364.8000 108.4000 365.4000 112.2000 ;
	    RECT 369.2000 111.6000 369.8000 115.0000 ;
	    RECT 373.4000 112.8000 374.2000 119.8000 ;
	    RECT 373.4000 112.2000 375.0000 112.8000 ;
	    RECT 366.0000 109.6000 366.8000 111.2000 ;
	    RECT 369.2000 111.0000 373.0000 111.6000 ;
	    RECT 369.2000 108.8000 370.0000 110.4000 ;
	    RECT 370.8000 108.8000 371.6000 110.4000 ;
	    RECT 372.4000 109.0000 373.0000 111.0000 ;
	    RECT 362.8000 107.8000 363.8000 108.2000 ;
	    RECT 334.0000 106.6000 337.8000 107.2000 ;
	    RECT 334.0000 102.2000 334.8000 106.6000 ;
	    RECT 337.0000 106.4000 337.8000 106.6000 ;
	    RECT 346.8000 105.6000 347.4000 107.6000 ;
	    RECT 354.0000 107.2000 354.8000 107.6000 ;
	    RECT 345.0000 105.4000 345.8000 105.6000 ;
	    RECT 338.8000 104.2000 339.6000 105.0000 ;
	    RECT 343.0000 104.8000 345.8000 105.4000 ;
	    RECT 346.8000 104.8000 347.6000 105.6000 ;
	    RECT 343.0000 104.2000 343.6000 104.8000 ;
	    RECT 348.4000 104.2000 349.2000 105.0000 ;
	    RECT 338.2000 103.6000 339.6000 104.2000 ;
	    RECT 338.2000 102.2000 339.4000 103.6000 ;
	    RECT 342.8000 102.2000 343.6000 104.2000 ;
	    RECT 347.2000 103.6000 349.2000 104.2000 ;
	    RECT 347.2000 102.2000 348.0000 103.6000 ;
	    RECT 351.6000 102.2000 352.4000 107.0000 ;
	    RECT 353.4000 106.2000 357.0000 106.6000 ;
	    RECT 358.0000 106.2000 358.6000 107.6000 ;
	    RECT 359.6000 107.2000 363.8000 107.8000 ;
	    RECT 364.8000 107.6000 366.8000 108.4000 ;
	    RECT 372.4000 108.2000 373.8000 109.0000 ;
	    RECT 374.4000 108.4000 375.0000 112.2000 ;
	    RECT 378.8000 111.2000 379.6000 119.8000 ;
	    RECT 383.0000 115.8000 384.2000 119.8000 ;
	    RECT 387.6000 115.8000 388.4000 119.8000 ;
	    RECT 392.0000 116.4000 392.8000 119.8000 ;
	    RECT 392.0000 115.8000 394.0000 116.4000 ;
	    RECT 383.6000 115.0000 384.4000 115.8000 ;
	    RECT 387.8000 115.2000 388.4000 115.8000 ;
	    RECT 387.0000 114.6000 390.6000 115.2000 ;
	    RECT 393.2000 115.0000 394.0000 115.8000 ;
	    RECT 387.0000 114.4000 387.8000 114.6000 ;
	    RECT 389.8000 114.4000 390.6000 114.6000 ;
	    RECT 382.8000 113.2000 384.2000 114.0000 ;
	    RECT 383.6000 112.2000 384.2000 113.2000 ;
	    RECT 385.8000 113.0000 388.0000 113.6000 ;
	    RECT 385.8000 112.8000 386.6000 113.0000 ;
	    RECT 383.6000 111.6000 386.0000 112.2000 ;
	    RECT 375.6000 109.6000 376.4000 111.2000 ;
	    RECT 378.8000 110.6000 383.0000 111.2000 ;
	    RECT 372.4000 107.8000 373.4000 108.2000 ;
	    RECT 353.2000 106.0000 357.2000 106.2000 ;
	    RECT 353.2000 102.2000 354.0000 106.0000 ;
	    RECT 356.4000 102.2000 357.2000 106.0000 ;
	    RECT 358.0000 102.2000 358.8000 106.2000 ;
	    RECT 359.6000 105.0000 360.2000 107.2000 ;
	    RECT 364.8000 107.0000 365.4000 107.6000 ;
	    RECT 364.6000 106.6000 365.4000 107.0000 ;
	    RECT 363.8000 106.0000 365.4000 106.6000 ;
	    RECT 369.2000 107.2000 373.4000 107.8000 ;
	    RECT 374.4000 107.6000 376.4000 108.4000 ;
	    RECT 359.6000 103.0000 360.4000 105.0000 ;
	    RECT 363.8000 104.4000 364.6000 106.0000 ;
	    RECT 362.8000 103.6000 364.6000 104.4000 ;
	    RECT 363.8000 103.0000 364.6000 103.6000 ;
	    RECT 369.2000 105.0000 369.8000 107.2000 ;
	    RECT 374.4000 107.0000 375.0000 107.6000 ;
	    RECT 374.2000 106.6000 375.0000 107.0000 ;
	    RECT 373.4000 106.4000 375.0000 106.6000 ;
	    RECT 372.4000 106.0000 375.0000 106.4000 ;
	    RECT 378.8000 107.2000 379.6000 110.6000 ;
	    RECT 382.2000 110.4000 383.0000 110.6000 ;
	    RECT 380.6000 109.8000 381.4000 110.0000 ;
	    RECT 380.6000 109.2000 384.4000 109.8000 ;
	    RECT 383.6000 109.0000 384.4000 109.2000 ;
	    RECT 385.4000 108.4000 386.0000 111.6000 ;
	    RECT 387.4000 111.8000 388.0000 113.0000 ;
	    RECT 388.6000 113.0000 389.4000 113.2000 ;
	    RECT 393.2000 113.0000 394.0000 113.2000 ;
	    RECT 388.6000 112.4000 394.0000 113.0000 ;
	    RECT 387.4000 111.4000 392.2000 111.8000 ;
	    RECT 396.4000 111.4000 397.2000 119.8000 ;
	    RECT 398.8000 113.6000 399.6000 114.4000 ;
	    RECT 398.8000 112.4000 399.4000 113.6000 ;
	    RECT 400.2000 112.4000 401.0000 119.8000 ;
	    RECT 404.4000 118.3000 405.2000 118.4000 ;
	    RECT 410.8000 118.3000 411.6000 119.8000 ;
	    RECT 404.4000 117.7000 411.6000 118.3000 ;
	    RECT 404.4000 117.6000 405.2000 117.7000 ;
	    RECT 398.0000 111.8000 399.4000 112.4000 ;
	    RECT 400.0000 111.8000 401.0000 112.4000 ;
	    RECT 398.0000 111.6000 398.8000 111.8000 ;
	    RECT 387.4000 111.2000 397.2000 111.4000 ;
	    RECT 391.4000 111.0000 397.2000 111.2000 ;
	    RECT 391.6000 110.8000 397.2000 111.0000 ;
	    RECT 390.0000 110.2000 390.8000 110.4000 ;
	    RECT 390.0000 109.6000 395.0000 110.2000 ;
	    RECT 394.2000 109.4000 395.0000 109.6000 ;
	    RECT 392.6000 108.4000 393.4000 108.6000 ;
	    RECT 400.0000 108.4000 400.6000 111.8000 ;
	    RECT 410.8000 111.2000 411.6000 117.7000 ;
	    RECT 415.0000 115.8000 416.2000 119.8000 ;
	    RECT 419.6000 115.8000 420.4000 119.8000 ;
	    RECT 424.0000 116.4000 424.8000 119.8000 ;
	    RECT 424.0000 115.8000 426.0000 116.4000 ;
	    RECT 415.6000 115.0000 416.4000 115.8000 ;
	    RECT 419.8000 115.2000 420.4000 115.8000 ;
	    RECT 419.0000 114.6000 422.6000 115.2000 ;
	    RECT 425.2000 115.0000 426.0000 115.8000 ;
	    RECT 419.0000 114.4000 419.8000 114.6000 ;
	    RECT 421.8000 114.4000 422.6000 114.6000 ;
	    RECT 414.8000 113.2000 416.2000 114.0000 ;
	    RECT 415.6000 112.2000 416.2000 113.2000 ;
	    RECT 417.8000 113.0000 420.0000 113.6000 ;
	    RECT 417.8000 112.8000 418.6000 113.0000 ;
	    RECT 415.6000 111.6000 418.0000 112.2000 ;
	    RECT 410.8000 110.6000 415.0000 111.2000 ;
	    RECT 401.2000 108.8000 402.0000 110.4000 ;
	    RECT 385.4000 107.8000 396.4000 108.4000 ;
	    RECT 385.8000 107.6000 386.6000 107.8000 ;
	    RECT 391.6000 107.6000 392.4000 107.8000 ;
	    RECT 394.8000 107.6000 396.4000 107.8000 ;
	    RECT 398.0000 107.6000 400.6000 108.4000 ;
	    RECT 402.8000 108.3000 403.6000 108.4000 ;
	    RECT 407.6000 108.3000 408.4000 108.4000 ;
	    RECT 402.8000 108.2000 408.4000 108.3000 ;
	    RECT 402.0000 107.7000 408.4000 108.2000 ;
	    RECT 402.0000 107.6000 403.6000 107.7000 ;
	    RECT 407.6000 107.6000 408.4000 107.7000 ;
	    RECT 378.8000 106.6000 382.6000 107.2000 ;
	    RECT 372.4000 105.6000 374.2000 106.0000 ;
	    RECT 369.2000 103.0000 370.0000 105.0000 ;
	    RECT 373.4000 103.0000 374.2000 105.6000 ;
	    RECT 378.8000 102.2000 379.6000 106.6000 ;
	    RECT 381.8000 106.4000 382.6000 106.6000 ;
	    RECT 391.6000 105.6000 392.2000 107.6000 ;
	    RECT 389.8000 105.4000 390.6000 105.6000 ;
	    RECT 383.6000 104.2000 384.4000 105.0000 ;
	    RECT 387.8000 104.8000 390.6000 105.4000 ;
	    RECT 391.6000 104.8000 392.4000 105.6000 ;
	    RECT 387.8000 104.2000 388.4000 104.8000 ;
	    RECT 393.2000 104.2000 394.0000 105.0000 ;
	    RECT 383.0000 103.6000 384.4000 104.2000 ;
	    RECT 383.0000 102.2000 384.2000 103.6000 ;
	    RECT 387.6000 102.2000 388.4000 104.2000 ;
	    RECT 392.0000 103.6000 394.0000 104.2000 ;
	    RECT 392.0000 102.2000 392.8000 103.6000 ;
	    RECT 396.4000 102.2000 397.2000 107.0000 ;
	    RECT 398.2000 106.2000 398.8000 107.6000 ;
	    RECT 402.0000 107.2000 402.8000 107.6000 ;
	    RECT 410.8000 107.2000 411.6000 110.6000 ;
	    RECT 414.2000 110.4000 415.0000 110.6000 ;
	    RECT 412.6000 109.8000 413.4000 110.0000 ;
	    RECT 412.6000 109.2000 416.4000 109.8000 ;
	    RECT 415.6000 109.0000 416.4000 109.2000 ;
	    RECT 417.4000 108.4000 418.0000 111.6000 ;
	    RECT 419.4000 111.8000 420.0000 113.0000 ;
	    RECT 420.6000 113.0000 421.4000 113.2000 ;
	    RECT 425.2000 113.0000 426.0000 113.2000 ;
	    RECT 420.6000 112.4000 426.0000 113.0000 ;
	    RECT 419.4000 111.4000 424.2000 111.8000 ;
	    RECT 428.4000 111.4000 429.2000 119.8000 ;
	    RECT 419.4000 111.2000 429.2000 111.4000 ;
	    RECT 423.4000 111.0000 429.2000 111.2000 ;
	    RECT 423.6000 110.8000 429.2000 111.0000 ;
	    RECT 422.0000 110.2000 422.8000 110.4000 ;
	    RECT 422.0000 109.6000 427.0000 110.2000 ;
	    RECT 426.2000 109.4000 427.0000 109.6000 ;
	    RECT 424.6000 108.4000 425.4000 108.6000 ;
	    RECT 417.4000 107.8000 428.4000 108.4000 ;
	    RECT 417.8000 107.6000 418.6000 107.8000 ;
	    RECT 410.8000 106.6000 414.6000 107.2000 ;
	    RECT 399.8000 106.2000 403.4000 106.6000 ;
	    RECT 398.0000 102.2000 398.8000 106.2000 ;
	    RECT 399.6000 106.0000 403.6000 106.2000 ;
	    RECT 399.6000 102.2000 400.4000 106.0000 ;
	    RECT 402.8000 102.2000 403.6000 106.0000 ;
	    RECT 410.8000 102.2000 411.6000 106.6000 ;
	    RECT 413.8000 106.4000 414.6000 106.6000 ;
	    RECT 423.6000 106.4000 424.2000 107.8000 ;
	    RECT 426.8000 107.6000 428.4000 107.8000 ;
	    RECT 421.8000 105.4000 422.6000 105.6000 ;
	    RECT 415.6000 104.2000 416.4000 105.0000 ;
	    RECT 419.8000 104.8000 422.6000 105.4000 ;
	    RECT 423.6000 104.8000 424.4000 106.4000 ;
	    RECT 419.8000 104.2000 420.4000 104.8000 ;
	    RECT 425.2000 104.2000 426.0000 105.0000 ;
	    RECT 415.0000 103.6000 416.4000 104.2000 ;
	    RECT 415.0000 102.2000 416.2000 103.6000 ;
	    RECT 419.6000 102.2000 420.4000 104.2000 ;
	    RECT 424.0000 103.6000 426.0000 104.2000 ;
	    RECT 424.0000 102.2000 424.8000 103.6000 ;
	    RECT 428.4000 102.2000 429.2000 107.0000 ;
	    RECT 430.0000 106.8000 430.8000 108.4000 ;
	    RECT 431.6000 106.2000 432.4000 119.8000 ;
	    RECT 433.2000 111.6000 434.0000 113.2000 ;
	    RECT 434.8000 111.2000 435.6000 119.8000 ;
	    RECT 439.0000 115.8000 440.2000 119.8000 ;
	    RECT 443.6000 115.8000 444.4000 119.8000 ;
	    RECT 448.0000 116.4000 448.8000 119.8000 ;
	    RECT 448.0000 115.8000 450.0000 116.4000 ;
	    RECT 439.6000 115.0000 440.4000 115.8000 ;
	    RECT 443.8000 115.2000 444.4000 115.8000 ;
	    RECT 443.0000 114.6000 446.6000 115.2000 ;
	    RECT 449.2000 115.0000 450.0000 115.8000 ;
	    RECT 443.0000 114.4000 443.8000 114.6000 ;
	    RECT 445.8000 114.4000 446.6000 114.6000 ;
	    RECT 438.8000 113.2000 440.2000 114.0000 ;
	    RECT 439.6000 112.2000 440.2000 113.2000 ;
	    RECT 441.8000 113.0000 444.0000 113.6000 ;
	    RECT 441.8000 112.8000 442.6000 113.0000 ;
	    RECT 439.6000 111.6000 442.0000 112.2000 ;
	    RECT 434.8000 110.6000 439.0000 111.2000 ;
	    RECT 434.8000 107.2000 435.6000 110.6000 ;
	    RECT 438.2000 110.4000 439.0000 110.6000 ;
	    RECT 436.6000 109.8000 437.4000 110.0000 ;
	    RECT 436.6000 109.2000 440.4000 109.8000 ;
	    RECT 439.6000 109.0000 440.4000 109.2000 ;
	    RECT 441.4000 108.4000 442.0000 111.6000 ;
	    RECT 443.4000 111.8000 444.0000 113.0000 ;
	    RECT 444.6000 113.0000 445.4000 113.2000 ;
	    RECT 449.2000 113.0000 450.0000 113.2000 ;
	    RECT 444.6000 112.4000 450.0000 113.0000 ;
	    RECT 443.4000 111.4000 448.2000 111.8000 ;
	    RECT 452.4000 111.4000 453.2000 119.8000 ;
	    RECT 443.4000 111.2000 453.2000 111.4000 ;
	    RECT 447.4000 111.0000 453.2000 111.2000 ;
	    RECT 447.6000 110.8000 453.2000 111.0000 ;
	    RECT 446.0000 110.2000 446.8000 110.4000 ;
	    RECT 455.6000 110.3000 456.4000 119.8000 ;
	    RECT 459.6000 113.6000 460.4000 114.4000 ;
	    RECT 457.2000 111.6000 458.0000 113.2000 ;
	    RECT 459.6000 112.4000 460.2000 113.6000 ;
	    RECT 461.0000 112.4000 461.8000 119.8000 ;
	    RECT 458.8000 111.8000 460.2000 112.4000 ;
	    RECT 460.8000 111.8000 461.8000 112.4000 ;
	    RECT 458.8000 111.6000 459.6000 111.8000 ;
	    RECT 458.9000 110.3000 459.5000 111.6000 ;
	    RECT 446.0000 109.6000 451.0000 110.2000 ;
	    RECT 447.6000 109.4000 448.4000 109.6000 ;
	    RECT 450.2000 109.4000 451.0000 109.6000 ;
	    RECT 455.6000 109.7000 459.5000 110.3000 ;
	    RECT 448.6000 108.4000 449.4000 108.6000 ;
	    RECT 441.4000 107.8000 452.4000 108.4000 ;
	    RECT 441.8000 107.6000 442.6000 107.8000 ;
	    RECT 434.8000 106.6000 438.6000 107.2000 ;
	    RECT 431.6000 105.6000 433.4000 106.2000 ;
	    RECT 432.6000 104.4000 433.4000 105.6000 ;
	    RECT 432.6000 103.6000 434.0000 104.4000 ;
	    RECT 432.6000 102.2000 433.4000 103.6000 ;
	    RECT 434.8000 102.2000 435.6000 106.6000 ;
	    RECT 437.8000 106.4000 438.6000 106.6000 ;
	    RECT 447.6000 106.4000 448.2000 107.8000 ;
	    RECT 450.8000 107.6000 452.4000 107.8000 ;
	    RECT 445.8000 105.4000 446.6000 105.6000 ;
	    RECT 439.6000 104.2000 440.4000 105.0000 ;
	    RECT 443.8000 104.8000 446.6000 105.4000 ;
	    RECT 447.6000 104.8000 448.4000 106.4000 ;
	    RECT 443.8000 104.2000 444.4000 104.8000 ;
	    RECT 449.2000 104.2000 450.0000 105.0000 ;
	    RECT 439.0000 103.6000 440.4000 104.2000 ;
	    RECT 439.0000 102.2000 440.2000 103.6000 ;
	    RECT 443.6000 102.2000 444.4000 104.2000 ;
	    RECT 448.0000 103.6000 450.0000 104.2000 ;
	    RECT 448.0000 102.2000 448.8000 103.6000 ;
	    RECT 452.4000 102.2000 453.2000 107.0000 ;
	    RECT 454.0000 106.8000 454.8000 108.4000 ;
	    RECT 455.6000 106.2000 456.4000 109.7000 ;
	    RECT 460.8000 108.4000 461.4000 111.8000 ;
	    RECT 462.0000 108.8000 462.8000 110.4000 ;
	    RECT 457.2000 108.3000 458.0000 108.4000 ;
	    RECT 458.8000 108.3000 461.4000 108.4000 ;
	    RECT 457.2000 107.7000 461.4000 108.3000 ;
	    RECT 463.6000 108.2000 464.4000 108.4000 ;
	    RECT 457.2000 107.6000 458.0000 107.7000 ;
	    RECT 458.8000 107.6000 461.4000 107.7000 ;
	    RECT 462.8000 107.6000 464.4000 108.2000 ;
	    RECT 459.0000 106.2000 459.6000 107.6000 ;
	    RECT 462.8000 107.2000 463.6000 107.6000 ;
	    RECT 460.6000 106.2000 464.2000 106.6000 ;
	    RECT 455.6000 105.6000 457.4000 106.2000 ;
	    RECT 456.6000 102.2000 457.4000 105.6000 ;
	    RECT 458.8000 102.2000 459.6000 106.2000 ;
	    RECT 460.4000 106.0000 464.4000 106.2000 ;
	    RECT 460.4000 102.2000 461.2000 106.0000 ;
	    RECT 463.6000 102.2000 464.4000 106.0000 ;
	    RECT 465.2000 102.2000 466.0000 119.8000 ;
	    RECT 468.4000 102.2000 469.2000 119.8000 ;
	    RECT 471.6000 111.2000 472.4000 119.8000 ;
	    RECT 475.8000 115.8000 477.0000 119.8000 ;
	    RECT 480.4000 115.8000 481.2000 119.8000 ;
	    RECT 484.8000 116.4000 485.6000 119.8000 ;
	    RECT 484.8000 115.8000 486.8000 116.4000 ;
	    RECT 476.4000 115.0000 477.2000 115.8000 ;
	    RECT 480.6000 115.2000 481.2000 115.8000 ;
	    RECT 479.8000 114.6000 483.4000 115.2000 ;
	    RECT 486.0000 115.0000 486.8000 115.8000 ;
	    RECT 479.8000 114.4000 480.6000 114.6000 ;
	    RECT 482.6000 114.4000 483.4000 114.6000 ;
	    RECT 475.6000 113.2000 477.0000 114.0000 ;
	    RECT 476.4000 112.2000 477.0000 113.2000 ;
	    RECT 478.6000 113.0000 480.8000 113.6000 ;
	    RECT 478.6000 112.8000 479.4000 113.0000 ;
	    RECT 476.4000 111.6000 478.8000 112.2000 ;
	    RECT 471.6000 110.6000 475.8000 111.2000 ;
	    RECT 471.6000 107.2000 472.4000 110.6000 ;
	    RECT 475.0000 110.4000 475.8000 110.6000 ;
	    RECT 473.4000 109.8000 474.2000 110.0000 ;
	    RECT 473.4000 109.2000 477.2000 109.8000 ;
	    RECT 476.4000 109.0000 477.2000 109.2000 ;
	    RECT 478.2000 108.4000 478.8000 111.6000 ;
	    RECT 480.2000 111.8000 480.8000 113.0000 ;
	    RECT 481.4000 113.0000 482.2000 113.2000 ;
	    RECT 486.0000 113.0000 486.8000 113.2000 ;
	    RECT 481.4000 112.4000 486.8000 113.0000 ;
	    RECT 480.2000 111.4000 485.0000 111.8000 ;
	    RECT 489.2000 111.4000 490.0000 119.8000 ;
	    RECT 480.2000 111.2000 490.0000 111.4000 ;
	    RECT 484.2000 111.0000 490.0000 111.2000 ;
	    RECT 484.4000 110.8000 490.0000 111.0000 ;
	    RECT 482.8000 110.2000 483.6000 110.4000 ;
	    RECT 482.8000 109.6000 487.8000 110.2000 ;
	    RECT 484.4000 109.4000 485.2000 109.6000 ;
	    RECT 487.0000 109.4000 487.8000 109.6000 ;
	    RECT 485.4000 108.4000 486.2000 108.6000 ;
	    RECT 478.2000 107.8000 489.2000 108.4000 ;
	    RECT 478.6000 107.6000 479.4000 107.8000 ;
	    RECT 471.6000 106.6000 475.4000 107.2000 ;
	    RECT 471.6000 102.2000 472.4000 106.6000 ;
	    RECT 474.6000 106.4000 475.4000 106.6000 ;
	    RECT 484.4000 106.4000 485.0000 107.8000 ;
	    RECT 487.6000 107.6000 489.2000 107.8000 ;
	    RECT 492.4000 108.3000 493.2000 119.8000 ;
	    RECT 496.6000 112.4000 497.4000 119.8000 ;
	    RECT 502.0000 115.8000 502.8000 119.8000 ;
	    RECT 502.2000 115.6000 502.8000 115.8000 ;
	    RECT 505.2000 115.8000 506.0000 119.8000 ;
	    RECT 508.4000 115.8000 509.2000 119.8000 ;
	    RECT 505.2000 115.6000 505.8000 115.8000 ;
	    RECT 502.2000 115.0000 505.8000 115.6000 ;
	    RECT 508.6000 115.6000 509.2000 115.8000 ;
	    RECT 511.6000 115.8000 512.4000 119.8000 ;
	    RECT 511.6000 115.6000 512.2000 115.8000 ;
	    RECT 508.6000 115.0000 512.2000 115.6000 ;
	    RECT 498.0000 113.6000 498.8000 114.4000 ;
	    RECT 498.2000 112.4000 498.8000 113.6000 ;
	    RECT 503.6000 112.8000 504.4000 114.4000 ;
	    RECT 505.2000 112.4000 505.8000 115.0000 ;
	    RECT 510.0000 112.8000 510.8000 114.4000 ;
	    RECT 511.6000 112.4000 512.2000 115.0000 ;
	    RECT 495.6000 111.6000 497.6000 112.4000 ;
	    RECT 498.2000 111.8000 499.6000 112.4000 ;
	    RECT 498.8000 111.6000 499.6000 111.8000 ;
	    RECT 505.2000 111.6000 506.0000 112.4000 ;
	    RECT 511.6000 111.6000 512.4000 112.4000 ;
	    RECT 494.0000 110.3000 494.8000 110.4000 ;
	    RECT 495.6000 110.3000 496.4000 110.4000 ;
	    RECT 494.0000 109.7000 496.4000 110.3000 ;
	    RECT 494.0000 109.6000 494.8000 109.7000 ;
	    RECT 495.6000 108.8000 496.4000 109.7000 ;
	    RECT 497.0000 108.4000 497.6000 111.6000 ;
	    RECT 502.0000 109.6000 503.6000 110.4000 ;
	    RECT 505.2000 108.4000 505.8000 111.6000 ;
	    RECT 508.4000 109.6000 510.0000 110.4000 ;
	    RECT 511.6000 108.4000 512.2000 111.6000 ;
	    RECT 494.0000 108.3000 494.8000 108.4000 ;
	    RECT 492.4000 108.2000 494.8000 108.3000 ;
	    RECT 492.4000 107.7000 495.6000 108.2000 ;
	    RECT 482.6000 105.4000 483.4000 105.6000 ;
	    RECT 476.4000 104.2000 477.2000 105.0000 ;
	    RECT 480.6000 104.8000 483.4000 105.4000 ;
	    RECT 484.4000 104.8000 485.2000 106.4000 ;
	    RECT 480.6000 104.2000 481.2000 104.8000 ;
	    RECT 486.0000 104.2000 486.8000 105.0000 ;
	    RECT 475.8000 103.6000 477.2000 104.2000 ;
	    RECT 475.8000 102.2000 477.0000 103.6000 ;
	    RECT 480.4000 102.2000 481.2000 104.2000 ;
	    RECT 484.8000 103.6000 486.8000 104.2000 ;
	    RECT 484.8000 102.2000 485.6000 103.6000 ;
	    RECT 489.2000 102.2000 490.0000 107.0000 ;
	    RECT 490.8000 104.8000 491.6000 106.4000 ;
	    RECT 492.4000 102.2000 493.2000 107.7000 ;
	    RECT 494.0000 107.6000 495.6000 107.7000 ;
	    RECT 497.0000 107.6000 499.6000 108.4000 ;
	    RECT 504.2000 108.2000 505.8000 108.4000 ;
	    RECT 510.6000 108.2000 512.2000 108.4000 ;
	    RECT 504.0000 107.8000 505.8000 108.2000 ;
	    RECT 510.4000 107.8000 512.2000 108.2000 ;
	    RECT 494.8000 107.2000 495.6000 107.6000 ;
	    RECT 494.2000 106.2000 497.8000 106.6000 ;
	    RECT 498.8000 106.2000 499.4000 107.6000 ;
	    RECT 494.0000 106.0000 498.0000 106.2000 ;
	    RECT 494.0000 102.2000 494.8000 106.0000 ;
	    RECT 497.2000 102.2000 498.0000 106.0000 ;
	    RECT 498.8000 102.2000 499.6000 106.2000 ;
	    RECT 504.0000 102.2000 504.8000 107.8000 ;
	    RECT 510.4000 102.2000 511.2000 107.8000 ;
	    RECT 4.4000 95.2000 5.2000 99.8000 ;
	    RECT 9.2000 95.2000 10.0000 99.8000 ;
	    RECT 10.8000 95.8000 11.6000 99.8000 ;
	    RECT 12.4000 96.0000 13.2000 99.8000 ;
	    RECT 15.6000 96.0000 16.4000 99.8000 ;
	    RECT 12.4000 95.8000 16.4000 96.0000 ;
	    RECT 17.2000 95.8000 18.0000 99.8000 ;
	    RECT 18.8000 96.0000 19.6000 99.8000 ;
	    RECT 22.0000 96.0000 22.8000 99.8000 ;
	    RECT 18.8000 95.8000 22.8000 96.0000 ;
	    RECT 23.6000 96.0000 24.4000 99.8000 ;
	    RECT 26.8000 96.0000 27.6000 99.8000 ;
	    RECT 23.6000 95.8000 27.6000 96.0000 ;
	    RECT 28.4000 95.8000 29.2000 99.8000 ;
	    RECT 3.0000 94.6000 5.2000 95.2000 ;
	    RECT 7.8000 94.6000 10.0000 95.2000 ;
	    RECT 3.0000 91.6000 3.6000 94.6000 ;
	    RECT 4.4000 91.6000 5.2000 93.2000 ;
	    RECT 7.8000 91.6000 8.4000 94.6000 ;
	    RECT 11.0000 94.4000 11.6000 95.8000 ;
	    RECT 12.6000 95.4000 16.2000 95.8000 ;
	    RECT 14.8000 94.4000 15.6000 94.8000 ;
	    RECT 17.4000 94.4000 18.0000 95.8000 ;
	    RECT 19.0000 95.4000 22.6000 95.8000 ;
	    RECT 23.8000 95.4000 27.4000 95.8000 ;
	    RECT 21.2000 94.4000 22.0000 94.8000 ;
	    RECT 24.4000 94.4000 25.2000 94.8000 ;
	    RECT 28.4000 94.4000 29.0000 95.8000 ;
	    RECT 30.0000 95.4000 30.8000 99.8000 ;
	    RECT 34.2000 98.4000 35.4000 99.8000 ;
	    RECT 34.2000 97.8000 35.6000 98.4000 ;
	    RECT 38.8000 97.8000 39.6000 99.8000 ;
	    RECT 43.2000 98.4000 44.0000 99.8000 ;
	    RECT 43.2000 97.8000 45.2000 98.4000 ;
	    RECT 34.8000 97.0000 35.6000 97.8000 ;
	    RECT 39.0000 97.2000 39.6000 97.8000 ;
	    RECT 39.0000 96.6000 41.8000 97.2000 ;
	    RECT 41.0000 96.4000 41.8000 96.6000 ;
	    RECT 42.8000 96.4000 43.6000 97.2000 ;
	    RECT 44.4000 97.0000 45.2000 97.8000 ;
	    RECT 33.0000 95.4000 33.8000 95.6000 ;
	    RECT 30.0000 94.8000 33.8000 95.4000 ;
	    RECT 10.8000 93.6000 13.4000 94.4000 ;
	    RECT 14.8000 93.8000 16.4000 94.4000 ;
	    RECT 15.6000 93.6000 16.4000 93.8000 ;
	    RECT 17.2000 93.6000 19.8000 94.4000 ;
	    RECT 21.2000 93.8000 22.8000 94.4000 ;
	    RECT 22.0000 93.6000 22.8000 93.8000 ;
	    RECT 23.6000 93.8000 25.2000 94.4000 ;
	    RECT 23.6000 93.6000 24.4000 93.8000 ;
	    RECT 26.6000 93.6000 29.2000 94.4000 ;
	    RECT 9.2000 91.6000 10.0000 93.2000 ;
	    RECT 2.4000 90.8000 3.6000 91.6000 ;
	    RECT 7.2000 90.8000 8.4000 91.6000 ;
	    RECT 3.0000 90.2000 3.6000 90.8000 ;
	    RECT 7.8000 90.2000 8.4000 90.8000 ;
	    RECT 10.8000 90.2000 11.6000 90.4000 ;
	    RECT 12.8000 90.2000 13.4000 93.6000 ;
	    RECT 14.0000 91.6000 14.8000 93.2000 ;
	    RECT 17.2000 90.2000 18.0000 90.4000 ;
	    RECT 19.2000 90.2000 19.8000 93.6000 ;
	    RECT 20.4000 92.3000 21.2000 93.2000 ;
	    RECT 22.0000 92.3000 22.8000 92.4000 ;
	    RECT 20.4000 91.7000 22.8000 92.3000 ;
	    RECT 20.4000 91.6000 21.2000 91.7000 ;
	    RECT 22.0000 91.6000 22.8000 91.7000 ;
	    RECT 25.2000 91.6000 26.0000 93.2000 ;
	    RECT 26.6000 92.3000 27.2000 93.6000 ;
	    RECT 28.4000 92.3000 29.2000 92.4000 ;
	    RECT 26.6000 91.7000 29.2000 92.3000 ;
	    RECT 26.6000 90.2000 27.2000 91.7000 ;
	    RECT 28.4000 91.6000 29.2000 91.7000 ;
	    RECT 30.0000 91.4000 30.8000 94.8000 ;
	    RECT 37.0000 94.2000 37.8000 94.4000 ;
	    RECT 42.8000 94.2000 43.4000 96.4000 ;
	    RECT 47.6000 95.0000 48.4000 99.8000 ;
	    RECT 49.2000 95.8000 50.0000 99.8000 ;
	    RECT 50.8000 96.0000 51.6000 99.8000 ;
	    RECT 54.0000 96.0000 54.8000 99.8000 ;
	    RECT 57.2000 97.8000 58.0000 99.8000 ;
	    RECT 62.0000 97.8000 62.8000 99.8000 ;
	    RECT 66.8000 97.8000 67.6000 99.8000 ;
	    RECT 71.6000 97.8000 72.4000 99.8000 ;
	    RECT 50.8000 95.8000 54.8000 96.0000 ;
	    RECT 49.4000 94.4000 50.0000 95.8000 ;
	    RECT 51.0000 95.4000 54.6000 95.8000 ;
	    RECT 55.6000 95.6000 56.4000 97.2000 ;
	    RECT 53.2000 94.4000 54.0000 94.8000 ;
	    RECT 57.4000 94.4000 58.0000 97.8000 ;
	    RECT 60.4000 95.6000 61.2000 97.2000 ;
	    RECT 62.2000 94.4000 62.8000 97.8000 ;
	    RECT 65.2000 95.6000 66.0000 97.2000 ;
	    RECT 67.0000 94.4000 67.6000 97.8000 ;
	    RECT 70.0000 95.6000 70.8000 97.2000 ;
	    RECT 71.8000 94.4000 72.4000 97.8000 ;
	    RECT 74.8000 95.8000 75.6000 99.8000 ;
	    RECT 76.4000 96.0000 77.2000 99.8000 ;
	    RECT 79.6000 96.0000 80.4000 99.8000 ;
	    RECT 76.4000 95.8000 80.4000 96.0000 ;
	    RECT 75.0000 94.4000 75.6000 95.8000 ;
	    RECT 76.6000 95.4000 80.2000 95.8000 ;
	    RECT 81.2000 95.0000 82.0000 99.8000 ;
	    RECT 85.6000 98.4000 86.4000 99.8000 ;
	    RECT 84.4000 97.8000 86.4000 98.4000 ;
	    RECT 90.0000 97.8000 90.8000 99.8000 ;
	    RECT 94.2000 98.4000 95.4000 99.8000 ;
	    RECT 94.0000 97.8000 95.4000 98.4000 ;
	    RECT 84.4000 97.0000 85.2000 97.8000 ;
	    RECT 90.0000 97.2000 90.6000 97.8000 ;
	    RECT 86.0000 96.4000 86.8000 97.2000 ;
	    RECT 87.8000 96.6000 90.6000 97.2000 ;
	    RECT 94.0000 97.0000 94.8000 97.8000 ;
	    RECT 87.8000 96.4000 88.6000 96.6000 ;
	    RECT 78.8000 94.4000 79.6000 94.8000 ;
	    RECT 46.0000 94.2000 47.6000 94.4000 ;
	    RECT 36.6000 93.6000 47.6000 94.2000 ;
	    RECT 49.2000 93.6000 51.8000 94.4000 ;
	    RECT 53.2000 94.3000 54.8000 94.4000 ;
	    RECT 57.2000 94.3000 58.0000 94.4000 ;
	    RECT 53.2000 93.8000 58.0000 94.3000 ;
	    RECT 54.0000 93.7000 58.0000 93.8000 ;
	    RECT 54.0000 93.6000 54.8000 93.7000 ;
	    RECT 57.2000 93.6000 58.0000 93.7000 ;
	    RECT 62.0000 93.6000 62.8000 94.4000 ;
	    RECT 63.6000 94.3000 64.4000 94.4000 ;
	    RECT 66.8000 94.3000 67.6000 94.4000 ;
	    RECT 63.6000 93.7000 67.6000 94.3000 ;
	    RECT 63.6000 93.6000 64.4000 93.7000 ;
	    RECT 66.8000 93.6000 67.6000 93.7000 ;
	    RECT 71.6000 93.6000 72.4000 94.4000 ;
	    RECT 73.2000 94.3000 74.0000 94.4000 ;
	    RECT 74.8000 94.3000 77.4000 94.4000 ;
	    RECT 73.2000 93.7000 77.4000 94.3000 ;
	    RECT 78.8000 93.8000 80.4000 94.4000 ;
	    RECT 73.2000 93.6000 74.0000 93.7000 ;
	    RECT 74.8000 93.6000 77.4000 93.7000 ;
	    RECT 79.6000 93.6000 80.4000 93.8000 ;
	    RECT 82.0000 94.2000 83.6000 94.4000 ;
	    RECT 86.2000 94.2000 86.8000 96.4000 ;
	    RECT 95.8000 95.4000 96.6000 95.6000 ;
	    RECT 98.8000 95.4000 99.6000 99.8000 ;
	    RECT 100.4000 96.0000 101.2000 99.8000 ;
	    RECT 103.6000 96.0000 104.4000 99.8000 ;
	    RECT 100.4000 95.8000 104.4000 96.0000 ;
	    RECT 105.2000 95.8000 106.0000 99.8000 ;
	    RECT 113.2000 95.8000 114.0000 99.8000 ;
	    RECT 114.8000 96.0000 115.6000 99.8000 ;
	    RECT 118.0000 96.0000 118.8000 99.8000 ;
	    RECT 114.8000 95.8000 118.8000 96.0000 ;
	    RECT 119.6000 95.8000 120.4000 99.8000 ;
	    RECT 121.2000 96.0000 122.0000 99.8000 ;
	    RECT 124.4000 96.0000 125.2000 99.8000 ;
	    RECT 121.2000 95.8000 125.2000 96.0000 ;
	    RECT 126.0000 95.8000 126.8000 99.8000 ;
	    RECT 127.6000 96.0000 128.4000 99.8000 ;
	    RECT 130.8000 96.0000 131.6000 99.8000 ;
	    RECT 134.0000 97.8000 134.8000 99.8000 ;
	    RECT 127.6000 95.8000 131.6000 96.0000 ;
	    RECT 100.6000 95.4000 104.2000 95.8000 ;
	    RECT 95.8000 94.8000 99.6000 95.4000 ;
	    RECT 87.6000 94.2000 88.4000 94.4000 ;
	    RECT 91.8000 94.2000 92.6000 94.4000 ;
	    RECT 82.0000 93.6000 93.0000 94.2000 ;
	    RECT 34.8000 92.8000 35.6000 93.0000 ;
	    RECT 31.8000 92.2000 35.6000 92.8000 ;
	    RECT 36.6000 92.4000 37.2000 93.6000 ;
	    RECT 43.8000 93.4000 44.6000 93.6000 ;
	    RECT 42.8000 92.4000 43.6000 92.6000 ;
	    RECT 45.4000 92.4000 46.2000 92.6000 ;
	    RECT 31.8000 92.0000 32.6000 92.2000 ;
	    RECT 36.4000 91.6000 37.2000 92.4000 ;
	    RECT 41.2000 91.8000 46.2000 92.4000 ;
	    RECT 41.2000 91.6000 42.0000 91.8000 ;
	    RECT 33.4000 91.4000 34.2000 91.6000 ;
	    RECT 30.0000 90.8000 34.2000 91.4000 ;
	    RECT 28.4000 90.2000 29.2000 90.4000 ;
	    RECT 3.0000 89.6000 5.2000 90.2000 ;
	    RECT 7.8000 89.6000 10.0000 90.2000 ;
	    RECT 10.8000 89.6000 12.2000 90.2000 ;
	    RECT 12.8000 89.6000 13.8000 90.2000 ;
	    RECT 17.2000 89.6000 18.6000 90.2000 ;
	    RECT 19.2000 89.6000 20.2000 90.2000 ;
	    RECT 4.4000 82.2000 5.2000 89.6000 ;
	    RECT 9.2000 82.2000 10.0000 89.6000 ;
	    RECT 11.6000 88.4000 12.2000 89.6000 ;
	    RECT 13.0000 88.4000 13.8000 89.6000 ;
	    RECT 18.0000 88.4000 18.6000 89.6000 ;
	    RECT 11.6000 87.6000 12.4000 88.4000 ;
	    RECT 13.0000 87.6000 14.8000 88.4000 ;
	    RECT 18.0000 87.6000 18.8000 88.4000 ;
	    RECT 13.0000 82.2000 13.8000 87.6000 ;
	    RECT 19.4000 82.2000 20.2000 89.6000 ;
	    RECT 26.2000 89.6000 27.2000 90.2000 ;
	    RECT 27.8000 89.6000 29.2000 90.2000 ;
	    RECT 26.2000 82.2000 27.0000 89.6000 ;
	    RECT 27.8000 88.4000 28.4000 89.6000 ;
	    RECT 27.6000 88.3000 28.4000 88.4000 ;
	    RECT 30.0000 88.3000 30.8000 90.8000 ;
	    RECT 36.6000 90.4000 37.2000 91.6000 ;
	    RECT 42.8000 91.0000 48.4000 91.2000 ;
	    RECT 42.6000 90.8000 48.4000 91.0000 ;
	    RECT 34.8000 89.8000 37.2000 90.4000 ;
	    RECT 38.6000 90.6000 48.4000 90.8000 ;
	    RECT 38.6000 90.2000 43.4000 90.6000 ;
	    RECT 34.8000 88.8000 35.4000 89.8000 ;
	    RECT 27.6000 87.7000 30.8000 88.3000 ;
	    RECT 34.0000 88.0000 35.4000 88.8000 ;
	    RECT 37.0000 89.0000 37.8000 89.2000 ;
	    RECT 38.6000 89.0000 39.2000 90.2000 ;
	    RECT 37.0000 88.4000 39.2000 89.0000 ;
	    RECT 39.8000 89.0000 45.2000 89.6000 ;
	    RECT 39.8000 88.8000 40.6000 89.0000 ;
	    RECT 44.4000 88.8000 45.2000 89.0000 ;
	    RECT 27.6000 87.6000 28.4000 87.7000 ;
	    RECT 30.0000 82.2000 30.8000 87.7000 ;
	    RECT 38.2000 87.4000 39.0000 87.6000 ;
	    RECT 41.0000 87.4000 41.8000 87.6000 ;
	    RECT 34.8000 86.2000 35.6000 87.0000 ;
	    RECT 38.2000 86.8000 41.8000 87.4000 ;
	    RECT 39.0000 86.2000 39.6000 86.8000 ;
	    RECT 44.4000 86.2000 45.2000 87.0000 ;
	    RECT 34.2000 82.2000 35.4000 86.2000 ;
	    RECT 38.8000 82.2000 39.6000 86.2000 ;
	    RECT 43.2000 85.6000 45.2000 86.2000 ;
	    RECT 43.2000 82.2000 44.0000 85.6000 ;
	    RECT 47.6000 82.2000 48.4000 90.6000 ;
	    RECT 49.2000 90.2000 50.0000 90.4000 ;
	    RECT 51.2000 90.2000 51.8000 93.6000 ;
	    RECT 52.4000 91.6000 53.2000 93.2000 ;
	    RECT 57.4000 90.2000 58.0000 93.6000 ;
	    RECT 58.8000 90.8000 59.6000 92.4000 ;
	    RECT 62.2000 90.2000 62.8000 93.6000 ;
	    RECT 63.6000 90.8000 64.4000 92.4000 ;
	    RECT 67.0000 90.2000 67.6000 93.6000 ;
	    RECT 68.4000 90.8000 69.2000 92.4000 ;
	    RECT 71.8000 90.2000 72.4000 93.6000 ;
	    RECT 73.2000 90.8000 74.0000 92.4000 ;
	    RECT 74.8000 90.2000 75.6000 90.4000 ;
	    RECT 76.8000 90.2000 77.4000 93.6000 ;
	    RECT 85.0000 93.4000 85.8000 93.6000 ;
	    RECT 78.0000 91.6000 78.8000 93.2000 ;
	    RECT 83.4000 92.4000 84.2000 92.6000 ;
	    RECT 83.4000 92.3000 88.4000 92.4000 ;
	    RECT 89.2000 92.3000 90.0000 92.4000 ;
	    RECT 83.4000 91.8000 90.0000 92.3000 ;
	    RECT 87.6000 91.7000 90.0000 91.8000 ;
	    RECT 87.6000 91.6000 88.4000 91.7000 ;
	    RECT 89.2000 91.6000 90.0000 91.7000 ;
	    RECT 81.2000 91.0000 86.8000 91.2000 ;
	    RECT 81.2000 90.8000 87.0000 91.0000 ;
	    RECT 81.2000 90.6000 91.0000 90.8000 ;
	    RECT 49.2000 89.6000 50.6000 90.2000 ;
	    RECT 51.2000 89.6000 52.2000 90.2000 ;
	    RECT 50.0000 88.4000 50.6000 89.6000 ;
	    RECT 50.0000 87.6000 50.8000 88.4000 ;
	    RECT 51.4000 82.2000 52.2000 89.6000 ;
	    RECT 57.2000 89.4000 59.0000 90.2000 ;
	    RECT 62.0000 89.4000 63.8000 90.2000 ;
	    RECT 66.8000 89.4000 68.6000 90.2000 ;
	    RECT 71.6000 89.4000 73.4000 90.2000 ;
	    RECT 74.8000 89.6000 76.2000 90.2000 ;
	    RECT 76.8000 89.6000 77.8000 90.2000 ;
	    RECT 58.2000 82.2000 59.0000 89.4000 ;
	    RECT 63.0000 84.4000 63.8000 89.4000 ;
	    RECT 62.0000 83.6000 63.8000 84.4000 ;
	    RECT 63.0000 82.2000 63.8000 83.6000 ;
	    RECT 67.8000 82.2000 68.6000 89.4000 ;
	    RECT 72.6000 84.4000 73.4000 89.4000 ;
	    RECT 75.6000 88.4000 76.2000 89.6000 ;
	    RECT 75.6000 87.6000 76.4000 88.4000 ;
	    RECT 71.6000 83.6000 73.4000 84.4000 ;
	    RECT 72.6000 82.2000 73.4000 83.6000 ;
	    RECT 77.0000 82.2000 77.8000 89.6000 ;
	    RECT 81.2000 82.2000 82.0000 90.6000 ;
	    RECT 86.2000 90.2000 91.0000 90.6000 ;
	    RECT 84.4000 89.0000 89.8000 89.6000 ;
	    RECT 84.4000 88.8000 85.2000 89.0000 ;
	    RECT 89.0000 88.8000 89.8000 89.0000 ;
	    RECT 90.4000 89.0000 91.0000 90.2000 ;
	    RECT 92.4000 90.4000 93.0000 93.6000 ;
	    RECT 94.0000 92.8000 94.8000 93.0000 ;
	    RECT 94.0000 92.2000 97.8000 92.8000 ;
	    RECT 97.0000 92.0000 97.8000 92.2000 ;
	    RECT 95.4000 91.4000 96.2000 91.6000 ;
	    RECT 98.8000 91.4000 99.6000 94.8000 ;
	    RECT 101.2000 94.4000 102.0000 94.8000 ;
	    RECT 105.2000 94.4000 105.8000 95.8000 ;
	    RECT 113.4000 94.4000 114.0000 95.8000 ;
	    RECT 115.0000 95.4000 118.6000 95.8000 ;
	    RECT 117.2000 94.4000 118.0000 94.8000 ;
	    RECT 119.8000 94.4000 120.4000 95.8000 ;
	    RECT 121.4000 95.4000 125.0000 95.8000 ;
	    RECT 123.6000 94.4000 124.4000 94.8000 ;
	    RECT 126.2000 94.4000 126.8000 95.8000 ;
	    RECT 127.8000 95.4000 131.4000 95.8000 ;
	    RECT 132.4000 95.6000 133.2000 97.2000 ;
	    RECT 130.0000 94.4000 130.8000 94.8000 ;
	    RECT 134.2000 94.4000 134.8000 97.8000 ;
	    RECT 137.2000 99.2000 141.2000 99.8000 ;
	    RECT 137.2000 95.8000 138.0000 99.2000 ;
	    RECT 138.8000 95.6000 139.6000 98.6000 ;
	    RECT 140.4000 96.0000 141.2000 99.2000 ;
	    RECT 143.6000 96.0000 144.4000 99.8000 ;
	    RECT 140.4000 95.8000 144.4000 96.0000 ;
	    RECT 145.2000 95.8000 146.0000 99.8000 ;
	    RECT 146.8000 96.0000 147.6000 99.8000 ;
	    RECT 150.0000 96.0000 150.8000 99.8000 ;
	    RECT 146.8000 95.8000 150.8000 96.0000 ;
	    RECT 151.6000 99.2000 155.6000 99.8000 ;
	    RECT 151.6000 95.8000 152.4000 99.2000 ;
	    RECT 153.2000 95.8000 154.0000 98.6000 ;
	    RECT 154.8000 96.0000 155.6000 99.2000 ;
	    RECT 158.0000 96.0000 158.8000 99.8000 ;
	    RECT 154.8000 95.8000 158.8000 96.0000 ;
	    RECT 159.6000 95.8000 160.4000 99.8000 ;
	    RECT 161.2000 96.0000 162.0000 99.8000 ;
	    RECT 164.4000 96.0000 165.2000 99.8000 ;
	    RECT 167.6000 97.8000 168.4000 99.8000 ;
	    RECT 161.2000 95.8000 165.2000 96.0000 ;
	    RECT 138.8000 94.4000 139.4000 95.6000 ;
	    RECT 140.6000 95.4000 144.2000 95.8000 ;
	    RECT 142.8000 94.4000 143.6000 94.8000 ;
	    RECT 145.4000 94.4000 146.0000 95.8000 ;
	    RECT 147.0000 95.4000 150.6000 95.8000 ;
	    RECT 149.2000 94.4000 150.0000 94.8000 ;
	    RECT 153.2000 94.4000 153.8000 95.8000 ;
	    RECT 155.0000 95.4000 158.6000 95.8000 ;
	    RECT 157.2000 94.4000 158.0000 94.8000 ;
	    RECT 159.8000 94.4000 160.4000 95.8000 ;
	    RECT 161.4000 95.4000 165.0000 95.8000 ;
	    RECT 166.0000 95.6000 166.8000 97.2000 ;
	    RECT 163.6000 94.4000 164.4000 94.8000 ;
	    RECT 167.8000 94.4000 168.4000 97.8000 ;
	    RECT 170.8000 95.8000 171.6000 99.8000 ;
	    RECT 172.4000 96.0000 173.2000 99.8000 ;
	    RECT 175.6000 96.0000 176.4000 99.8000 ;
	    RECT 172.4000 95.8000 176.4000 96.0000 ;
	    RECT 177.2000 96.0000 178.0000 99.8000 ;
	    RECT 180.4000 99.2000 184.4000 99.8000 ;
	    RECT 180.4000 96.0000 181.2000 99.2000 ;
	    RECT 177.2000 95.8000 181.2000 96.0000 ;
	    RECT 182.0000 95.8000 182.8000 98.6000 ;
	    RECT 183.6000 95.8000 184.4000 99.2000 ;
	    RECT 185.2000 99.2000 189.2000 99.8000 ;
	    RECT 185.2000 95.8000 186.0000 99.2000 ;
	    RECT 186.8000 95.8000 187.6000 98.6000 ;
	    RECT 188.4000 96.0000 189.2000 99.2000 ;
	    RECT 191.6000 96.0000 192.4000 99.8000 ;
	    RECT 188.4000 95.8000 192.4000 96.0000 ;
	    RECT 193.2000 95.8000 194.0000 99.8000 ;
	    RECT 194.8000 96.0000 195.6000 99.8000 ;
	    RECT 198.0000 96.0000 198.8000 99.8000 ;
	    RECT 194.8000 95.8000 198.8000 96.0000 ;
	    RECT 199.6000 95.8000 200.4000 99.8000 ;
	    RECT 201.2000 96.0000 202.0000 99.8000 ;
	    RECT 204.4000 96.0000 205.2000 99.8000 ;
	    RECT 201.2000 95.8000 205.2000 96.0000 ;
	    RECT 206.0000 97.0000 206.8000 99.0000 ;
	    RECT 171.0000 94.4000 171.6000 95.8000 ;
	    RECT 172.6000 95.4000 176.2000 95.8000 ;
	    RECT 177.4000 95.4000 181.0000 95.8000 ;
	    RECT 174.8000 94.4000 175.6000 94.8000 ;
	    RECT 178.0000 94.4000 178.8000 94.8000 ;
	    RECT 182.2000 94.4000 182.8000 95.8000 ;
	    RECT 186.8000 94.4000 187.4000 95.8000 ;
	    RECT 188.6000 95.4000 192.2000 95.8000 ;
	    RECT 190.8000 94.4000 191.6000 94.8000 ;
	    RECT 193.4000 94.4000 194.0000 95.8000 ;
	    RECT 195.0000 95.4000 198.6000 95.8000 ;
	    RECT 197.2000 94.4000 198.0000 94.8000 ;
	    RECT 199.8000 94.4000 200.4000 95.8000 ;
	    RECT 201.4000 95.4000 205.0000 95.8000 ;
	    RECT 206.0000 94.8000 206.6000 97.0000 ;
	    RECT 210.2000 96.4000 211.0000 99.0000 ;
	    RECT 209.2000 96.0000 211.0000 96.4000 ;
	    RECT 219.4000 96.0000 220.2000 99.0000 ;
	    RECT 223.6000 97.0000 224.4000 99.0000 ;
	    RECT 226.8000 97.8000 227.6000 99.8000 ;
	    RECT 209.2000 95.6000 211.8000 96.0000 ;
	    RECT 210.2000 95.4000 211.8000 95.6000 ;
	    RECT 211.0000 95.0000 211.8000 95.4000 ;
	    RECT 203.6000 94.4000 204.4000 94.8000 ;
	    RECT 100.4000 93.8000 102.0000 94.4000 ;
	    RECT 100.4000 93.6000 101.2000 93.8000 ;
	    RECT 103.4000 93.6000 106.0000 94.4000 ;
	    RECT 113.2000 93.6000 115.8000 94.4000 ;
	    RECT 117.2000 93.8000 118.8000 94.4000 ;
	    RECT 118.0000 93.6000 118.8000 93.8000 ;
	    RECT 119.6000 93.6000 122.2000 94.4000 ;
	    RECT 123.6000 93.8000 125.2000 94.4000 ;
	    RECT 124.4000 93.6000 125.2000 93.8000 ;
	    RECT 126.0000 93.6000 128.6000 94.4000 ;
	    RECT 130.0000 94.3000 131.6000 94.4000 ;
	    RECT 132.4000 94.3000 133.2000 94.4000 ;
	    RECT 130.0000 93.8000 133.2000 94.3000 ;
	    RECT 130.8000 93.7000 133.2000 93.8000 ;
	    RECT 130.8000 93.6000 131.6000 93.7000 ;
	    RECT 132.4000 93.6000 133.2000 93.7000 ;
	    RECT 134.0000 93.6000 134.8000 94.4000 ;
	    RECT 102.0000 91.6000 102.8000 93.2000 ;
	    RECT 95.4000 90.8000 99.6000 91.4000 ;
	    RECT 92.4000 89.8000 94.8000 90.4000 ;
	    RECT 91.8000 89.0000 92.6000 89.2000 ;
	    RECT 90.4000 88.4000 92.6000 89.0000 ;
	    RECT 94.2000 88.8000 94.8000 89.8000 ;
	    RECT 94.2000 88.0000 95.6000 88.8000 ;
	    RECT 87.8000 87.4000 88.6000 87.6000 ;
	    RECT 90.6000 87.4000 91.4000 87.6000 ;
	    RECT 84.4000 86.2000 85.2000 87.0000 ;
	    RECT 87.8000 86.8000 91.4000 87.4000 ;
	    RECT 90.0000 86.2000 90.6000 86.8000 ;
	    RECT 94.0000 86.2000 94.8000 87.0000 ;
	    RECT 84.4000 85.6000 86.4000 86.2000 ;
	    RECT 85.6000 82.2000 86.4000 85.6000 ;
	    RECT 90.0000 82.2000 90.8000 86.2000 ;
	    RECT 94.2000 82.2000 95.4000 86.2000 ;
	    RECT 98.8000 82.2000 99.6000 90.8000 ;
	    RECT 103.4000 90.2000 104.0000 93.6000 ;
	    RECT 115.2000 92.3000 115.8000 93.6000 ;
	    RECT 105.3000 91.7000 115.8000 92.3000 ;
	    RECT 105.3000 90.4000 105.9000 91.7000 ;
	    RECT 105.2000 90.2000 106.0000 90.4000 ;
	    RECT 103.0000 89.6000 104.0000 90.2000 ;
	    RECT 104.6000 89.6000 106.0000 90.2000 ;
	    RECT 111.6000 90.3000 112.4000 90.4000 ;
	    RECT 113.2000 90.3000 114.0000 90.4000 ;
	    RECT 111.6000 90.2000 114.0000 90.3000 ;
	    RECT 115.2000 90.2000 115.8000 91.7000 ;
	    RECT 116.4000 91.6000 117.2000 93.2000 ;
	    RECT 119.6000 90.2000 120.4000 90.4000 ;
	    RECT 121.6000 90.2000 122.2000 93.6000 ;
	    RECT 122.8000 92.3000 123.6000 93.2000 ;
	    RECT 128.0000 92.3000 128.6000 93.6000 ;
	    RECT 122.8000 91.7000 128.6000 92.3000 ;
	    RECT 122.8000 91.6000 123.6000 91.7000 ;
	    RECT 126.0000 90.2000 126.8000 90.4000 ;
	    RECT 128.0000 90.2000 128.6000 91.7000 ;
	    RECT 129.2000 91.6000 130.0000 93.2000 ;
	    RECT 134.2000 90.2000 134.8000 93.6000 ;
	    RECT 137.2000 92.8000 138.0000 94.4000 ;
	    RECT 138.8000 93.8000 141.2000 94.4000 ;
	    RECT 142.8000 94.3000 144.4000 94.4000 ;
	    RECT 145.2000 94.3000 147.8000 94.4000 ;
	    RECT 142.8000 93.8000 147.8000 94.3000 ;
	    RECT 149.2000 93.8000 150.8000 94.4000 ;
	    RECT 140.4000 93.6000 141.2000 93.8000 ;
	    RECT 143.6000 93.7000 147.8000 93.8000 ;
	    RECT 143.6000 93.6000 144.4000 93.7000 ;
	    RECT 145.2000 93.6000 147.8000 93.7000 ;
	    RECT 150.0000 93.6000 150.8000 93.8000 ;
	    RECT 135.6000 90.8000 136.4000 92.4000 ;
	    RECT 138.8000 91.6000 139.6000 93.2000 ;
	    RECT 140.6000 90.2000 141.2000 93.6000 ;
	    RECT 142.0000 91.6000 142.8000 93.2000 ;
	    RECT 145.2000 90.2000 146.0000 90.4000 ;
	    RECT 147.2000 90.2000 147.8000 93.6000 ;
	    RECT 148.4000 91.6000 149.2000 93.2000 ;
	    RECT 151.6000 92.8000 152.4000 94.4000 ;
	    RECT 153.2000 93.8000 155.6000 94.4000 ;
	    RECT 157.2000 94.3000 158.8000 94.4000 ;
	    RECT 159.6000 94.3000 162.2000 94.4000 ;
	    RECT 157.2000 93.8000 162.2000 94.3000 ;
	    RECT 163.6000 93.8000 165.2000 94.4000 ;
	    RECT 154.8000 93.6000 155.6000 93.8000 ;
	    RECT 158.0000 93.7000 162.2000 93.8000 ;
	    RECT 158.0000 93.6000 158.8000 93.7000 ;
	    RECT 159.6000 93.6000 162.2000 93.7000 ;
	    RECT 164.4000 93.6000 165.2000 93.8000 ;
	    RECT 167.6000 93.6000 168.4000 94.4000 ;
	    RECT 170.8000 93.6000 173.4000 94.4000 ;
	    RECT 174.8000 93.8000 176.4000 94.4000 ;
	    RECT 175.6000 93.6000 176.4000 93.8000 ;
	    RECT 177.2000 93.8000 178.8000 94.4000 ;
	    RECT 180.4000 93.8000 182.8000 94.4000 ;
	    RECT 177.2000 93.6000 178.0000 93.8000 ;
	    RECT 180.4000 93.6000 181.2000 93.8000 ;
	    RECT 153.2000 91.6000 154.0000 93.2000 ;
	    RECT 155.0000 90.2000 155.6000 93.6000 ;
	    RECT 156.4000 92.3000 157.2000 93.2000 ;
	    RECT 158.0000 92.3000 158.8000 92.4000 ;
	    RECT 156.4000 91.7000 158.8000 92.3000 ;
	    RECT 156.4000 91.6000 157.2000 91.7000 ;
	    RECT 158.0000 91.6000 158.8000 91.7000 ;
	    RECT 159.6000 90.2000 160.4000 90.4000 ;
	    RECT 161.6000 90.2000 162.2000 93.6000 ;
	    RECT 162.8000 91.6000 163.6000 93.2000 ;
	    RECT 167.8000 90.2000 168.4000 93.6000 ;
	    RECT 169.2000 92.3000 170.0000 92.4000 ;
	    RECT 170.8000 92.3000 171.6000 92.4000 ;
	    RECT 169.2000 91.7000 171.6000 92.3000 ;
	    RECT 169.2000 90.8000 170.0000 91.7000 ;
	    RECT 170.8000 91.6000 171.6000 91.7000 ;
	    RECT 170.8000 90.2000 171.6000 90.4000 ;
	    RECT 172.8000 90.2000 173.4000 93.6000 ;
	    RECT 174.0000 91.6000 174.8000 93.2000 ;
	    RECT 178.8000 91.6000 179.6000 93.2000 ;
	    RECT 180.4000 90.4000 181.0000 93.6000 ;
	    RECT 182.0000 91.6000 182.8000 93.2000 ;
	    RECT 183.6000 92.8000 184.4000 94.4000 ;
	    RECT 185.2000 92.8000 186.0000 94.4000 ;
	    RECT 186.8000 93.8000 189.2000 94.4000 ;
	    RECT 190.8000 94.3000 192.4000 94.4000 ;
	    RECT 193.2000 94.3000 195.8000 94.4000 ;
	    RECT 190.8000 93.8000 195.8000 94.3000 ;
	    RECT 197.2000 93.8000 198.8000 94.4000 ;
	    RECT 188.4000 93.6000 189.2000 93.8000 ;
	    RECT 191.6000 93.7000 195.8000 93.8000 ;
	    RECT 191.6000 93.6000 192.4000 93.7000 ;
	    RECT 193.2000 93.6000 195.8000 93.7000 ;
	    RECT 198.0000 93.6000 198.8000 93.8000 ;
	    RECT 199.6000 93.6000 202.2000 94.4000 ;
	    RECT 203.6000 93.8000 205.2000 94.4000 ;
	    RECT 206.0000 94.2000 210.2000 94.8000 ;
	    RECT 204.4000 93.6000 205.2000 93.8000 ;
	    RECT 209.2000 93.8000 210.2000 94.2000 ;
	    RECT 211.2000 94.4000 211.8000 95.0000 ;
	    RECT 218.6000 95.4000 220.2000 96.0000 ;
	    RECT 218.6000 95.0000 219.4000 95.4000 ;
	    RECT 218.6000 94.4000 219.2000 95.0000 ;
	    RECT 223.8000 94.8000 224.4000 97.0000 ;
	    RECT 225.2000 95.6000 226.0000 97.2000 ;
	    RECT 186.8000 91.6000 187.6000 93.2000 ;
	    RECT 188.6000 90.4000 189.2000 93.6000 ;
	    RECT 190.0000 91.6000 190.8000 93.2000 ;
	    RECT 178.8000 90.2000 181.0000 90.4000 ;
	    RECT 186.8000 90.2000 189.2000 90.4000 ;
	    RECT 193.2000 90.2000 194.0000 90.4000 ;
	    RECT 195.2000 90.2000 195.8000 93.6000 ;
	    RECT 196.4000 91.6000 197.2000 93.2000 ;
	    RECT 199.6000 90.2000 200.4000 90.4000 ;
	    RECT 201.6000 90.2000 202.2000 93.6000 ;
	    RECT 202.8000 91.6000 203.6000 93.2000 ;
	    RECT 206.0000 91.6000 206.8000 93.2000 ;
	    RECT 207.6000 91.6000 208.4000 93.2000 ;
	    RECT 209.2000 93.0000 210.6000 93.8000 ;
	    RECT 211.2000 93.6000 213.2000 94.4000 ;
	    RECT 217.2000 93.6000 219.2000 94.4000 ;
	    RECT 220.2000 94.2000 224.4000 94.8000 ;
	    RECT 227.0000 94.4000 227.6000 97.8000 ;
	    RECT 232.6000 96.4000 233.4000 99.8000 ;
	    RECT 231.6000 95.8000 233.4000 96.4000 ;
	    RECT 234.8000 95.8000 235.6000 99.8000 ;
	    RECT 236.4000 96.0000 237.2000 99.8000 ;
	    RECT 239.6000 96.0000 240.4000 99.8000 ;
	    RECT 236.4000 95.8000 240.4000 96.0000 ;
	    RECT 220.2000 93.8000 221.2000 94.2000 ;
	    RECT 209.2000 91.0000 209.8000 93.0000 ;
	    RECT 206.0000 90.4000 209.8000 91.0000 ;
	    RECT 111.6000 89.7000 114.6000 90.2000 ;
	    RECT 111.6000 89.6000 112.4000 89.7000 ;
	    RECT 113.2000 89.6000 114.6000 89.7000 ;
	    RECT 115.2000 89.6000 116.2000 90.2000 ;
	    RECT 119.6000 89.6000 121.0000 90.2000 ;
	    RECT 121.6000 89.6000 122.6000 90.2000 ;
	    RECT 126.0000 89.6000 127.4000 90.2000 ;
	    RECT 128.0000 89.6000 129.0000 90.2000 ;
	    RECT 103.0000 82.2000 103.8000 89.6000 ;
	    RECT 104.6000 88.4000 105.2000 89.6000 ;
	    RECT 104.4000 87.6000 105.2000 88.4000 ;
	    RECT 114.0000 88.4000 114.6000 89.6000 ;
	    RECT 114.0000 87.6000 114.8000 88.4000 ;
	    RECT 115.4000 82.2000 116.2000 89.6000 ;
	    RECT 120.4000 88.4000 121.0000 89.6000 ;
	    RECT 120.4000 87.6000 121.2000 88.4000 ;
	    RECT 121.8000 82.2000 122.6000 89.6000 ;
	    RECT 126.8000 88.4000 127.4000 89.6000 ;
	    RECT 126.8000 87.6000 127.6000 88.4000 ;
	    RECT 128.2000 82.2000 129.0000 89.6000 ;
	    RECT 134.0000 89.4000 135.8000 90.2000 ;
	    RECT 135.0000 84.4000 135.8000 89.4000 ;
	    RECT 134.0000 83.6000 135.8000 84.4000 ;
	    RECT 135.0000 82.2000 135.8000 83.6000 ;
	    RECT 139.8000 82.2000 141.8000 90.2000 ;
	    RECT 145.2000 89.6000 146.6000 90.2000 ;
	    RECT 147.2000 89.6000 148.2000 90.2000 ;
	    RECT 146.0000 88.4000 146.6000 89.6000 ;
	    RECT 146.0000 87.6000 146.8000 88.4000 ;
	    RECT 147.4000 82.2000 148.2000 89.6000 ;
	    RECT 154.2000 82.2000 156.2000 90.2000 ;
	    RECT 159.6000 89.6000 161.0000 90.2000 ;
	    RECT 161.6000 89.6000 162.6000 90.2000 ;
	    RECT 160.4000 88.4000 161.0000 89.6000 ;
	    RECT 160.4000 87.6000 161.2000 88.4000 ;
	    RECT 161.8000 82.2000 162.6000 89.6000 ;
	    RECT 167.6000 89.4000 169.4000 90.2000 ;
	    RECT 170.8000 89.6000 172.2000 90.2000 ;
	    RECT 172.8000 89.6000 173.8000 90.2000 ;
	    RECT 178.8000 89.6000 181.8000 90.2000 ;
	    RECT 186.8000 89.6000 189.8000 90.2000 ;
	    RECT 193.2000 89.6000 194.6000 90.2000 ;
	    RECT 195.2000 89.6000 196.2000 90.2000 ;
	    RECT 199.6000 89.6000 201.0000 90.2000 ;
	    RECT 201.6000 89.6000 202.6000 90.2000 ;
	    RECT 168.6000 84.4000 169.4000 89.4000 ;
	    RECT 171.6000 88.4000 172.2000 89.6000 ;
	    RECT 171.6000 87.6000 172.4000 88.4000 ;
	    RECT 167.6000 83.6000 169.4000 84.4000 ;
	    RECT 168.6000 82.2000 169.4000 83.6000 ;
	    RECT 173.0000 84.4000 173.8000 89.6000 ;
	    RECT 173.0000 83.6000 174.8000 84.4000 ;
	    RECT 173.0000 82.2000 173.8000 83.6000 ;
	    RECT 179.8000 82.2000 181.8000 89.6000 ;
	    RECT 187.8000 82.2000 189.8000 89.6000 ;
	    RECT 194.0000 88.4000 194.6000 89.6000 ;
	    RECT 194.0000 87.6000 194.8000 88.4000 ;
	    RECT 195.4000 82.2000 196.2000 89.6000 ;
	    RECT 200.4000 88.4000 201.0000 89.6000 ;
	    RECT 200.4000 87.6000 201.2000 88.4000 ;
	    RECT 201.8000 84.4000 202.6000 89.6000 ;
	    RECT 206.0000 87.0000 206.6000 90.4000 ;
	    RECT 211.2000 89.8000 211.8000 93.6000 ;
	    RECT 212.4000 92.3000 213.2000 92.4000 ;
	    RECT 215.6000 92.3000 216.4000 92.4000 ;
	    RECT 217.2000 92.3000 218.0000 92.4000 ;
	    RECT 212.4000 91.7000 218.0000 92.3000 ;
	    RECT 212.4000 90.8000 213.2000 91.7000 ;
	    RECT 215.6000 91.6000 216.4000 91.7000 ;
	    RECT 217.2000 90.8000 218.0000 91.7000 ;
	    RECT 210.2000 89.2000 211.8000 89.8000 ;
	    RECT 218.6000 90.4000 219.2000 93.6000 ;
	    RECT 219.8000 93.0000 221.2000 93.8000 ;
	    RECT 226.8000 93.6000 227.6000 94.4000 ;
	    RECT 230.0000 93.6000 230.8000 95.2000 ;
	    RECT 220.6000 91.0000 221.2000 93.0000 ;
	    RECT 222.0000 91.6000 222.8000 93.2000 ;
	    RECT 223.6000 91.6000 224.4000 93.2000 ;
	    RECT 220.6000 90.4000 224.4000 91.0000 ;
	    RECT 218.6000 89.8000 219.6000 90.4000 ;
	    RECT 218.6000 89.2000 220.2000 89.8000 ;
	    RECT 201.8000 83.6000 203.6000 84.4000 ;
	    RECT 201.8000 82.2000 202.6000 83.6000 ;
	    RECT 206.0000 83.0000 206.8000 87.0000 ;
	    RECT 210.2000 82.2000 211.0000 89.2000 ;
	    RECT 219.4000 82.2000 220.2000 89.2000 ;
	    RECT 223.8000 87.0000 224.4000 90.4000 ;
	    RECT 227.0000 90.2000 227.6000 93.6000 ;
	    RECT 228.4000 90.8000 229.2000 92.4000 ;
	    RECT 231.6000 92.3000 232.4000 95.8000 ;
	    RECT 235.0000 94.4000 235.6000 95.8000 ;
	    RECT 236.6000 95.4000 240.2000 95.8000 ;
	    RECT 241.2000 95.4000 242.0000 99.8000 ;
	    RECT 245.4000 98.4000 246.6000 99.8000 ;
	    RECT 245.4000 97.8000 246.8000 98.4000 ;
	    RECT 250.0000 97.8000 250.8000 99.8000 ;
	    RECT 254.4000 98.4000 255.2000 99.8000 ;
	    RECT 254.4000 97.8000 256.4000 98.4000 ;
	    RECT 246.0000 97.0000 246.8000 97.8000 ;
	    RECT 250.2000 97.2000 250.8000 97.8000 ;
	    RECT 250.2000 96.6000 253.0000 97.2000 ;
	    RECT 252.2000 96.4000 253.0000 96.6000 ;
	    RECT 254.0000 96.4000 254.8000 97.2000 ;
	    RECT 255.6000 97.0000 256.4000 97.8000 ;
	    RECT 244.2000 95.4000 245.0000 95.6000 ;
	    RECT 241.2000 94.8000 245.0000 95.4000 ;
	    RECT 238.8000 94.4000 239.6000 94.8000 ;
	    RECT 234.8000 93.6000 237.4000 94.4000 ;
	    RECT 238.8000 93.8000 240.4000 94.4000 ;
	    RECT 239.6000 93.6000 240.4000 93.8000 ;
	    RECT 231.6000 91.7000 235.5000 92.3000 ;
	    RECT 226.8000 89.4000 228.6000 90.2000 ;
	    RECT 223.6000 83.0000 224.4000 87.0000 ;
	    RECT 227.8000 86.4000 228.6000 89.4000 ;
	    RECT 226.8000 85.6000 228.6000 86.4000 ;
	    RECT 227.8000 82.2000 228.6000 85.6000 ;
	    RECT 231.6000 82.2000 232.4000 91.7000 ;
	    RECT 234.9000 90.4000 235.5000 91.7000 ;
	    RECT 236.8000 90.4000 237.4000 93.6000 ;
	    RECT 238.0000 91.6000 238.8000 93.2000 ;
	    RECT 241.2000 91.4000 242.0000 94.8000 ;
	    RECT 254.0000 94.4000 254.6000 96.4000 ;
	    RECT 258.8000 95.0000 259.6000 99.8000 ;
	    RECT 263.6000 98.3000 264.4000 98.4000 ;
	    RECT 267.4000 98.3000 268.2000 99.8000 ;
	    RECT 263.6000 97.7000 268.2000 98.3000 ;
	    RECT 263.6000 97.6000 264.4000 97.7000 ;
	    RECT 267.4000 96.4000 268.2000 97.7000 ;
	    RECT 267.4000 95.8000 269.2000 96.4000 ;
	    RECT 248.2000 94.2000 249.0000 94.4000 ;
	    RECT 254.0000 94.2000 254.8000 94.4000 ;
	    RECT 257.2000 94.2000 258.8000 94.4000 ;
	    RECT 247.8000 93.6000 258.8000 94.2000 ;
	    RECT 260.4000 94.3000 261.2000 94.4000 ;
	    RECT 266.8000 94.3000 267.6000 94.4000 ;
	    RECT 260.4000 93.7000 267.6000 94.3000 ;
	    RECT 260.4000 93.6000 261.2000 93.7000 ;
	    RECT 266.8000 93.6000 267.6000 93.7000 ;
	    RECT 246.0000 92.8000 246.8000 93.0000 ;
	    RECT 243.0000 92.2000 246.8000 92.8000 ;
	    RECT 243.0000 92.0000 243.8000 92.2000 ;
	    RECT 244.6000 91.4000 245.4000 91.6000 ;
	    RECT 241.2000 90.8000 245.4000 91.4000 ;
	    RECT 233.2000 88.8000 234.0000 90.4000 ;
	    RECT 234.8000 90.2000 235.6000 90.4000 ;
	    RECT 234.8000 89.6000 236.2000 90.2000 ;
	    RECT 236.8000 89.6000 238.8000 90.4000 ;
	    RECT 235.6000 88.4000 236.2000 89.6000 ;
	    RECT 235.6000 87.6000 236.4000 88.4000 ;
	    RECT 237.0000 82.2000 237.8000 89.6000 ;
	    RECT 241.2000 82.2000 242.0000 90.8000 ;
	    RECT 247.8000 90.4000 248.4000 93.6000 ;
	    RECT 255.0000 93.4000 255.8000 93.6000 ;
	    RECT 256.6000 92.4000 257.4000 92.6000 ;
	    RECT 252.4000 91.8000 257.4000 92.4000 ;
	    RECT 252.4000 91.6000 253.2000 91.8000 ;
	    RECT 254.0000 91.0000 259.6000 91.2000 ;
	    RECT 253.8000 90.8000 259.6000 91.0000 ;
	    RECT 246.0000 89.8000 248.4000 90.4000 ;
	    RECT 249.8000 90.6000 259.6000 90.8000 ;
	    RECT 249.8000 90.2000 254.6000 90.6000 ;
	    RECT 246.0000 88.8000 246.6000 89.8000 ;
	    RECT 245.2000 88.0000 246.6000 88.8000 ;
	    RECT 248.2000 89.0000 249.0000 89.2000 ;
	    RECT 249.8000 89.0000 250.4000 90.2000 ;
	    RECT 248.2000 88.4000 250.4000 89.0000 ;
	    RECT 251.0000 89.0000 256.4000 89.6000 ;
	    RECT 251.0000 88.8000 251.8000 89.0000 ;
	    RECT 255.6000 88.8000 256.4000 89.0000 ;
	    RECT 249.4000 87.4000 250.2000 87.6000 ;
	    RECT 252.2000 87.4000 253.0000 87.6000 ;
	    RECT 246.0000 86.2000 246.8000 87.0000 ;
	    RECT 249.4000 86.8000 253.0000 87.4000 ;
	    RECT 250.2000 86.2000 250.8000 86.8000 ;
	    RECT 255.6000 86.2000 256.4000 87.0000 ;
	    RECT 245.4000 82.2000 246.6000 86.2000 ;
	    RECT 250.0000 82.2000 250.8000 86.2000 ;
	    RECT 254.4000 85.6000 256.4000 86.2000 ;
	    RECT 254.4000 82.2000 255.2000 85.6000 ;
	    RECT 258.8000 82.2000 259.6000 90.6000 ;
	    RECT 266.8000 88.8000 267.6000 90.4000 ;
	    RECT 268.4000 82.2000 269.2000 95.8000 ;
	    RECT 270.0000 93.6000 270.8000 95.2000 ;
	    RECT 271.6000 92.4000 272.4000 99.8000 ;
	    RECT 274.8000 95.2000 275.6000 99.8000 ;
	    RECT 273.4000 94.6000 275.6000 95.2000 ;
	    RECT 271.6000 90.2000 272.2000 92.4000 ;
	    RECT 273.4000 91.6000 274.0000 94.6000 ;
	    RECT 274.8000 91.6000 275.6000 93.2000 ;
	    RECT 276.4000 92.4000 277.2000 99.8000 ;
	    RECT 279.6000 95.2000 280.4000 99.8000 ;
	    RECT 281.2000 99.2000 285.2000 99.8000 ;
	    RECT 281.2000 95.8000 282.0000 99.2000 ;
	    RECT 282.8000 95.8000 283.6000 98.6000 ;
	    RECT 284.4000 96.0000 285.2000 99.2000 ;
	    RECT 287.6000 96.0000 288.4000 99.8000 ;
	    RECT 284.4000 95.8000 288.4000 96.0000 ;
	    RECT 278.2000 94.6000 280.4000 95.2000 ;
	    RECT 272.8000 90.8000 274.0000 91.6000 ;
	    RECT 273.4000 90.2000 274.0000 90.8000 ;
	    RECT 276.4000 90.2000 277.0000 92.4000 ;
	    RECT 278.2000 91.6000 278.8000 94.6000 ;
	    RECT 282.8000 94.4000 283.4000 95.8000 ;
	    RECT 284.6000 95.4000 288.2000 95.8000 ;
	    RECT 289.2000 95.2000 290.0000 99.8000 ;
	    RECT 286.8000 94.4000 287.6000 94.8000 ;
	    RECT 289.2000 94.6000 291.4000 95.2000 ;
	    RECT 281.2000 92.8000 282.0000 94.4000 ;
	    RECT 282.8000 93.8000 285.2000 94.4000 ;
	    RECT 286.8000 93.8000 288.4000 94.4000 ;
	    RECT 284.4000 93.6000 285.2000 93.8000 ;
	    RECT 287.6000 93.6000 288.4000 93.8000 ;
	    RECT 282.8000 91.6000 283.6000 93.2000 ;
	    RECT 277.6000 90.8000 278.8000 91.6000 ;
	    RECT 278.2000 90.2000 278.8000 90.8000 ;
	    RECT 284.6000 90.2000 285.2000 93.6000 ;
	    RECT 286.0000 91.6000 286.8000 93.2000 ;
	    RECT 290.8000 91.6000 291.4000 94.6000 ;
	    RECT 292.4000 94.3000 293.2000 99.8000 ;
	    RECT 294.0000 96.0000 294.8000 99.8000 ;
	    RECT 297.2000 96.0000 298.0000 99.8000 ;
	    RECT 294.0000 95.8000 298.0000 96.0000 ;
	    RECT 298.8000 95.8000 299.6000 99.8000 ;
	    RECT 300.4000 99.2000 304.4000 99.8000 ;
	    RECT 300.4000 95.8000 301.2000 99.2000 ;
	    RECT 302.0000 95.8000 302.8000 98.6000 ;
	    RECT 303.6000 96.0000 304.4000 99.2000 ;
	    RECT 306.8000 96.0000 307.6000 99.8000 ;
	    RECT 303.6000 95.8000 307.6000 96.0000 ;
	    RECT 308.4000 95.8000 309.2000 99.8000 ;
	    RECT 310.0000 96.0000 310.8000 99.8000 ;
	    RECT 313.2000 96.0000 314.0000 99.8000 ;
	    RECT 310.0000 95.8000 314.0000 96.0000 ;
	    RECT 316.4000 97.8000 317.2000 99.8000 ;
	    RECT 294.2000 95.4000 297.8000 95.8000 ;
	    RECT 294.8000 94.4000 295.6000 94.8000 ;
	    RECT 298.8000 94.4000 299.4000 95.8000 ;
	    RECT 302.0000 94.4000 302.6000 95.8000 ;
	    RECT 303.8000 95.4000 307.4000 95.8000 ;
	    RECT 306.0000 94.4000 306.8000 94.8000 ;
	    RECT 308.6000 94.4000 309.2000 95.8000 ;
	    RECT 310.2000 95.4000 313.8000 95.8000 ;
	    RECT 312.4000 94.4000 313.2000 94.8000 ;
	    RECT 316.4000 94.4000 317.0000 97.8000 ;
	    RECT 318.0000 95.6000 318.8000 97.2000 ;
	    RECT 319.6000 96.0000 320.4000 99.8000 ;
	    RECT 322.8000 99.2000 326.8000 99.8000 ;
	    RECT 322.8000 96.0000 323.6000 99.2000 ;
	    RECT 319.6000 95.8000 323.6000 96.0000 ;
	    RECT 324.4000 95.8000 325.2000 98.6000 ;
	    RECT 326.0000 95.8000 326.8000 99.2000 ;
	    RECT 319.8000 95.4000 323.4000 95.8000 ;
	    RECT 320.4000 94.4000 321.2000 94.8000 ;
	    RECT 324.6000 94.4000 325.2000 95.8000 ;
	    RECT 327.6000 95.2000 328.4000 99.8000 ;
	    RECT 327.6000 94.6000 329.8000 95.2000 ;
	    RECT 294.0000 94.3000 295.6000 94.4000 ;
	    RECT 292.4000 93.8000 295.6000 94.3000 ;
	    RECT 292.4000 93.7000 294.8000 93.8000 ;
	    RECT 292.4000 92.4000 293.2000 93.7000 ;
	    RECT 294.0000 93.6000 294.8000 93.7000 ;
	    RECT 297.0000 93.6000 299.6000 94.4000 ;
	    RECT 290.8000 90.8000 292.0000 91.6000 ;
	    RECT 290.8000 90.2000 291.4000 90.8000 ;
	    RECT 292.6000 90.2000 293.2000 92.4000 ;
	    RECT 295.6000 91.6000 296.4000 93.2000 ;
	    RECT 297.0000 90.4000 297.6000 93.6000 ;
	    RECT 300.4000 92.8000 301.2000 94.4000 ;
	    RECT 302.0000 93.8000 304.4000 94.4000 ;
	    RECT 306.0000 94.3000 307.6000 94.4000 ;
	    RECT 308.4000 94.3000 311.0000 94.4000 ;
	    RECT 306.0000 93.8000 311.0000 94.3000 ;
	    RECT 312.4000 93.8000 314.0000 94.4000 ;
	    RECT 303.6000 93.6000 304.4000 93.8000 ;
	    RECT 306.8000 93.7000 311.0000 93.8000 ;
	    RECT 306.8000 93.6000 307.6000 93.7000 ;
	    RECT 308.4000 93.6000 311.0000 93.7000 ;
	    RECT 313.2000 93.6000 314.0000 93.8000 ;
	    RECT 316.4000 93.6000 317.2000 94.4000 ;
	    RECT 319.6000 93.8000 321.2000 94.4000 ;
	    RECT 322.8000 93.8000 325.2000 94.4000 ;
	    RECT 319.6000 93.6000 320.4000 93.8000 ;
	    RECT 322.8000 93.6000 323.6000 93.8000 ;
	    RECT 302.0000 91.6000 302.8000 93.2000 ;
	    RECT 271.6000 82.2000 272.4000 90.2000 ;
	    RECT 273.4000 89.6000 275.6000 90.2000 ;
	    RECT 274.8000 82.2000 275.6000 89.6000 ;
	    RECT 276.4000 82.2000 277.2000 90.2000 ;
	    RECT 278.2000 89.6000 280.4000 90.2000 ;
	    RECT 279.6000 82.2000 280.4000 89.6000 ;
	    RECT 283.8000 82.2000 285.8000 90.2000 ;
	    RECT 289.2000 89.6000 291.4000 90.2000 ;
	    RECT 289.2000 82.2000 290.0000 89.6000 ;
	    RECT 292.4000 82.2000 293.2000 90.2000 ;
	    RECT 295.6000 89.6000 297.6000 90.4000 ;
	    RECT 298.8000 90.2000 299.6000 90.4000 ;
	    RECT 303.8000 90.2000 304.4000 93.6000 ;
	    RECT 305.2000 92.3000 306.0000 93.2000 ;
	    RECT 308.4000 92.3000 309.2000 92.4000 ;
	    RECT 305.2000 91.7000 309.2000 92.3000 ;
	    RECT 305.2000 91.6000 306.0000 91.7000 ;
	    RECT 308.4000 91.6000 309.2000 91.7000 ;
	    RECT 308.4000 90.2000 309.2000 90.4000 ;
	    RECT 310.4000 90.2000 311.0000 93.6000 ;
	    RECT 311.6000 91.6000 312.4000 93.2000 ;
	    RECT 314.8000 90.8000 315.6000 92.4000 ;
	    RECT 316.4000 92.3000 317.0000 93.6000 ;
	    RECT 321.2000 92.3000 322.0000 93.2000 ;
	    RECT 316.4000 91.7000 322.0000 92.3000 ;
	    RECT 316.4000 90.2000 317.0000 91.7000 ;
	    RECT 321.2000 91.6000 322.0000 91.7000 ;
	    RECT 322.8000 92.4000 323.4000 93.6000 ;
	    RECT 322.8000 91.6000 323.6000 92.4000 ;
	    RECT 324.4000 91.6000 325.2000 93.2000 ;
	    RECT 326.0000 92.8000 326.8000 94.4000 ;
	    RECT 329.2000 91.6000 329.8000 94.6000 ;
	    RECT 330.8000 92.4000 331.6000 99.8000 ;
	    RECT 332.4000 97.0000 333.2000 99.0000 ;
	    RECT 332.4000 94.8000 333.0000 97.0000 ;
	    RECT 336.6000 96.4000 337.4000 99.0000 ;
	    RECT 345.8000 98.4000 346.6000 99.0000 ;
	    RECT 345.2000 97.6000 346.6000 98.4000 ;
	    RECT 335.6000 96.0000 337.4000 96.4000 ;
	    RECT 345.8000 96.0000 346.6000 97.6000 ;
	    RECT 350.0000 97.0000 350.8000 99.0000 ;
	    RECT 335.6000 95.6000 338.2000 96.0000 ;
	    RECT 336.6000 95.4000 338.2000 95.6000 ;
	    RECT 337.4000 95.0000 338.2000 95.4000 ;
	    RECT 332.4000 94.2000 336.6000 94.8000 ;
	    RECT 335.6000 93.8000 336.6000 94.2000 ;
	    RECT 337.6000 94.4000 338.2000 95.0000 ;
	    RECT 345.0000 95.4000 346.6000 96.0000 ;
	    RECT 345.0000 95.0000 345.8000 95.4000 ;
	    RECT 345.0000 94.4000 345.6000 95.0000 ;
	    RECT 350.2000 94.8000 350.8000 97.0000 ;
	    RECT 322.8000 90.2000 323.4000 91.6000 ;
	    RECT 329.2000 90.8000 330.4000 91.6000 ;
	    RECT 329.2000 90.2000 329.8000 90.8000 ;
	    RECT 331.0000 90.2000 331.6000 92.4000 ;
	    RECT 332.4000 91.6000 333.2000 93.2000 ;
	    RECT 334.0000 91.6000 334.8000 93.2000 ;
	    RECT 335.6000 93.0000 337.0000 93.8000 ;
	    RECT 337.6000 93.6000 339.6000 94.4000 ;
	    RECT 343.6000 93.6000 345.6000 94.4000 ;
	    RECT 346.6000 94.2000 350.8000 94.8000 ;
	    RECT 353.2000 97.8000 354.0000 99.8000 ;
	    RECT 353.2000 94.4000 353.8000 97.8000 ;
	    RECT 354.8000 95.6000 355.6000 97.2000 ;
	    RECT 356.4000 96.0000 357.2000 99.8000 ;
	    RECT 359.6000 99.2000 363.6000 99.8000 ;
	    RECT 359.6000 96.0000 360.4000 99.2000 ;
	    RECT 356.4000 95.8000 360.4000 96.0000 ;
	    RECT 361.2000 95.8000 362.0000 98.6000 ;
	    RECT 362.8000 95.8000 363.6000 99.2000 ;
	    RECT 364.4000 95.8000 365.2000 99.8000 ;
	    RECT 366.0000 96.0000 366.8000 99.8000 ;
	    RECT 369.2000 96.0000 370.0000 99.8000 ;
	    RECT 366.0000 95.8000 370.0000 96.0000 ;
	    RECT 356.6000 95.4000 360.2000 95.8000 ;
	    RECT 357.2000 94.4000 358.0000 94.8000 ;
	    RECT 361.4000 94.4000 362.0000 95.8000 ;
	    RECT 364.6000 94.4000 365.2000 95.8000 ;
	    RECT 366.2000 95.4000 369.8000 95.8000 ;
	    RECT 368.4000 94.4000 369.2000 94.8000 ;
	    RECT 346.6000 93.8000 347.6000 94.2000 ;
	    RECT 335.6000 91.0000 336.2000 93.0000 ;
	    RECT 298.2000 89.6000 299.6000 90.2000 ;
	    RECT 296.6000 82.2000 297.4000 89.6000 ;
	    RECT 298.2000 88.4000 298.8000 89.6000 ;
	    RECT 298.0000 87.6000 298.8000 88.4000 ;
	    RECT 303.0000 84.4000 305.0000 90.2000 ;
	    RECT 308.4000 89.6000 309.8000 90.2000 ;
	    RECT 310.4000 89.6000 311.4000 90.2000 ;
	    RECT 309.2000 88.4000 309.8000 89.6000 ;
	    RECT 309.2000 87.6000 310.0000 88.4000 ;
	    RECT 302.0000 83.6000 305.0000 84.4000 ;
	    RECT 303.0000 82.2000 305.0000 83.6000 ;
	    RECT 310.6000 82.2000 311.4000 89.6000 ;
	    RECT 315.4000 89.4000 317.2000 90.2000 ;
	    RECT 315.4000 82.2000 316.2000 89.4000 ;
	    RECT 322.2000 82.2000 324.2000 90.2000 ;
	    RECT 327.6000 89.6000 329.8000 90.2000 ;
	    RECT 327.6000 82.2000 328.4000 89.6000 ;
	    RECT 330.8000 82.2000 331.6000 90.2000 ;
	    RECT 332.4000 90.4000 336.2000 91.0000 ;
	    RECT 332.4000 87.0000 333.0000 90.4000 ;
	    RECT 337.6000 89.8000 338.2000 93.6000 ;
	    RECT 338.8000 92.3000 339.6000 92.4000 ;
	    RECT 343.6000 92.3000 344.4000 92.4000 ;
	    RECT 338.8000 91.7000 344.4000 92.3000 ;
	    RECT 338.8000 90.8000 339.6000 91.7000 ;
	    RECT 343.6000 90.8000 344.4000 91.7000 ;
	    RECT 336.6000 89.2000 338.2000 89.8000 ;
	    RECT 345.0000 89.8000 345.6000 93.6000 ;
	    RECT 346.2000 93.0000 347.6000 93.8000 ;
	    RECT 353.2000 93.6000 354.0000 94.4000 ;
	    RECT 356.4000 93.8000 358.0000 94.4000 ;
	    RECT 359.6000 93.8000 362.0000 94.4000 ;
	    RECT 356.4000 93.6000 357.2000 93.8000 ;
	    RECT 359.6000 93.6000 360.4000 93.8000 ;
	    RECT 347.0000 91.0000 347.6000 93.0000 ;
	    RECT 348.4000 91.6000 349.2000 93.2000 ;
	    RECT 350.0000 91.6000 350.8000 93.2000 ;
	    RECT 347.0000 90.4000 350.8000 91.0000 ;
	    RECT 351.6000 90.8000 352.4000 92.4000 ;
	    RECT 353.2000 92.3000 353.8000 93.6000 ;
	    RECT 358.0000 92.3000 358.8000 93.2000 ;
	    RECT 353.2000 91.7000 358.8000 92.3000 ;
	    RECT 345.0000 89.2000 346.6000 89.8000 ;
	    RECT 332.4000 83.0000 333.2000 87.0000 ;
	    RECT 336.6000 82.2000 337.4000 89.2000 ;
	    RECT 345.8000 82.2000 346.6000 89.2000 ;
	    RECT 350.2000 87.0000 350.8000 90.4000 ;
	    RECT 353.2000 90.2000 353.8000 91.7000 ;
	    RECT 358.0000 91.6000 358.8000 91.7000 ;
	    RECT 359.6000 90.2000 360.2000 93.6000 ;
	    RECT 361.2000 91.6000 362.0000 93.2000 ;
	    RECT 362.8000 92.3000 363.6000 94.4000 ;
	    RECT 364.4000 93.6000 367.0000 94.4000 ;
	    RECT 368.4000 93.8000 370.0000 94.4000 ;
	    RECT 369.2000 93.6000 370.0000 93.8000 ;
	    RECT 362.8000 91.7000 365.1000 92.3000 ;
	    RECT 364.5000 90.4000 365.1000 91.7000 ;
	    RECT 364.4000 90.2000 365.2000 90.4000 ;
	    RECT 366.4000 90.2000 367.0000 93.6000 ;
	    RECT 367.6000 91.6000 368.4000 93.2000 ;
	    RECT 370.8000 92.4000 371.6000 99.8000 ;
	    RECT 374.0000 95.2000 374.8000 99.8000 ;
	    RECT 375.6000 96.0000 376.4000 99.8000 ;
	    RECT 378.8000 96.0000 379.6000 99.8000 ;
	    RECT 375.6000 95.8000 379.6000 96.0000 ;
	    RECT 380.4000 95.8000 381.2000 99.8000 ;
	    RECT 382.0000 95.8000 382.8000 99.8000 ;
	    RECT 383.6000 96.0000 384.4000 99.8000 ;
	    RECT 386.8000 96.0000 387.6000 99.8000 ;
	    RECT 383.6000 95.8000 387.6000 96.0000 ;
	    RECT 375.8000 95.4000 379.4000 95.8000 ;
	    RECT 372.6000 94.6000 374.8000 95.2000 ;
	    RECT 370.8000 90.2000 371.4000 92.4000 ;
	    RECT 372.6000 91.6000 373.2000 94.6000 ;
	    RECT 376.4000 94.4000 377.2000 94.8000 ;
	    RECT 380.4000 94.4000 381.0000 95.8000 ;
	    RECT 382.2000 94.4000 382.8000 95.8000 ;
	    RECT 383.8000 95.4000 387.4000 95.8000 ;
	    RECT 388.4000 95.4000 389.2000 99.8000 ;
	    RECT 392.6000 98.4000 393.8000 99.8000 ;
	    RECT 392.6000 97.8000 394.0000 98.4000 ;
	    RECT 397.2000 97.8000 398.0000 99.8000 ;
	    RECT 401.6000 98.4000 402.4000 99.8000 ;
	    RECT 401.6000 97.8000 403.6000 98.4000 ;
	    RECT 393.2000 97.0000 394.0000 97.8000 ;
	    RECT 397.4000 97.2000 398.0000 97.8000 ;
	    RECT 397.4000 96.6000 400.2000 97.2000 ;
	    RECT 399.4000 96.4000 400.2000 96.6000 ;
	    RECT 401.2000 96.4000 402.0000 97.2000 ;
	    RECT 402.8000 97.0000 403.6000 97.8000 ;
	    RECT 391.4000 95.4000 392.2000 95.6000 ;
	    RECT 388.4000 94.8000 392.2000 95.4000 ;
	    RECT 386.0000 94.4000 386.8000 94.8000 ;
	    RECT 375.6000 93.8000 377.2000 94.4000 ;
	    RECT 375.6000 93.6000 376.4000 93.8000 ;
	    RECT 378.6000 93.6000 381.2000 94.4000 ;
	    RECT 382.0000 93.6000 384.6000 94.4000 ;
	    RECT 386.0000 93.8000 387.6000 94.4000 ;
	    RECT 386.8000 93.6000 387.6000 93.8000 ;
	    RECT 374.0000 91.6000 374.8000 93.2000 ;
	    RECT 377.2000 91.6000 378.0000 93.2000 ;
	    RECT 378.6000 92.3000 379.2000 93.6000 ;
	    RECT 384.0000 92.4000 384.6000 93.6000 ;
	    RECT 378.6000 91.7000 382.7000 92.3000 ;
	    RECT 372.0000 90.8000 373.2000 91.6000 ;
	    RECT 372.6000 90.2000 373.2000 90.8000 ;
	    RECT 378.6000 90.2000 379.2000 91.7000 ;
	    RECT 382.1000 90.4000 382.7000 91.7000 ;
	    RECT 383.6000 91.6000 384.6000 92.4000 ;
	    RECT 385.2000 91.6000 386.0000 93.2000 ;
	    RECT 380.4000 90.2000 381.2000 90.4000 ;
	    RECT 350.0000 83.0000 350.8000 87.0000 ;
	    RECT 352.2000 89.4000 354.0000 90.2000 ;
	    RECT 352.2000 82.2000 353.0000 89.4000 ;
	    RECT 359.0000 84.4000 361.0000 90.2000 ;
	    RECT 364.4000 89.6000 365.8000 90.2000 ;
	    RECT 366.4000 89.6000 367.4000 90.2000 ;
	    RECT 365.2000 88.4000 365.8000 89.6000 ;
	    RECT 365.2000 87.6000 366.0000 88.4000 ;
	    RECT 358.0000 83.6000 361.0000 84.4000 ;
	    RECT 359.0000 82.2000 361.0000 83.6000 ;
	    RECT 366.6000 82.2000 367.4000 89.6000 ;
	    RECT 370.8000 82.2000 371.6000 90.2000 ;
	    RECT 372.6000 89.6000 374.8000 90.2000 ;
	    RECT 374.0000 82.2000 374.8000 89.6000 ;
	    RECT 378.2000 89.6000 379.2000 90.2000 ;
	    RECT 379.8000 89.6000 381.2000 90.2000 ;
	    RECT 382.0000 90.2000 382.8000 90.4000 ;
	    RECT 384.0000 90.2000 384.6000 91.6000 ;
	    RECT 388.4000 91.4000 389.2000 94.8000 ;
	    RECT 395.4000 94.2000 396.2000 94.4000 ;
	    RECT 401.2000 94.2000 401.8000 96.4000 ;
	    RECT 406.0000 95.0000 406.8000 99.8000 ;
	    RECT 414.0000 95.4000 414.8000 99.8000 ;
	    RECT 418.2000 98.4000 419.4000 99.8000 ;
	    RECT 418.2000 97.8000 419.6000 98.4000 ;
	    RECT 422.8000 97.8000 423.6000 99.8000 ;
	    RECT 427.2000 98.4000 428.0000 99.8000 ;
	    RECT 427.2000 97.8000 429.2000 98.4000 ;
	    RECT 418.8000 97.0000 419.6000 97.8000 ;
	    RECT 423.0000 97.2000 423.6000 97.8000 ;
	    RECT 423.0000 96.6000 425.8000 97.2000 ;
	    RECT 425.0000 96.4000 425.8000 96.6000 ;
	    RECT 426.8000 96.4000 427.6000 97.2000 ;
	    RECT 428.4000 97.0000 429.2000 97.8000 ;
	    RECT 417.0000 95.4000 417.8000 95.6000 ;
	    RECT 414.0000 94.8000 417.8000 95.4000 ;
	    RECT 404.4000 94.2000 406.0000 94.4000 ;
	    RECT 395.0000 93.6000 406.0000 94.2000 ;
	    RECT 393.2000 92.8000 394.0000 93.0000 ;
	    RECT 390.2000 92.2000 394.0000 92.8000 ;
	    RECT 390.2000 92.0000 391.0000 92.2000 ;
	    RECT 391.8000 91.4000 392.6000 91.6000 ;
	    RECT 388.4000 90.8000 392.6000 91.4000 ;
	    RECT 382.0000 89.6000 383.4000 90.2000 ;
	    RECT 384.0000 89.6000 385.0000 90.2000 ;
	    RECT 378.2000 82.2000 379.0000 89.6000 ;
	    RECT 379.8000 88.4000 380.4000 89.6000 ;
	    RECT 379.6000 87.6000 380.4000 88.4000 ;
	    RECT 382.8000 88.4000 383.4000 89.6000 ;
	    RECT 382.8000 87.6000 383.6000 88.4000 ;
	    RECT 384.2000 82.2000 385.0000 89.6000 ;
	    RECT 388.4000 82.2000 389.2000 90.8000 ;
	    RECT 395.0000 90.4000 395.6000 93.6000 ;
	    RECT 402.2000 93.4000 403.0000 93.6000 ;
	    RECT 403.8000 92.4000 404.6000 92.6000 ;
	    RECT 396.4000 92.3000 397.2000 92.4000 ;
	    RECT 399.6000 92.3000 404.6000 92.4000 ;
	    RECT 396.4000 91.8000 404.6000 92.3000 ;
	    RECT 396.4000 91.7000 400.4000 91.8000 ;
	    RECT 396.4000 91.6000 397.2000 91.7000 ;
	    RECT 399.6000 91.6000 400.4000 91.7000 ;
	    RECT 414.0000 91.4000 414.8000 94.8000 ;
	    RECT 421.0000 94.2000 421.8000 94.4000 ;
	    RECT 423.6000 94.2000 424.4000 94.4000 ;
	    RECT 426.8000 94.2000 427.4000 96.4000 ;
	    RECT 431.6000 95.0000 432.4000 99.8000 ;
	    RECT 433.2000 95.8000 434.0000 99.8000 ;
	    RECT 434.8000 96.0000 435.6000 99.8000 ;
	    RECT 438.0000 96.0000 438.8000 99.8000 ;
	    RECT 434.8000 95.8000 438.8000 96.0000 ;
	    RECT 433.4000 94.4000 434.0000 95.8000 ;
	    RECT 435.0000 95.4000 438.6000 95.8000 ;
	    RECT 439.6000 95.4000 440.4000 99.8000 ;
	    RECT 443.8000 98.4000 445.0000 99.8000 ;
	    RECT 443.8000 97.8000 445.2000 98.4000 ;
	    RECT 448.4000 97.8000 449.2000 99.8000 ;
	    RECT 452.8000 98.4000 453.6000 99.8000 ;
	    RECT 452.8000 97.8000 454.8000 98.4000 ;
	    RECT 444.4000 97.0000 445.2000 97.8000 ;
	    RECT 448.6000 97.2000 449.2000 97.8000 ;
	    RECT 448.6000 96.6000 451.4000 97.2000 ;
	    RECT 450.6000 96.4000 451.4000 96.6000 ;
	    RECT 452.4000 96.4000 453.2000 97.2000 ;
	    RECT 454.0000 97.0000 454.8000 97.8000 ;
	    RECT 442.6000 95.4000 443.4000 95.6000 ;
	    RECT 439.6000 94.8000 443.4000 95.4000 ;
	    RECT 437.2000 94.4000 438.0000 94.8000 ;
	    RECT 430.0000 94.2000 431.6000 94.4000 ;
	    RECT 420.6000 93.6000 431.6000 94.2000 ;
	    RECT 433.2000 93.6000 435.8000 94.4000 ;
	    RECT 437.2000 93.8000 438.8000 94.4000 ;
	    RECT 438.0000 93.6000 438.8000 93.8000 ;
	    RECT 418.8000 92.8000 419.6000 93.0000 ;
	    RECT 415.8000 92.2000 419.6000 92.8000 ;
	    RECT 415.8000 92.0000 416.6000 92.2000 ;
	    RECT 417.4000 91.4000 418.2000 91.6000 ;
	    RECT 401.2000 91.0000 406.8000 91.2000 ;
	    RECT 401.0000 90.8000 406.8000 91.0000 ;
	    RECT 393.2000 89.8000 395.6000 90.4000 ;
	    RECT 397.0000 90.6000 406.8000 90.8000 ;
	    RECT 397.0000 90.2000 401.8000 90.6000 ;
	    RECT 393.2000 88.8000 393.8000 89.8000 ;
	    RECT 392.4000 88.0000 393.8000 88.8000 ;
	    RECT 395.4000 89.0000 396.2000 89.2000 ;
	    RECT 397.0000 89.0000 397.6000 90.2000 ;
	    RECT 395.4000 88.4000 397.6000 89.0000 ;
	    RECT 398.2000 89.0000 403.6000 89.6000 ;
	    RECT 398.2000 88.8000 399.0000 89.0000 ;
	    RECT 402.8000 88.8000 403.6000 89.0000 ;
	    RECT 396.6000 87.4000 397.4000 87.6000 ;
	    RECT 399.4000 87.4000 400.2000 87.6000 ;
	    RECT 393.2000 86.2000 394.0000 87.0000 ;
	    RECT 396.6000 86.8000 400.2000 87.4000 ;
	    RECT 397.4000 86.2000 398.0000 86.8000 ;
	    RECT 402.8000 86.2000 403.6000 87.0000 ;
	    RECT 392.6000 82.2000 393.8000 86.2000 ;
	    RECT 397.2000 82.2000 398.0000 86.2000 ;
	    RECT 401.6000 85.6000 403.6000 86.2000 ;
	    RECT 401.6000 82.2000 402.4000 85.6000 ;
	    RECT 406.0000 82.2000 406.8000 90.6000 ;
	    RECT 414.0000 90.8000 418.2000 91.4000 ;
	    RECT 414.0000 82.2000 414.8000 90.8000 ;
	    RECT 420.6000 90.4000 421.2000 93.6000 ;
	    RECT 427.8000 93.4000 428.6000 93.6000 ;
	    RECT 426.8000 92.4000 427.6000 92.6000 ;
	    RECT 429.4000 92.4000 430.2000 92.6000 ;
	    RECT 435.2000 92.4000 435.8000 93.6000 ;
	    RECT 425.2000 91.8000 430.2000 92.4000 ;
	    RECT 425.2000 91.6000 426.0000 91.8000 ;
	    RECT 434.8000 91.6000 435.8000 92.4000 ;
	    RECT 436.4000 92.3000 437.2000 93.2000 ;
	    RECT 438.0000 92.3000 438.8000 92.4000 ;
	    RECT 436.4000 91.7000 438.8000 92.3000 ;
	    RECT 436.4000 91.6000 437.2000 91.7000 ;
	    RECT 438.0000 91.6000 438.8000 91.7000 ;
	    RECT 426.8000 91.0000 432.4000 91.2000 ;
	    RECT 426.6000 90.8000 432.4000 91.0000 ;
	    RECT 418.8000 89.8000 421.2000 90.4000 ;
	    RECT 422.6000 90.6000 432.4000 90.8000 ;
	    RECT 422.6000 90.2000 427.4000 90.6000 ;
	    RECT 418.8000 88.8000 419.4000 89.8000 ;
	    RECT 418.0000 88.0000 419.4000 88.8000 ;
	    RECT 421.0000 89.0000 421.8000 89.2000 ;
	    RECT 422.6000 89.0000 423.2000 90.2000 ;
	    RECT 421.0000 88.4000 423.2000 89.0000 ;
	    RECT 423.8000 89.0000 429.2000 89.6000 ;
	    RECT 423.8000 88.8000 424.6000 89.0000 ;
	    RECT 428.4000 88.8000 429.2000 89.0000 ;
	    RECT 422.2000 87.4000 423.0000 87.6000 ;
	    RECT 425.0000 87.4000 425.8000 87.6000 ;
	    RECT 418.8000 86.2000 419.6000 87.0000 ;
	    RECT 422.2000 86.8000 425.8000 87.4000 ;
	    RECT 423.0000 86.2000 423.6000 86.8000 ;
	    RECT 428.4000 86.2000 429.2000 87.0000 ;
	    RECT 418.2000 82.2000 419.4000 86.2000 ;
	    RECT 422.8000 82.2000 423.6000 86.2000 ;
	    RECT 427.2000 85.6000 429.2000 86.2000 ;
	    RECT 427.2000 82.2000 428.0000 85.6000 ;
	    RECT 431.6000 82.2000 432.4000 90.6000 ;
	    RECT 433.2000 90.2000 434.0000 90.4000 ;
	    RECT 435.2000 90.2000 435.8000 91.6000 ;
	    RECT 439.6000 91.4000 440.4000 94.8000 ;
	    RECT 446.6000 94.2000 448.4000 94.4000 ;
	    RECT 452.4000 94.2000 453.0000 96.4000 ;
	    RECT 457.2000 95.0000 458.0000 99.8000 ;
	    RECT 458.8000 95.6000 459.6000 97.2000 ;
	    RECT 455.6000 94.2000 457.2000 94.4000 ;
	    RECT 446.2000 93.6000 457.2000 94.2000 ;
	    RECT 460.4000 94.3000 461.2000 99.8000 ;
	    RECT 462.0000 96.0000 462.8000 99.8000 ;
	    RECT 465.2000 96.0000 466.0000 99.8000 ;
	    RECT 462.0000 95.8000 466.0000 96.0000 ;
	    RECT 466.8000 95.8000 467.6000 99.8000 ;
	    RECT 462.2000 95.4000 465.8000 95.8000 ;
	    RECT 462.8000 94.4000 463.6000 94.8000 ;
	    RECT 466.8000 94.4000 467.4000 95.8000 ;
	    RECT 468.4000 95.4000 469.2000 99.8000 ;
	    RECT 472.6000 98.4000 473.8000 99.8000 ;
	    RECT 472.6000 97.8000 474.0000 98.4000 ;
	    RECT 477.2000 97.8000 478.0000 99.8000 ;
	    RECT 481.6000 98.4000 482.4000 99.8000 ;
	    RECT 481.6000 97.8000 483.6000 98.4000 ;
	    RECT 473.2000 97.0000 474.0000 97.8000 ;
	    RECT 477.4000 97.2000 478.0000 97.8000 ;
	    RECT 477.4000 96.6000 480.2000 97.2000 ;
	    RECT 479.4000 96.4000 480.2000 96.6000 ;
	    RECT 481.2000 96.4000 482.0000 97.2000 ;
	    RECT 482.8000 97.0000 483.6000 97.8000 ;
	    RECT 471.4000 95.4000 472.2000 95.6000 ;
	    RECT 468.4000 94.8000 472.2000 95.4000 ;
	    RECT 462.0000 94.3000 463.6000 94.4000 ;
	    RECT 460.4000 93.8000 463.6000 94.3000 ;
	    RECT 460.4000 93.7000 462.8000 93.8000 ;
	    RECT 444.4000 92.8000 445.2000 93.0000 ;
	    RECT 441.4000 92.2000 445.2000 92.8000 ;
	    RECT 441.4000 92.0000 442.2000 92.2000 ;
	    RECT 443.0000 91.4000 443.8000 91.6000 ;
	    RECT 439.6000 90.8000 443.8000 91.4000 ;
	    RECT 433.2000 89.6000 434.6000 90.2000 ;
	    RECT 435.2000 89.6000 436.2000 90.2000 ;
	    RECT 434.0000 88.4000 434.6000 89.6000 ;
	    RECT 434.0000 87.6000 434.8000 88.4000 ;
	    RECT 435.4000 82.2000 436.2000 89.6000 ;
	    RECT 439.6000 82.2000 440.4000 90.8000 ;
	    RECT 446.2000 90.4000 446.8000 93.6000 ;
	    RECT 453.4000 93.4000 454.2000 93.6000 ;
	    RECT 452.4000 92.4000 453.2000 92.6000 ;
	    RECT 455.0000 92.4000 455.8000 92.6000 ;
	    RECT 450.8000 91.8000 455.8000 92.4000 ;
	    RECT 450.8000 91.6000 451.6000 91.8000 ;
	    RECT 452.4000 91.0000 458.0000 91.2000 ;
	    RECT 452.2000 90.8000 458.0000 91.0000 ;
	    RECT 444.4000 89.8000 446.8000 90.4000 ;
	    RECT 448.2000 90.6000 458.0000 90.8000 ;
	    RECT 448.2000 90.2000 453.0000 90.6000 ;
	    RECT 444.4000 88.8000 445.0000 89.8000 ;
	    RECT 443.6000 88.0000 445.0000 88.8000 ;
	    RECT 446.6000 89.0000 447.4000 89.2000 ;
	    RECT 448.2000 89.0000 448.8000 90.2000 ;
	    RECT 446.6000 88.4000 448.8000 89.0000 ;
	    RECT 449.4000 89.0000 454.8000 89.6000 ;
	    RECT 449.4000 88.8000 450.2000 89.0000 ;
	    RECT 454.0000 88.8000 454.8000 89.0000 ;
	    RECT 447.8000 87.4000 448.6000 87.6000 ;
	    RECT 450.6000 87.4000 451.4000 87.6000 ;
	    RECT 444.4000 86.2000 445.2000 87.0000 ;
	    RECT 447.8000 86.8000 451.4000 87.4000 ;
	    RECT 448.6000 86.2000 449.2000 86.8000 ;
	    RECT 454.0000 86.2000 454.8000 87.0000 ;
	    RECT 443.8000 82.2000 445.0000 86.2000 ;
	    RECT 448.4000 82.2000 449.2000 86.2000 ;
	    RECT 452.8000 85.6000 454.8000 86.2000 ;
	    RECT 452.8000 82.2000 453.6000 85.6000 ;
	    RECT 457.2000 82.2000 458.0000 90.6000 ;
	    RECT 460.4000 82.2000 461.2000 93.7000 ;
	    RECT 462.0000 93.6000 462.8000 93.7000 ;
	    RECT 465.0000 93.6000 467.6000 94.4000 ;
	    RECT 463.6000 91.6000 464.4000 93.2000 ;
	    RECT 465.0000 90.2000 465.6000 93.6000 ;
	    RECT 468.4000 91.4000 469.2000 94.8000 ;
	    RECT 475.4000 94.2000 476.2000 94.4000 ;
	    RECT 481.2000 94.2000 481.8000 96.4000 ;
	    RECT 486.0000 95.0000 486.8000 99.8000 ;
	    RECT 487.6000 95.6000 488.4000 99.8000 ;
	    RECT 489.2000 96.0000 490.0000 99.8000 ;
	    RECT 492.4000 96.0000 493.2000 99.8000 ;
	    RECT 489.2000 95.8000 493.2000 96.0000 ;
	    RECT 487.8000 94.4000 488.4000 95.6000 ;
	    RECT 489.4000 95.4000 493.0000 95.8000 ;
	    RECT 494.0000 95.6000 494.8000 97.2000 ;
	    RECT 491.6000 94.4000 492.4000 94.8000 ;
	    RECT 484.4000 94.2000 486.0000 94.4000 ;
	    RECT 475.0000 93.6000 486.0000 94.2000 ;
	    RECT 487.6000 93.6000 490.2000 94.4000 ;
	    RECT 491.6000 94.3000 493.2000 94.4000 ;
	    RECT 495.6000 94.3000 496.4000 99.8000 ;
	    RECT 491.6000 93.8000 496.4000 94.3000 ;
	    RECT 500.8000 94.2000 501.6000 99.8000 ;
	    RECT 504.8000 94.2000 505.6000 99.8000 ;
	    RECT 500.8000 93.8000 502.6000 94.2000 ;
	    RECT 492.4000 93.7000 496.4000 93.8000 ;
	    RECT 492.4000 93.6000 493.2000 93.7000 ;
	    RECT 473.2000 92.8000 474.0000 93.0000 ;
	    RECT 470.2000 92.2000 474.0000 92.8000 ;
	    RECT 475.0000 92.4000 475.6000 93.6000 ;
	    RECT 482.2000 93.4000 483.0000 93.6000 ;
	    RECT 481.2000 92.4000 482.0000 92.6000 ;
	    RECT 483.8000 92.4000 484.6000 92.6000 ;
	    RECT 470.2000 92.0000 471.0000 92.2000 ;
	    RECT 474.8000 91.6000 475.6000 92.4000 ;
	    RECT 479.6000 91.8000 484.6000 92.4000 ;
	    RECT 479.6000 91.6000 480.4000 91.8000 ;
	    RECT 471.8000 91.4000 472.6000 91.6000 ;
	    RECT 468.4000 90.8000 472.6000 91.4000 ;
	    RECT 466.8000 90.2000 467.6000 90.4000 ;
	    RECT 464.6000 89.6000 465.6000 90.2000 ;
	    RECT 466.2000 89.6000 467.6000 90.2000 ;
	    RECT 464.6000 82.2000 465.4000 89.6000 ;
	    RECT 466.2000 88.4000 466.8000 89.6000 ;
	    RECT 466.0000 87.6000 466.8000 88.4000 ;
	    RECT 468.4000 82.2000 469.2000 90.8000 ;
	    RECT 475.0000 90.4000 475.6000 91.6000 ;
	    RECT 481.2000 91.0000 486.8000 91.2000 ;
	    RECT 481.0000 90.8000 486.8000 91.0000 ;
	    RECT 473.2000 89.8000 475.6000 90.4000 ;
	    RECT 477.0000 90.6000 486.8000 90.8000 ;
	    RECT 477.0000 90.2000 481.8000 90.6000 ;
	    RECT 473.2000 88.8000 473.8000 89.8000 ;
	    RECT 472.4000 88.0000 473.8000 88.8000 ;
	    RECT 475.4000 89.0000 476.2000 89.2000 ;
	    RECT 477.0000 89.0000 477.6000 90.2000 ;
	    RECT 475.4000 88.4000 477.6000 89.0000 ;
	    RECT 478.2000 89.0000 483.6000 89.6000 ;
	    RECT 478.2000 88.8000 479.0000 89.0000 ;
	    RECT 482.8000 88.8000 483.6000 89.0000 ;
	    RECT 476.6000 87.4000 477.4000 87.6000 ;
	    RECT 479.4000 87.4000 480.2000 87.6000 ;
	    RECT 473.2000 86.2000 474.0000 87.0000 ;
	    RECT 476.6000 86.8000 480.2000 87.4000 ;
	    RECT 477.4000 86.2000 478.0000 86.8000 ;
	    RECT 482.8000 86.2000 483.6000 87.0000 ;
	    RECT 472.6000 82.2000 473.8000 86.2000 ;
	    RECT 477.2000 82.2000 478.0000 86.2000 ;
	    RECT 481.6000 85.6000 483.6000 86.2000 ;
	    RECT 481.6000 82.2000 482.4000 85.6000 ;
	    RECT 486.0000 82.2000 486.8000 90.6000 ;
	    RECT 487.6000 90.2000 488.4000 90.4000 ;
	    RECT 489.6000 90.2000 490.2000 93.6000 ;
	    RECT 490.8000 92.3000 491.6000 93.2000 ;
	    RECT 492.4000 92.3000 493.2000 92.4000 ;
	    RECT 490.8000 91.7000 493.2000 92.3000 ;
	    RECT 490.8000 91.6000 491.6000 91.7000 ;
	    RECT 492.4000 91.6000 493.2000 91.7000 ;
	    RECT 487.6000 89.6000 489.0000 90.2000 ;
	    RECT 489.6000 89.6000 490.6000 90.2000 ;
	    RECT 488.4000 88.4000 489.0000 89.6000 ;
	    RECT 488.4000 87.6000 489.2000 88.4000 ;
	    RECT 489.8000 82.2000 490.6000 89.6000 ;
	    RECT 495.6000 82.2000 496.4000 93.7000 ;
	    RECT 501.0000 93.6000 502.6000 93.8000 ;
	    RECT 498.8000 91.6000 500.4000 92.4000 ;
	    RECT 502.0000 90.4000 502.6000 93.6000 ;
	    RECT 503.8000 93.8000 505.6000 94.2000 ;
	    RECT 503.8000 93.6000 505.4000 93.8000 ;
	    RECT 503.8000 90.4000 504.4000 93.6000 ;
	    RECT 506.0000 91.6000 507.6000 92.4000 ;
	    RECT 502.0000 89.6000 502.8000 90.4000 ;
	    RECT 503.6000 89.6000 504.4000 90.4000 ;
	    RECT 500.4000 87.6000 501.2000 89.2000 ;
	    RECT 502.0000 87.0000 502.6000 89.6000 ;
	    RECT 499.0000 86.4000 502.6000 87.0000 ;
	    RECT 498.8000 82.2000 499.6000 86.4000 ;
	    RECT 502.0000 86.2000 502.6000 86.4000 ;
	    RECT 503.8000 87.0000 504.4000 89.6000 ;
	    RECT 505.2000 87.6000 506.0000 89.2000 ;
	    RECT 503.8000 86.4000 507.4000 87.0000 ;
	    RECT 503.8000 86.2000 504.4000 86.4000 ;
	    RECT 502.0000 82.2000 502.8000 86.2000 ;
	    RECT 503.6000 82.2000 504.4000 86.2000 ;
	    RECT 506.8000 86.2000 507.4000 86.4000 ;
	    RECT 506.8000 82.2000 507.6000 86.2000 ;
	    RECT 4.4000 72.4000 5.2000 79.8000 ;
	    RECT 3.0000 71.8000 5.2000 72.4000 ;
	    RECT 6.0000 72.4000 6.8000 79.8000 ;
	    RECT 6.0000 71.8000 8.2000 72.4000 ;
	    RECT 9.2000 71.8000 10.0000 79.8000 ;
	    RECT 10.8000 72.4000 11.6000 79.8000 ;
	    RECT 10.8000 71.8000 13.0000 72.4000 ;
	    RECT 14.0000 71.8000 14.8000 79.8000 ;
	    RECT 3.0000 71.2000 3.6000 71.8000 ;
	    RECT 2.4000 70.4000 3.6000 71.2000 ;
	    RECT 7.6000 71.2000 8.2000 71.8000 ;
	    RECT 7.6000 70.4000 8.8000 71.2000 ;
	    RECT 3.0000 67.4000 3.6000 70.4000 ;
	    RECT 4.4000 68.8000 5.2000 70.4000 ;
	    RECT 7.6000 67.4000 8.2000 70.4000 ;
	    RECT 9.4000 69.6000 10.0000 71.8000 ;
	    RECT 3.0000 66.8000 5.2000 67.4000 ;
	    RECT 4.4000 62.2000 5.2000 66.8000 ;
	    RECT 6.0000 66.8000 8.2000 67.4000 ;
	    RECT 6.0000 62.2000 6.8000 66.8000 ;
	    RECT 9.2000 62.2000 10.0000 69.6000 ;
	    RECT 12.4000 71.2000 13.0000 71.8000 ;
	    RECT 12.4000 70.4000 13.6000 71.2000 ;
	    RECT 12.4000 67.4000 13.0000 70.4000 ;
	    RECT 14.2000 69.6000 14.8000 71.8000 ;
	    RECT 10.8000 66.8000 13.0000 67.4000 ;
	    RECT 10.8000 62.2000 11.6000 66.8000 ;
	    RECT 14.0000 62.2000 14.8000 69.6000 ;
	    RECT 15.6000 71.2000 16.4000 79.8000 ;
	    RECT 19.8000 75.8000 21.0000 79.8000 ;
	    RECT 24.4000 75.8000 25.2000 79.8000 ;
	    RECT 28.8000 76.4000 29.6000 79.8000 ;
	    RECT 28.8000 75.8000 30.8000 76.4000 ;
	    RECT 20.4000 75.0000 21.2000 75.8000 ;
	    RECT 24.6000 75.2000 25.2000 75.8000 ;
	    RECT 23.8000 74.6000 27.4000 75.2000 ;
	    RECT 30.0000 75.0000 30.8000 75.8000 ;
	    RECT 23.8000 74.4000 24.6000 74.6000 ;
	    RECT 26.6000 74.4000 27.4000 74.6000 ;
	    RECT 19.6000 73.2000 21.0000 74.0000 ;
	    RECT 20.4000 72.2000 21.0000 73.2000 ;
	    RECT 22.6000 73.0000 24.8000 73.6000 ;
	    RECT 22.6000 72.8000 23.4000 73.0000 ;
	    RECT 20.4000 71.6000 22.8000 72.2000 ;
	    RECT 15.6000 70.6000 19.8000 71.2000 ;
	    RECT 15.6000 67.2000 16.4000 70.6000 ;
	    RECT 19.0000 70.4000 19.8000 70.6000 ;
	    RECT 17.4000 69.8000 18.2000 70.0000 ;
	    RECT 17.4000 69.2000 21.2000 69.8000 ;
	    RECT 20.4000 69.0000 21.2000 69.2000 ;
	    RECT 22.2000 68.4000 22.8000 71.6000 ;
	    RECT 24.2000 71.8000 24.8000 73.0000 ;
	    RECT 25.4000 73.0000 26.2000 73.2000 ;
	    RECT 30.0000 73.0000 30.8000 73.2000 ;
	    RECT 25.4000 72.4000 30.8000 73.0000 ;
	    RECT 24.2000 71.4000 29.0000 71.8000 ;
	    RECT 33.2000 71.4000 34.0000 79.8000 ;
	    RECT 34.8000 72.4000 35.6000 79.8000 ;
	    RECT 34.8000 71.8000 37.0000 72.4000 ;
	    RECT 38.0000 71.8000 38.8000 79.8000 ;
	    RECT 41.8000 74.4000 42.6000 79.8000 ;
	    RECT 40.4000 73.6000 41.2000 74.4000 ;
	    RECT 41.8000 73.6000 43.6000 74.4000 ;
	    RECT 40.4000 72.4000 41.0000 73.6000 ;
	    RECT 41.8000 72.4000 42.6000 73.6000 ;
	    RECT 24.2000 71.2000 34.0000 71.4000 ;
	    RECT 28.2000 71.0000 34.0000 71.2000 ;
	    RECT 28.4000 70.8000 34.0000 71.0000 ;
	    RECT 36.4000 71.2000 37.0000 71.8000 ;
	    RECT 36.4000 70.4000 37.6000 71.2000 ;
	    RECT 26.8000 70.2000 27.6000 70.4000 ;
	    RECT 26.8000 69.6000 31.8000 70.2000 ;
	    RECT 28.4000 69.4000 29.2000 69.6000 ;
	    RECT 31.0000 69.4000 31.8000 69.6000 ;
	    RECT 34.8000 68.8000 35.6000 70.4000 ;
	    RECT 29.4000 68.4000 30.2000 68.6000 ;
	    RECT 22.2000 67.8000 33.2000 68.4000 ;
	    RECT 22.6000 67.6000 23.4000 67.8000 ;
	    RECT 26.8000 67.6000 27.6000 67.8000 ;
	    RECT 15.6000 66.6000 19.4000 67.2000 ;
	    RECT 15.6000 62.2000 16.4000 66.6000 ;
	    RECT 18.6000 66.4000 19.4000 66.6000 ;
	    RECT 28.4000 65.6000 29.0000 67.8000 ;
	    RECT 31.6000 67.6000 33.2000 67.8000 ;
	    RECT 36.4000 67.4000 37.0000 70.4000 ;
	    RECT 38.2000 69.6000 38.8000 71.8000 ;
	    RECT 39.6000 71.8000 41.0000 72.4000 ;
	    RECT 41.6000 71.8000 42.6000 72.4000 ;
	    RECT 46.0000 72.4000 46.8000 79.8000 ;
	    RECT 46.0000 71.8000 48.2000 72.4000 ;
	    RECT 49.2000 71.8000 50.0000 79.8000 ;
	    RECT 51.6000 73.6000 52.4000 74.4000 ;
	    RECT 51.6000 72.4000 52.2000 73.6000 ;
	    RECT 53.0000 72.4000 53.8000 79.8000 ;
	    RECT 39.6000 71.6000 40.4000 71.8000 ;
	    RECT 26.6000 65.4000 27.4000 65.6000 ;
	    RECT 20.4000 64.2000 21.2000 65.0000 ;
	    RECT 24.6000 64.8000 27.4000 65.4000 ;
	    RECT 28.4000 64.8000 29.2000 65.6000 ;
	    RECT 24.6000 64.2000 25.2000 64.8000 ;
	    RECT 30.0000 64.2000 30.8000 65.0000 ;
	    RECT 19.8000 63.6000 21.2000 64.2000 ;
	    RECT 19.8000 62.2000 21.0000 63.6000 ;
	    RECT 24.4000 62.2000 25.2000 64.2000 ;
	    RECT 28.8000 63.6000 30.8000 64.2000 ;
	    RECT 28.8000 62.2000 29.6000 63.6000 ;
	    RECT 33.2000 62.2000 34.0000 67.0000 ;
	    RECT 34.8000 66.8000 37.0000 67.4000 ;
	    RECT 34.8000 62.2000 35.6000 66.8000 ;
	    RECT 38.0000 62.2000 38.8000 69.6000 ;
	    RECT 41.6000 68.4000 42.2000 71.8000 ;
	    RECT 47.6000 71.2000 48.2000 71.8000 ;
	    RECT 47.6000 70.4000 48.8000 71.2000 ;
	    RECT 42.8000 68.8000 43.6000 70.4000 ;
	    RECT 46.0000 68.8000 46.8000 70.4000 ;
	    RECT 39.6000 67.6000 42.2000 68.4000 ;
	    RECT 44.4000 68.2000 45.2000 68.4000 ;
	    RECT 43.6000 67.6000 45.2000 68.2000 ;
	    RECT 39.8000 66.2000 40.4000 67.6000 ;
	    RECT 43.6000 67.2000 44.4000 67.6000 ;
	    RECT 47.6000 67.4000 48.2000 70.4000 ;
	    RECT 49.4000 69.6000 50.0000 71.8000 ;
	    RECT 50.8000 71.8000 52.2000 72.4000 ;
	    RECT 52.8000 71.8000 53.8000 72.4000 ;
	    RECT 50.8000 71.6000 51.6000 71.8000 ;
	    RECT 52.8000 70.4000 53.4000 71.8000 ;
	    RECT 58.8000 71.2000 59.6000 79.8000 ;
	    RECT 62.0000 71.2000 62.8000 79.8000 ;
	    RECT 65.2000 71.2000 66.0000 79.8000 ;
	    RECT 68.4000 71.2000 69.2000 79.8000 ;
	    RECT 73.8000 78.4000 74.6000 79.8000 ;
	    RECT 73.8000 77.6000 75.6000 78.4000 ;
	    RECT 72.4000 73.6000 73.2000 74.4000 ;
	    RECT 72.4000 72.4000 73.0000 73.6000 ;
	    RECT 73.8000 72.4000 74.6000 77.6000 ;
	    RECT 71.6000 71.8000 73.0000 72.4000 ;
	    RECT 73.6000 71.8000 74.6000 72.4000 ;
	    RECT 78.0000 72.4000 78.8000 79.8000 ;
	    RECT 78.0000 71.8000 80.2000 72.4000 ;
	    RECT 81.2000 71.8000 82.0000 79.8000 ;
	    RECT 71.6000 71.6000 72.4000 71.8000 ;
	    RECT 58.8000 70.4000 60.6000 71.2000 ;
	    RECT 62.0000 70.4000 64.2000 71.2000 ;
	    RECT 65.2000 70.4000 67.4000 71.2000 ;
	    RECT 68.4000 70.4000 70.8000 71.2000 ;
	    RECT 52.4000 69.6000 53.4000 70.4000 ;
	    RECT 46.0000 66.8000 48.2000 67.4000 ;
	    RECT 41.4000 66.2000 45.0000 66.6000 ;
	    RECT 39.6000 62.2000 40.4000 66.2000 ;
	    RECT 41.2000 66.0000 45.2000 66.2000 ;
	    RECT 41.2000 62.2000 42.0000 66.0000 ;
	    RECT 44.4000 62.2000 45.2000 66.0000 ;
	    RECT 46.0000 62.2000 46.8000 66.8000 ;
	    RECT 49.2000 62.2000 50.0000 69.6000 ;
	    RECT 52.8000 68.4000 53.4000 69.6000 ;
	    RECT 54.0000 70.3000 54.8000 70.4000 ;
	    RECT 57.2000 70.3000 58.0000 70.4000 ;
	    RECT 54.0000 69.7000 58.0000 70.3000 ;
	    RECT 54.0000 68.8000 54.8000 69.7000 ;
	    RECT 57.2000 69.6000 58.0000 69.7000 ;
	    RECT 59.8000 69.0000 60.6000 70.4000 ;
	    RECT 63.4000 69.0000 64.2000 70.4000 ;
	    RECT 66.6000 69.0000 67.4000 70.4000 ;
	    RECT 50.8000 67.6000 53.4000 68.4000 ;
	    RECT 55.6000 68.2000 56.4000 68.4000 ;
	    RECT 54.8000 67.6000 56.4000 68.2000 ;
	    RECT 59.8000 68.2000 62.4000 69.0000 ;
	    RECT 63.4000 68.2000 65.8000 69.0000 ;
	    RECT 66.6000 68.2000 69.2000 69.0000 ;
	    RECT 59.8000 67.6000 60.6000 68.2000 ;
	    RECT 63.4000 67.6000 64.2000 68.2000 ;
	    RECT 66.6000 67.6000 67.4000 68.2000 ;
	    RECT 70.0000 67.6000 70.8000 70.4000 ;
	    RECT 73.6000 68.4000 74.2000 71.8000 ;
	    RECT 79.6000 71.2000 80.2000 71.8000 ;
	    RECT 79.6000 70.4000 80.8000 71.2000 ;
	    RECT 74.8000 68.8000 75.6000 70.4000 ;
	    RECT 71.6000 67.6000 74.2000 68.4000 ;
	    RECT 76.4000 68.2000 77.2000 68.4000 ;
	    RECT 75.6000 67.6000 77.2000 68.2000 ;
	    RECT 51.0000 66.2000 51.6000 67.6000 ;
	    RECT 54.8000 67.2000 55.6000 67.6000 ;
	    RECT 58.8000 66.8000 60.6000 67.6000 ;
	    RECT 62.0000 66.8000 64.2000 67.6000 ;
	    RECT 65.2000 66.8000 67.4000 67.6000 ;
	    RECT 68.4000 66.8000 70.8000 67.6000 ;
	    RECT 52.6000 66.2000 56.2000 66.6000 ;
	    RECT 50.8000 62.2000 51.6000 66.2000 ;
	    RECT 52.4000 66.0000 56.4000 66.2000 ;
	    RECT 52.4000 62.2000 53.2000 66.0000 ;
	    RECT 55.6000 62.2000 56.4000 66.0000 ;
	    RECT 58.8000 62.2000 59.6000 66.8000 ;
	    RECT 62.0000 62.2000 62.8000 66.8000 ;
	    RECT 65.2000 62.2000 66.0000 66.8000 ;
	    RECT 68.4000 62.2000 69.2000 66.8000 ;
	    RECT 71.8000 66.2000 72.4000 67.6000 ;
	    RECT 75.6000 67.2000 76.4000 67.6000 ;
	    RECT 79.6000 67.4000 80.2000 70.4000 ;
	    RECT 81.4000 69.6000 82.0000 71.8000 ;
	    RECT 82.8000 71.4000 83.6000 79.8000 ;
	    RECT 87.2000 76.4000 88.0000 79.8000 ;
	    RECT 86.0000 75.8000 88.0000 76.4000 ;
	    RECT 91.6000 75.8000 92.4000 79.8000 ;
	    RECT 95.8000 75.8000 97.0000 79.8000 ;
	    RECT 86.0000 75.0000 86.8000 75.8000 ;
	    RECT 91.6000 75.2000 92.2000 75.8000 ;
	    RECT 89.4000 74.6000 93.0000 75.2000 ;
	    RECT 95.6000 75.0000 96.4000 75.8000 ;
	    RECT 89.4000 74.4000 90.2000 74.6000 ;
	    RECT 92.2000 74.4000 93.0000 74.6000 ;
	    RECT 86.0000 73.0000 86.8000 73.2000 ;
	    RECT 90.6000 73.0000 91.4000 73.2000 ;
	    RECT 86.0000 72.4000 91.4000 73.0000 ;
	    RECT 92.0000 73.0000 94.2000 73.6000 ;
	    RECT 92.0000 71.8000 92.6000 73.0000 ;
	    RECT 93.4000 72.8000 94.2000 73.0000 ;
	    RECT 95.8000 73.2000 97.2000 74.0000 ;
	    RECT 95.8000 72.2000 96.4000 73.2000 ;
	    RECT 87.8000 71.4000 92.6000 71.8000 ;
	    RECT 82.8000 71.2000 92.6000 71.4000 ;
	    RECT 94.0000 71.6000 96.4000 72.2000 ;
	    RECT 82.8000 71.0000 88.6000 71.2000 ;
	    RECT 82.8000 70.8000 88.4000 71.0000 ;
	    RECT 89.2000 70.3000 90.0000 70.4000 ;
	    RECT 92.4000 70.3000 93.2000 70.4000 ;
	    RECT 89.2000 70.2000 93.2000 70.3000 ;
	    RECT 78.0000 66.8000 80.2000 67.4000 ;
	    RECT 73.4000 66.2000 77.0000 66.6000 ;
	    RECT 71.6000 62.2000 72.4000 66.2000 ;
	    RECT 73.2000 66.0000 77.2000 66.2000 ;
	    RECT 73.2000 62.2000 74.0000 66.0000 ;
	    RECT 76.4000 62.2000 77.2000 66.0000 ;
	    RECT 78.0000 62.2000 78.8000 66.8000 ;
	    RECT 81.2000 62.2000 82.0000 69.6000 ;
	    RECT 85.0000 69.7000 93.2000 70.2000 ;
	    RECT 85.0000 69.6000 90.0000 69.7000 ;
	    RECT 92.4000 69.6000 93.2000 69.7000 ;
	    RECT 85.0000 69.4000 85.8000 69.6000 ;
	    RECT 86.6000 68.4000 87.4000 68.6000 ;
	    RECT 94.0000 68.4000 94.6000 71.6000 ;
	    RECT 100.4000 71.2000 101.2000 79.8000 ;
	    RECT 104.6000 72.4000 105.4000 79.8000 ;
	    RECT 106.0000 73.6000 106.8000 74.4000 ;
	    RECT 106.2000 72.4000 106.8000 73.6000 ;
	    RECT 104.6000 71.8000 105.6000 72.4000 ;
	    RECT 106.2000 71.8000 107.6000 72.4000 ;
	    RECT 97.0000 70.6000 101.2000 71.2000 ;
	    RECT 97.0000 70.4000 97.8000 70.6000 ;
	    RECT 98.6000 69.8000 99.4000 70.0000 ;
	    RECT 95.6000 69.2000 99.4000 69.8000 ;
	    RECT 95.6000 69.0000 96.4000 69.2000 ;
	    RECT 83.6000 67.8000 94.6000 68.4000 ;
	    RECT 83.6000 67.6000 85.2000 67.8000 ;
	    RECT 87.6000 67.6000 88.4000 67.8000 ;
	    RECT 93.4000 67.6000 94.2000 67.8000 ;
	    RECT 82.8000 62.2000 83.6000 67.0000 ;
	    RECT 87.8000 65.6000 88.4000 67.6000 ;
	    RECT 100.4000 67.2000 101.2000 70.6000 ;
	    RECT 105.0000 70.4000 105.6000 71.8000 ;
	    RECT 106.8000 71.6000 107.6000 71.8000 ;
	    RECT 113.2000 72.3000 114.0000 72.4000 ;
	    RECT 114.8000 72.3000 115.6000 73.2000 ;
	    RECT 113.2000 71.7000 115.6000 72.3000 ;
	    RECT 113.2000 71.6000 114.0000 71.7000 ;
	    RECT 114.8000 71.6000 115.6000 71.7000 ;
	    RECT 103.6000 68.8000 104.4000 70.4000 ;
	    RECT 105.0000 69.6000 106.0000 70.4000 ;
	    RECT 106.9000 70.3000 107.5000 71.6000 ;
	    RECT 116.4000 70.3000 117.2000 79.8000 ;
	    RECT 119.6000 72.4000 120.4000 79.8000 ;
	    RECT 119.6000 71.8000 121.8000 72.4000 ;
	    RECT 122.8000 71.8000 123.6000 79.8000 ;
	    RECT 106.9000 69.7000 117.2000 70.3000 ;
	    RECT 105.0000 68.4000 105.6000 69.6000 ;
	    RECT 102.0000 68.2000 102.8000 68.4000 ;
	    RECT 102.0000 67.6000 103.6000 68.2000 ;
	    RECT 105.0000 67.6000 107.6000 68.4000 ;
	    RECT 102.8000 67.2000 103.6000 67.6000 ;
	    RECT 97.4000 66.6000 101.2000 67.2000 ;
	    RECT 97.4000 66.4000 98.2000 66.6000 ;
	    RECT 86.0000 64.2000 86.8000 65.0000 ;
	    RECT 87.6000 64.8000 88.4000 65.6000 ;
	    RECT 89.4000 65.4000 90.2000 65.6000 ;
	    RECT 89.4000 64.8000 92.2000 65.4000 ;
	    RECT 91.6000 64.2000 92.2000 64.8000 ;
	    RECT 95.6000 64.2000 96.4000 65.0000 ;
	    RECT 86.0000 63.6000 88.0000 64.2000 ;
	    RECT 87.2000 62.2000 88.0000 63.6000 ;
	    RECT 91.6000 62.2000 92.4000 64.2000 ;
	    RECT 95.6000 63.6000 97.0000 64.2000 ;
	    RECT 95.8000 62.2000 97.0000 63.6000 ;
	    RECT 100.4000 62.2000 101.2000 66.6000 ;
	    RECT 102.2000 66.2000 105.8000 66.6000 ;
	    RECT 106.8000 66.2000 107.4000 67.6000 ;
	    RECT 116.4000 66.2000 117.2000 69.7000 ;
	    RECT 121.2000 71.2000 121.8000 71.8000 ;
	    RECT 121.2000 70.4000 122.4000 71.2000 ;
	    RECT 118.0000 66.8000 118.8000 68.4000 ;
	    RECT 121.2000 67.4000 121.8000 70.4000 ;
	    RECT 123.0000 69.6000 123.6000 71.8000 ;
	    RECT 124.4000 75.0000 125.2000 79.0000 ;
	    RECT 128.6000 78.4000 129.4000 79.8000 ;
	    RECT 128.6000 77.6000 130.0000 78.4000 ;
	    RECT 124.4000 71.6000 125.0000 75.0000 ;
	    RECT 128.6000 72.8000 129.4000 77.6000 ;
	    RECT 134.0000 75.0000 134.8000 79.0000 ;
	    RECT 138.2000 78.4000 139.0000 79.8000 ;
	    RECT 138.2000 77.6000 139.6000 78.4000 ;
	    RECT 128.6000 72.2000 130.2000 72.8000 ;
	    RECT 124.4000 71.0000 128.2000 71.6000 ;
	    RECT 119.6000 66.8000 121.8000 67.4000 ;
	    RECT 102.0000 66.0000 106.0000 66.2000 ;
	    RECT 102.0000 62.2000 102.8000 66.0000 ;
	    RECT 105.2000 62.2000 106.0000 66.0000 ;
	    RECT 106.8000 62.2000 107.6000 66.2000 ;
	    RECT 115.4000 65.6000 117.2000 66.2000 ;
	    RECT 115.4000 62.2000 116.2000 65.6000 ;
	    RECT 119.6000 62.2000 120.4000 66.8000 ;
	    RECT 122.8000 62.2000 123.6000 69.6000 ;
	    RECT 124.4000 68.8000 125.2000 70.4000 ;
	    RECT 126.0000 68.8000 126.8000 70.4000 ;
	    RECT 127.6000 69.0000 128.2000 71.0000 ;
	    RECT 127.6000 68.2000 129.0000 69.0000 ;
	    RECT 129.6000 68.4000 130.2000 72.2000 ;
	    RECT 134.0000 71.6000 134.6000 75.0000 ;
	    RECT 138.2000 72.8000 139.0000 77.6000 ;
	    RECT 138.2000 72.2000 139.8000 72.8000 ;
	    RECT 130.8000 69.6000 131.6000 71.2000 ;
	    RECT 134.0000 71.0000 137.8000 71.6000 ;
	    RECT 134.0000 68.8000 134.8000 70.4000 ;
	    RECT 135.6000 68.8000 136.4000 70.4000 ;
	    RECT 137.2000 69.0000 137.8000 71.0000 ;
	    RECT 127.6000 67.8000 128.6000 68.2000 ;
	    RECT 124.4000 67.2000 128.6000 67.8000 ;
	    RECT 129.6000 67.6000 131.6000 68.4000 ;
	    RECT 137.2000 68.2000 138.6000 69.0000 ;
	    RECT 139.2000 68.4000 139.8000 72.2000 ;
	    RECT 140.4000 69.6000 141.2000 71.2000 ;
	    RECT 145.2000 70.3000 146.0000 79.8000 ;
	    RECT 149.2000 73.6000 150.0000 74.4000 ;
	    RECT 146.8000 71.6000 147.6000 73.2000 ;
	    RECT 149.2000 72.4000 149.8000 73.6000 ;
	    RECT 150.6000 72.4000 151.4000 79.8000 ;
	    RECT 148.4000 71.8000 149.8000 72.4000 ;
	    RECT 150.4000 71.8000 151.4000 72.4000 ;
	    RECT 154.8000 72.4000 155.6000 79.8000 ;
	    RECT 154.8000 71.8000 157.0000 72.4000 ;
	    RECT 158.0000 71.8000 158.8000 79.8000 ;
	    RECT 160.4000 73.6000 161.2000 74.4000 ;
	    RECT 160.4000 72.4000 161.0000 73.6000 ;
	    RECT 161.8000 72.4000 162.6000 79.8000 ;
	    RECT 166.8000 73.6000 167.6000 74.4000 ;
	    RECT 166.8000 72.4000 167.4000 73.6000 ;
	    RECT 168.2000 72.4000 169.0000 79.8000 ;
	    RECT 175.0000 76.4000 175.8000 79.8000 ;
	    RECT 174.0000 75.6000 175.8000 76.4000 ;
	    RECT 148.4000 71.6000 149.2000 71.8000 ;
	    RECT 148.5000 70.3000 149.1000 71.6000 ;
	    RECT 145.2000 69.7000 149.1000 70.3000 ;
	    RECT 137.2000 67.8000 138.2000 68.2000 ;
	    RECT 124.4000 65.0000 125.0000 67.2000 ;
	    RECT 129.6000 67.0000 130.2000 67.6000 ;
	    RECT 129.4000 66.6000 130.2000 67.0000 ;
	    RECT 128.6000 66.0000 130.2000 66.6000 ;
	    RECT 134.0000 67.2000 138.2000 67.8000 ;
	    RECT 139.2000 67.6000 141.2000 68.4000 ;
	    RECT 142.0000 68.3000 142.8000 68.4000 ;
	    RECT 143.6000 68.3000 144.4000 68.4000 ;
	    RECT 142.0000 67.7000 144.4000 68.3000 ;
	    RECT 142.0000 67.6000 142.8000 67.7000 ;
	    RECT 124.4000 63.0000 125.2000 65.0000 ;
	    RECT 128.6000 63.0000 129.4000 66.0000 ;
	    RECT 134.0000 65.0000 134.6000 67.2000 ;
	    RECT 139.2000 67.0000 139.8000 67.6000 ;
	    RECT 139.0000 66.6000 139.8000 67.0000 ;
	    RECT 143.6000 66.8000 144.4000 67.7000 ;
	    RECT 138.2000 66.0000 139.8000 66.6000 ;
	    RECT 145.2000 66.2000 146.0000 69.7000 ;
	    RECT 150.4000 68.4000 151.0000 71.8000 ;
	    RECT 156.4000 71.2000 157.0000 71.8000 ;
	    RECT 156.4000 70.4000 157.6000 71.2000 ;
	    RECT 151.6000 68.8000 152.4000 70.4000 ;
	    RECT 154.8000 68.8000 155.6000 70.4000 ;
	    RECT 148.4000 67.6000 151.0000 68.4000 ;
	    RECT 153.2000 68.2000 154.0000 68.4000 ;
	    RECT 152.4000 67.6000 154.0000 68.2000 ;
	    RECT 148.6000 66.2000 149.2000 67.6000 ;
	    RECT 152.4000 67.2000 153.2000 67.6000 ;
	    RECT 156.4000 67.4000 157.0000 70.4000 ;
	    RECT 158.2000 69.6000 158.8000 71.8000 ;
	    RECT 159.6000 71.8000 161.0000 72.4000 ;
	    RECT 161.6000 71.8000 162.6000 72.4000 ;
	    RECT 166.0000 71.8000 167.4000 72.4000 ;
	    RECT 168.0000 71.8000 169.0000 72.4000 ;
	    RECT 175.0000 72.4000 175.8000 75.6000 ;
	    RECT 176.4000 73.6000 177.2000 74.4000 ;
	    RECT 176.6000 72.4000 177.2000 73.6000 ;
	    RECT 179.6000 73.6000 180.4000 74.4000 ;
	    RECT 179.6000 72.4000 180.2000 73.6000 ;
	    RECT 181.0000 72.4000 181.8000 79.8000 ;
	    RECT 175.0000 71.8000 176.0000 72.4000 ;
	    RECT 176.6000 72.3000 178.0000 72.4000 ;
	    RECT 178.8000 72.3000 180.2000 72.4000 ;
	    RECT 176.6000 71.8000 180.2000 72.3000 ;
	    RECT 180.8000 71.8000 181.8000 72.4000 ;
	    RECT 159.6000 71.6000 160.4000 71.8000 ;
	    RECT 154.8000 66.8000 157.0000 67.4000 ;
	    RECT 150.2000 66.2000 153.8000 66.6000 ;
	    RECT 134.0000 63.0000 134.8000 65.0000 ;
	    RECT 138.2000 63.0000 139.0000 66.0000 ;
	    RECT 145.2000 65.6000 147.0000 66.2000 ;
	    RECT 146.2000 62.2000 147.0000 65.6000 ;
	    RECT 148.4000 62.2000 149.2000 66.2000 ;
	    RECT 150.0000 66.0000 154.0000 66.2000 ;
	    RECT 150.0000 62.2000 150.8000 66.0000 ;
	    RECT 153.2000 62.2000 154.0000 66.0000 ;
	    RECT 154.8000 62.2000 155.6000 66.8000 ;
	    RECT 158.0000 62.2000 158.8000 69.6000 ;
	    RECT 161.6000 68.4000 162.2000 71.8000 ;
	    RECT 166.0000 71.6000 166.8000 71.8000 ;
	    RECT 162.8000 68.8000 163.6000 70.4000 ;
	    RECT 168.0000 68.4000 168.6000 71.8000 ;
	    RECT 169.2000 68.8000 170.0000 70.4000 ;
	    RECT 174.0000 68.8000 174.8000 70.4000 ;
	    RECT 175.4000 68.4000 176.0000 71.8000 ;
	    RECT 177.2000 71.7000 179.6000 71.8000 ;
	    RECT 177.2000 71.6000 178.0000 71.7000 ;
	    RECT 178.8000 71.6000 179.6000 71.7000 ;
	    RECT 178.8000 70.3000 179.6000 70.4000 ;
	    RECT 180.8000 70.3000 181.4000 71.8000 ;
	    RECT 185.2000 71.2000 186.0000 79.8000 ;
	    RECT 189.4000 75.8000 190.6000 79.8000 ;
	    RECT 194.0000 75.8000 194.8000 79.8000 ;
	    RECT 198.4000 76.4000 199.2000 79.8000 ;
	    RECT 198.4000 75.8000 200.4000 76.4000 ;
	    RECT 190.0000 75.0000 190.8000 75.8000 ;
	    RECT 194.2000 75.2000 194.8000 75.8000 ;
	    RECT 193.4000 74.6000 197.0000 75.2000 ;
	    RECT 199.6000 75.0000 200.4000 75.8000 ;
	    RECT 193.4000 74.4000 194.2000 74.6000 ;
	    RECT 196.2000 74.4000 197.0000 74.6000 ;
	    RECT 189.2000 73.2000 190.6000 74.0000 ;
	    RECT 190.0000 72.2000 190.6000 73.2000 ;
	    RECT 192.2000 73.0000 194.4000 73.6000 ;
	    RECT 192.2000 72.8000 193.0000 73.0000 ;
	    RECT 190.0000 71.6000 192.4000 72.2000 ;
	    RECT 185.2000 70.6000 189.4000 71.2000 ;
	    RECT 178.8000 69.7000 181.4000 70.3000 ;
	    RECT 178.8000 69.6000 179.6000 69.7000 ;
	    RECT 180.8000 68.4000 181.4000 69.7000 ;
	    RECT 182.0000 68.8000 182.8000 70.4000 ;
	    RECT 159.6000 67.6000 162.2000 68.4000 ;
	    RECT 164.4000 68.2000 165.2000 68.4000 ;
	    RECT 163.6000 67.6000 165.2000 68.2000 ;
	    RECT 166.0000 67.6000 168.6000 68.4000 ;
	    RECT 170.8000 68.2000 171.6000 68.4000 ;
	    RECT 170.0000 67.6000 171.6000 68.2000 ;
	    RECT 172.4000 68.2000 173.2000 68.4000 ;
	    RECT 172.4000 67.6000 174.0000 68.2000 ;
	    RECT 175.4000 67.6000 178.0000 68.4000 ;
	    RECT 178.8000 67.6000 181.4000 68.4000 ;
	    RECT 183.6000 68.2000 184.4000 68.4000 ;
	    RECT 182.8000 67.6000 184.4000 68.2000 ;
	    RECT 159.8000 66.2000 160.4000 67.6000 ;
	    RECT 163.6000 67.2000 164.4000 67.6000 ;
	    RECT 161.4000 66.2000 165.0000 66.6000 ;
	    RECT 166.2000 66.2000 166.8000 67.6000 ;
	    RECT 170.0000 67.2000 170.8000 67.6000 ;
	    RECT 173.2000 67.2000 174.0000 67.6000 ;
	    RECT 167.8000 66.2000 171.4000 66.6000 ;
	    RECT 172.6000 66.2000 176.2000 66.6000 ;
	    RECT 177.2000 66.2000 177.8000 67.6000 ;
	    RECT 179.0000 66.2000 179.6000 67.6000 ;
	    RECT 182.8000 67.2000 183.6000 67.6000 ;
	    RECT 185.2000 67.2000 186.0000 70.6000 ;
	    RECT 188.6000 70.4000 189.4000 70.6000 ;
	    RECT 187.0000 69.8000 187.8000 70.0000 ;
	    RECT 187.0000 69.2000 190.8000 69.8000 ;
	    RECT 190.0000 69.0000 190.8000 69.2000 ;
	    RECT 191.8000 68.4000 192.4000 71.6000 ;
	    RECT 193.8000 71.8000 194.4000 73.0000 ;
	    RECT 195.0000 73.0000 195.8000 73.2000 ;
	    RECT 199.6000 73.0000 200.4000 73.2000 ;
	    RECT 195.0000 72.4000 200.4000 73.0000 ;
	    RECT 193.8000 71.4000 198.6000 71.8000 ;
	    RECT 202.8000 71.4000 203.6000 79.8000 ;
	    RECT 205.2000 73.6000 206.0000 74.4000 ;
	    RECT 205.2000 72.4000 205.8000 73.6000 ;
	    RECT 206.6000 72.4000 207.4000 79.8000 ;
	    RECT 204.4000 71.8000 205.8000 72.4000 ;
	    RECT 206.4000 71.8000 207.4000 72.4000 ;
	    RECT 210.8000 72.4000 211.6000 79.8000 ;
	    RECT 210.8000 71.8000 213.0000 72.4000 ;
	    RECT 214.0000 71.8000 214.8000 79.8000 ;
	    RECT 218.2000 71.8000 220.2000 79.8000 ;
	    RECT 224.4000 73.6000 225.2000 74.4000 ;
	    RECT 224.4000 72.4000 225.0000 73.6000 ;
	    RECT 225.8000 72.4000 226.6000 79.8000 ;
	    RECT 232.6000 72.6000 233.4000 79.8000 ;
	    RECT 237.4000 76.4000 239.4000 79.8000 ;
	    RECT 236.4000 75.6000 239.4000 76.4000 ;
	    RECT 223.6000 71.8000 225.0000 72.4000 ;
	    RECT 225.6000 71.8000 226.6000 72.4000 ;
	    RECT 231.6000 71.8000 233.4000 72.6000 ;
	    RECT 237.4000 71.8000 239.4000 75.6000 ;
	    RECT 245.4000 72.4000 246.2000 79.8000 ;
	    RECT 246.8000 73.6000 247.6000 74.4000 ;
	    RECT 247.0000 72.4000 247.6000 73.6000 ;
	    RECT 250.0000 73.6000 250.8000 74.4000 ;
	    RECT 250.0000 72.4000 250.6000 73.6000 ;
	    RECT 251.4000 72.4000 252.2000 79.8000 ;
	    RECT 245.4000 71.8000 246.4000 72.4000 ;
	    RECT 247.0000 71.8000 248.4000 72.4000 ;
	    RECT 204.4000 71.6000 205.2000 71.8000 ;
	    RECT 193.8000 71.2000 203.6000 71.4000 ;
	    RECT 197.8000 71.0000 203.6000 71.2000 ;
	    RECT 198.0000 70.8000 203.6000 71.0000 ;
	    RECT 206.4000 70.4000 207.0000 71.8000 ;
	    RECT 212.4000 71.2000 213.0000 71.8000 ;
	    RECT 212.4000 70.4000 213.6000 71.2000 ;
	    RECT 196.4000 70.2000 197.2000 70.4000 ;
	    RECT 196.4000 69.6000 201.4000 70.2000 ;
	    RECT 206.0000 69.6000 207.0000 70.4000 ;
	    RECT 198.0000 69.4000 198.8000 69.6000 ;
	    RECT 200.6000 69.4000 201.4000 69.6000 ;
	    RECT 199.0000 68.4000 199.8000 68.6000 ;
	    RECT 206.4000 68.4000 207.0000 69.6000 ;
	    RECT 207.6000 68.8000 208.4000 70.4000 ;
	    RECT 191.8000 67.8000 202.8000 68.4000 ;
	    RECT 192.2000 67.6000 193.0000 67.8000 ;
	    RECT 185.2000 66.6000 189.0000 67.2000 ;
	    RECT 180.6000 66.2000 184.2000 66.6000 ;
	    RECT 159.6000 62.2000 160.4000 66.2000 ;
	    RECT 161.2000 66.0000 165.2000 66.2000 ;
	    RECT 161.2000 62.2000 162.0000 66.0000 ;
	    RECT 164.4000 62.2000 165.2000 66.0000 ;
	    RECT 166.0000 62.2000 166.8000 66.2000 ;
	    RECT 167.6000 66.0000 171.6000 66.2000 ;
	    RECT 167.6000 62.2000 168.4000 66.0000 ;
	    RECT 170.8000 62.2000 171.6000 66.0000 ;
	    RECT 172.4000 66.0000 176.4000 66.2000 ;
	    RECT 172.4000 62.2000 173.2000 66.0000 ;
	    RECT 175.6000 62.2000 176.4000 66.0000 ;
	    RECT 177.2000 62.2000 178.0000 66.2000 ;
	    RECT 178.8000 62.2000 179.6000 66.2000 ;
	    RECT 180.4000 66.0000 184.4000 66.2000 ;
	    RECT 180.4000 62.2000 181.2000 66.0000 ;
	    RECT 183.6000 62.2000 184.4000 66.0000 ;
	    RECT 185.2000 62.2000 186.0000 66.6000 ;
	    RECT 188.2000 66.4000 189.0000 66.6000 ;
	    RECT 198.0000 65.6000 198.6000 67.8000 ;
	    RECT 201.2000 67.6000 202.8000 67.8000 ;
	    RECT 204.4000 67.6000 207.0000 68.4000 ;
	    RECT 209.2000 68.2000 210.0000 68.4000 ;
	    RECT 208.4000 67.6000 210.0000 68.2000 ;
	    RECT 196.2000 65.4000 197.0000 65.6000 ;
	    RECT 190.0000 64.2000 190.8000 65.0000 ;
	    RECT 194.2000 64.8000 197.0000 65.4000 ;
	    RECT 198.0000 64.8000 198.8000 65.6000 ;
	    RECT 194.2000 64.2000 194.8000 64.8000 ;
	    RECT 199.6000 64.2000 200.4000 65.0000 ;
	    RECT 189.4000 63.6000 190.8000 64.2000 ;
	    RECT 189.4000 62.2000 190.6000 63.6000 ;
	    RECT 194.0000 62.2000 194.8000 64.2000 ;
	    RECT 198.4000 63.6000 200.4000 64.2000 ;
	    RECT 198.4000 62.2000 199.2000 63.6000 ;
	    RECT 202.8000 62.2000 203.6000 67.0000 ;
	    RECT 204.6000 66.2000 205.2000 67.6000 ;
	    RECT 208.4000 67.2000 209.2000 67.6000 ;
	    RECT 212.4000 67.4000 213.0000 70.4000 ;
	    RECT 214.2000 69.6000 214.8000 71.8000 ;
	    RECT 210.8000 66.8000 213.0000 67.4000 ;
	    RECT 214.0000 68.3000 214.8000 69.6000 ;
	    RECT 215.6000 68.3000 216.4000 70.4000 ;
	    RECT 217.2000 68.8000 218.0000 70.4000 ;
	    RECT 219.0000 68.4000 219.6000 71.8000 ;
	    RECT 223.6000 71.6000 224.4000 71.8000 ;
	    RECT 220.4000 70.3000 221.2000 70.4000 ;
	    RECT 223.6000 70.3000 224.4000 70.4000 ;
	    RECT 220.4000 69.7000 224.4000 70.3000 ;
	    RECT 220.4000 68.8000 221.2000 69.7000 ;
	    RECT 223.6000 69.6000 224.4000 69.7000 ;
	    RECT 225.6000 68.4000 226.2000 71.8000 ;
	    RECT 226.8000 68.8000 227.6000 70.4000 ;
	    RECT 228.4000 70.3000 229.2000 70.4000 ;
	    RECT 231.8000 70.3000 232.4000 71.8000 ;
	    RECT 228.4000 69.7000 232.4000 70.3000 ;
	    RECT 228.4000 69.6000 229.2000 69.7000 ;
	    RECT 231.8000 68.4000 232.4000 69.7000 ;
	    RECT 233.2000 69.6000 234.0000 71.2000 ;
	    RECT 214.0000 67.7000 216.4000 68.3000 ;
	    RECT 218.8000 68.2000 219.6000 68.4000 ;
	    RECT 222.0000 68.3000 222.8000 68.4000 ;
	    RECT 223.6000 68.3000 226.2000 68.4000 ;
	    RECT 222.0000 68.2000 226.2000 68.3000 ;
	    RECT 228.4000 68.3000 229.2000 68.4000 ;
	    RECT 230.0000 68.3000 230.8000 68.4000 ;
	    RECT 228.4000 68.2000 230.8000 68.3000 ;
	    RECT 206.2000 66.2000 209.8000 66.6000 ;
	    RECT 204.4000 62.2000 205.2000 66.2000 ;
	    RECT 206.0000 66.0000 210.0000 66.2000 ;
	    RECT 206.0000 62.2000 206.8000 66.0000 ;
	    RECT 209.2000 62.2000 210.0000 66.0000 ;
	    RECT 210.8000 62.2000 211.6000 66.8000 ;
	    RECT 214.0000 62.2000 214.8000 67.7000 ;
	    RECT 215.6000 67.6000 216.4000 67.7000 ;
	    RECT 217.2000 67.6000 219.6000 68.2000 ;
	    RECT 221.2000 67.7000 226.2000 68.2000 ;
	    RECT 221.2000 67.6000 222.8000 67.7000 ;
	    RECT 223.6000 67.6000 226.2000 67.7000 ;
	    RECT 227.6000 67.7000 230.8000 68.2000 ;
	    RECT 227.6000 67.6000 229.2000 67.7000 ;
	    RECT 230.0000 67.6000 230.8000 67.7000 ;
	    RECT 231.6000 67.6000 232.4000 68.4000 ;
	    RECT 234.8000 67.6000 235.6000 69.2000 ;
	    RECT 236.4000 68.8000 237.2000 70.4000 ;
	    RECT 238.2000 68.4000 238.8000 71.8000 ;
	    RECT 239.6000 68.8000 240.4000 70.4000 ;
	    RECT 244.4000 68.8000 245.2000 70.4000 ;
	    RECT 245.8000 68.4000 246.4000 71.8000 ;
	    RECT 247.6000 71.6000 248.4000 71.8000 ;
	    RECT 249.2000 71.8000 250.6000 72.4000 ;
	    RECT 251.2000 71.8000 252.2000 72.4000 ;
	    RECT 262.6000 72.6000 263.4000 79.8000 ;
	    RECT 267.6000 73.6000 268.4000 74.4000 ;
	    RECT 262.6000 71.8000 264.4000 72.6000 ;
	    RECT 267.6000 72.4000 268.2000 73.6000 ;
	    RECT 269.0000 72.4000 269.8000 79.8000 ;
	    RECT 275.8000 72.4000 277.8000 79.8000 ;
	    RECT 283.8000 72.6000 284.6000 79.8000 ;
	    RECT 266.8000 71.8000 268.2000 72.4000 ;
	    RECT 268.8000 71.8000 269.8000 72.4000 ;
	    RECT 274.8000 71.8000 277.8000 72.4000 ;
	    RECT 282.8000 71.8000 284.6000 72.6000 ;
	    RECT 249.2000 71.6000 250.0000 71.8000 ;
	    RECT 251.2000 68.4000 251.8000 71.8000 ;
	    RECT 252.4000 70.3000 253.2000 70.4000 ;
	    RECT 257.2000 70.3000 258.0000 70.4000 ;
	    RECT 252.4000 69.7000 258.0000 70.3000 ;
	    RECT 252.4000 68.8000 253.2000 69.7000 ;
	    RECT 257.2000 69.6000 258.0000 69.7000 ;
	    RECT 262.0000 69.6000 262.8000 71.2000 ;
	    RECT 263.6000 68.4000 264.2000 71.8000 ;
	    RECT 266.8000 71.6000 267.6000 71.8000 ;
	    RECT 268.8000 68.4000 269.4000 71.8000 ;
	    RECT 274.8000 71.6000 277.2000 71.8000 ;
	    RECT 270.0000 68.8000 270.8000 70.4000 ;
	    RECT 238.0000 68.2000 238.8000 68.4000 ;
	    RECT 241.2000 68.2000 242.0000 68.4000 ;
	    RECT 236.4000 67.6000 238.8000 68.2000 ;
	    RECT 240.4000 67.6000 242.0000 68.2000 ;
	    RECT 242.8000 68.2000 243.6000 68.4000 ;
	    RECT 242.8000 67.6000 244.4000 68.2000 ;
	    RECT 245.8000 67.6000 248.4000 68.4000 ;
	    RECT 249.2000 67.6000 251.8000 68.4000 ;
	    RECT 254.0000 68.3000 254.8000 68.4000 ;
	    RECT 255.6000 68.3000 256.4000 68.4000 ;
	    RECT 254.0000 68.2000 256.4000 68.3000 ;
	    RECT 253.2000 67.7000 256.4000 68.2000 ;
	    RECT 253.2000 67.6000 254.8000 67.7000 ;
	    RECT 255.6000 67.6000 256.4000 67.7000 ;
	    RECT 258.8000 68.3000 259.6000 68.4000 ;
	    RECT 263.6000 68.3000 264.4000 68.4000 ;
	    RECT 258.8000 67.7000 264.4000 68.3000 ;
	    RECT 258.8000 67.6000 259.6000 67.7000 ;
	    RECT 263.6000 67.6000 264.4000 67.7000 ;
	    RECT 266.8000 67.6000 269.4000 68.4000 ;
	    RECT 271.6000 68.2000 272.4000 68.4000 ;
	    RECT 270.8000 67.6000 272.4000 68.2000 ;
	    RECT 273.2000 67.6000 274.0000 69.2000 ;
	    RECT 274.8000 68.8000 275.6000 70.4000 ;
	    RECT 276.6000 68.4000 277.2000 71.6000 ;
	    RECT 278.0000 70.3000 278.8000 70.4000 ;
	    RECT 283.0000 70.3000 283.6000 71.8000 ;
	    RECT 286.0000 71.4000 286.8000 79.8000 ;
	    RECT 290.4000 76.4000 291.2000 79.8000 ;
	    RECT 289.2000 75.8000 291.2000 76.4000 ;
	    RECT 294.8000 75.8000 295.6000 79.8000 ;
	    RECT 299.0000 75.8000 300.2000 79.8000 ;
	    RECT 289.2000 75.0000 290.0000 75.8000 ;
	    RECT 294.8000 75.2000 295.4000 75.8000 ;
	    RECT 292.6000 74.6000 296.2000 75.2000 ;
	    RECT 298.8000 75.0000 299.6000 75.8000 ;
	    RECT 292.6000 74.4000 293.4000 74.6000 ;
	    RECT 295.4000 74.4000 296.2000 74.6000 ;
	    RECT 289.2000 73.0000 290.0000 73.2000 ;
	    RECT 293.8000 73.0000 294.6000 73.2000 ;
	    RECT 289.2000 72.4000 294.6000 73.0000 ;
	    RECT 295.2000 73.0000 297.4000 73.6000 ;
	    RECT 295.2000 71.8000 295.8000 73.0000 ;
	    RECT 296.6000 72.8000 297.4000 73.0000 ;
	    RECT 299.0000 73.2000 300.4000 74.0000 ;
	    RECT 299.0000 72.2000 299.6000 73.2000 ;
	    RECT 291.0000 71.4000 295.8000 71.8000 ;
	    RECT 286.0000 71.2000 295.8000 71.4000 ;
	    RECT 297.2000 71.6000 299.6000 72.2000 ;
	    RECT 278.0000 69.7000 283.6000 70.3000 ;
	    RECT 278.0000 68.8000 278.8000 69.7000 ;
	    RECT 283.0000 68.4000 283.6000 69.7000 ;
	    RECT 284.4000 69.6000 285.2000 71.2000 ;
	    RECT 286.0000 71.0000 291.8000 71.2000 ;
	    RECT 286.0000 70.8000 291.6000 71.0000 ;
	    RECT 292.4000 70.2000 293.2000 70.4000 ;
	    RECT 288.2000 69.6000 293.2000 70.2000 ;
	    RECT 288.2000 69.4000 289.0000 69.6000 ;
	    RECT 290.8000 69.4000 291.6000 69.6000 ;
	    RECT 289.8000 68.4000 290.6000 68.6000 ;
	    RECT 297.2000 68.4000 297.8000 71.6000 ;
	    RECT 303.6000 71.2000 304.4000 79.8000 ;
	    RECT 309.0000 72.8000 309.8000 79.8000 ;
	    RECT 313.2000 75.0000 314.0000 79.0000 ;
	    RECT 318.6000 76.4000 319.4000 79.8000 ;
	    RECT 318.0000 75.6000 319.4000 76.4000 ;
	    RECT 308.2000 72.2000 309.8000 72.8000 ;
	    RECT 300.2000 70.6000 304.4000 71.2000 ;
	    RECT 300.2000 70.4000 301.0000 70.6000 ;
	    RECT 301.8000 69.8000 302.6000 70.0000 ;
	    RECT 298.8000 69.2000 302.6000 69.8000 ;
	    RECT 298.8000 69.0000 299.6000 69.2000 ;
	    RECT 276.4000 68.2000 277.2000 68.4000 ;
	    RECT 279.6000 68.2000 280.4000 68.4000 ;
	    RECT 274.8000 67.6000 277.2000 68.2000 ;
	    RECT 278.8000 67.6000 280.4000 68.2000 ;
	    RECT 282.8000 67.6000 283.6000 68.4000 ;
	    RECT 286.8000 67.8000 297.8000 68.4000 ;
	    RECT 286.8000 67.6000 288.4000 67.8000 ;
	    RECT 217.2000 66.4000 217.8000 67.6000 ;
	    RECT 221.2000 67.2000 222.0000 67.6000 ;
	    RECT 215.6000 62.8000 216.4000 66.2000 ;
	    RECT 217.2000 63.4000 218.0000 66.4000 ;
	    RECT 219.0000 66.2000 222.6000 66.6000 ;
	    RECT 223.8000 66.2000 224.4000 67.6000 ;
	    RECT 227.6000 67.2000 228.4000 67.6000 ;
	    RECT 225.4000 66.2000 229.0000 66.6000 ;
	    RECT 218.8000 66.0000 222.8000 66.2000 ;
	    RECT 218.8000 62.8000 219.6000 66.0000 ;
	    RECT 215.6000 62.2000 219.6000 62.8000 ;
	    RECT 222.0000 62.2000 222.8000 66.0000 ;
	    RECT 223.6000 62.2000 224.4000 66.2000 ;
	    RECT 225.2000 66.0000 229.2000 66.2000 ;
	    RECT 225.2000 62.2000 226.0000 66.0000 ;
	    RECT 228.4000 62.2000 229.2000 66.0000 ;
	    RECT 230.0000 64.8000 230.8000 66.4000 ;
	    RECT 231.8000 64.2000 232.4000 67.6000 ;
	    RECT 236.4000 66.2000 237.0000 67.6000 ;
	    RECT 240.4000 67.2000 241.2000 67.6000 ;
	    RECT 243.6000 67.2000 244.4000 67.6000 ;
	    RECT 238.2000 66.2000 241.8000 66.6000 ;
	    RECT 243.0000 66.2000 246.6000 66.6000 ;
	    RECT 247.6000 66.2000 248.2000 67.6000 ;
	    RECT 249.4000 66.2000 250.0000 67.6000 ;
	    RECT 253.2000 67.2000 254.0000 67.6000 ;
	    RECT 251.0000 66.2000 254.6000 66.6000 ;
	    RECT 231.6000 62.2000 232.4000 64.2000 ;
	    RECT 234.8000 62.8000 235.6000 66.2000 ;
	    RECT 236.4000 63.4000 237.2000 66.2000 ;
	    RECT 238.0000 66.0000 242.0000 66.2000 ;
	    RECT 238.0000 62.8000 238.8000 66.0000 ;
	    RECT 234.8000 62.2000 238.8000 62.8000 ;
	    RECT 241.2000 62.2000 242.0000 66.0000 ;
	    RECT 242.8000 66.0000 246.8000 66.2000 ;
	    RECT 242.8000 62.2000 243.6000 66.0000 ;
	    RECT 246.0000 62.2000 246.8000 66.0000 ;
	    RECT 247.6000 62.2000 248.4000 66.2000 ;
	    RECT 249.2000 62.2000 250.0000 66.2000 ;
	    RECT 250.8000 66.0000 254.8000 66.2000 ;
	    RECT 250.8000 62.2000 251.6000 66.0000 ;
	    RECT 254.0000 62.2000 254.8000 66.0000 ;
	    RECT 263.6000 64.2000 264.2000 67.6000 ;
	    RECT 265.2000 64.8000 266.0000 66.4000 ;
	    RECT 267.0000 66.2000 267.6000 67.6000 ;
	    RECT 270.8000 67.2000 271.6000 67.6000 ;
	    RECT 268.6000 66.2000 272.2000 66.6000 ;
	    RECT 274.8000 66.2000 275.4000 67.6000 ;
	    RECT 278.8000 67.2000 279.6000 67.6000 ;
	    RECT 276.6000 66.2000 280.2000 66.6000 ;
	    RECT 263.6000 62.2000 264.4000 64.2000 ;
	    RECT 266.8000 62.2000 267.6000 66.2000 ;
	    RECT 268.4000 66.0000 272.4000 66.2000 ;
	    RECT 268.4000 62.2000 269.2000 66.0000 ;
	    RECT 271.6000 62.2000 272.4000 66.0000 ;
	    RECT 273.2000 62.8000 274.0000 66.2000 ;
	    RECT 274.8000 63.4000 275.6000 66.2000 ;
	    RECT 276.4000 66.0000 280.4000 66.2000 ;
	    RECT 276.4000 62.8000 277.2000 66.0000 ;
	    RECT 273.2000 62.2000 277.2000 62.8000 ;
	    RECT 279.6000 62.2000 280.4000 66.0000 ;
	    RECT 281.2000 64.8000 282.0000 66.4000 ;
	    RECT 283.0000 64.2000 283.6000 67.6000 ;
	    RECT 282.8000 62.2000 283.6000 64.2000 ;
	    RECT 286.0000 62.2000 286.8000 67.0000 ;
	    RECT 291.0000 65.6000 291.6000 67.8000 ;
	    RECT 294.0000 67.6000 294.8000 67.8000 ;
	    RECT 296.6000 67.6000 297.4000 67.8000 ;
	    RECT 303.6000 67.2000 304.4000 70.6000 ;
	    RECT 306.8000 69.6000 307.6000 71.2000 ;
	    RECT 308.2000 68.4000 308.8000 72.2000 ;
	    RECT 313.4000 71.6000 314.0000 75.0000 ;
	    RECT 318.6000 72.8000 319.4000 75.6000 ;
	    RECT 322.8000 75.0000 323.6000 79.0000 ;
	    RECT 310.2000 71.0000 314.0000 71.6000 ;
	    RECT 317.8000 72.2000 319.4000 72.8000 ;
	    RECT 310.2000 69.0000 310.8000 71.0000 ;
	    RECT 305.2000 68.3000 306.0000 68.4000 ;
	    RECT 306.8000 68.3000 308.8000 68.4000 ;
	    RECT 305.2000 67.7000 308.8000 68.3000 ;
	    RECT 309.4000 68.2000 310.8000 69.0000 ;
	    RECT 311.6000 68.8000 312.4000 70.4000 ;
	    RECT 313.2000 68.8000 314.0000 70.4000 ;
	    RECT 314.8000 70.3000 315.6000 70.4000 ;
	    RECT 316.4000 70.3000 317.2000 71.2000 ;
	    RECT 314.8000 69.7000 317.2000 70.3000 ;
	    RECT 314.8000 69.6000 315.6000 69.7000 ;
	    RECT 316.4000 69.6000 317.2000 69.7000 ;
	    RECT 317.8000 68.4000 318.4000 72.2000 ;
	    RECT 323.0000 71.6000 323.6000 75.0000 ;
	    RECT 327.0000 72.4000 327.8000 79.8000 ;
	    RECT 328.4000 73.6000 329.2000 74.4000 ;
	    RECT 328.6000 72.4000 329.2000 73.6000 ;
	    RECT 327.0000 71.8000 328.0000 72.4000 ;
	    RECT 328.6000 71.8000 330.0000 72.4000 ;
	    RECT 319.8000 71.0000 323.6000 71.6000 ;
	    RECT 319.8000 69.0000 320.4000 71.0000 ;
	    RECT 305.2000 67.6000 306.0000 67.7000 ;
	    RECT 306.8000 67.6000 308.8000 67.7000 ;
	    RECT 300.6000 66.6000 304.4000 67.2000 ;
	    RECT 300.6000 66.4000 301.4000 66.6000 ;
	    RECT 289.2000 64.2000 290.0000 65.0000 ;
	    RECT 290.8000 64.8000 291.6000 65.6000 ;
	    RECT 292.6000 65.4000 293.4000 65.6000 ;
	    RECT 292.6000 64.8000 295.4000 65.4000 ;
	    RECT 294.8000 64.2000 295.4000 64.8000 ;
	    RECT 298.8000 64.2000 299.6000 65.0000 ;
	    RECT 289.2000 63.6000 291.2000 64.2000 ;
	    RECT 290.4000 62.2000 291.2000 63.6000 ;
	    RECT 294.8000 62.2000 295.6000 64.2000 ;
	    RECT 298.8000 63.6000 300.2000 64.2000 ;
	    RECT 299.0000 62.2000 300.2000 63.6000 ;
	    RECT 303.6000 62.2000 304.4000 66.6000 ;
	    RECT 308.2000 67.0000 308.8000 67.6000 ;
	    RECT 309.8000 67.8000 310.8000 68.2000 ;
	    RECT 309.8000 67.2000 314.0000 67.8000 ;
	    RECT 316.4000 67.6000 318.4000 68.4000 ;
	    RECT 319.0000 68.2000 320.4000 69.0000 ;
	    RECT 321.2000 68.8000 322.0000 70.4000 ;
	    RECT 322.8000 68.8000 323.6000 70.4000 ;
	    RECT 326.0000 68.8000 326.8000 70.4000 ;
	    RECT 327.4000 68.4000 328.0000 71.8000 ;
	    RECT 329.2000 71.6000 330.0000 71.8000 ;
	    RECT 330.8000 71.6000 331.6000 73.2000 ;
	    RECT 329.3000 70.3000 329.9000 71.6000 ;
	    RECT 332.4000 70.3000 333.2000 79.8000 ;
	    RECT 329.3000 69.7000 333.2000 70.3000 ;
	    RECT 308.2000 66.6000 309.0000 67.0000 ;
	    RECT 308.2000 66.0000 309.8000 66.6000 ;
	    RECT 309.0000 63.0000 309.8000 66.0000 ;
	    RECT 313.4000 65.0000 314.0000 67.2000 ;
	    RECT 317.8000 67.0000 318.4000 67.6000 ;
	    RECT 319.4000 67.8000 320.4000 68.2000 ;
	    RECT 324.4000 68.2000 325.2000 68.4000 ;
	    RECT 319.4000 67.2000 323.6000 67.8000 ;
	    RECT 324.4000 67.6000 326.0000 68.2000 ;
	    RECT 327.4000 67.6000 330.0000 68.4000 ;
	    RECT 325.2000 67.2000 326.0000 67.6000 ;
	    RECT 317.8000 66.6000 318.6000 67.0000 ;
	    RECT 317.8000 66.0000 319.4000 66.6000 ;
	    RECT 313.2000 63.0000 314.0000 65.0000 ;
	    RECT 318.6000 63.0000 319.4000 66.0000 ;
	    RECT 323.0000 65.0000 323.6000 67.2000 ;
	    RECT 324.6000 66.2000 328.2000 66.6000 ;
	    RECT 329.2000 66.4000 329.8000 67.6000 ;
	    RECT 322.8000 63.0000 323.6000 65.0000 ;
	    RECT 324.4000 66.0000 328.4000 66.2000 ;
	    RECT 324.4000 62.2000 325.2000 66.0000 ;
	    RECT 327.6000 62.2000 328.4000 66.0000 ;
	    RECT 329.2000 62.2000 330.0000 66.4000 ;
	    RECT 332.4000 66.2000 333.2000 69.7000 ;
	    RECT 335.6000 71.2000 336.4000 79.8000 ;
	    RECT 339.8000 75.8000 341.0000 79.8000 ;
	    RECT 344.4000 75.8000 345.2000 79.8000 ;
	    RECT 348.8000 76.4000 349.6000 79.8000 ;
	    RECT 348.8000 75.8000 350.8000 76.4000 ;
	    RECT 340.4000 75.0000 341.2000 75.8000 ;
	    RECT 344.6000 75.2000 345.2000 75.8000 ;
	    RECT 343.8000 74.6000 347.4000 75.2000 ;
	    RECT 350.0000 75.0000 350.8000 75.8000 ;
	    RECT 343.8000 74.4000 344.6000 74.6000 ;
	    RECT 346.6000 74.4000 347.4000 74.6000 ;
	    RECT 339.6000 73.2000 341.0000 74.0000 ;
	    RECT 340.4000 72.2000 341.0000 73.2000 ;
	    RECT 342.6000 73.0000 344.8000 73.6000 ;
	    RECT 342.6000 72.8000 343.4000 73.0000 ;
	    RECT 340.4000 71.6000 342.8000 72.2000 ;
	    RECT 335.6000 70.6000 339.8000 71.2000 ;
	    RECT 334.0000 68.3000 334.8000 68.4000 ;
	    RECT 335.6000 68.3000 336.4000 70.6000 ;
	    RECT 339.0000 70.4000 339.8000 70.6000 ;
	    RECT 337.4000 69.8000 338.2000 70.0000 ;
	    RECT 337.4000 69.2000 341.2000 69.8000 ;
	    RECT 340.4000 69.0000 341.2000 69.2000 ;
	    RECT 334.0000 67.7000 336.4000 68.3000 ;
	    RECT 342.2000 68.4000 342.8000 71.6000 ;
	    RECT 344.2000 71.8000 344.8000 73.0000 ;
	    RECT 345.4000 73.0000 346.2000 73.2000 ;
	    RECT 350.0000 73.0000 350.8000 73.2000 ;
	    RECT 345.4000 72.4000 350.8000 73.0000 ;
	    RECT 344.2000 71.4000 349.0000 71.8000 ;
	    RECT 353.2000 71.4000 354.0000 79.8000 ;
	    RECT 354.8000 72.4000 355.6000 79.8000 ;
	    RECT 358.0000 74.3000 358.8000 79.8000 ;
	    RECT 359.6000 74.3000 360.4000 74.4000 ;
	    RECT 358.0000 73.7000 360.4000 74.3000 ;
	    RECT 354.8000 71.8000 357.0000 72.4000 ;
	    RECT 358.0000 71.8000 358.8000 73.7000 ;
	    RECT 359.6000 73.6000 360.4000 73.7000 ;
	    RECT 344.2000 71.2000 354.0000 71.4000 ;
	    RECT 348.2000 71.0000 354.0000 71.2000 ;
	    RECT 348.4000 70.8000 354.0000 71.0000 ;
	    RECT 356.4000 71.2000 357.0000 71.8000 ;
	    RECT 356.4000 70.4000 357.6000 71.2000 ;
	    RECT 343.6000 70.3000 344.4000 70.4000 ;
	    RECT 346.8000 70.3000 347.6000 70.4000 ;
	    RECT 343.6000 70.2000 347.6000 70.3000 ;
	    RECT 343.6000 69.7000 351.8000 70.2000 ;
	    RECT 343.6000 69.6000 344.4000 69.7000 ;
	    RECT 346.8000 69.6000 351.8000 69.7000 ;
	    RECT 351.0000 69.4000 351.8000 69.6000 ;
	    RECT 354.8000 68.8000 355.6000 70.4000 ;
	    RECT 349.4000 68.4000 350.2000 68.6000 ;
	    RECT 342.2000 67.8000 353.2000 68.4000 ;
	    RECT 334.0000 66.8000 334.8000 67.7000 ;
	    RECT 335.6000 67.2000 336.4000 67.7000 ;
	    RECT 342.6000 67.6000 343.4000 67.8000 ;
	    RECT 346.8000 67.6000 347.6000 67.8000 ;
	    RECT 331.4000 65.6000 333.2000 66.2000 ;
	    RECT 335.6000 66.6000 339.4000 67.2000 ;
	    RECT 331.4000 62.2000 332.2000 65.6000 ;
	    RECT 335.6000 62.2000 336.4000 66.6000 ;
	    RECT 338.6000 66.4000 339.4000 66.6000 ;
	    RECT 348.4000 65.6000 349.0000 67.8000 ;
	    RECT 351.6000 67.6000 353.2000 67.8000 ;
	    RECT 356.4000 67.4000 357.0000 70.4000 ;
	    RECT 358.2000 69.6000 358.8000 71.8000 ;
	    RECT 346.6000 65.4000 347.4000 65.6000 ;
	    RECT 340.4000 64.2000 341.2000 65.0000 ;
	    RECT 344.6000 64.8000 347.4000 65.4000 ;
	    RECT 348.4000 64.8000 349.2000 65.6000 ;
	    RECT 344.6000 64.2000 345.2000 64.8000 ;
	    RECT 350.0000 64.2000 350.8000 65.0000 ;
	    RECT 339.8000 63.6000 341.2000 64.2000 ;
	    RECT 339.8000 62.2000 341.0000 63.6000 ;
	    RECT 344.4000 62.2000 345.2000 64.2000 ;
	    RECT 348.8000 63.6000 350.8000 64.2000 ;
	    RECT 348.8000 62.2000 349.6000 63.6000 ;
	    RECT 353.2000 62.2000 354.0000 67.0000 ;
	    RECT 354.8000 66.8000 357.0000 67.4000 ;
	    RECT 354.8000 62.2000 355.6000 66.8000 ;
	    RECT 358.0000 62.2000 358.8000 69.6000 ;
	    RECT 359.6000 66.8000 360.4000 68.4000 ;
	    RECT 361.2000 68.3000 362.0000 79.8000 ;
	    RECT 362.8000 71.6000 363.6000 73.2000 ;
	    RECT 364.4000 71.2000 365.2000 79.8000 ;
	    RECT 368.6000 75.8000 369.8000 79.8000 ;
	    RECT 373.2000 75.8000 374.0000 79.8000 ;
	    RECT 377.6000 76.4000 378.4000 79.8000 ;
	    RECT 377.6000 75.8000 379.6000 76.4000 ;
	    RECT 369.2000 75.0000 370.0000 75.8000 ;
	    RECT 373.4000 75.2000 374.0000 75.8000 ;
	    RECT 372.6000 74.6000 376.2000 75.2000 ;
	    RECT 378.8000 75.0000 379.6000 75.8000 ;
	    RECT 372.6000 74.4000 373.4000 74.6000 ;
	    RECT 375.4000 74.4000 376.2000 74.6000 ;
	    RECT 368.4000 73.2000 369.8000 74.0000 ;
	    RECT 369.2000 72.2000 369.8000 73.2000 ;
	    RECT 371.4000 73.0000 373.6000 73.6000 ;
	    RECT 371.4000 72.8000 372.2000 73.0000 ;
	    RECT 369.2000 71.6000 371.6000 72.2000 ;
	    RECT 364.4000 70.6000 368.6000 71.2000 ;
	    RECT 362.8000 68.3000 363.6000 68.4000 ;
	    RECT 361.2000 67.7000 363.6000 68.3000 ;
	    RECT 361.2000 66.2000 362.0000 67.7000 ;
	    RECT 362.8000 67.6000 363.6000 67.7000 ;
	    RECT 364.4000 67.2000 365.2000 70.6000 ;
	    RECT 367.8000 70.4000 368.6000 70.6000 ;
	    RECT 366.2000 69.8000 367.0000 70.0000 ;
	    RECT 366.2000 69.2000 370.0000 69.8000 ;
	    RECT 369.2000 69.0000 370.0000 69.2000 ;
	    RECT 371.0000 68.4000 371.6000 71.6000 ;
	    RECT 373.0000 71.8000 373.6000 73.0000 ;
	    RECT 374.2000 73.0000 375.0000 73.2000 ;
	    RECT 378.8000 73.0000 379.6000 73.2000 ;
	    RECT 374.2000 72.4000 379.6000 73.0000 ;
	    RECT 373.0000 71.4000 377.8000 71.8000 ;
	    RECT 382.0000 71.4000 382.8000 79.8000 ;
	    RECT 384.4000 73.6000 385.2000 74.4000 ;
	    RECT 384.4000 72.4000 385.0000 73.6000 ;
	    RECT 385.8000 72.4000 386.6000 79.8000 ;
	    RECT 383.6000 71.8000 385.0000 72.4000 ;
	    RECT 385.6000 71.8000 386.6000 72.4000 ;
	    RECT 390.0000 71.8000 390.8000 79.8000 ;
	    RECT 393.2000 72.4000 394.0000 79.8000 ;
	    RECT 391.8000 71.8000 394.0000 72.4000 ;
	    RECT 383.6000 71.6000 384.4000 71.8000 ;
	    RECT 373.0000 71.2000 382.8000 71.4000 ;
	    RECT 377.0000 71.0000 382.8000 71.2000 ;
	    RECT 377.2000 70.8000 382.8000 71.0000 ;
	    RECT 385.6000 70.4000 386.2000 71.8000 ;
	    RECT 375.6000 70.2000 376.4000 70.4000 ;
	    RECT 375.6000 69.6000 380.6000 70.2000 ;
	    RECT 385.2000 69.6000 386.2000 70.4000 ;
	    RECT 377.2000 69.4000 378.0000 69.6000 ;
	    RECT 379.8000 69.4000 380.6000 69.6000 ;
	    RECT 378.2000 68.4000 379.0000 68.6000 ;
	    RECT 385.6000 68.4000 386.2000 69.6000 ;
	    RECT 386.8000 70.3000 387.6000 70.4000 ;
	    RECT 388.4000 70.3000 389.2000 70.4000 ;
	    RECT 386.8000 69.7000 389.2000 70.3000 ;
	    RECT 386.8000 68.8000 387.6000 69.7000 ;
	    RECT 388.4000 69.6000 389.2000 69.7000 ;
	    RECT 390.0000 69.6000 390.6000 71.8000 ;
	    RECT 391.8000 71.2000 392.4000 71.8000 ;
	    RECT 391.2000 70.4000 392.4000 71.2000 ;
	    RECT 394.8000 71.2000 395.6000 79.8000 ;
	    RECT 399.0000 75.8000 400.2000 79.8000 ;
	    RECT 403.6000 75.8000 404.4000 79.8000 ;
	    RECT 408.0000 76.4000 408.8000 79.8000 ;
	    RECT 408.0000 75.8000 410.0000 76.4000 ;
	    RECT 399.6000 75.0000 400.4000 75.8000 ;
	    RECT 403.8000 75.2000 404.4000 75.8000 ;
	    RECT 403.0000 74.6000 406.6000 75.2000 ;
	    RECT 409.2000 75.0000 410.0000 75.8000 ;
	    RECT 403.0000 74.4000 403.8000 74.6000 ;
	    RECT 405.8000 74.4000 406.6000 74.6000 ;
	    RECT 398.8000 73.2000 400.2000 74.0000 ;
	    RECT 399.6000 72.2000 400.2000 73.2000 ;
	    RECT 401.8000 73.0000 404.0000 73.6000 ;
	    RECT 401.8000 72.8000 402.6000 73.0000 ;
	    RECT 399.6000 71.6000 402.0000 72.2000 ;
	    RECT 394.8000 70.6000 399.0000 71.2000 ;
	    RECT 371.0000 67.8000 382.0000 68.4000 ;
	    RECT 371.4000 67.6000 372.2000 67.8000 ;
	    RECT 364.4000 66.6000 368.2000 67.2000 ;
	    RECT 361.2000 65.6000 363.0000 66.2000 ;
	    RECT 362.2000 62.2000 363.0000 65.6000 ;
	    RECT 364.4000 62.2000 365.2000 66.6000 ;
	    RECT 367.4000 66.4000 368.2000 66.6000 ;
	    RECT 377.2000 66.4000 377.8000 67.8000 ;
	    RECT 380.4000 67.6000 382.0000 67.8000 ;
	    RECT 383.6000 67.6000 386.2000 68.4000 ;
	    RECT 388.4000 68.2000 389.2000 68.4000 ;
	    RECT 387.6000 67.6000 389.2000 68.2000 ;
	    RECT 375.4000 65.4000 376.2000 65.6000 ;
	    RECT 369.2000 64.2000 370.0000 65.0000 ;
	    RECT 373.4000 64.8000 376.2000 65.4000 ;
	    RECT 377.2000 64.8000 378.0000 66.4000 ;
	    RECT 373.4000 64.2000 374.0000 64.8000 ;
	    RECT 378.8000 64.2000 379.6000 65.0000 ;
	    RECT 368.6000 63.6000 370.0000 64.2000 ;
	    RECT 368.6000 62.2000 369.8000 63.6000 ;
	    RECT 373.2000 62.2000 374.0000 64.2000 ;
	    RECT 377.6000 63.6000 379.6000 64.2000 ;
	    RECT 377.6000 62.2000 378.4000 63.6000 ;
	    RECT 382.0000 62.2000 382.8000 67.0000 ;
	    RECT 383.8000 66.2000 384.4000 67.6000 ;
	    RECT 387.6000 67.2000 388.4000 67.6000 ;
	    RECT 385.4000 66.2000 389.0000 66.6000 ;
	    RECT 383.6000 62.2000 384.4000 66.2000 ;
	    RECT 385.2000 66.0000 389.2000 66.2000 ;
	    RECT 385.2000 62.2000 386.0000 66.0000 ;
	    RECT 388.4000 62.2000 389.2000 66.0000 ;
	    RECT 390.0000 62.2000 390.8000 69.6000 ;
	    RECT 391.8000 67.4000 392.4000 70.4000 ;
	    RECT 393.2000 68.8000 394.0000 70.4000 ;
	    RECT 391.8000 66.8000 394.0000 67.4000 ;
	    RECT 393.2000 62.2000 394.0000 66.8000 ;
	    RECT 394.8000 67.2000 395.6000 70.6000 ;
	    RECT 398.2000 70.4000 399.0000 70.6000 ;
	    RECT 396.6000 69.8000 397.4000 70.0000 ;
	    RECT 396.6000 69.2000 400.4000 69.8000 ;
	    RECT 399.6000 69.0000 400.4000 69.2000 ;
	    RECT 401.4000 68.4000 402.0000 71.6000 ;
	    RECT 403.4000 71.8000 404.0000 73.0000 ;
	    RECT 404.6000 73.0000 405.4000 73.2000 ;
	    RECT 409.2000 73.0000 410.0000 73.2000 ;
	    RECT 404.6000 72.4000 410.0000 73.0000 ;
	    RECT 403.4000 71.4000 408.2000 71.8000 ;
	    RECT 412.4000 71.4000 413.2000 79.8000 ;
	    RECT 403.4000 71.2000 413.2000 71.4000 ;
	    RECT 407.4000 71.0000 413.2000 71.2000 ;
	    RECT 407.6000 70.8000 413.2000 71.0000 ;
	    RECT 406.0000 70.2000 406.8000 70.4000 ;
	    RECT 422.0000 70.3000 422.8000 79.8000 ;
	    RECT 426.0000 73.6000 426.8000 74.4000 ;
	    RECT 423.6000 71.6000 424.4000 73.2000 ;
	    RECT 426.0000 72.4000 426.6000 73.6000 ;
	    RECT 427.4000 72.4000 428.2000 79.8000 ;
	    RECT 425.2000 71.8000 426.6000 72.4000 ;
	    RECT 427.2000 71.8000 428.2000 72.4000 ;
	    RECT 425.2000 71.6000 426.0000 71.8000 ;
	    RECT 425.3000 70.3000 425.9000 71.6000 ;
	    RECT 406.0000 69.6000 411.0000 70.2000 ;
	    RECT 407.6000 69.4000 408.4000 69.6000 ;
	    RECT 410.2000 69.4000 411.0000 69.6000 ;
	    RECT 422.0000 69.7000 425.9000 70.3000 ;
	    RECT 408.6000 68.4000 409.4000 68.6000 ;
	    RECT 401.4000 67.8000 412.4000 68.4000 ;
	    RECT 401.8000 67.6000 402.6000 67.8000 ;
	    RECT 394.8000 66.6000 398.6000 67.2000 ;
	    RECT 394.8000 62.2000 395.6000 66.6000 ;
	    RECT 397.8000 66.4000 398.6000 66.6000 ;
	    RECT 407.6000 65.6000 408.2000 67.8000 ;
	    RECT 410.8000 67.6000 412.4000 67.8000 ;
	    RECT 414.0000 68.3000 414.8000 68.4000 ;
	    RECT 420.4000 68.3000 421.2000 68.4000 ;
	    RECT 414.0000 67.7000 421.2000 68.3000 ;
	    RECT 414.0000 67.6000 414.8000 67.7000 ;
	    RECT 405.8000 65.4000 406.6000 65.6000 ;
	    RECT 399.6000 64.2000 400.4000 65.0000 ;
	    RECT 403.8000 64.8000 406.6000 65.4000 ;
	    RECT 407.6000 64.8000 408.4000 65.6000 ;
	    RECT 403.8000 64.2000 404.4000 64.8000 ;
	    RECT 409.2000 64.2000 410.0000 65.0000 ;
	    RECT 399.0000 63.6000 400.4000 64.2000 ;
	    RECT 399.0000 62.2000 400.2000 63.6000 ;
	    RECT 403.6000 62.2000 404.4000 64.2000 ;
	    RECT 408.0000 63.6000 410.0000 64.2000 ;
	    RECT 408.0000 62.2000 408.8000 63.6000 ;
	    RECT 412.4000 62.2000 413.2000 67.0000 ;
	    RECT 420.4000 66.8000 421.2000 67.7000 ;
	    RECT 422.0000 66.2000 422.8000 69.7000 ;
	    RECT 427.2000 68.4000 427.8000 71.8000 ;
	    RECT 433.2000 71.2000 434.0000 79.8000 ;
	    RECT 436.4000 71.2000 437.2000 79.8000 ;
	    RECT 439.6000 71.2000 440.4000 79.8000 ;
	    RECT 442.8000 71.2000 443.6000 79.8000 ;
	    RECT 431.6000 70.4000 434.0000 71.2000 ;
	    RECT 435.0000 70.4000 437.2000 71.2000 ;
	    RECT 438.2000 70.4000 440.4000 71.2000 ;
	    RECT 441.8000 70.4000 443.6000 71.2000 ;
	    RECT 428.4000 68.8000 429.2000 70.4000 ;
	    RECT 425.2000 67.6000 427.8000 68.4000 ;
	    RECT 430.0000 68.2000 430.8000 68.4000 ;
	    RECT 429.2000 67.6000 430.8000 68.2000 ;
	    RECT 431.6000 67.6000 432.4000 70.4000 ;
	    RECT 435.0000 69.0000 435.8000 70.4000 ;
	    RECT 438.2000 69.0000 439.0000 70.4000 ;
	    RECT 441.8000 69.0000 442.6000 70.4000 ;
	    RECT 433.2000 68.2000 435.8000 69.0000 ;
	    RECT 436.6000 68.2000 439.0000 69.0000 ;
	    RECT 440.0000 68.2000 442.6000 69.0000 ;
	    RECT 435.0000 67.6000 435.8000 68.2000 ;
	    RECT 438.2000 67.6000 439.0000 68.2000 ;
	    RECT 441.8000 67.6000 442.6000 68.2000 ;
	    RECT 447.6000 68.3000 448.4000 79.8000 ;
	    RECT 451.8000 72.4000 452.6000 79.8000 ;
	    RECT 453.2000 73.6000 454.0000 74.4000 ;
	    RECT 453.4000 72.4000 454.0000 73.6000 ;
	    RECT 451.8000 71.8000 452.8000 72.4000 ;
	    RECT 453.4000 71.8000 454.8000 72.4000 ;
	    RECT 450.8000 68.8000 451.6000 70.4000 ;
	    RECT 452.2000 68.4000 452.8000 71.8000 ;
	    RECT 454.0000 71.6000 454.8000 71.8000 ;
	    RECT 455.6000 71.2000 456.4000 79.8000 ;
	    RECT 459.8000 75.8000 461.0000 79.8000 ;
	    RECT 464.4000 75.8000 465.2000 79.8000 ;
	    RECT 468.8000 76.4000 469.6000 79.8000 ;
	    RECT 468.8000 75.8000 470.8000 76.4000 ;
	    RECT 460.4000 75.0000 461.2000 75.8000 ;
	    RECT 464.6000 75.2000 465.2000 75.8000 ;
	    RECT 463.8000 74.6000 467.4000 75.2000 ;
	    RECT 470.0000 75.0000 470.8000 75.8000 ;
	    RECT 463.8000 74.4000 464.6000 74.6000 ;
	    RECT 466.6000 74.4000 467.4000 74.6000 ;
	    RECT 459.6000 73.2000 461.0000 74.0000 ;
	    RECT 460.4000 72.2000 461.0000 73.2000 ;
	    RECT 462.6000 73.0000 464.8000 73.6000 ;
	    RECT 462.6000 72.8000 463.4000 73.0000 ;
	    RECT 460.4000 71.6000 462.8000 72.2000 ;
	    RECT 455.6000 70.6000 459.8000 71.2000 ;
	    RECT 449.2000 68.3000 450.0000 68.4000 ;
	    RECT 447.6000 68.2000 450.0000 68.3000 ;
	    RECT 447.6000 67.7000 450.8000 68.2000 ;
	    RECT 425.4000 66.2000 426.0000 67.6000 ;
	    RECT 429.2000 67.2000 430.0000 67.6000 ;
	    RECT 431.6000 66.8000 434.0000 67.6000 ;
	    RECT 435.0000 66.8000 437.2000 67.6000 ;
	    RECT 438.2000 66.8000 440.4000 67.6000 ;
	    RECT 441.8000 66.8000 443.6000 67.6000 ;
	    RECT 427.0000 66.2000 430.6000 66.6000 ;
	    RECT 422.0000 65.6000 423.8000 66.2000 ;
	    RECT 423.0000 62.2000 423.8000 65.6000 ;
	    RECT 425.2000 62.2000 426.0000 66.2000 ;
	    RECT 426.8000 66.0000 430.8000 66.2000 ;
	    RECT 426.8000 62.2000 427.6000 66.0000 ;
	    RECT 430.0000 62.2000 430.8000 66.0000 ;
	    RECT 433.2000 62.2000 434.0000 66.8000 ;
	    RECT 436.4000 62.2000 437.2000 66.8000 ;
	    RECT 439.6000 62.2000 440.4000 66.8000 ;
	    RECT 442.8000 62.2000 443.6000 66.8000 ;
	    RECT 446.0000 64.8000 446.8000 66.4000 ;
	    RECT 447.6000 62.2000 448.4000 67.7000 ;
	    RECT 449.2000 67.6000 450.8000 67.7000 ;
	    RECT 452.2000 67.6000 454.8000 68.4000 ;
	    RECT 450.0000 67.2000 450.8000 67.6000 ;
	    RECT 449.4000 66.2000 453.0000 66.6000 ;
	    RECT 454.0000 66.2000 454.6000 67.6000 ;
	    RECT 455.6000 67.2000 456.4000 70.6000 ;
	    RECT 459.0000 70.4000 459.8000 70.6000 ;
	    RECT 462.2000 70.4000 462.8000 71.6000 ;
	    RECT 464.2000 71.8000 464.8000 73.0000 ;
	    RECT 465.4000 73.0000 466.2000 73.2000 ;
	    RECT 470.0000 73.0000 470.8000 73.2000 ;
	    RECT 465.4000 72.4000 470.8000 73.0000 ;
	    RECT 464.2000 71.4000 469.0000 71.8000 ;
	    RECT 473.2000 71.4000 474.0000 79.8000 ;
	    RECT 464.2000 71.2000 474.0000 71.4000 ;
	    RECT 468.2000 71.0000 474.0000 71.2000 ;
	    RECT 468.4000 70.8000 474.0000 71.0000 ;
	    RECT 457.4000 69.8000 458.2000 70.0000 ;
	    RECT 457.4000 69.2000 461.2000 69.8000 ;
	    RECT 462.0000 69.6000 462.8000 70.4000 ;
	    RECT 466.8000 70.2000 467.6000 70.4000 ;
	    RECT 466.8000 69.6000 471.8000 70.2000 ;
	    RECT 460.4000 69.0000 461.2000 69.2000 ;
	    RECT 462.2000 68.4000 462.8000 69.6000 ;
	    RECT 468.4000 69.4000 469.2000 69.6000 ;
	    RECT 471.0000 69.4000 471.8000 69.6000 ;
	    RECT 469.4000 68.4000 470.2000 68.6000 ;
	    RECT 462.2000 67.8000 473.2000 68.4000 ;
	    RECT 462.6000 67.6000 463.4000 67.8000 ;
	    RECT 455.6000 66.6000 459.4000 67.2000 ;
	    RECT 449.2000 66.0000 453.2000 66.2000 ;
	    RECT 449.2000 62.2000 450.0000 66.0000 ;
	    RECT 452.4000 62.2000 453.2000 66.0000 ;
	    RECT 454.0000 62.2000 454.8000 66.2000 ;
	    RECT 455.6000 62.2000 456.4000 66.6000 ;
	    RECT 458.6000 66.4000 459.4000 66.6000 ;
	    RECT 468.4000 65.6000 469.0000 67.8000 ;
	    RECT 471.6000 67.6000 473.2000 67.8000 ;
	    RECT 476.4000 68.3000 477.2000 79.8000 ;
	    RECT 480.6000 72.4000 481.4000 79.8000 ;
	    RECT 484.4000 75.8000 485.2000 79.8000 ;
	    RECT 484.6000 75.6000 485.2000 75.8000 ;
	    RECT 487.6000 75.8000 488.4000 79.8000 ;
	    RECT 487.6000 75.6000 488.2000 75.8000 ;
	    RECT 484.6000 75.0000 488.2000 75.6000 ;
	    RECT 482.0000 73.6000 482.8000 74.4000 ;
	    RECT 482.2000 72.4000 482.8000 73.6000 ;
	    RECT 484.6000 72.4000 485.2000 75.0000 ;
	    RECT 486.0000 72.8000 486.8000 74.4000 ;
	    RECT 479.6000 71.6000 481.6000 72.4000 ;
	    RECT 482.2000 71.8000 483.6000 72.4000 ;
	    RECT 482.8000 71.6000 483.6000 71.8000 ;
	    RECT 484.4000 71.6000 485.2000 72.4000 ;
	    RECT 478.0000 70.3000 478.8000 70.4000 ;
	    RECT 479.6000 70.3000 480.4000 70.4000 ;
	    RECT 478.0000 69.7000 480.4000 70.3000 ;
	    RECT 478.0000 69.6000 478.8000 69.7000 ;
	    RECT 479.6000 68.8000 480.4000 69.7000 ;
	    RECT 481.0000 68.4000 481.6000 71.6000 ;
	    RECT 484.6000 68.4000 485.2000 71.6000 ;
	    RECT 486.8000 69.6000 488.4000 70.4000 ;
	    RECT 478.0000 68.3000 478.8000 68.4000 ;
	    RECT 476.4000 68.2000 478.8000 68.3000 ;
	    RECT 476.4000 67.7000 479.6000 68.2000 ;
	    RECT 466.6000 65.4000 467.4000 65.6000 ;
	    RECT 460.4000 64.2000 461.2000 65.0000 ;
	    RECT 464.6000 64.8000 467.4000 65.4000 ;
	    RECT 468.4000 64.8000 469.2000 65.6000 ;
	    RECT 464.6000 64.2000 465.2000 64.8000 ;
	    RECT 470.0000 64.2000 470.8000 65.0000 ;
	    RECT 459.8000 63.6000 461.2000 64.2000 ;
	    RECT 459.8000 62.2000 461.0000 63.6000 ;
	    RECT 464.4000 62.2000 465.2000 64.2000 ;
	    RECT 468.8000 63.6000 470.8000 64.2000 ;
	    RECT 468.8000 62.2000 469.6000 63.6000 ;
	    RECT 473.2000 62.2000 474.0000 67.0000 ;
	    RECT 474.8000 64.8000 475.6000 66.4000 ;
	    RECT 476.4000 62.2000 477.2000 67.7000 ;
	    RECT 478.0000 67.6000 479.6000 67.7000 ;
	    RECT 481.0000 67.6000 483.6000 68.4000 ;
	    RECT 484.6000 68.2000 486.2000 68.4000 ;
	    RECT 492.4000 68.3000 493.2000 79.8000 ;
	    RECT 496.6000 72.4000 497.4000 79.8000 ;
	    RECT 498.0000 73.6000 498.8000 74.4000 ;
	    RECT 498.2000 72.4000 498.8000 73.6000 ;
	    RECT 496.6000 71.8000 497.6000 72.4000 ;
	    RECT 498.2000 71.8000 499.6000 72.4000 ;
	    RECT 495.6000 68.8000 496.4000 70.4000 ;
	    RECT 497.0000 68.4000 497.6000 71.8000 ;
	    RECT 498.8000 71.6000 499.6000 71.8000 ;
	    RECT 502.0000 71.2000 502.8000 79.8000 ;
	    RECT 505.2000 71.2000 506.0000 79.8000 ;
	    RECT 508.4000 71.2000 509.2000 79.8000 ;
	    RECT 511.6000 71.2000 512.4000 79.8000 ;
	    RECT 500.4000 70.4000 502.8000 71.2000 ;
	    RECT 503.8000 70.4000 506.0000 71.2000 ;
	    RECT 507.0000 70.4000 509.2000 71.2000 ;
	    RECT 510.6000 70.4000 512.4000 71.2000 ;
	    RECT 494.0000 68.3000 494.8000 68.4000 ;
	    RECT 492.4000 68.2000 494.8000 68.3000 ;
	    RECT 484.6000 67.8000 486.4000 68.2000 ;
	    RECT 478.8000 67.2000 479.6000 67.6000 ;
	    RECT 478.2000 66.2000 481.8000 66.6000 ;
	    RECT 482.8000 66.2000 483.4000 67.6000 ;
	    RECT 478.0000 66.0000 482.0000 66.2000 ;
	    RECT 478.0000 62.2000 478.8000 66.0000 ;
	    RECT 481.2000 62.2000 482.0000 66.0000 ;
	    RECT 482.8000 62.2000 483.6000 66.2000 ;
	    RECT 485.6000 62.2000 486.4000 67.8000 ;
	    RECT 492.4000 67.7000 495.6000 68.2000 ;
	    RECT 490.8000 64.8000 491.6000 66.4000 ;
	    RECT 492.4000 62.2000 493.2000 67.7000 ;
	    RECT 494.0000 67.6000 495.6000 67.7000 ;
	    RECT 497.0000 67.6000 499.6000 68.4000 ;
	    RECT 500.4000 67.6000 501.2000 70.4000 ;
	    RECT 503.8000 69.0000 504.6000 70.4000 ;
	    RECT 507.0000 69.0000 507.8000 70.4000 ;
	    RECT 510.6000 69.0000 511.4000 70.4000 ;
	    RECT 502.0000 68.2000 504.6000 69.0000 ;
	    RECT 505.4000 68.2000 507.8000 69.0000 ;
	    RECT 508.8000 68.2000 511.4000 69.0000 ;
	    RECT 503.8000 67.6000 504.6000 68.2000 ;
	    RECT 507.0000 67.6000 507.8000 68.2000 ;
	    RECT 510.6000 67.6000 511.4000 68.2000 ;
	    RECT 494.8000 67.2000 495.6000 67.6000 ;
	    RECT 494.2000 66.2000 497.8000 66.6000 ;
	    RECT 498.8000 66.2000 499.4000 67.6000 ;
	    RECT 500.4000 66.8000 502.8000 67.6000 ;
	    RECT 503.8000 66.8000 506.0000 67.6000 ;
	    RECT 507.0000 66.8000 509.2000 67.6000 ;
	    RECT 510.6000 66.8000 512.4000 67.6000 ;
	    RECT 494.0000 66.0000 498.0000 66.2000 ;
	    RECT 494.0000 62.2000 494.8000 66.0000 ;
	    RECT 497.2000 62.2000 498.0000 66.0000 ;
	    RECT 498.8000 62.2000 499.6000 66.2000 ;
	    RECT 502.0000 62.2000 502.8000 66.8000 ;
	    RECT 505.2000 62.2000 506.0000 66.8000 ;
	    RECT 508.4000 62.2000 509.2000 66.8000 ;
	    RECT 511.6000 62.2000 512.4000 66.8000 ;
	    RECT 4.4000 55.2000 5.2000 59.8000 ;
	    RECT 3.0000 54.6000 5.2000 55.2000 ;
	    RECT 7.6000 55.2000 8.4000 59.8000 ;
	    RECT 10.8000 55.2000 11.6000 59.8000 ;
	    RECT 14.0000 55.2000 14.8000 59.8000 ;
	    RECT 17.2000 55.2000 18.0000 59.8000 ;
	    RECT 20.4000 55.4000 21.2000 59.8000 ;
	    RECT 24.6000 58.4000 25.8000 59.8000 ;
	    RECT 24.6000 57.8000 26.0000 58.4000 ;
	    RECT 29.2000 57.8000 30.0000 59.8000 ;
	    RECT 33.6000 58.4000 34.4000 59.8000 ;
	    RECT 33.6000 57.8000 35.6000 58.4000 ;
	    RECT 25.2000 57.0000 26.0000 57.8000 ;
	    RECT 29.4000 57.2000 30.0000 57.8000 ;
	    RECT 29.4000 56.6000 32.2000 57.2000 ;
	    RECT 31.4000 56.4000 32.2000 56.6000 ;
	    RECT 33.2000 56.4000 34.0000 57.2000 ;
	    RECT 34.8000 57.0000 35.6000 57.8000 ;
	    RECT 23.4000 55.4000 24.2000 55.6000 ;
	    RECT 3.0000 51.6000 3.6000 54.6000 ;
	    RECT 7.6000 54.4000 9.4000 55.2000 ;
	    RECT 10.8000 54.4000 13.0000 55.2000 ;
	    RECT 14.0000 54.4000 16.2000 55.2000 ;
	    RECT 17.2000 54.4000 19.6000 55.2000 ;
	    RECT 8.6000 53.8000 9.4000 54.4000 ;
	    RECT 12.2000 53.8000 13.0000 54.4000 ;
	    RECT 15.4000 53.8000 16.2000 54.4000 ;
	    RECT 4.4000 51.6000 5.2000 53.2000 ;
	    RECT 8.6000 53.0000 11.2000 53.8000 ;
	    RECT 12.2000 53.0000 14.6000 53.8000 ;
	    RECT 15.4000 53.0000 18.0000 53.8000 ;
	    RECT 8.6000 51.6000 9.4000 53.0000 ;
	    RECT 12.2000 51.6000 13.0000 53.0000 ;
	    RECT 15.4000 51.6000 16.2000 53.0000 ;
	    RECT 18.8000 51.6000 19.6000 54.4000 ;
	    RECT 2.4000 50.8000 3.6000 51.6000 ;
	    RECT 3.0000 50.2000 3.6000 50.8000 ;
	    RECT 7.6000 50.8000 9.4000 51.6000 ;
	    RECT 10.8000 50.8000 13.0000 51.6000 ;
	    RECT 14.0000 50.8000 16.2000 51.6000 ;
	    RECT 17.2000 50.8000 19.6000 51.6000 ;
	    RECT 20.4000 54.8000 24.2000 55.4000 ;
	    RECT 20.4000 51.4000 21.2000 54.8000 ;
	    RECT 27.4000 54.2000 28.2000 54.4000 ;
	    RECT 33.2000 54.2000 33.8000 56.4000 ;
	    RECT 38.0000 55.0000 38.8000 59.8000 ;
	    RECT 39.6000 55.8000 40.4000 59.8000 ;
	    RECT 41.2000 56.0000 42.0000 59.8000 ;
	    RECT 44.4000 56.0000 45.2000 59.8000 ;
	    RECT 41.2000 55.8000 45.2000 56.0000 ;
	    RECT 46.0000 55.8000 46.8000 59.8000 ;
	    RECT 47.6000 56.0000 48.4000 59.8000 ;
	    RECT 50.8000 56.0000 51.6000 59.8000 ;
	    RECT 47.6000 55.8000 51.6000 56.0000 ;
	    RECT 39.8000 54.4000 40.4000 55.8000 ;
	    RECT 41.4000 55.4000 45.0000 55.8000 ;
	    RECT 43.6000 54.4000 44.4000 54.8000 ;
	    RECT 46.2000 54.4000 46.8000 55.8000 ;
	    RECT 47.8000 55.4000 51.4000 55.8000 ;
	    RECT 52.4000 55.6000 53.2000 59.8000 ;
	    RECT 54.0000 56.0000 54.8000 59.8000 ;
	    RECT 57.2000 56.0000 58.0000 59.8000 ;
	    RECT 54.0000 55.8000 58.0000 56.0000 ;
	    RECT 58.8000 55.8000 59.6000 59.8000 ;
	    RECT 60.4000 56.0000 61.2000 59.8000 ;
	    RECT 63.6000 56.0000 64.4000 59.8000 ;
	    RECT 60.4000 55.8000 64.4000 56.0000 ;
	    RECT 50.0000 54.4000 50.8000 54.8000 ;
	    RECT 52.6000 54.4000 53.2000 55.6000 ;
	    RECT 54.2000 55.4000 57.8000 55.8000 ;
	    RECT 56.4000 54.4000 57.2000 54.8000 ;
	    RECT 59.0000 54.4000 59.6000 55.8000 ;
	    RECT 60.6000 55.4000 64.2000 55.8000 ;
	    RECT 65.2000 55.4000 66.0000 59.8000 ;
	    RECT 69.4000 58.4000 70.6000 59.8000 ;
	    RECT 69.4000 57.8000 70.8000 58.4000 ;
	    RECT 74.0000 57.8000 74.8000 59.8000 ;
	    RECT 78.4000 58.4000 79.2000 59.8000 ;
	    RECT 78.4000 57.8000 80.4000 58.4000 ;
	    RECT 70.0000 57.0000 70.8000 57.8000 ;
	    RECT 74.2000 57.2000 74.8000 57.8000 ;
	    RECT 74.2000 56.6000 77.0000 57.2000 ;
	    RECT 76.2000 56.4000 77.0000 56.6000 ;
	    RECT 78.0000 56.4000 78.8000 57.2000 ;
	    RECT 79.6000 57.0000 80.4000 57.8000 ;
	    RECT 71.6000 56.3000 72.4000 56.4000 ;
	    RECT 68.4000 55.7000 72.4000 56.3000 ;
	    RECT 68.4000 55.6000 69.2000 55.7000 ;
	    RECT 71.6000 55.6000 72.4000 55.7000 ;
	    RECT 68.2000 55.4000 69.2000 55.6000 ;
	    RECT 65.2000 54.8000 69.2000 55.4000 ;
	    RECT 62.8000 54.4000 63.6000 54.8000 ;
	    RECT 36.4000 54.2000 38.0000 54.4000 ;
	    RECT 27.0000 53.6000 38.0000 54.2000 ;
	    RECT 39.6000 53.6000 42.2000 54.4000 ;
	    RECT 43.6000 53.8000 45.2000 54.4000 ;
	    RECT 44.4000 53.6000 45.2000 53.8000 ;
	    RECT 46.0000 53.6000 48.6000 54.4000 ;
	    RECT 50.0000 53.8000 51.6000 54.4000 ;
	    RECT 50.8000 53.6000 51.6000 53.8000 ;
	    RECT 52.4000 53.6000 55.0000 54.4000 ;
	    RECT 56.4000 53.8000 58.0000 54.4000 ;
	    RECT 57.2000 53.6000 58.0000 53.8000 ;
	    RECT 58.8000 53.6000 61.4000 54.4000 ;
	    RECT 62.8000 53.8000 64.4000 54.4000 ;
	    RECT 63.6000 53.6000 64.4000 53.8000 ;
	    RECT 25.2000 52.8000 26.0000 53.0000 ;
	    RECT 22.2000 52.2000 26.0000 52.8000 ;
	    RECT 27.0000 52.4000 27.6000 53.6000 ;
	    RECT 34.2000 53.4000 35.0000 53.6000 ;
	    RECT 33.2000 52.4000 34.0000 52.6000 ;
	    RECT 35.8000 52.4000 36.6000 52.6000 ;
	    RECT 22.2000 52.0000 23.0000 52.2000 ;
	    RECT 26.8000 51.6000 27.6000 52.4000 ;
	    RECT 31.6000 51.8000 36.6000 52.4000 ;
	    RECT 31.6000 51.6000 32.4000 51.8000 ;
	    RECT 23.8000 51.4000 24.6000 51.6000 ;
	    RECT 20.4000 50.8000 24.6000 51.4000 ;
	    RECT 3.0000 49.6000 5.2000 50.2000 ;
	    RECT 4.4000 42.2000 5.2000 49.6000 ;
	    RECT 7.6000 42.2000 8.4000 50.8000 ;
	    RECT 10.8000 42.2000 11.6000 50.8000 ;
	    RECT 14.0000 42.2000 14.8000 50.8000 ;
	    RECT 17.2000 42.2000 18.0000 50.8000 ;
	    RECT 20.4000 42.2000 21.2000 50.8000 ;
	    RECT 27.0000 50.4000 27.6000 51.6000 ;
	    RECT 33.2000 51.0000 38.8000 51.2000 ;
	    RECT 33.0000 50.8000 38.8000 51.0000 ;
	    RECT 25.2000 49.8000 27.6000 50.4000 ;
	    RECT 29.0000 50.6000 38.8000 50.8000 ;
	    RECT 29.0000 50.2000 33.8000 50.6000 ;
	    RECT 25.2000 48.8000 25.8000 49.8000 ;
	    RECT 24.4000 48.0000 25.8000 48.8000 ;
	    RECT 27.4000 49.0000 28.2000 49.2000 ;
	    RECT 29.0000 49.0000 29.6000 50.2000 ;
	    RECT 27.4000 48.4000 29.6000 49.0000 ;
	    RECT 30.2000 49.0000 35.6000 49.6000 ;
	    RECT 30.2000 48.8000 31.0000 49.0000 ;
	    RECT 34.8000 48.8000 35.6000 49.0000 ;
	    RECT 28.6000 47.4000 29.4000 47.6000 ;
	    RECT 31.4000 47.4000 32.2000 47.6000 ;
	    RECT 25.2000 46.2000 26.0000 47.0000 ;
	    RECT 28.6000 46.8000 32.2000 47.4000 ;
	    RECT 29.4000 46.2000 30.0000 46.8000 ;
	    RECT 34.8000 46.2000 35.6000 47.0000 ;
	    RECT 24.6000 42.2000 25.8000 46.2000 ;
	    RECT 29.2000 42.2000 30.0000 46.2000 ;
	    RECT 33.6000 45.6000 35.6000 46.2000 ;
	    RECT 33.6000 42.2000 34.4000 45.6000 ;
	    RECT 38.0000 42.2000 38.8000 50.6000 ;
	    RECT 41.6000 50.4000 42.2000 53.6000 ;
	    RECT 42.8000 51.6000 43.6000 53.2000 ;
	    RECT 46.0000 52.3000 46.8000 52.4000 ;
	    RECT 48.0000 52.3000 48.6000 53.6000 ;
	    RECT 46.0000 51.7000 48.6000 52.3000 ;
	    RECT 46.0000 51.6000 46.8000 51.7000 ;
	    RECT 39.6000 50.2000 40.4000 50.4000 ;
	    RECT 39.6000 49.6000 41.0000 50.2000 ;
	    RECT 41.6000 49.6000 43.6000 50.4000 ;
	    RECT 46.0000 50.2000 46.8000 50.4000 ;
	    RECT 48.0000 50.2000 48.6000 51.7000 ;
	    RECT 49.2000 52.3000 50.0000 53.2000 ;
	    RECT 50.8000 52.3000 51.6000 52.4000 ;
	    RECT 49.2000 51.7000 51.6000 52.3000 ;
	    RECT 49.2000 51.6000 50.0000 51.7000 ;
	    RECT 50.8000 51.6000 51.6000 51.7000 ;
	    RECT 52.4000 50.2000 53.2000 50.4000 ;
	    RECT 54.4000 50.2000 55.0000 53.6000 ;
	    RECT 55.6000 51.6000 56.4000 53.2000 ;
	    RECT 58.8000 50.2000 59.6000 50.4000 ;
	    RECT 60.8000 50.2000 61.4000 53.6000 ;
	    RECT 62.0000 51.6000 62.8000 53.2000 ;
	    RECT 65.2000 51.4000 66.0000 54.8000 ;
	    RECT 72.2000 54.2000 73.0000 54.4000 ;
	    RECT 78.0000 54.2000 78.6000 56.4000 ;
	    RECT 82.8000 55.0000 83.6000 59.8000 ;
	    RECT 81.2000 54.2000 82.8000 54.4000 ;
	    RECT 71.8000 53.6000 82.8000 54.2000 ;
	    RECT 70.0000 52.8000 70.8000 53.0000 ;
	    RECT 67.0000 52.2000 70.8000 52.8000 ;
	    RECT 67.0000 52.0000 67.8000 52.2000 ;
	    RECT 68.6000 51.4000 69.4000 51.6000 ;
	    RECT 65.2000 50.8000 69.4000 51.4000 ;
	    RECT 46.0000 49.6000 47.4000 50.2000 ;
	    RECT 48.0000 49.6000 49.0000 50.2000 ;
	    RECT 52.4000 49.6000 53.8000 50.2000 ;
	    RECT 54.4000 49.6000 55.4000 50.2000 ;
	    RECT 58.8000 49.6000 60.2000 50.2000 ;
	    RECT 60.8000 49.6000 61.8000 50.2000 ;
	    RECT 40.4000 48.4000 41.0000 49.6000 ;
	    RECT 39.6000 47.6000 41.2000 48.4000 ;
	    RECT 41.8000 42.2000 42.6000 49.6000 ;
	    RECT 46.8000 48.4000 47.4000 49.6000 ;
	    RECT 46.8000 47.6000 47.6000 48.4000 ;
	    RECT 48.2000 42.2000 49.0000 49.6000 ;
	    RECT 53.2000 48.4000 53.8000 49.6000 ;
	    RECT 53.2000 47.6000 54.0000 48.4000 ;
	    RECT 54.6000 42.2000 55.4000 49.6000 ;
	    RECT 59.6000 48.4000 60.2000 49.6000 ;
	    RECT 59.6000 47.6000 60.4000 48.4000 ;
	    RECT 61.0000 42.2000 61.8000 49.6000 ;
	    RECT 65.2000 42.2000 66.0000 50.8000 ;
	    RECT 71.8000 50.4000 72.4000 53.6000 ;
	    RECT 79.0000 53.4000 79.8000 53.6000 ;
	    RECT 78.0000 52.4000 78.8000 52.6000 ;
	    RECT 80.6000 52.4000 81.4000 52.6000 ;
	    RECT 76.4000 51.8000 81.4000 52.4000 ;
	    RECT 84.4000 52.4000 85.2000 59.8000 ;
	    RECT 87.6000 55.2000 88.4000 59.8000 ;
	    RECT 89.2000 55.8000 90.0000 59.8000 ;
	    RECT 90.8000 56.0000 91.6000 59.8000 ;
	    RECT 94.0000 56.0000 94.8000 59.8000 ;
	    RECT 90.8000 55.8000 94.8000 56.0000 ;
	    RECT 95.6000 55.8000 96.4000 59.8000 ;
	    RECT 97.2000 56.0000 98.0000 59.8000 ;
	    RECT 100.4000 56.0000 101.2000 59.8000 ;
	    RECT 97.2000 55.8000 101.2000 56.0000 ;
	    RECT 86.2000 54.6000 88.4000 55.2000 ;
	    RECT 76.4000 51.6000 77.2000 51.8000 ;
	    RECT 78.0000 51.0000 83.6000 51.2000 ;
	    RECT 77.8000 50.8000 83.6000 51.0000 ;
	    RECT 70.0000 49.8000 72.4000 50.4000 ;
	    RECT 73.8000 50.6000 83.6000 50.8000 ;
	    RECT 73.8000 50.2000 78.6000 50.6000 ;
	    RECT 70.0000 48.8000 70.6000 49.8000 ;
	    RECT 69.2000 48.0000 70.6000 48.8000 ;
	    RECT 72.2000 49.0000 73.0000 49.2000 ;
	    RECT 73.8000 49.0000 74.4000 50.2000 ;
	    RECT 72.2000 48.4000 74.4000 49.0000 ;
	    RECT 75.0000 49.0000 80.4000 49.6000 ;
	    RECT 75.0000 48.8000 75.8000 49.0000 ;
	    RECT 79.6000 48.8000 80.4000 49.0000 ;
	    RECT 73.4000 47.4000 74.2000 47.6000 ;
	    RECT 76.2000 47.4000 77.0000 47.6000 ;
	    RECT 70.0000 46.2000 70.8000 47.0000 ;
	    RECT 73.4000 46.8000 77.0000 47.4000 ;
	    RECT 74.2000 46.2000 74.8000 46.8000 ;
	    RECT 79.6000 46.2000 80.4000 47.0000 ;
	    RECT 69.4000 42.2000 70.6000 46.2000 ;
	    RECT 74.0000 42.2000 74.8000 46.2000 ;
	    RECT 78.4000 45.6000 80.4000 46.2000 ;
	    RECT 78.4000 42.2000 79.2000 45.6000 ;
	    RECT 82.8000 42.2000 83.6000 50.6000 ;
	    RECT 84.4000 50.2000 85.0000 52.4000 ;
	    RECT 86.2000 51.6000 86.8000 54.6000 ;
	    RECT 89.4000 54.4000 90.0000 55.8000 ;
	    RECT 91.0000 55.4000 94.6000 55.8000 ;
	    RECT 93.2000 54.4000 94.0000 54.8000 ;
	    RECT 95.8000 54.4000 96.4000 55.8000 ;
	    RECT 97.4000 55.4000 101.0000 55.8000 ;
	    RECT 99.6000 54.4000 100.4000 54.8000 ;
	    RECT 89.2000 53.6000 91.8000 54.4000 ;
	    RECT 93.2000 53.8000 94.8000 54.4000 ;
	    RECT 94.0000 53.6000 94.8000 53.8000 ;
	    RECT 95.6000 53.6000 98.2000 54.4000 ;
	    RECT 99.6000 53.8000 101.2000 54.4000 ;
	    RECT 100.4000 53.6000 101.2000 53.8000 ;
	    RECT 87.6000 51.6000 88.4000 53.2000 ;
	    RECT 85.6000 50.8000 86.8000 51.6000 ;
	    RECT 86.2000 50.2000 86.8000 50.8000 ;
	    RECT 89.2000 50.2000 90.0000 50.4000 ;
	    RECT 91.2000 50.2000 91.8000 53.6000 ;
	    RECT 92.4000 52.3000 93.2000 53.2000 ;
	    RECT 97.6000 52.4000 98.2000 53.6000 ;
	    RECT 94.0000 52.3000 94.8000 52.4000 ;
	    RECT 92.4000 51.7000 94.8000 52.3000 ;
	    RECT 92.4000 51.6000 93.2000 51.7000 ;
	    RECT 94.0000 51.6000 94.8000 51.7000 ;
	    RECT 97.2000 51.6000 98.2000 52.4000 ;
	    RECT 98.8000 51.6000 99.6000 53.2000 ;
	    RECT 102.0000 52.4000 102.8000 59.8000 ;
	    RECT 105.2000 55.2000 106.0000 59.8000 ;
	    RECT 113.2000 55.8000 114.0000 59.8000 ;
	    RECT 114.8000 56.0000 115.6000 59.8000 ;
	    RECT 118.0000 56.0000 118.8000 59.8000 ;
	    RECT 114.8000 55.8000 118.8000 56.0000 ;
	    RECT 103.8000 54.6000 106.0000 55.2000 ;
	    RECT 95.6000 50.2000 96.4000 50.4000 ;
	    RECT 97.6000 50.2000 98.2000 51.6000 ;
	    RECT 102.0000 50.2000 102.6000 52.4000 ;
	    RECT 103.8000 51.6000 104.4000 54.6000 ;
	    RECT 113.4000 54.4000 114.0000 55.8000 ;
	    RECT 115.0000 55.4000 118.6000 55.8000 ;
	    RECT 117.2000 54.4000 118.0000 54.8000 ;
	    RECT 113.2000 53.6000 115.8000 54.4000 ;
	    RECT 117.2000 54.3000 118.8000 54.4000 ;
	    RECT 119.6000 54.3000 120.4000 59.8000 ;
	    RECT 122.8000 55.2000 123.6000 59.8000 ;
	    RECT 117.2000 53.8000 120.4000 54.3000 ;
	    RECT 118.0000 53.7000 120.4000 53.8000 ;
	    RECT 118.0000 53.6000 118.8000 53.7000 ;
	    RECT 105.2000 51.6000 106.0000 53.2000 ;
	    RECT 106.8000 52.3000 107.6000 52.4000 ;
	    RECT 115.2000 52.3000 115.8000 53.6000 ;
	    RECT 106.8000 51.7000 115.8000 52.3000 ;
	    RECT 106.8000 51.6000 107.6000 51.7000 ;
	    RECT 103.2000 50.8000 104.4000 51.6000 ;
	    RECT 103.8000 50.2000 104.4000 50.8000 ;
	    RECT 113.2000 50.2000 114.0000 50.4000 ;
	    RECT 115.2000 50.2000 115.8000 51.7000 ;
	    RECT 116.4000 51.6000 117.2000 53.2000 ;
	    RECT 119.6000 52.4000 120.4000 53.7000 ;
	    RECT 121.4000 54.6000 123.6000 55.2000 ;
	    RECT 124.4000 55.2000 125.2000 59.8000 ;
	    RECT 124.4000 54.6000 126.6000 55.2000 ;
	    RECT 119.6000 50.2000 120.2000 52.4000 ;
	    RECT 121.4000 51.6000 122.0000 54.6000 ;
	    RECT 120.8000 50.8000 122.0000 51.6000 ;
	    RECT 121.4000 50.2000 122.0000 50.8000 ;
	    RECT 126.0000 51.6000 126.6000 54.6000 ;
	    RECT 127.6000 52.4000 128.4000 59.8000 ;
	    RECT 129.2000 55.8000 130.0000 59.8000 ;
	    RECT 130.8000 56.0000 131.6000 59.8000 ;
	    RECT 134.0000 56.0000 134.8000 59.8000 ;
	    RECT 130.8000 55.8000 134.8000 56.0000 ;
	    RECT 129.4000 54.4000 130.0000 55.8000 ;
	    RECT 131.0000 55.4000 134.6000 55.8000 ;
	    RECT 135.6000 55.4000 136.4000 59.8000 ;
	    RECT 139.8000 58.4000 141.0000 59.8000 ;
	    RECT 139.8000 57.8000 141.2000 58.4000 ;
	    RECT 144.4000 57.8000 145.2000 59.8000 ;
	    RECT 148.8000 58.4000 149.6000 59.8000 ;
	    RECT 148.8000 57.8000 150.8000 58.4000 ;
	    RECT 140.4000 57.0000 141.2000 57.8000 ;
	    RECT 144.6000 57.2000 145.2000 57.8000 ;
	    RECT 144.6000 56.6000 147.4000 57.2000 ;
	    RECT 146.6000 56.4000 147.4000 56.6000 ;
	    RECT 148.4000 56.4000 149.2000 57.2000 ;
	    RECT 150.0000 57.0000 150.8000 57.8000 ;
	    RECT 138.6000 55.4000 139.4000 55.6000 ;
	    RECT 135.6000 54.8000 139.4000 55.4000 ;
	    RECT 133.2000 54.4000 134.0000 54.8000 ;
	    RECT 129.2000 53.6000 131.8000 54.4000 ;
	    RECT 133.2000 53.8000 134.8000 54.4000 ;
	    RECT 134.0000 53.6000 134.8000 53.8000 ;
	    RECT 126.0000 50.8000 127.2000 51.6000 ;
	    RECT 126.0000 50.2000 126.6000 50.8000 ;
	    RECT 127.8000 50.2000 128.4000 52.4000 ;
	    RECT 84.4000 42.2000 85.2000 50.2000 ;
	    RECT 86.2000 49.6000 88.4000 50.2000 ;
	    RECT 89.2000 49.6000 90.6000 50.2000 ;
	    RECT 91.2000 49.6000 92.2000 50.2000 ;
	    RECT 95.6000 49.6000 97.0000 50.2000 ;
	    RECT 97.6000 49.6000 98.6000 50.2000 ;
	    RECT 87.6000 42.2000 88.4000 49.6000 ;
	    RECT 90.0000 48.4000 90.6000 49.6000 ;
	    RECT 90.0000 47.6000 90.8000 48.4000 ;
	    RECT 91.4000 42.2000 92.2000 49.6000 ;
	    RECT 96.4000 48.4000 97.0000 49.6000 ;
	    RECT 96.4000 47.6000 97.2000 48.4000 ;
	    RECT 97.8000 42.2000 98.6000 49.6000 ;
	    RECT 102.0000 42.2000 102.8000 50.2000 ;
	    RECT 103.8000 49.6000 106.0000 50.2000 ;
	    RECT 113.2000 49.6000 114.6000 50.2000 ;
	    RECT 115.2000 49.6000 116.2000 50.2000 ;
	    RECT 105.2000 42.2000 106.0000 49.6000 ;
	    RECT 114.0000 48.4000 114.6000 49.6000 ;
	    RECT 114.0000 47.6000 114.8000 48.4000 ;
	    RECT 115.4000 42.2000 116.2000 49.6000 ;
	    RECT 119.6000 42.2000 120.4000 50.2000 ;
	    RECT 121.4000 49.6000 123.6000 50.2000 ;
	    RECT 122.8000 42.2000 123.6000 49.6000 ;
	    RECT 124.4000 49.6000 126.6000 50.2000 ;
	    RECT 124.4000 42.2000 125.2000 49.6000 ;
	    RECT 127.6000 42.2000 128.4000 50.2000 ;
	    RECT 129.2000 50.2000 130.0000 50.4000 ;
	    RECT 131.2000 50.2000 131.8000 53.6000 ;
	    RECT 132.4000 52.3000 133.2000 53.2000 ;
	    RECT 134.0000 52.3000 134.8000 52.4000 ;
	    RECT 132.4000 51.7000 134.8000 52.3000 ;
	    RECT 132.4000 51.6000 133.2000 51.7000 ;
	    RECT 134.0000 51.6000 134.8000 51.7000 ;
	    RECT 135.6000 51.4000 136.4000 54.8000 ;
	    RECT 142.6000 54.2000 144.4000 54.4000 ;
	    RECT 145.2000 54.2000 146.0000 54.4000 ;
	    RECT 148.4000 54.2000 149.0000 56.4000 ;
	    RECT 153.2000 55.0000 154.0000 59.8000 ;
	    RECT 154.8000 55.8000 155.6000 59.8000 ;
	    RECT 156.4000 56.0000 157.2000 59.8000 ;
	    RECT 159.6000 56.0000 160.4000 59.8000 ;
	    RECT 156.4000 55.8000 160.4000 56.0000 ;
	    RECT 161.2000 55.8000 162.0000 59.8000 ;
	    RECT 162.8000 56.0000 163.6000 59.8000 ;
	    RECT 166.0000 56.0000 166.8000 59.8000 ;
	    RECT 162.8000 55.8000 166.8000 56.0000 ;
	    RECT 167.6000 55.8000 168.4000 59.8000 ;
	    RECT 169.2000 56.0000 170.0000 59.8000 ;
	    RECT 172.4000 56.0000 173.2000 59.8000 ;
	    RECT 169.2000 55.8000 173.2000 56.0000 ;
	    RECT 174.0000 55.8000 174.8000 59.8000 ;
	    RECT 175.6000 56.0000 176.4000 59.8000 ;
	    RECT 178.8000 56.0000 179.6000 59.8000 ;
	    RECT 175.6000 55.8000 179.6000 56.0000 ;
	    RECT 180.4000 55.8000 181.2000 59.8000 ;
	    RECT 182.0000 56.0000 182.8000 59.8000 ;
	    RECT 185.2000 56.0000 186.0000 59.8000 ;
	    RECT 182.0000 55.8000 186.0000 56.0000 ;
	    RECT 186.8000 56.0000 187.6000 59.8000 ;
	    RECT 190.0000 56.0000 190.8000 59.8000 ;
	    RECT 186.8000 55.8000 190.8000 56.0000 ;
	    RECT 191.6000 55.8000 192.4000 59.8000 ;
	    RECT 193.2000 55.8000 194.0000 59.8000 ;
	    RECT 194.8000 56.0000 195.6000 59.8000 ;
	    RECT 198.0000 56.0000 198.8000 59.8000 ;
	    RECT 194.8000 55.8000 198.8000 56.0000 ;
	    RECT 199.6000 55.8000 200.4000 59.8000 ;
	    RECT 201.2000 56.0000 202.0000 59.8000 ;
	    RECT 204.4000 56.0000 205.2000 59.8000 ;
	    RECT 201.2000 55.8000 205.2000 56.0000 ;
	    RECT 206.0000 55.8000 206.8000 59.8000 ;
	    RECT 207.6000 56.0000 208.4000 59.8000 ;
	    RECT 210.8000 56.0000 211.6000 59.8000 ;
	    RECT 207.6000 55.8000 211.6000 56.0000 ;
	    RECT 155.0000 54.4000 155.6000 55.8000 ;
	    RECT 156.6000 55.4000 160.2000 55.8000 ;
	    RECT 158.8000 54.4000 159.6000 54.8000 ;
	    RECT 161.4000 54.4000 162.0000 55.8000 ;
	    RECT 163.0000 55.4000 166.6000 55.8000 ;
	    RECT 165.2000 54.4000 166.0000 54.8000 ;
	    RECT 167.8000 54.4000 168.4000 55.8000 ;
	    RECT 169.4000 55.4000 173.0000 55.8000 ;
	    RECT 171.6000 54.4000 172.4000 54.8000 ;
	    RECT 174.2000 54.4000 174.8000 55.8000 ;
	    RECT 175.8000 55.4000 179.4000 55.8000 ;
	    RECT 178.0000 54.4000 178.8000 54.8000 ;
	    RECT 180.6000 54.4000 181.2000 55.8000 ;
	    RECT 182.2000 55.4000 185.8000 55.8000 ;
	    RECT 187.0000 55.4000 190.6000 55.8000 ;
	    RECT 184.4000 54.4000 185.2000 54.8000 ;
	    RECT 187.6000 54.4000 188.4000 54.8000 ;
	    RECT 191.6000 54.4000 192.2000 55.8000 ;
	    RECT 193.4000 54.4000 194.0000 55.8000 ;
	    RECT 195.0000 55.4000 198.6000 55.8000 ;
	    RECT 197.2000 54.4000 198.0000 54.8000 ;
	    RECT 199.8000 54.4000 200.4000 55.8000 ;
	    RECT 201.4000 55.4000 205.0000 55.8000 ;
	    RECT 203.6000 54.4000 204.4000 54.8000 ;
	    RECT 206.2000 54.4000 206.8000 55.8000 ;
	    RECT 207.8000 55.4000 211.4000 55.8000 ;
	    RECT 212.4000 55.6000 213.2000 59.8000 ;
	    RECT 214.0000 56.0000 214.8000 59.8000 ;
	    RECT 217.2000 56.0000 218.0000 59.8000 ;
	    RECT 214.0000 55.8000 218.0000 56.0000 ;
	    RECT 218.8000 55.8000 219.6000 59.8000 ;
	    RECT 220.4000 56.0000 221.2000 59.8000 ;
	    RECT 223.6000 56.0000 224.4000 59.8000 ;
	    RECT 220.4000 55.8000 224.4000 56.0000 ;
	    RECT 225.2000 59.2000 229.2000 59.8000 ;
	    RECT 225.2000 55.8000 226.0000 59.2000 ;
	    RECT 210.0000 54.4000 210.8000 54.8000 ;
	    RECT 212.6000 54.4000 213.2000 55.6000 ;
	    RECT 214.2000 55.4000 217.8000 55.8000 ;
	    RECT 216.4000 54.4000 217.2000 54.8000 ;
	    RECT 219.0000 54.4000 219.6000 55.8000 ;
	    RECT 220.6000 55.4000 224.2000 55.8000 ;
	    RECT 226.8000 55.6000 227.6000 58.6000 ;
	    RECT 228.4000 56.0000 229.2000 59.2000 ;
	    RECT 231.6000 56.0000 232.4000 59.8000 ;
	    RECT 228.4000 55.8000 232.4000 56.0000 ;
	    RECT 233.2000 55.8000 234.0000 59.8000 ;
	    RECT 234.8000 56.0000 235.6000 59.8000 ;
	    RECT 238.0000 56.0000 238.8000 59.8000 ;
	    RECT 241.2000 57.8000 242.0000 59.8000 ;
	    RECT 234.8000 55.8000 238.8000 56.0000 ;
	    RECT 222.8000 54.4000 223.6000 54.8000 ;
	    RECT 226.8000 54.4000 227.4000 55.6000 ;
	    RECT 228.6000 55.4000 232.2000 55.8000 ;
	    RECT 230.8000 54.4000 231.6000 54.8000 ;
	    RECT 233.4000 54.4000 234.0000 55.8000 ;
	    RECT 235.0000 55.4000 238.6000 55.8000 ;
	    RECT 239.6000 55.6000 240.4000 57.2000 ;
	    RECT 237.2000 54.4000 238.0000 54.8000 ;
	    RECT 241.4000 54.4000 242.0000 57.8000 ;
	    RECT 244.4000 55.2000 245.2000 59.8000 ;
	    RECT 244.4000 54.6000 246.6000 55.2000 ;
	    RECT 151.6000 54.2000 153.2000 54.4000 ;
	    RECT 142.2000 53.6000 153.2000 54.2000 ;
	    RECT 154.8000 53.6000 157.4000 54.4000 ;
	    RECT 158.8000 53.8000 160.4000 54.4000 ;
	    RECT 159.6000 53.6000 160.4000 53.8000 ;
	    RECT 161.2000 53.6000 163.8000 54.4000 ;
	    RECT 165.2000 53.8000 166.8000 54.4000 ;
	    RECT 166.0000 53.6000 166.8000 53.8000 ;
	    RECT 167.6000 53.6000 170.2000 54.4000 ;
	    RECT 171.6000 53.8000 173.2000 54.4000 ;
	    RECT 172.4000 53.6000 173.2000 53.8000 ;
	    RECT 174.0000 53.6000 176.6000 54.4000 ;
	    RECT 178.0000 53.8000 179.6000 54.4000 ;
	    RECT 178.8000 53.6000 179.6000 53.8000 ;
	    RECT 180.4000 53.6000 183.0000 54.4000 ;
	    RECT 184.4000 53.8000 186.0000 54.4000 ;
	    RECT 185.2000 53.6000 186.0000 53.8000 ;
	    RECT 186.8000 53.8000 188.4000 54.4000 ;
	    RECT 186.8000 53.6000 187.6000 53.8000 ;
	    RECT 189.8000 53.6000 192.4000 54.4000 ;
	    RECT 193.2000 53.6000 195.8000 54.4000 ;
	    RECT 197.2000 53.8000 198.8000 54.4000 ;
	    RECT 198.0000 53.6000 198.8000 53.8000 ;
	    RECT 199.6000 53.6000 202.2000 54.4000 ;
	    RECT 203.6000 53.8000 205.2000 54.4000 ;
	    RECT 204.4000 53.6000 205.2000 53.8000 ;
	    RECT 206.0000 53.6000 208.6000 54.4000 ;
	    RECT 210.0000 53.8000 211.6000 54.4000 ;
	    RECT 210.8000 53.6000 211.6000 53.8000 ;
	    RECT 212.4000 53.6000 215.0000 54.4000 ;
	    RECT 216.4000 53.8000 218.0000 54.4000 ;
	    RECT 217.2000 53.6000 218.0000 53.8000 ;
	    RECT 218.8000 53.6000 221.4000 54.4000 ;
	    RECT 222.8000 53.8000 224.4000 54.4000 ;
	    RECT 223.6000 53.6000 224.4000 53.8000 ;
	    RECT 140.4000 52.8000 141.2000 53.0000 ;
	    RECT 137.4000 52.2000 141.2000 52.8000 ;
	    RECT 142.2000 52.4000 142.8000 53.6000 ;
	    RECT 149.4000 53.4000 150.2000 53.6000 ;
	    RECT 148.4000 52.4000 149.2000 52.6000 ;
	    RECT 151.0000 52.4000 151.8000 52.6000 ;
	    RECT 137.4000 52.0000 138.2000 52.2000 ;
	    RECT 142.0000 51.6000 142.8000 52.4000 ;
	    RECT 146.8000 51.8000 151.8000 52.4000 ;
	    RECT 146.8000 51.6000 147.6000 51.8000 ;
	    RECT 139.0000 51.4000 139.8000 51.6000 ;
	    RECT 135.6000 50.8000 139.8000 51.4000 ;
	    RECT 129.2000 49.6000 130.6000 50.2000 ;
	    RECT 131.2000 49.6000 132.2000 50.2000 ;
	    RECT 130.0000 48.4000 130.6000 49.6000 ;
	    RECT 130.0000 47.6000 130.8000 48.4000 ;
	    RECT 131.4000 44.4000 132.2000 49.6000 ;
	    RECT 131.4000 43.6000 133.2000 44.4000 ;
	    RECT 131.4000 42.2000 132.2000 43.6000 ;
	    RECT 135.6000 42.2000 136.4000 50.8000 ;
	    RECT 142.2000 50.4000 142.8000 51.6000 ;
	    RECT 148.4000 51.0000 154.0000 51.2000 ;
	    RECT 148.2000 50.8000 154.0000 51.0000 ;
	    RECT 140.4000 49.8000 142.8000 50.4000 ;
	    RECT 144.2000 50.6000 154.0000 50.8000 ;
	    RECT 144.2000 50.2000 149.0000 50.6000 ;
	    RECT 140.4000 48.8000 141.0000 49.8000 ;
	    RECT 139.6000 48.0000 141.0000 48.8000 ;
	    RECT 142.6000 49.0000 143.4000 49.2000 ;
	    RECT 144.2000 49.0000 144.8000 50.2000 ;
	    RECT 142.6000 48.4000 144.8000 49.0000 ;
	    RECT 145.4000 49.0000 150.8000 49.6000 ;
	    RECT 145.4000 48.8000 146.2000 49.0000 ;
	    RECT 150.0000 48.8000 150.8000 49.0000 ;
	    RECT 143.8000 47.4000 144.6000 47.6000 ;
	    RECT 146.6000 47.4000 147.4000 47.6000 ;
	    RECT 140.4000 46.2000 141.2000 47.0000 ;
	    RECT 143.8000 46.8000 147.4000 47.4000 ;
	    RECT 144.6000 46.2000 145.2000 46.8000 ;
	    RECT 150.0000 46.2000 150.8000 47.0000 ;
	    RECT 139.8000 42.2000 141.0000 46.2000 ;
	    RECT 144.4000 42.2000 145.2000 46.2000 ;
	    RECT 148.8000 45.6000 150.8000 46.2000 ;
	    RECT 148.8000 42.2000 149.6000 45.6000 ;
	    RECT 153.2000 42.2000 154.0000 50.6000 ;
	    RECT 154.8000 50.2000 155.6000 50.4000 ;
	    RECT 156.8000 50.2000 157.4000 53.6000 ;
	    RECT 158.0000 52.3000 158.8000 53.2000 ;
	    RECT 159.6000 52.3000 160.4000 52.4000 ;
	    RECT 158.0000 51.7000 160.4000 52.3000 ;
	    RECT 158.0000 51.6000 158.8000 51.7000 ;
	    RECT 159.6000 51.6000 160.4000 51.7000 ;
	    RECT 161.2000 50.2000 162.0000 50.4000 ;
	    RECT 163.2000 50.2000 163.8000 53.6000 ;
	    RECT 164.4000 52.3000 165.2000 53.2000 ;
	    RECT 169.6000 52.3000 170.2000 53.6000 ;
	    RECT 164.4000 51.7000 170.2000 52.3000 ;
	    RECT 164.4000 51.6000 165.2000 51.7000 ;
	    RECT 167.6000 50.2000 168.4000 50.4000 ;
	    RECT 169.6000 50.2000 170.2000 51.7000 ;
	    RECT 170.8000 51.6000 171.6000 53.2000 ;
	    RECT 172.4000 52.3000 173.2000 52.4000 ;
	    RECT 176.0000 52.3000 176.6000 53.6000 ;
	    RECT 172.4000 51.7000 176.6000 52.3000 ;
	    RECT 172.4000 51.6000 173.2000 51.7000 ;
	    RECT 174.0000 50.2000 174.8000 50.4000 ;
	    RECT 176.0000 50.2000 176.6000 51.7000 ;
	    RECT 177.2000 52.3000 178.0000 53.2000 ;
	    RECT 182.4000 52.3000 183.0000 53.6000 ;
	    RECT 177.2000 51.7000 183.0000 52.3000 ;
	    RECT 177.2000 51.6000 178.0000 51.7000 ;
	    RECT 180.4000 50.2000 181.2000 50.4000 ;
	    RECT 182.4000 50.2000 183.0000 51.7000 ;
	    RECT 183.6000 52.3000 184.4000 53.2000 ;
	    RECT 185.2000 52.3000 186.0000 52.4000 ;
	    RECT 183.6000 51.7000 186.0000 52.3000 ;
	    RECT 183.6000 51.6000 184.4000 51.7000 ;
	    RECT 185.2000 51.6000 186.0000 51.7000 ;
	    RECT 186.8000 52.3000 187.6000 52.4000 ;
	    RECT 188.4000 52.3000 189.2000 53.2000 ;
	    RECT 186.8000 51.7000 189.2000 52.3000 ;
	    RECT 186.8000 51.6000 187.6000 51.7000 ;
	    RECT 188.4000 51.6000 189.2000 51.7000 ;
	    RECT 189.8000 50.2000 190.4000 53.6000 ;
	    RECT 195.2000 52.4000 195.8000 53.6000 ;
	    RECT 194.8000 51.6000 195.8000 52.4000 ;
	    RECT 196.4000 51.6000 197.2000 53.2000 ;
	    RECT 191.6000 50.2000 192.4000 50.4000 ;
	    RECT 154.8000 49.6000 156.2000 50.2000 ;
	    RECT 156.8000 49.6000 157.8000 50.2000 ;
	    RECT 161.2000 49.6000 162.6000 50.2000 ;
	    RECT 163.2000 49.6000 164.2000 50.2000 ;
	    RECT 167.6000 49.6000 169.0000 50.2000 ;
	    RECT 169.6000 49.6000 170.6000 50.2000 ;
	    RECT 174.0000 49.6000 175.4000 50.2000 ;
	    RECT 176.0000 49.6000 177.0000 50.2000 ;
	    RECT 180.4000 49.6000 181.8000 50.2000 ;
	    RECT 182.4000 49.6000 183.4000 50.2000 ;
	    RECT 155.6000 48.4000 156.2000 49.6000 ;
	    RECT 157.0000 48.4000 157.8000 49.6000 ;
	    RECT 162.0000 48.4000 162.6000 49.6000 ;
	    RECT 155.6000 47.6000 156.4000 48.4000 ;
	    RECT 157.0000 47.6000 158.8000 48.4000 ;
	    RECT 162.0000 47.6000 162.8000 48.4000 ;
	    RECT 157.0000 42.2000 157.8000 47.6000 ;
	    RECT 163.4000 42.2000 164.2000 49.6000 ;
	    RECT 168.4000 48.4000 169.0000 49.6000 ;
	    RECT 168.4000 47.6000 169.2000 48.4000 ;
	    RECT 169.8000 42.2000 170.6000 49.6000 ;
	    RECT 174.8000 48.4000 175.4000 49.6000 ;
	    RECT 174.8000 47.6000 175.6000 48.4000 ;
	    RECT 176.2000 42.2000 177.0000 49.6000 ;
	    RECT 181.2000 48.4000 181.8000 49.6000 ;
	    RECT 181.2000 47.6000 182.0000 48.4000 ;
	    RECT 182.6000 42.2000 183.4000 49.6000 ;
	    RECT 189.4000 49.6000 190.4000 50.2000 ;
	    RECT 191.0000 49.6000 192.4000 50.2000 ;
	    RECT 193.2000 50.2000 194.0000 50.4000 ;
	    RECT 195.2000 50.2000 195.8000 51.6000 ;
	    RECT 199.6000 50.2000 200.4000 50.4000 ;
	    RECT 201.6000 50.2000 202.2000 53.6000 ;
	    RECT 202.8000 51.6000 203.6000 53.2000 ;
	    RECT 204.4000 52.3000 205.2000 52.4000 ;
	    RECT 208.0000 52.3000 208.6000 53.6000 ;
	    RECT 204.4000 51.7000 208.6000 52.3000 ;
	    RECT 204.4000 51.6000 205.2000 51.7000 ;
	    RECT 206.0000 50.2000 206.8000 50.4000 ;
	    RECT 208.0000 50.2000 208.6000 51.7000 ;
	    RECT 209.2000 52.3000 210.0000 53.2000 ;
	    RECT 210.8000 52.3000 211.6000 52.4000 ;
	    RECT 209.2000 51.7000 211.6000 52.3000 ;
	    RECT 209.2000 51.6000 210.0000 51.7000 ;
	    RECT 210.8000 51.6000 211.6000 51.7000 ;
	    RECT 212.4000 50.2000 213.2000 50.4000 ;
	    RECT 214.4000 50.2000 215.0000 53.6000 ;
	    RECT 215.6000 51.6000 216.4000 53.2000 ;
	    RECT 218.8000 50.2000 219.6000 50.4000 ;
	    RECT 220.8000 50.2000 221.4000 53.6000 ;
	    RECT 222.0000 51.6000 222.8000 53.2000 ;
	    RECT 225.2000 52.8000 226.0000 54.4000 ;
	    RECT 226.8000 53.8000 229.2000 54.4000 ;
	    RECT 230.8000 54.3000 232.4000 54.4000 ;
	    RECT 233.2000 54.3000 235.8000 54.4000 ;
	    RECT 230.8000 53.8000 235.8000 54.3000 ;
	    RECT 237.2000 53.8000 238.8000 54.4000 ;
	    RECT 228.4000 53.6000 229.2000 53.8000 ;
	    RECT 231.6000 53.7000 235.8000 53.8000 ;
	    RECT 231.6000 53.6000 232.4000 53.7000 ;
	    RECT 233.2000 53.6000 235.8000 53.7000 ;
	    RECT 238.0000 53.6000 238.8000 53.8000 ;
	    RECT 241.2000 53.6000 242.0000 54.4000 ;
	    RECT 226.8000 51.6000 227.6000 53.2000 ;
	    RECT 228.6000 50.2000 229.2000 53.6000 ;
	    RECT 230.0000 52.3000 230.8000 53.2000 ;
	    RECT 233.2000 52.3000 234.0000 52.4000 ;
	    RECT 230.0000 51.7000 234.0000 52.3000 ;
	    RECT 230.0000 51.6000 230.8000 51.7000 ;
	    RECT 233.2000 51.6000 234.0000 51.7000 ;
	    RECT 233.2000 50.2000 234.0000 50.4000 ;
	    RECT 235.2000 50.2000 235.8000 53.6000 ;
	    RECT 236.4000 51.6000 237.2000 53.2000 ;
	    RECT 239.6000 52.3000 240.4000 52.4000 ;
	    RECT 241.4000 52.3000 242.0000 53.6000 ;
	    RECT 239.6000 51.7000 242.0000 52.3000 ;
	    RECT 239.6000 51.6000 240.4000 51.7000 ;
	    RECT 241.4000 50.2000 242.0000 51.7000 ;
	    RECT 242.8000 50.8000 243.6000 52.4000 ;
	    RECT 246.0000 51.6000 246.6000 54.6000 ;
	    RECT 247.6000 52.4000 248.4000 59.8000 ;
	    RECT 249.8000 58.4000 250.6000 59.8000 ;
	    RECT 263.0000 58.4000 263.8000 59.8000 ;
	    RECT 265.2000 59.2000 269.2000 59.8000 ;
	    RECT 249.8000 57.6000 251.6000 58.4000 ;
	    RECT 263.0000 57.6000 264.4000 58.4000 ;
	    RECT 249.8000 56.4000 250.6000 57.6000 ;
	    RECT 263.0000 56.4000 263.8000 57.6000 ;
	    RECT 249.8000 55.8000 251.6000 56.4000 ;
	    RECT 246.0000 50.8000 247.2000 51.6000 ;
	    RECT 246.0000 50.2000 246.6000 50.8000 ;
	    RECT 247.8000 50.2000 248.4000 52.4000 ;
	    RECT 193.2000 49.6000 194.6000 50.2000 ;
	    RECT 195.2000 49.6000 196.2000 50.2000 ;
	    RECT 199.6000 49.6000 201.0000 50.2000 ;
	    RECT 201.6000 49.6000 202.6000 50.2000 ;
	    RECT 206.0000 49.6000 207.4000 50.2000 ;
	    RECT 208.0000 49.6000 209.0000 50.2000 ;
	    RECT 212.4000 49.6000 213.8000 50.2000 ;
	    RECT 214.4000 49.6000 215.4000 50.2000 ;
	    RECT 218.8000 49.6000 220.2000 50.2000 ;
	    RECT 220.8000 49.6000 221.8000 50.2000 ;
	    RECT 189.4000 42.2000 190.2000 49.6000 ;
	    RECT 191.0000 48.4000 191.6000 49.6000 ;
	    RECT 194.0000 48.4000 194.6000 49.6000 ;
	    RECT 190.8000 47.6000 192.4000 48.4000 ;
	    RECT 194.0000 47.6000 194.8000 48.4000 ;
	    RECT 195.4000 42.2000 196.2000 49.6000 ;
	    RECT 200.4000 48.4000 201.0000 49.6000 ;
	    RECT 201.8000 48.4000 202.6000 49.6000 ;
	    RECT 206.8000 48.4000 207.4000 49.6000 ;
	    RECT 200.4000 47.6000 201.2000 48.4000 ;
	    RECT 201.8000 47.6000 203.6000 48.4000 ;
	    RECT 206.8000 47.6000 207.6000 48.4000 ;
	    RECT 201.8000 42.2000 202.6000 47.6000 ;
	    RECT 208.2000 42.2000 209.0000 49.6000 ;
	    RECT 213.2000 48.4000 213.8000 49.6000 ;
	    RECT 213.2000 47.6000 214.0000 48.4000 ;
	    RECT 214.6000 42.2000 215.4000 49.6000 ;
	    RECT 219.6000 48.4000 220.2000 49.6000 ;
	    RECT 219.6000 47.6000 220.4000 48.4000 ;
	    RECT 221.0000 42.2000 221.8000 49.6000 ;
	    RECT 227.8000 42.2000 229.8000 50.2000 ;
	    RECT 233.2000 49.6000 234.6000 50.2000 ;
	    RECT 235.2000 49.6000 236.2000 50.2000 ;
	    RECT 234.0000 48.4000 234.6000 49.6000 ;
	    RECT 234.0000 47.6000 234.8000 48.4000 ;
	    RECT 235.4000 42.2000 236.2000 49.6000 ;
	    RECT 241.2000 49.4000 243.0000 50.2000 ;
	    RECT 242.2000 42.2000 243.0000 49.4000 ;
	    RECT 244.4000 49.6000 246.6000 50.2000 ;
	    RECT 244.4000 42.2000 245.2000 49.6000 ;
	    RECT 247.6000 42.2000 248.4000 50.2000 ;
	    RECT 249.2000 48.8000 250.0000 50.4000 ;
	    RECT 250.8000 42.2000 251.6000 55.8000 ;
	    RECT 262.0000 55.8000 263.8000 56.4000 ;
	    RECT 265.2000 55.8000 266.0000 59.2000 ;
	    RECT 266.8000 55.8000 267.6000 58.6000 ;
	    RECT 268.4000 56.0000 269.2000 59.2000 ;
	    RECT 271.6000 56.0000 272.4000 59.8000 ;
	    RECT 268.4000 55.8000 272.4000 56.0000 ;
	    RECT 273.2000 55.8000 274.0000 59.8000 ;
	    RECT 274.8000 56.0000 275.6000 59.8000 ;
	    RECT 278.0000 56.0000 278.8000 59.8000 ;
	    RECT 274.8000 55.8000 278.8000 56.0000 ;
	    RECT 279.6000 55.8000 280.4000 59.8000 ;
	    RECT 281.2000 56.0000 282.0000 59.8000 ;
	    RECT 284.4000 56.0000 285.2000 59.8000 ;
	    RECT 281.2000 55.8000 285.2000 56.0000 ;
	    RECT 287.6000 57.8000 288.4000 59.8000 ;
	    RECT 290.8000 59.2000 294.8000 59.8000 ;
	    RECT 252.4000 54.3000 253.2000 55.2000 ;
	    RECT 254.0000 54.3000 254.8000 54.4000 ;
	    RECT 252.4000 53.7000 254.8000 54.3000 ;
	    RECT 252.4000 53.6000 253.2000 53.7000 ;
	    RECT 254.0000 53.6000 254.8000 53.7000 ;
	    RECT 260.4000 53.6000 261.2000 55.2000 ;
	    RECT 262.0000 42.2000 262.8000 55.8000 ;
	    RECT 266.8000 54.4000 267.4000 55.8000 ;
	    RECT 268.6000 55.4000 272.2000 55.8000 ;
	    RECT 270.8000 54.4000 271.6000 54.8000 ;
	    RECT 273.4000 54.4000 274.0000 55.8000 ;
	    RECT 275.0000 55.4000 278.6000 55.8000 ;
	    RECT 277.2000 54.4000 278.0000 54.8000 ;
	    RECT 279.8000 54.4000 280.4000 55.8000 ;
	    RECT 281.4000 55.4000 285.0000 55.8000 ;
	    RECT 283.6000 54.4000 284.4000 54.8000 ;
	    RECT 287.6000 54.4000 288.2000 57.8000 ;
	    RECT 289.2000 55.6000 290.0000 57.2000 ;
	    RECT 290.8000 55.8000 291.6000 59.2000 ;
	    RECT 292.4000 55.8000 293.2000 58.6000 ;
	    RECT 294.0000 56.0000 294.8000 59.2000 ;
	    RECT 297.2000 56.0000 298.0000 59.8000 ;
	    RECT 294.0000 55.8000 298.0000 56.0000 ;
	    RECT 298.8000 55.8000 299.6000 59.8000 ;
	    RECT 300.4000 56.0000 301.2000 59.8000 ;
	    RECT 303.6000 56.0000 304.4000 59.8000 ;
	    RECT 300.4000 55.8000 304.4000 56.0000 ;
	    RECT 306.8000 57.6000 307.6000 59.8000 ;
	    RECT 292.4000 54.4000 293.0000 55.8000 ;
	    RECT 294.2000 55.4000 297.8000 55.8000 ;
	    RECT 296.4000 54.4000 297.2000 54.8000 ;
	    RECT 299.0000 54.4000 299.6000 55.8000 ;
	    RECT 300.6000 55.4000 304.2000 55.8000 ;
	    RECT 302.8000 54.4000 303.6000 54.8000 ;
	    RECT 306.8000 54.4000 307.4000 57.6000 ;
	    RECT 308.4000 55.6000 309.2000 57.2000 ;
	    RECT 310.0000 56.0000 310.8000 59.8000 ;
	    RECT 313.2000 56.0000 314.0000 59.8000 ;
	    RECT 310.0000 55.8000 314.0000 56.0000 ;
	    RECT 314.8000 55.8000 315.6000 59.8000 ;
	    RECT 316.4000 56.0000 317.2000 59.8000 ;
	    RECT 319.6000 59.2000 323.6000 59.8000 ;
	    RECT 319.6000 56.0000 320.4000 59.2000 ;
	    RECT 316.4000 55.8000 320.4000 56.0000 ;
	    RECT 321.2000 55.8000 322.0000 58.6000 ;
	    RECT 322.8000 55.8000 323.6000 59.2000 ;
	    RECT 326.0000 57.8000 326.8000 59.8000 ;
	    RECT 310.2000 55.4000 313.8000 55.8000 ;
	    RECT 310.8000 54.4000 311.6000 54.8000 ;
	    RECT 314.8000 54.4000 315.4000 55.8000 ;
	    RECT 316.6000 55.4000 320.2000 55.8000 ;
	    RECT 317.2000 54.4000 318.0000 54.8000 ;
	    RECT 321.4000 54.4000 322.0000 55.8000 ;
	    RECT 324.4000 55.6000 325.2000 57.2000 ;
	    RECT 326.2000 56.4000 326.8000 57.8000 ;
	    RECT 326.0000 55.6000 326.8000 56.4000 ;
	    RECT 326.2000 54.4000 326.8000 55.6000 ;
	    RECT 265.2000 52.8000 266.0000 54.4000 ;
	    RECT 266.8000 53.8000 269.2000 54.4000 ;
	    RECT 270.8000 54.3000 272.4000 54.4000 ;
	    RECT 273.2000 54.3000 275.8000 54.4000 ;
	    RECT 270.8000 53.8000 275.8000 54.3000 ;
	    RECT 277.2000 53.8000 278.8000 54.4000 ;
	    RECT 268.4000 53.6000 269.2000 53.8000 ;
	    RECT 271.6000 53.7000 275.8000 53.8000 ;
	    RECT 271.6000 53.6000 272.4000 53.7000 ;
	    RECT 273.2000 53.6000 275.8000 53.7000 ;
	    RECT 278.0000 53.6000 278.8000 53.8000 ;
	    RECT 279.6000 53.6000 282.2000 54.4000 ;
	    RECT 283.6000 54.3000 285.2000 54.4000 ;
	    RECT 286.0000 54.3000 286.8000 54.4000 ;
	    RECT 283.6000 53.8000 286.8000 54.3000 ;
	    RECT 284.4000 53.7000 286.8000 53.8000 ;
	    RECT 284.4000 53.6000 285.2000 53.7000 ;
	    RECT 286.0000 53.6000 286.8000 53.7000 ;
	    RECT 287.6000 53.6000 288.4000 54.4000 ;
	    RECT 266.8000 51.6000 267.6000 53.2000 ;
	    RECT 268.6000 50.4000 269.2000 53.6000 ;
	    RECT 270.0000 51.6000 270.8000 53.2000 ;
	    RECT 263.6000 48.8000 264.4000 50.4000 ;
	    RECT 268.4000 50.2000 269.2000 50.4000 ;
	    RECT 273.2000 50.2000 274.0000 50.4000 ;
	    RECT 275.2000 50.2000 275.8000 53.6000 ;
	    RECT 276.4000 51.6000 277.2000 53.2000 ;
	    RECT 279.6000 50.2000 280.4000 50.4000 ;
	    RECT 281.6000 50.2000 282.2000 53.6000 ;
	    RECT 282.8000 51.6000 283.6000 53.2000 ;
	    RECT 286.0000 50.8000 286.8000 52.4000 ;
	    RECT 287.6000 50.2000 288.2000 53.6000 ;
	    RECT 290.8000 52.8000 291.6000 54.4000 ;
	    RECT 292.4000 53.8000 294.8000 54.4000 ;
	    RECT 296.4000 54.3000 298.0000 54.4000 ;
	    RECT 298.8000 54.3000 301.4000 54.4000 ;
	    RECT 296.4000 53.8000 301.4000 54.3000 ;
	    RECT 302.8000 54.3000 304.4000 54.4000 ;
	    RECT 305.2000 54.3000 306.0000 54.4000 ;
	    RECT 302.8000 53.8000 306.0000 54.3000 ;
	    RECT 294.0000 53.6000 294.8000 53.8000 ;
	    RECT 297.2000 53.7000 301.4000 53.8000 ;
	    RECT 297.2000 53.6000 298.0000 53.7000 ;
	    RECT 298.8000 53.6000 301.4000 53.7000 ;
	    RECT 303.6000 53.7000 306.0000 53.8000 ;
	    RECT 303.6000 53.6000 304.4000 53.7000 ;
	    RECT 305.2000 53.6000 306.0000 53.7000 ;
	    RECT 306.8000 53.6000 307.6000 54.4000 ;
	    RECT 310.0000 53.8000 311.6000 54.4000 ;
	    RECT 313.0000 54.3000 315.6000 54.4000 ;
	    RECT 316.4000 54.3000 318.0000 54.4000 ;
	    RECT 313.0000 53.8000 318.0000 54.3000 ;
	    RECT 319.6000 53.8000 322.0000 54.4000 ;
	    RECT 322.8000 54.3000 323.6000 54.4000 ;
	    RECT 324.4000 54.3000 325.2000 54.4000 ;
	    RECT 310.0000 53.6000 310.8000 53.8000 ;
	    RECT 313.0000 53.7000 317.2000 53.8000 ;
	    RECT 313.0000 53.6000 315.6000 53.7000 ;
	    RECT 316.4000 53.6000 317.2000 53.7000 ;
	    RECT 319.6000 53.6000 320.4000 53.8000 ;
	    RECT 322.8000 53.7000 325.2000 54.3000 ;
	    RECT 292.4000 51.6000 293.2000 53.2000 ;
	    RECT 294.2000 50.2000 294.8000 53.6000 ;
	    RECT 295.6000 51.6000 296.4000 53.2000 ;
	    RECT 298.8000 50.2000 299.6000 50.4000 ;
	    RECT 300.8000 50.2000 301.4000 53.6000 ;
	    RECT 302.0000 51.6000 302.8000 53.2000 ;
	    RECT 303.6000 52.3000 304.4000 52.4000 ;
	    RECT 305.2000 52.3000 306.0000 52.4000 ;
	    RECT 303.6000 51.7000 306.0000 52.3000 ;
	    RECT 303.6000 51.6000 304.4000 51.7000 ;
	    RECT 305.2000 50.8000 306.0000 51.7000 ;
	    RECT 306.8000 50.2000 307.4000 53.6000 ;
	    RECT 311.6000 51.6000 312.4000 53.2000 ;
	    RECT 313.0000 50.2000 313.6000 53.6000 ;
	    RECT 318.0000 51.6000 318.8000 53.2000 ;
	    RECT 319.6000 50.4000 320.2000 53.6000 ;
	    RECT 321.2000 51.6000 322.0000 53.2000 ;
	    RECT 322.8000 52.8000 323.6000 53.7000 ;
	    RECT 324.4000 53.6000 325.2000 53.7000 ;
	    RECT 326.0000 53.6000 326.8000 54.4000 ;
	    RECT 314.8000 50.2000 315.6000 50.4000 ;
	    RECT 267.8000 42.2000 269.8000 50.2000 ;
	    RECT 273.2000 49.6000 274.6000 50.2000 ;
	    RECT 275.2000 49.6000 276.2000 50.2000 ;
	    RECT 279.6000 49.6000 281.0000 50.2000 ;
	    RECT 281.6000 49.6000 282.6000 50.2000 ;
	    RECT 274.0000 48.4000 274.6000 49.6000 ;
	    RECT 274.0000 47.6000 274.8000 48.4000 ;
	    RECT 275.4000 42.2000 276.2000 49.6000 ;
	    RECT 280.4000 48.4000 281.0000 49.6000 ;
	    RECT 280.4000 47.6000 281.2000 48.4000 ;
	    RECT 281.8000 42.2000 282.6000 49.6000 ;
	    RECT 286.6000 49.4000 288.4000 50.2000 ;
	    RECT 286.6000 48.4000 287.4000 49.4000 ;
	    RECT 286.0000 47.6000 287.4000 48.4000 ;
	    RECT 286.6000 42.2000 287.4000 47.6000 ;
	    RECT 293.4000 44.4000 295.4000 50.2000 ;
	    RECT 298.8000 49.6000 300.2000 50.2000 ;
	    RECT 300.8000 49.6000 301.8000 50.2000 ;
	    RECT 299.6000 48.4000 300.2000 49.6000 ;
	    RECT 299.6000 47.6000 300.4000 48.4000 ;
	    RECT 292.4000 43.6000 295.4000 44.4000 ;
	    RECT 293.4000 42.2000 295.4000 43.6000 ;
	    RECT 301.0000 42.2000 301.8000 49.6000 ;
	    RECT 305.8000 49.4000 307.6000 50.2000 ;
	    RECT 312.6000 49.6000 313.6000 50.2000 ;
	    RECT 314.2000 49.6000 315.6000 50.2000 ;
	    RECT 318.0000 50.2000 320.2000 50.4000 ;
	    RECT 326.2000 50.2000 326.8000 53.6000 ;
	    RECT 330.8000 57.8000 331.6000 59.8000 ;
	    RECT 330.8000 54.4000 331.4000 57.8000 ;
	    RECT 332.4000 55.6000 333.2000 57.2000 ;
	    RECT 334.0000 57.0000 334.8000 59.0000 ;
	    RECT 338.2000 58.4000 339.0000 59.0000 ;
	    RECT 337.2000 57.6000 339.0000 58.4000 ;
	    RECT 334.0000 54.8000 334.6000 57.0000 ;
	    RECT 338.2000 56.0000 339.0000 57.6000 ;
	    RECT 347.4000 56.0000 348.2000 59.0000 ;
	    RECT 351.6000 57.0000 352.4000 59.0000 ;
	    RECT 338.2000 55.4000 339.8000 56.0000 ;
	    RECT 339.0000 55.0000 339.8000 55.4000 ;
	    RECT 330.8000 53.6000 331.6000 54.4000 ;
	    RECT 334.0000 54.2000 338.2000 54.8000 ;
	    RECT 337.2000 53.8000 338.2000 54.2000 ;
	    RECT 339.2000 54.4000 339.8000 55.0000 ;
	    RECT 346.6000 55.4000 348.2000 56.0000 ;
	    RECT 346.6000 55.0000 347.4000 55.4000 ;
	    RECT 346.6000 54.4000 347.2000 55.0000 ;
	    RECT 351.8000 54.8000 352.4000 57.0000 ;
	    RECT 353.2000 55.8000 354.0000 59.8000 ;
	    RECT 354.8000 56.0000 355.6000 59.8000 ;
	    RECT 358.0000 56.0000 358.8000 59.8000 ;
	    RECT 354.8000 55.8000 358.8000 56.0000 ;
	    RECT 359.6000 56.0000 360.4000 59.8000 ;
	    RECT 362.8000 56.0000 363.6000 59.8000 ;
	    RECT 359.6000 55.8000 363.6000 56.0000 ;
	    RECT 364.4000 55.8000 365.2000 59.8000 ;
	    RECT 327.6000 52.3000 328.4000 52.4000 ;
	    RECT 329.2000 52.3000 330.0000 52.4000 ;
	    RECT 327.6000 51.7000 330.0000 52.3000 ;
	    RECT 327.6000 50.8000 328.4000 51.7000 ;
	    RECT 329.2000 50.8000 330.0000 51.7000 ;
	    RECT 330.8000 50.2000 331.4000 53.6000 ;
	    RECT 334.0000 51.6000 334.8000 53.2000 ;
	    RECT 335.6000 51.6000 336.4000 53.2000 ;
	    RECT 337.2000 53.0000 338.6000 53.8000 ;
	    RECT 339.2000 53.6000 341.2000 54.4000 ;
	    RECT 342.0000 54.3000 342.8000 54.4000 ;
	    RECT 345.2000 54.3000 347.2000 54.4000 ;
	    RECT 342.0000 53.7000 347.2000 54.3000 ;
	    RECT 348.2000 54.2000 352.4000 54.8000 ;
	    RECT 353.4000 54.4000 354.0000 55.8000 ;
	    RECT 355.0000 55.4000 358.6000 55.8000 ;
	    RECT 359.8000 55.4000 363.4000 55.8000 ;
	    RECT 357.2000 54.4000 358.0000 54.8000 ;
	    RECT 360.4000 54.4000 361.2000 54.8000 ;
	    RECT 364.4000 54.4000 365.0000 55.8000 ;
	    RECT 366.0000 55.4000 366.8000 59.8000 ;
	    RECT 370.2000 58.4000 371.4000 59.8000 ;
	    RECT 370.2000 57.8000 371.6000 58.4000 ;
	    RECT 374.8000 57.8000 375.6000 59.8000 ;
	    RECT 379.2000 58.4000 380.0000 59.8000 ;
	    RECT 379.2000 57.8000 381.2000 58.4000 ;
	    RECT 370.8000 57.0000 371.6000 57.8000 ;
	    RECT 375.0000 57.2000 375.6000 57.8000 ;
	    RECT 375.0000 56.6000 377.8000 57.2000 ;
	    RECT 377.0000 56.4000 377.8000 56.6000 ;
	    RECT 378.8000 56.4000 379.6000 57.2000 ;
	    RECT 380.4000 57.0000 381.2000 57.8000 ;
	    RECT 369.0000 55.4000 369.8000 55.6000 ;
	    RECT 366.0000 54.8000 369.8000 55.4000 ;
	    RECT 348.2000 53.8000 349.2000 54.2000 ;
	    RECT 342.0000 53.6000 342.8000 53.7000 ;
	    RECT 345.2000 53.6000 347.2000 53.7000 ;
	    RECT 337.2000 51.0000 337.8000 53.0000 ;
	    RECT 334.0000 50.4000 337.8000 51.0000 ;
	    RECT 318.0000 49.6000 321.0000 50.2000 ;
	    RECT 305.8000 42.2000 306.6000 49.4000 ;
	    RECT 312.6000 42.2000 313.4000 49.6000 ;
	    RECT 314.2000 48.4000 314.8000 49.6000 ;
	    RECT 314.0000 47.6000 314.8000 48.4000 ;
	    RECT 319.0000 42.2000 321.0000 49.6000 ;
	    RECT 326.0000 49.4000 327.8000 50.2000 ;
	    RECT 327.0000 42.2000 327.8000 49.4000 ;
	    RECT 329.8000 49.4000 331.6000 50.2000 ;
	    RECT 329.8000 44.4000 330.6000 49.4000 ;
	    RECT 329.2000 43.6000 330.6000 44.4000 ;
	    RECT 329.8000 42.2000 330.6000 43.6000 ;
	    RECT 334.0000 47.0000 334.6000 50.4000 ;
	    RECT 339.2000 49.8000 339.8000 53.6000 ;
	    RECT 340.4000 52.3000 341.2000 52.4000 ;
	    RECT 345.2000 52.3000 346.0000 52.4000 ;
	    RECT 340.4000 51.7000 346.0000 52.3000 ;
	    RECT 340.4000 50.8000 341.2000 51.7000 ;
	    RECT 345.2000 50.8000 346.0000 51.7000 ;
	    RECT 338.2000 49.2000 339.8000 49.8000 ;
	    RECT 346.6000 49.8000 347.2000 53.6000 ;
	    RECT 347.8000 53.0000 349.2000 53.8000 ;
	    RECT 353.2000 53.6000 355.8000 54.4000 ;
	    RECT 357.2000 54.3000 358.8000 54.4000 ;
	    RECT 359.6000 54.3000 361.2000 54.4000 ;
	    RECT 357.2000 53.8000 361.2000 54.3000 ;
	    RECT 358.0000 53.7000 360.4000 53.8000 ;
	    RECT 358.0000 53.6000 358.8000 53.7000 ;
	    RECT 359.6000 53.6000 360.4000 53.7000 ;
	    RECT 362.6000 53.6000 365.2000 54.4000 ;
	    RECT 348.6000 51.0000 349.2000 53.0000 ;
	    RECT 350.0000 51.6000 350.8000 53.2000 ;
	    RECT 351.6000 51.6000 352.4000 53.2000 ;
	    RECT 348.6000 50.4000 352.4000 51.0000 ;
	    RECT 346.6000 49.2000 348.2000 49.8000 ;
	    RECT 334.0000 43.0000 334.8000 47.0000 ;
	    RECT 338.2000 42.2000 339.0000 49.2000 ;
	    RECT 347.4000 42.2000 348.2000 49.2000 ;
	    RECT 351.8000 47.0000 352.4000 50.4000 ;
	    RECT 353.2000 50.2000 354.0000 50.4000 ;
	    RECT 355.2000 50.2000 355.8000 53.6000 ;
	    RECT 356.4000 52.3000 357.2000 53.2000 ;
	    RECT 361.2000 52.3000 362.0000 53.2000 ;
	    RECT 356.4000 51.7000 362.0000 52.3000 ;
	    RECT 356.4000 51.6000 357.2000 51.7000 ;
	    RECT 361.2000 51.6000 362.0000 51.7000 ;
	    RECT 362.6000 50.2000 363.2000 53.6000 ;
	    RECT 366.0000 51.4000 366.8000 54.8000 ;
	    RECT 373.0000 54.2000 373.8000 54.4000 ;
	    RECT 377.2000 54.2000 378.0000 54.4000 ;
	    RECT 378.8000 54.2000 379.4000 56.4000 ;
	    RECT 383.6000 55.0000 384.4000 59.8000 ;
	    RECT 385.2000 55.8000 386.0000 59.8000 ;
	    RECT 386.8000 56.0000 387.6000 59.8000 ;
	    RECT 390.0000 56.0000 390.8000 59.8000 ;
	    RECT 394.2000 56.4000 395.0000 59.8000 ;
	    RECT 386.8000 55.8000 390.8000 56.0000 ;
	    RECT 393.2000 55.8000 395.0000 56.4000 ;
	    RECT 396.4000 56.0000 397.2000 59.8000 ;
	    RECT 399.6000 56.0000 400.4000 59.8000 ;
	    RECT 396.4000 55.8000 400.4000 56.0000 ;
	    RECT 401.2000 55.8000 402.0000 59.8000 ;
	    RECT 385.4000 54.4000 386.0000 55.8000 ;
	    RECT 387.0000 55.4000 390.6000 55.8000 ;
	    RECT 389.2000 54.4000 390.0000 54.8000 ;
	    RECT 382.0000 54.2000 383.6000 54.4000 ;
	    RECT 372.6000 53.6000 383.6000 54.2000 ;
	    RECT 385.2000 53.6000 387.8000 54.4000 ;
	    RECT 389.2000 53.8000 390.8000 54.4000 ;
	    RECT 390.0000 53.6000 390.8000 53.8000 ;
	    RECT 391.6000 53.6000 392.4000 55.2000 ;
	    RECT 370.8000 52.8000 371.6000 53.0000 ;
	    RECT 367.8000 52.2000 371.6000 52.8000 ;
	    RECT 367.8000 52.0000 368.6000 52.2000 ;
	    RECT 369.4000 51.4000 370.2000 51.6000 ;
	    RECT 366.0000 50.8000 370.2000 51.4000 ;
	    RECT 364.4000 50.2000 365.2000 50.4000 ;
	    RECT 353.2000 49.6000 354.6000 50.2000 ;
	    RECT 355.2000 49.6000 356.2000 50.2000 ;
	    RECT 354.0000 48.4000 354.6000 49.6000 ;
	    RECT 354.0000 47.6000 354.8000 48.4000 ;
	    RECT 351.6000 43.0000 352.4000 47.0000 ;
	    RECT 355.4000 44.4000 356.2000 49.6000 ;
	    RECT 362.2000 49.6000 363.2000 50.2000 ;
	    RECT 363.8000 49.6000 365.2000 50.2000 ;
	    RECT 362.2000 48.4000 363.0000 49.6000 ;
	    RECT 363.8000 48.4000 364.4000 49.6000 ;
	    RECT 361.2000 47.6000 363.0000 48.4000 ;
	    RECT 363.6000 48.3000 364.4000 48.4000 ;
	    RECT 366.0000 48.3000 366.8000 50.8000 ;
	    RECT 372.6000 50.4000 373.2000 53.6000 ;
	    RECT 379.8000 53.4000 380.6000 53.6000 ;
	    RECT 378.8000 52.4000 379.6000 52.6000 ;
	    RECT 381.4000 52.4000 382.2000 52.6000 ;
	    RECT 377.2000 51.8000 382.2000 52.4000 ;
	    RECT 377.2000 51.6000 378.0000 51.8000 ;
	    RECT 378.8000 51.0000 384.4000 51.2000 ;
	    RECT 378.6000 50.8000 384.4000 51.0000 ;
	    RECT 370.8000 49.8000 373.2000 50.4000 ;
	    RECT 374.6000 50.6000 384.4000 50.8000 ;
	    RECT 374.6000 50.2000 379.4000 50.6000 ;
	    RECT 370.8000 48.8000 371.4000 49.8000 ;
	    RECT 363.6000 47.7000 366.8000 48.3000 ;
	    RECT 370.0000 48.0000 371.4000 48.8000 ;
	    RECT 373.0000 49.0000 373.8000 49.2000 ;
	    RECT 374.6000 49.0000 375.2000 50.2000 ;
	    RECT 373.0000 48.4000 375.2000 49.0000 ;
	    RECT 375.8000 49.0000 381.2000 49.6000 ;
	    RECT 375.8000 48.8000 376.6000 49.0000 ;
	    RECT 380.4000 48.8000 381.2000 49.0000 ;
	    RECT 363.6000 47.6000 364.4000 47.7000 ;
	    RECT 355.4000 43.6000 357.2000 44.4000 ;
	    RECT 355.4000 42.2000 356.2000 43.6000 ;
	    RECT 362.2000 42.2000 363.0000 47.6000 ;
	    RECT 366.0000 42.2000 366.8000 47.7000 ;
	    RECT 374.2000 47.4000 375.0000 47.6000 ;
	    RECT 377.0000 47.4000 377.8000 47.6000 ;
	    RECT 370.8000 46.2000 371.6000 47.0000 ;
	    RECT 374.2000 46.8000 377.8000 47.4000 ;
	    RECT 375.0000 46.2000 375.6000 46.8000 ;
	    RECT 380.4000 46.2000 381.2000 47.0000 ;
	    RECT 370.2000 42.2000 371.4000 46.2000 ;
	    RECT 374.8000 42.2000 375.6000 46.2000 ;
	    RECT 379.2000 45.6000 381.2000 46.2000 ;
	    RECT 379.2000 42.2000 380.0000 45.6000 ;
	    RECT 383.6000 42.2000 384.4000 50.6000 ;
	    RECT 385.2000 50.2000 386.0000 50.4000 ;
	    RECT 387.2000 50.2000 387.8000 53.6000 ;
	    RECT 388.4000 51.6000 389.2000 53.2000 ;
	    RECT 385.2000 49.6000 386.6000 50.2000 ;
	    RECT 387.2000 49.6000 388.2000 50.2000 ;
	    RECT 386.0000 48.4000 386.6000 49.6000 ;
	    RECT 386.0000 47.6000 386.8000 48.4000 ;
	    RECT 387.4000 42.2000 388.2000 49.6000 ;
	    RECT 393.2000 42.2000 394.0000 55.8000 ;
	    RECT 396.6000 55.4000 400.2000 55.8000 ;
	    RECT 397.2000 54.4000 398.0000 54.8000 ;
	    RECT 401.2000 54.4000 401.8000 55.8000 ;
	    RECT 409.2000 55.4000 410.0000 59.8000 ;
	    RECT 413.4000 58.4000 414.6000 59.8000 ;
	    RECT 413.4000 57.8000 414.8000 58.4000 ;
	    RECT 418.0000 57.8000 418.8000 59.8000 ;
	    RECT 422.4000 58.4000 423.2000 59.8000 ;
	    RECT 422.4000 57.8000 424.4000 58.4000 ;
	    RECT 414.0000 57.0000 414.8000 57.8000 ;
	    RECT 418.2000 57.2000 418.8000 57.8000 ;
	    RECT 418.2000 56.6000 421.0000 57.2000 ;
	    RECT 420.2000 56.4000 421.0000 56.6000 ;
	    RECT 422.0000 56.4000 422.8000 57.2000 ;
	    RECT 423.6000 57.0000 424.4000 57.8000 ;
	    RECT 412.2000 55.4000 413.0000 55.6000 ;
	    RECT 409.2000 54.8000 413.0000 55.4000 ;
	    RECT 396.4000 53.8000 398.0000 54.4000 ;
	    RECT 396.4000 53.6000 397.2000 53.8000 ;
	    RECT 399.4000 53.6000 402.0000 54.4000 ;
	    RECT 394.8000 52.3000 395.6000 52.4000 ;
	    RECT 398.0000 52.3000 398.8000 53.2000 ;
	    RECT 394.8000 51.7000 398.8000 52.3000 ;
	    RECT 394.8000 51.6000 395.6000 51.7000 ;
	    RECT 398.0000 51.6000 398.8000 51.7000 ;
	    RECT 394.8000 48.8000 395.6000 50.4000 ;
	    RECT 399.4000 50.2000 400.0000 53.6000 ;
	    RECT 409.2000 51.4000 410.0000 54.8000 ;
	    RECT 416.2000 54.2000 417.0000 54.4000 ;
	    RECT 422.0000 54.2000 422.6000 56.4000 ;
	    RECT 426.8000 55.0000 427.6000 59.8000 ;
	    RECT 431.0000 56.4000 431.8000 59.8000 ;
	    RECT 430.0000 55.8000 431.8000 56.4000 ;
	    RECT 425.2000 54.2000 426.8000 54.4000 ;
	    RECT 415.8000 53.6000 426.8000 54.2000 ;
	    RECT 428.4000 53.6000 429.2000 55.2000 ;
	    RECT 414.0000 52.8000 414.8000 53.0000 ;
	    RECT 411.0000 52.2000 414.8000 52.8000 ;
	    RECT 411.0000 52.0000 411.8000 52.2000 ;
	    RECT 412.6000 51.4000 413.4000 51.6000 ;
	    RECT 409.2000 50.8000 413.4000 51.4000 ;
	    RECT 401.2000 50.2000 402.0000 50.4000 ;
	    RECT 399.0000 49.6000 400.0000 50.2000 ;
	    RECT 400.6000 49.6000 402.0000 50.2000 ;
	    RECT 399.0000 44.4000 399.8000 49.6000 ;
	    RECT 400.6000 48.4000 401.2000 49.6000 ;
	    RECT 400.4000 47.6000 401.2000 48.4000 ;
	    RECT 398.0000 43.6000 399.8000 44.4000 ;
	    RECT 399.0000 42.2000 399.8000 43.6000 ;
	    RECT 409.2000 42.2000 410.0000 50.8000 ;
	    RECT 415.8000 50.4000 416.4000 53.6000 ;
	    RECT 423.0000 53.4000 423.8000 53.6000 ;
	    RECT 422.0000 52.4000 422.8000 52.6000 ;
	    RECT 424.6000 52.4000 425.4000 52.6000 ;
	    RECT 420.4000 51.8000 425.4000 52.4000 ;
	    RECT 430.0000 52.3000 430.8000 55.8000 ;
	    RECT 433.2000 55.6000 434.0000 59.8000 ;
	    RECT 434.8000 56.0000 435.6000 59.8000 ;
	    RECT 438.0000 56.0000 438.8000 59.8000 ;
	    RECT 434.8000 55.8000 438.8000 56.0000 ;
	    RECT 433.4000 54.4000 434.0000 55.6000 ;
	    RECT 435.0000 55.4000 438.6000 55.8000 ;
	    RECT 439.6000 55.2000 440.4000 59.8000 ;
	    RECT 437.2000 54.4000 438.0000 54.8000 ;
	    RECT 439.6000 54.6000 441.8000 55.2000 ;
	    RECT 433.2000 53.6000 435.8000 54.4000 ;
	    RECT 437.2000 53.8000 438.8000 54.4000 ;
	    RECT 438.0000 53.6000 438.8000 53.8000 ;
	    RECT 420.4000 51.6000 421.2000 51.8000 ;
	    RECT 430.0000 51.7000 433.9000 52.3000 ;
	    RECT 422.0000 51.0000 427.6000 51.2000 ;
	    RECT 421.8000 50.8000 427.6000 51.0000 ;
	    RECT 414.0000 49.8000 416.4000 50.4000 ;
	    RECT 417.8000 50.6000 427.6000 50.8000 ;
	    RECT 417.8000 50.2000 422.6000 50.6000 ;
	    RECT 414.0000 48.8000 414.6000 49.8000 ;
	    RECT 413.2000 48.0000 414.6000 48.8000 ;
	    RECT 416.2000 49.0000 417.0000 49.2000 ;
	    RECT 417.8000 49.0000 418.4000 50.2000 ;
	    RECT 416.2000 48.4000 418.4000 49.0000 ;
	    RECT 419.0000 49.0000 424.4000 49.6000 ;
	    RECT 419.0000 48.8000 419.8000 49.0000 ;
	    RECT 423.6000 48.8000 424.4000 49.0000 ;
	    RECT 417.4000 47.4000 418.2000 47.6000 ;
	    RECT 420.2000 47.4000 421.0000 47.6000 ;
	    RECT 414.0000 46.2000 414.8000 47.0000 ;
	    RECT 417.4000 46.8000 421.0000 47.4000 ;
	    RECT 418.2000 46.2000 418.8000 46.8000 ;
	    RECT 423.6000 46.2000 424.4000 47.0000 ;
	    RECT 413.4000 42.2000 414.6000 46.2000 ;
	    RECT 418.0000 42.2000 418.8000 46.2000 ;
	    RECT 422.4000 45.6000 424.4000 46.2000 ;
	    RECT 422.4000 42.2000 423.2000 45.6000 ;
	    RECT 426.8000 42.2000 427.6000 50.6000 ;
	    RECT 430.0000 42.2000 430.8000 51.7000 ;
	    RECT 433.3000 50.4000 433.9000 51.7000 ;
	    RECT 431.6000 48.8000 432.4000 50.4000 ;
	    RECT 433.2000 50.2000 434.0000 50.4000 ;
	    RECT 435.2000 50.2000 435.8000 53.6000 ;
	    RECT 436.4000 51.6000 437.2000 53.2000 ;
	    RECT 439.6000 51.6000 440.4000 53.2000 ;
	    RECT 441.2000 51.6000 441.8000 54.6000 ;
	    RECT 442.8000 52.4000 443.6000 59.8000 ;
	    RECT 441.2000 50.8000 442.4000 51.6000 ;
	    RECT 441.2000 50.2000 441.8000 50.8000 ;
	    RECT 443.0000 50.2000 443.6000 52.4000 ;
	    RECT 433.2000 49.6000 434.6000 50.2000 ;
	    RECT 435.2000 49.6000 436.2000 50.2000 ;
	    RECT 434.0000 48.4000 434.6000 49.6000 ;
	    RECT 434.0000 47.6000 434.8000 48.4000 ;
	    RECT 435.4000 42.2000 436.2000 49.6000 ;
	    RECT 439.6000 49.6000 441.8000 50.2000 ;
	    RECT 439.6000 42.2000 440.4000 49.6000 ;
	    RECT 442.8000 42.2000 443.6000 50.2000 ;
	    RECT 444.4000 55.4000 445.2000 59.8000 ;
	    RECT 448.6000 58.4000 449.8000 59.8000 ;
	    RECT 448.6000 57.8000 450.0000 58.4000 ;
	    RECT 453.2000 57.8000 454.0000 59.8000 ;
	    RECT 457.6000 58.4000 458.4000 59.8000 ;
	    RECT 457.6000 57.8000 459.6000 58.4000 ;
	    RECT 449.2000 57.0000 450.0000 57.8000 ;
	    RECT 453.4000 57.2000 454.0000 57.8000 ;
	    RECT 453.4000 56.6000 456.2000 57.2000 ;
	    RECT 455.4000 56.4000 456.2000 56.6000 ;
	    RECT 457.2000 56.4000 458.0000 57.2000 ;
	    RECT 458.8000 57.0000 459.6000 57.8000 ;
	    RECT 447.4000 55.4000 448.2000 55.6000 ;
	    RECT 444.4000 54.8000 448.2000 55.4000 ;
	    RECT 444.4000 51.4000 445.2000 54.8000 ;
	    RECT 451.4000 54.2000 452.2000 54.4000 ;
	    RECT 457.2000 54.2000 457.8000 56.4000 ;
	    RECT 462.0000 55.0000 462.8000 59.8000 ;
	    RECT 460.4000 54.2000 462.0000 54.4000 ;
	    RECT 451.0000 53.6000 462.0000 54.2000 ;
	    RECT 449.2000 52.8000 450.0000 53.0000 ;
	    RECT 446.2000 52.2000 450.0000 52.8000 ;
	    RECT 451.0000 52.4000 451.6000 53.6000 ;
	    RECT 458.2000 53.4000 459.0000 53.6000 ;
	    RECT 459.8000 52.4000 460.6000 52.6000 ;
	    RECT 446.2000 52.0000 447.0000 52.2000 ;
	    RECT 450.8000 51.6000 451.6000 52.4000 ;
	    RECT 454.0000 52.3000 454.8000 52.4000 ;
	    RECT 455.6000 52.3000 460.6000 52.4000 ;
	    RECT 454.0000 51.8000 460.6000 52.3000 ;
	    RECT 454.0000 51.7000 456.4000 51.8000 ;
	    RECT 454.0000 51.6000 454.8000 51.7000 ;
	    RECT 455.6000 51.6000 456.4000 51.7000 ;
	    RECT 447.8000 51.4000 448.6000 51.6000 ;
	    RECT 444.4000 50.8000 448.6000 51.4000 ;
	    RECT 444.4000 42.2000 445.2000 50.8000 ;
	    RECT 451.0000 50.4000 451.6000 51.6000 ;
	    RECT 457.2000 51.0000 462.8000 51.2000 ;
	    RECT 457.0000 50.8000 462.8000 51.0000 ;
	    RECT 449.2000 49.8000 451.6000 50.4000 ;
	    RECT 453.0000 50.6000 462.8000 50.8000 ;
	    RECT 453.0000 50.2000 457.8000 50.6000 ;
	    RECT 449.2000 48.8000 449.8000 49.8000 ;
	    RECT 448.4000 48.0000 449.8000 48.8000 ;
	    RECT 451.4000 49.0000 452.2000 49.2000 ;
	    RECT 453.0000 49.0000 453.6000 50.2000 ;
	    RECT 451.4000 48.4000 453.6000 49.0000 ;
	    RECT 454.2000 49.0000 459.6000 49.6000 ;
	    RECT 454.2000 48.8000 455.0000 49.0000 ;
	    RECT 458.8000 48.8000 459.6000 49.0000 ;
	    RECT 452.6000 47.4000 453.4000 47.6000 ;
	    RECT 455.4000 47.4000 456.2000 47.6000 ;
	    RECT 449.2000 46.2000 450.0000 47.0000 ;
	    RECT 452.6000 46.8000 456.2000 47.4000 ;
	    RECT 453.4000 46.2000 454.0000 46.8000 ;
	    RECT 458.8000 46.2000 459.6000 47.0000 ;
	    RECT 448.6000 42.2000 449.8000 46.2000 ;
	    RECT 453.2000 42.2000 454.0000 46.2000 ;
	    RECT 457.6000 45.6000 459.6000 46.2000 ;
	    RECT 457.6000 42.2000 458.4000 45.6000 ;
	    RECT 462.0000 42.2000 462.8000 50.6000 ;
	    RECT 463.6000 42.2000 464.4000 59.8000 ;
	    RECT 468.0000 54.2000 468.8000 59.8000 ;
	    RECT 467.0000 53.8000 468.8000 54.2000 ;
	    RECT 467.0000 53.6000 468.6000 53.8000 ;
	    RECT 467.0000 50.4000 467.6000 53.6000 ;
	    RECT 469.2000 51.6000 470.8000 52.4000 ;
	    RECT 466.8000 49.6000 467.6000 50.4000 ;
	    RECT 467.0000 47.0000 467.6000 49.6000 ;
	    RECT 468.4000 47.6000 469.2000 49.2000 ;
	    RECT 467.0000 46.4000 470.6000 47.0000 ;
	    RECT 467.0000 46.2000 467.6000 46.4000 ;
	    RECT 466.8000 42.2000 467.6000 46.2000 ;
	    RECT 470.0000 46.2000 470.6000 46.4000 ;
	    RECT 470.0000 42.2000 470.8000 46.2000 ;
	    RECT 473.2000 42.2000 474.0000 59.8000 ;
	    RECT 480.0000 54.2000 480.8000 59.8000 ;
	    RECT 480.0000 53.8000 481.8000 54.2000 ;
	    RECT 480.2000 53.6000 481.8000 53.8000 ;
	    RECT 478.0000 51.6000 479.6000 52.4000 ;
	    RECT 481.2000 50.4000 481.8000 53.6000 ;
	    RECT 481.2000 49.6000 482.0000 50.4000 ;
	    RECT 479.6000 47.6000 480.4000 49.2000 ;
	    RECT 481.2000 47.0000 481.8000 49.6000 ;
	    RECT 478.2000 46.4000 481.8000 47.0000 ;
	    RECT 478.2000 46.2000 478.8000 46.4000 ;
	    RECT 478.0000 42.2000 478.8000 46.2000 ;
	    RECT 481.2000 46.2000 481.8000 46.4000 ;
	    RECT 481.2000 42.2000 482.0000 46.2000 ;
	    RECT 482.8000 42.2000 483.6000 59.8000 ;
	    RECT 487.2000 54.2000 488.0000 59.8000 ;
	    RECT 486.2000 53.8000 488.0000 54.2000 ;
	    RECT 492.4000 55.4000 493.2000 59.8000 ;
	    RECT 496.6000 58.4000 497.8000 59.8000 ;
	    RECT 496.6000 57.8000 498.0000 58.4000 ;
	    RECT 501.2000 57.8000 502.0000 59.8000 ;
	    RECT 505.6000 58.4000 506.4000 59.8000 ;
	    RECT 505.6000 57.8000 507.6000 58.4000 ;
	    RECT 497.2000 57.0000 498.0000 57.8000 ;
	    RECT 501.4000 57.2000 502.0000 57.8000 ;
	    RECT 501.4000 56.6000 504.2000 57.2000 ;
	    RECT 503.4000 56.4000 504.2000 56.6000 ;
	    RECT 505.2000 56.4000 506.0000 57.2000 ;
	    RECT 506.8000 57.0000 507.6000 57.8000 ;
	    RECT 495.4000 55.4000 496.2000 55.6000 ;
	    RECT 492.4000 54.8000 496.2000 55.4000 ;
	    RECT 486.2000 53.6000 487.8000 53.8000 ;
	    RECT 486.2000 50.4000 486.8000 53.6000 ;
	    RECT 488.4000 51.6000 490.0000 52.4000 ;
	    RECT 486.0000 49.6000 486.8000 50.4000 ;
	    RECT 486.2000 47.0000 486.8000 49.6000 ;
	    RECT 492.4000 51.4000 493.2000 54.8000 ;
	    RECT 499.4000 54.2000 500.2000 54.4000 ;
	    RECT 502.0000 54.2000 502.8000 54.4000 ;
	    RECT 505.2000 54.2000 505.8000 56.4000 ;
	    RECT 510.0000 55.0000 510.8000 59.8000 ;
	    RECT 508.4000 54.2000 510.0000 54.4000 ;
	    RECT 499.0000 53.6000 510.0000 54.2000 ;
	    RECT 497.2000 52.8000 498.0000 53.0000 ;
	    RECT 494.2000 52.2000 498.0000 52.8000 ;
	    RECT 494.2000 52.0000 495.0000 52.2000 ;
	    RECT 495.8000 51.4000 496.6000 51.6000 ;
	    RECT 492.4000 50.8000 496.6000 51.4000 ;
	    RECT 487.6000 47.6000 488.4000 49.2000 ;
	    RECT 486.2000 46.4000 489.8000 47.0000 ;
	    RECT 486.2000 46.2000 486.8000 46.4000 ;
	    RECT 486.0000 42.2000 486.8000 46.2000 ;
	    RECT 489.2000 46.2000 489.8000 46.4000 ;
	    RECT 489.2000 42.2000 490.0000 46.2000 ;
	    RECT 492.4000 42.2000 493.2000 50.8000 ;
	    RECT 499.0000 50.4000 499.6000 53.6000 ;
	    RECT 506.2000 53.4000 507.0000 53.6000 ;
	    RECT 507.8000 52.4000 508.6000 52.6000 ;
	    RECT 500.4000 52.3000 501.2000 52.4000 ;
	    RECT 503.6000 52.3000 508.6000 52.4000 ;
	    RECT 500.4000 51.8000 508.6000 52.3000 ;
	    RECT 500.4000 51.7000 504.4000 51.8000 ;
	    RECT 500.4000 51.6000 501.2000 51.7000 ;
	    RECT 503.6000 51.6000 504.4000 51.7000 ;
	    RECT 505.2000 51.0000 510.8000 51.2000 ;
	    RECT 505.0000 50.8000 510.8000 51.0000 ;
	    RECT 497.2000 49.8000 499.6000 50.4000 ;
	    RECT 501.0000 50.6000 510.8000 50.8000 ;
	    RECT 501.0000 50.2000 505.8000 50.6000 ;
	    RECT 497.2000 48.8000 497.8000 49.8000 ;
	    RECT 496.4000 48.0000 497.8000 48.8000 ;
	    RECT 499.4000 49.0000 500.2000 49.2000 ;
	    RECT 501.0000 49.0000 501.6000 50.2000 ;
	    RECT 499.4000 48.4000 501.6000 49.0000 ;
	    RECT 502.2000 49.0000 507.6000 49.6000 ;
	    RECT 502.2000 48.8000 503.0000 49.0000 ;
	    RECT 506.8000 48.8000 507.6000 49.0000 ;
	    RECT 500.6000 47.4000 501.4000 47.6000 ;
	    RECT 503.4000 47.4000 504.2000 47.6000 ;
	    RECT 497.2000 46.2000 498.0000 47.0000 ;
	    RECT 500.6000 46.8000 504.2000 47.4000 ;
	    RECT 501.4000 46.2000 502.0000 46.8000 ;
	    RECT 506.8000 46.2000 507.6000 47.0000 ;
	    RECT 496.6000 42.2000 497.8000 46.2000 ;
	    RECT 501.2000 42.2000 502.0000 46.2000 ;
	    RECT 505.6000 45.6000 507.6000 46.2000 ;
	    RECT 505.6000 42.2000 506.4000 45.6000 ;
	    RECT 510.0000 42.2000 510.8000 50.6000 ;
	    RECT 1.2000 31.2000 2.0000 39.8000 ;
	    RECT 5.4000 35.8000 6.6000 39.8000 ;
	    RECT 10.0000 35.8000 10.8000 39.8000 ;
	    RECT 14.4000 36.4000 15.2000 39.8000 ;
	    RECT 14.4000 35.8000 16.4000 36.4000 ;
	    RECT 6.0000 35.0000 6.8000 35.8000 ;
	    RECT 10.2000 35.2000 10.8000 35.8000 ;
	    RECT 9.4000 34.6000 13.0000 35.2000 ;
	    RECT 15.6000 35.0000 16.4000 35.8000 ;
	    RECT 9.4000 34.4000 10.2000 34.6000 ;
	    RECT 12.2000 34.4000 13.0000 34.6000 ;
	    RECT 5.2000 33.2000 6.6000 34.0000 ;
	    RECT 6.0000 32.2000 6.6000 33.2000 ;
	    RECT 8.2000 33.0000 10.4000 33.6000 ;
	    RECT 8.2000 32.8000 9.0000 33.0000 ;
	    RECT 6.0000 31.6000 8.4000 32.2000 ;
	    RECT 1.2000 30.6000 5.4000 31.2000 ;
	    RECT 1.2000 27.2000 2.0000 30.6000 ;
	    RECT 4.6000 30.4000 5.4000 30.6000 ;
	    RECT 3.0000 29.8000 3.8000 30.0000 ;
	    RECT 3.0000 29.2000 6.8000 29.8000 ;
	    RECT 6.0000 29.0000 6.8000 29.2000 ;
	    RECT 7.8000 28.4000 8.4000 31.6000 ;
	    RECT 9.8000 31.8000 10.4000 33.0000 ;
	    RECT 11.0000 33.0000 11.8000 33.2000 ;
	    RECT 15.6000 33.0000 16.4000 33.2000 ;
	    RECT 11.0000 32.4000 16.4000 33.0000 ;
	    RECT 9.8000 31.4000 14.6000 31.8000 ;
	    RECT 18.8000 31.4000 19.6000 39.8000 ;
	    RECT 9.8000 31.2000 19.6000 31.4000 ;
	    RECT 13.8000 31.0000 19.6000 31.2000 ;
	    RECT 14.0000 30.8000 19.6000 31.0000 ;
	    RECT 20.4000 31.4000 21.2000 39.8000 ;
	    RECT 24.8000 36.4000 25.6000 39.8000 ;
	    RECT 23.6000 35.8000 25.6000 36.4000 ;
	    RECT 29.2000 35.8000 30.0000 39.8000 ;
	    RECT 33.4000 35.8000 34.6000 39.8000 ;
	    RECT 23.6000 35.0000 24.4000 35.8000 ;
	    RECT 29.2000 35.2000 29.8000 35.8000 ;
	    RECT 27.0000 34.6000 30.6000 35.2000 ;
	    RECT 33.2000 35.0000 34.0000 35.8000 ;
	    RECT 27.0000 34.4000 27.8000 34.6000 ;
	    RECT 29.8000 34.4000 30.6000 34.6000 ;
	    RECT 38.0000 34.3000 38.8000 39.8000 ;
	    RECT 41.8000 38.4000 42.6000 39.8000 ;
	    RECT 41.8000 37.6000 43.6000 38.4000 ;
	    RECT 40.4000 34.3000 41.2000 34.4000 ;
	    RECT 23.6000 33.0000 24.4000 33.2000 ;
	    RECT 28.2000 33.0000 29.0000 33.2000 ;
	    RECT 23.6000 32.4000 29.0000 33.0000 ;
	    RECT 29.6000 33.0000 31.8000 33.6000 ;
	    RECT 29.6000 31.8000 30.2000 33.0000 ;
	    RECT 31.0000 32.8000 31.8000 33.0000 ;
	    RECT 33.4000 33.2000 34.8000 34.0000 ;
	    RECT 38.0000 33.7000 41.2000 34.3000 ;
	    RECT 33.4000 32.2000 34.0000 33.2000 ;
	    RECT 25.4000 31.4000 30.2000 31.8000 ;
	    RECT 20.4000 31.2000 30.2000 31.4000 ;
	    RECT 31.6000 31.6000 34.0000 32.2000 ;
	    RECT 20.4000 31.0000 26.2000 31.2000 ;
	    RECT 20.4000 30.8000 26.0000 31.0000 ;
	    RECT 12.4000 30.2000 13.2000 30.4000 ;
	    RECT 26.8000 30.3000 27.6000 30.4000 ;
	    RECT 28.4000 30.3000 29.2000 30.4000 ;
	    RECT 26.8000 30.2000 29.2000 30.3000 ;
	    RECT 12.4000 29.6000 17.4000 30.2000 ;
	    RECT 14.0000 29.4000 14.8000 29.6000 ;
	    RECT 16.6000 29.4000 17.4000 29.6000 ;
	    RECT 22.6000 29.7000 29.2000 30.2000 ;
	    RECT 22.6000 29.6000 27.6000 29.7000 ;
	    RECT 28.4000 29.6000 29.2000 29.7000 ;
	    RECT 22.6000 29.4000 23.4000 29.6000 ;
	    RECT 15.0000 28.4000 15.8000 28.6000 ;
	    RECT 24.2000 28.4000 25.0000 28.6000 ;
	    RECT 31.6000 28.4000 32.2000 31.6000 ;
	    RECT 38.0000 31.2000 38.8000 33.7000 ;
	    RECT 40.4000 33.6000 41.2000 33.7000 ;
	    RECT 40.4000 32.4000 41.0000 33.6000 ;
	    RECT 41.8000 32.4000 42.6000 37.6000 ;
	    RECT 46.0000 33.6000 47.6000 34.4000 ;
	    RECT 46.8000 32.4000 47.4000 33.6000 ;
	    RECT 48.2000 32.4000 49.0000 39.8000 ;
	    RECT 39.6000 31.8000 41.0000 32.4000 ;
	    RECT 41.6000 31.8000 42.6000 32.4000 ;
	    RECT 46.0000 31.8000 47.4000 32.4000 ;
	    RECT 48.0000 31.8000 49.0000 32.4000 ;
	    RECT 55.0000 32.4000 55.8000 39.8000 ;
	    RECT 56.4000 33.6000 57.2000 34.4000 ;
	    RECT 56.6000 32.4000 57.2000 33.6000 ;
	    RECT 59.6000 33.6000 60.4000 34.4000 ;
	    RECT 59.6000 32.4000 60.2000 33.6000 ;
	    RECT 61.0000 32.4000 61.8000 39.8000 ;
	    RECT 55.0000 31.8000 56.0000 32.4000 ;
	    RECT 56.6000 31.8000 58.0000 32.4000 ;
	    RECT 39.6000 31.6000 40.4000 31.8000 ;
	    RECT 34.6000 30.6000 38.8000 31.2000 ;
	    RECT 34.6000 30.4000 35.4000 30.6000 ;
	    RECT 36.2000 29.8000 37.0000 30.0000 ;
	    RECT 33.2000 29.2000 37.0000 29.8000 ;
	    RECT 33.2000 29.0000 34.0000 29.2000 ;
	    RECT 7.8000 27.8000 18.8000 28.4000 ;
	    RECT 8.2000 27.6000 9.0000 27.8000 ;
	    RECT 1.2000 26.6000 5.2000 27.2000 ;
	    RECT 1.2000 22.2000 2.0000 26.6000 ;
	    RECT 4.2000 26.4000 5.2000 26.6000 ;
	    RECT 4.4000 25.6000 5.2000 26.4000 ;
	    RECT 14.0000 25.6000 14.6000 27.8000 ;
	    RECT 17.2000 27.6000 18.8000 27.8000 ;
	    RECT 21.2000 27.8000 32.2000 28.4000 ;
	    RECT 21.2000 27.6000 22.8000 27.8000 ;
	    RECT 12.2000 25.4000 13.0000 25.6000 ;
	    RECT 6.0000 24.2000 6.8000 25.0000 ;
	    RECT 10.2000 24.8000 13.0000 25.4000 ;
	    RECT 14.0000 24.8000 14.8000 25.6000 ;
	    RECT 10.2000 24.2000 10.8000 24.8000 ;
	    RECT 15.6000 24.2000 16.4000 25.0000 ;
	    RECT 5.4000 23.6000 6.8000 24.2000 ;
	    RECT 5.4000 22.2000 6.6000 23.6000 ;
	    RECT 10.0000 22.2000 10.8000 24.2000 ;
	    RECT 14.4000 23.6000 16.4000 24.2000 ;
	    RECT 14.4000 22.2000 15.2000 23.6000 ;
	    RECT 18.8000 22.2000 19.6000 27.0000 ;
	    RECT 20.4000 22.2000 21.2000 27.0000 ;
	    RECT 25.4000 25.6000 26.0000 27.8000 ;
	    RECT 26.8000 27.6000 27.6000 27.8000 ;
	    RECT 31.0000 27.6000 31.8000 27.8000 ;
	    RECT 38.0000 27.2000 38.8000 30.6000 ;
	    RECT 41.6000 28.4000 42.2000 31.8000 ;
	    RECT 46.0000 31.6000 46.8000 31.8000 ;
	    RECT 48.0000 30.4000 48.6000 31.8000 ;
	    RECT 42.8000 28.8000 43.6000 30.4000 ;
	    RECT 47.6000 29.6000 48.6000 30.4000 ;
	    RECT 48.0000 28.4000 48.6000 29.6000 ;
	    RECT 49.2000 28.8000 50.0000 30.4000 ;
	    RECT 54.0000 28.8000 54.8000 30.4000 ;
	    RECT 55.4000 30.3000 56.0000 31.8000 ;
	    RECT 57.2000 31.6000 58.0000 31.8000 ;
	    RECT 58.8000 31.8000 60.2000 32.4000 ;
	    RECT 60.8000 31.8000 61.8000 32.4000 ;
	    RECT 65.2000 32.4000 66.0000 39.8000 ;
	    RECT 65.2000 31.8000 67.4000 32.4000 ;
	    RECT 58.8000 31.6000 59.6000 31.8000 ;
	    RECT 58.9000 30.3000 59.5000 31.6000 ;
	    RECT 55.4000 29.7000 59.5000 30.3000 ;
	    RECT 55.4000 28.4000 56.0000 29.7000 ;
	    RECT 60.8000 28.4000 61.4000 31.8000 ;
	    RECT 66.8000 31.2000 67.4000 31.8000 ;
	    RECT 70.0000 31.2000 70.8000 39.8000 ;
	    RECT 74.2000 35.8000 75.4000 39.8000 ;
	    RECT 78.8000 35.8000 79.6000 39.8000 ;
	    RECT 83.2000 36.4000 84.0000 39.8000 ;
	    RECT 83.2000 35.8000 85.2000 36.4000 ;
	    RECT 74.8000 35.0000 75.6000 35.8000 ;
	    RECT 79.0000 35.2000 79.6000 35.8000 ;
	    RECT 78.2000 34.6000 81.8000 35.2000 ;
	    RECT 84.4000 35.0000 85.2000 35.8000 ;
	    RECT 78.2000 34.4000 79.0000 34.6000 ;
	    RECT 81.0000 34.4000 81.8000 34.6000 ;
	    RECT 74.0000 33.2000 75.4000 34.0000 ;
	    RECT 74.8000 32.2000 75.4000 33.2000 ;
	    RECT 77.0000 33.0000 79.2000 33.6000 ;
	    RECT 77.0000 32.8000 77.8000 33.0000 ;
	    RECT 74.8000 31.6000 77.2000 32.2000 ;
	    RECT 66.8000 30.4000 68.0000 31.2000 ;
	    RECT 70.0000 30.6000 74.2000 31.2000 ;
	    RECT 62.0000 28.8000 62.8000 30.4000 ;
	    RECT 65.2000 28.8000 66.0000 30.4000 ;
	    RECT 39.6000 27.6000 42.2000 28.4000 ;
	    RECT 44.4000 28.2000 45.2000 28.4000 ;
	    RECT 43.6000 27.6000 45.2000 28.2000 ;
	    RECT 46.0000 27.6000 48.6000 28.4000 ;
	    RECT 50.8000 28.3000 51.6000 28.4000 ;
	    RECT 52.4000 28.3000 53.2000 28.4000 ;
	    RECT 50.8000 28.2000 53.2000 28.3000 ;
	    RECT 50.0000 27.7000 54.0000 28.2000 ;
	    RECT 50.0000 27.6000 51.6000 27.7000 ;
	    RECT 52.4000 27.6000 54.0000 27.7000 ;
	    RECT 55.4000 27.6000 58.0000 28.4000 ;
	    RECT 58.8000 27.6000 61.4000 28.4000 ;
	    RECT 63.6000 28.2000 64.4000 28.4000 ;
	    RECT 62.8000 27.6000 64.4000 28.2000 ;
	    RECT 35.0000 26.6000 38.8000 27.2000 ;
	    RECT 35.0000 26.4000 35.8000 26.6000 ;
	    RECT 23.6000 24.2000 24.4000 25.0000 ;
	    RECT 25.2000 24.8000 26.0000 25.6000 ;
	    RECT 27.0000 25.4000 27.8000 25.6000 ;
	    RECT 27.0000 24.8000 29.8000 25.4000 ;
	    RECT 29.2000 24.2000 29.8000 24.8000 ;
	    RECT 33.2000 24.2000 34.0000 25.0000 ;
	    RECT 23.6000 23.6000 25.6000 24.2000 ;
	    RECT 24.8000 22.2000 25.6000 23.6000 ;
	    RECT 29.2000 22.2000 30.0000 24.2000 ;
	    RECT 33.2000 23.6000 34.6000 24.2000 ;
	    RECT 33.4000 22.2000 34.6000 23.6000 ;
	    RECT 38.0000 22.2000 38.8000 26.6000 ;
	    RECT 39.8000 26.2000 40.4000 27.6000 ;
	    RECT 43.6000 27.2000 44.4000 27.6000 ;
	    RECT 41.4000 26.2000 45.0000 26.6000 ;
	    RECT 46.2000 26.2000 46.8000 27.6000 ;
	    RECT 50.0000 27.2000 50.8000 27.6000 ;
	    RECT 53.2000 27.2000 54.0000 27.6000 ;
	    RECT 47.8000 26.2000 51.4000 26.6000 ;
	    RECT 52.6000 26.2000 56.2000 26.6000 ;
	    RECT 57.2000 26.2000 57.8000 27.6000 ;
	    RECT 59.0000 26.2000 59.6000 27.6000 ;
	    RECT 62.8000 27.2000 63.6000 27.6000 ;
	    RECT 66.8000 27.4000 67.4000 30.4000 ;
	    RECT 65.2000 26.8000 67.4000 27.4000 ;
	    RECT 70.0000 27.2000 70.8000 30.6000 ;
	    RECT 73.4000 30.4000 74.2000 30.6000 ;
	    RECT 71.8000 29.8000 72.6000 30.0000 ;
	    RECT 71.8000 29.2000 75.6000 29.8000 ;
	    RECT 74.8000 29.0000 75.6000 29.2000 ;
	    RECT 76.6000 28.4000 77.2000 31.6000 ;
	    RECT 78.6000 31.8000 79.2000 33.0000 ;
	    RECT 79.8000 33.0000 80.6000 33.2000 ;
	    RECT 84.4000 33.0000 85.2000 33.2000 ;
	    RECT 79.8000 32.4000 85.2000 33.0000 ;
	    RECT 78.6000 31.4000 83.4000 31.8000 ;
	    RECT 87.6000 31.4000 88.4000 39.8000 ;
	    RECT 91.4000 38.4000 92.2000 39.8000 ;
	    RECT 91.4000 37.6000 93.2000 38.4000 ;
	    RECT 90.0000 33.6000 90.8000 34.4000 ;
	    RECT 90.0000 32.4000 90.6000 33.6000 ;
	    RECT 91.4000 32.4000 92.2000 37.6000 ;
	    RECT 97.8000 34.4000 98.6000 39.8000 ;
	    RECT 96.4000 33.6000 97.2000 34.4000 ;
	    RECT 97.8000 33.6000 99.6000 34.4000 ;
	    RECT 96.4000 32.4000 97.0000 33.6000 ;
	    RECT 97.8000 32.4000 98.6000 33.6000 ;
	    RECT 105.2000 32.4000 106.0000 39.8000 ;
	    RECT 111.6000 34.3000 112.4000 34.4000 ;
	    RECT 113.2000 34.3000 114.0000 39.8000 ;
	    RECT 117.4000 35.8000 118.6000 39.8000 ;
	    RECT 122.0000 35.8000 122.8000 39.8000 ;
	    RECT 126.4000 36.4000 127.2000 39.8000 ;
	    RECT 126.4000 35.8000 128.4000 36.4000 ;
	    RECT 118.0000 35.0000 118.8000 35.8000 ;
	    RECT 122.2000 35.2000 122.8000 35.8000 ;
	    RECT 121.4000 34.6000 125.0000 35.2000 ;
	    RECT 127.6000 35.0000 128.4000 35.8000 ;
	    RECT 121.4000 34.4000 122.2000 34.6000 ;
	    RECT 124.2000 34.4000 125.0000 34.6000 ;
	    RECT 111.6000 33.7000 114.0000 34.3000 ;
	    RECT 111.6000 33.6000 112.4000 33.7000 ;
	    RECT 89.2000 31.8000 90.6000 32.4000 ;
	    RECT 91.2000 31.8000 92.2000 32.4000 ;
	    RECT 95.6000 31.8000 97.0000 32.4000 ;
	    RECT 97.6000 31.8000 98.6000 32.4000 ;
	    RECT 103.8000 31.8000 106.0000 32.4000 ;
	    RECT 89.2000 31.6000 90.0000 31.8000 ;
	    RECT 78.6000 31.2000 88.4000 31.4000 ;
	    RECT 82.6000 31.0000 88.4000 31.2000 ;
	    RECT 82.8000 30.8000 88.4000 31.0000 ;
	    RECT 81.2000 30.2000 82.0000 30.4000 ;
	    RECT 81.2000 29.6000 86.2000 30.2000 ;
	    RECT 82.8000 29.4000 83.6000 29.6000 ;
	    RECT 85.4000 29.4000 86.2000 29.6000 ;
	    RECT 83.8000 28.4000 84.6000 28.6000 ;
	    RECT 91.2000 28.4000 91.8000 31.8000 ;
	    RECT 95.6000 31.6000 96.4000 31.8000 ;
	    RECT 92.4000 30.3000 93.2000 30.4000 ;
	    RECT 94.0000 30.3000 94.8000 30.4000 ;
	    RECT 92.4000 29.7000 94.8000 30.3000 ;
	    RECT 92.4000 28.8000 93.2000 29.7000 ;
	    RECT 94.0000 29.6000 94.8000 29.7000 ;
	    RECT 97.6000 28.4000 98.2000 31.8000 ;
	    RECT 103.8000 31.2000 104.4000 31.8000 ;
	    RECT 103.2000 30.4000 104.4000 31.2000 ;
	    RECT 113.2000 31.2000 114.0000 33.7000 ;
	    RECT 117.2000 33.2000 118.6000 34.0000 ;
	    RECT 118.0000 32.2000 118.6000 33.2000 ;
	    RECT 120.2000 33.0000 122.4000 33.6000 ;
	    RECT 120.2000 32.8000 121.0000 33.0000 ;
	    RECT 118.0000 31.6000 120.4000 32.2000 ;
	    RECT 113.2000 30.6000 117.4000 31.2000 ;
	    RECT 98.8000 28.8000 99.6000 30.4000 ;
	    RECT 76.6000 27.8000 87.6000 28.4000 ;
	    RECT 77.0000 27.6000 77.8000 27.8000 ;
	    RECT 81.2000 27.6000 82.0000 27.8000 ;
	    RECT 60.6000 26.2000 64.2000 26.6000 ;
	    RECT 39.6000 22.2000 40.4000 26.2000 ;
	    RECT 41.2000 26.0000 45.2000 26.2000 ;
	    RECT 41.2000 22.2000 42.0000 26.0000 ;
	    RECT 44.4000 22.2000 45.2000 26.0000 ;
	    RECT 46.0000 22.2000 46.8000 26.2000 ;
	    RECT 47.6000 26.0000 51.6000 26.2000 ;
	    RECT 47.6000 22.2000 48.4000 26.0000 ;
	    RECT 50.8000 22.2000 51.6000 26.0000 ;
	    RECT 52.4000 26.0000 56.4000 26.2000 ;
	    RECT 52.4000 22.2000 53.2000 26.0000 ;
	    RECT 55.6000 22.2000 56.4000 26.0000 ;
	    RECT 57.2000 22.2000 58.0000 26.2000 ;
	    RECT 58.8000 22.2000 59.6000 26.2000 ;
	    RECT 60.4000 26.0000 64.4000 26.2000 ;
	    RECT 60.4000 22.2000 61.2000 26.0000 ;
	    RECT 63.6000 22.2000 64.4000 26.0000 ;
	    RECT 65.2000 22.2000 66.0000 26.8000 ;
	    RECT 70.0000 26.6000 73.8000 27.2000 ;
	    RECT 70.0000 22.2000 70.8000 26.6000 ;
	    RECT 73.0000 26.4000 73.8000 26.6000 ;
	    RECT 82.8000 25.6000 83.4000 27.8000 ;
	    RECT 86.0000 27.6000 87.6000 27.8000 ;
	    RECT 89.2000 27.6000 91.8000 28.4000 ;
	    RECT 94.0000 28.2000 94.8000 28.4000 ;
	    RECT 93.2000 27.6000 94.8000 28.2000 ;
	    RECT 95.6000 27.6000 98.2000 28.4000 ;
	    RECT 100.4000 28.2000 101.2000 28.4000 ;
	    RECT 99.6000 27.6000 101.2000 28.2000 ;
	    RECT 81.0000 25.4000 81.8000 25.6000 ;
	    RECT 74.8000 24.2000 75.6000 25.0000 ;
	    RECT 79.0000 24.8000 81.8000 25.4000 ;
	    RECT 82.8000 24.8000 83.6000 25.6000 ;
	    RECT 79.0000 24.2000 79.6000 24.8000 ;
	    RECT 84.4000 24.2000 85.2000 25.0000 ;
	    RECT 74.2000 23.6000 75.6000 24.2000 ;
	    RECT 74.2000 22.2000 75.4000 23.6000 ;
	    RECT 78.8000 22.2000 79.6000 24.2000 ;
	    RECT 83.2000 23.6000 85.2000 24.2000 ;
	    RECT 83.2000 22.2000 84.0000 23.6000 ;
	    RECT 87.6000 22.2000 88.4000 27.0000 ;
	    RECT 89.4000 26.2000 90.0000 27.6000 ;
	    RECT 93.2000 27.2000 94.0000 27.6000 ;
	    RECT 91.0000 26.2000 94.6000 26.6000 ;
	    RECT 95.8000 26.2000 96.4000 27.6000 ;
	    RECT 99.6000 27.2000 100.4000 27.6000 ;
	    RECT 103.8000 27.4000 104.4000 30.4000 ;
	    RECT 105.2000 30.3000 106.0000 30.4000 ;
	    RECT 111.6000 30.3000 112.4000 30.4000 ;
	    RECT 105.2000 29.7000 112.4000 30.3000 ;
	    RECT 105.2000 28.8000 106.0000 29.7000 ;
	    RECT 111.6000 29.6000 112.4000 29.7000 ;
	    RECT 103.8000 26.8000 106.0000 27.4000 ;
	    RECT 97.4000 26.2000 101.0000 26.6000 ;
	    RECT 89.2000 22.2000 90.0000 26.2000 ;
	    RECT 90.8000 26.0000 94.8000 26.2000 ;
	    RECT 90.8000 22.2000 91.6000 26.0000 ;
	    RECT 94.0000 22.2000 94.8000 26.0000 ;
	    RECT 95.6000 22.2000 96.4000 26.2000 ;
	    RECT 97.2000 26.0000 101.2000 26.2000 ;
	    RECT 97.2000 22.2000 98.0000 26.0000 ;
	    RECT 100.4000 22.2000 101.2000 26.0000 ;
	    RECT 105.2000 22.2000 106.0000 26.8000 ;
	    RECT 113.2000 27.2000 114.0000 30.6000 ;
	    RECT 116.6000 30.4000 117.4000 30.6000 ;
	    RECT 115.0000 29.8000 115.8000 30.0000 ;
	    RECT 115.0000 29.2000 118.8000 29.8000 ;
	    RECT 118.0000 29.0000 118.8000 29.2000 ;
	    RECT 119.8000 28.4000 120.4000 31.6000 ;
	    RECT 121.8000 31.8000 122.4000 33.0000 ;
	    RECT 123.0000 33.0000 123.8000 33.2000 ;
	    RECT 127.6000 33.0000 128.4000 33.2000 ;
	    RECT 123.0000 32.4000 128.4000 33.0000 ;
	    RECT 121.8000 31.4000 126.6000 31.8000 ;
	    RECT 130.8000 31.4000 131.6000 39.8000 ;
	    RECT 135.0000 38.4000 135.8000 39.8000 ;
	    RECT 134.0000 37.6000 135.8000 38.4000 ;
	    RECT 135.0000 32.4000 135.8000 37.6000 ;
	    RECT 136.4000 33.6000 137.2000 34.4000 ;
	    RECT 136.6000 32.4000 137.2000 33.6000 ;
	    RECT 135.0000 31.8000 136.0000 32.4000 ;
	    RECT 136.6000 31.8000 138.0000 32.4000 ;
	    RECT 121.8000 31.2000 131.6000 31.4000 ;
	    RECT 125.8000 31.0000 131.6000 31.2000 ;
	    RECT 126.0000 30.8000 131.6000 31.0000 ;
	    RECT 124.4000 30.2000 125.2000 30.4000 ;
	    RECT 124.4000 29.6000 129.4000 30.2000 ;
	    RECT 128.6000 29.4000 129.4000 29.6000 ;
	    RECT 134.0000 28.8000 134.8000 30.4000 ;
	    RECT 127.0000 28.4000 127.8000 28.6000 ;
	    RECT 135.4000 28.4000 136.0000 31.8000 ;
	    RECT 137.2000 31.6000 138.0000 31.8000 ;
	    RECT 138.8000 31.2000 139.6000 39.8000 ;
	    RECT 143.0000 35.8000 144.2000 39.8000 ;
	    RECT 147.6000 35.8000 148.4000 39.8000 ;
	    RECT 152.0000 36.4000 152.8000 39.8000 ;
	    RECT 152.0000 35.8000 154.0000 36.4000 ;
	    RECT 143.6000 35.0000 144.4000 35.8000 ;
	    RECT 147.8000 35.2000 148.4000 35.8000 ;
	    RECT 147.0000 34.6000 150.6000 35.2000 ;
	    RECT 153.2000 35.0000 154.0000 35.8000 ;
	    RECT 147.0000 34.4000 147.8000 34.6000 ;
	    RECT 149.8000 34.4000 150.6000 34.6000 ;
	    RECT 142.8000 33.2000 144.2000 34.0000 ;
	    RECT 143.6000 32.2000 144.2000 33.2000 ;
	    RECT 145.8000 33.0000 148.0000 33.6000 ;
	    RECT 145.8000 32.8000 146.6000 33.0000 ;
	    RECT 143.6000 31.6000 146.0000 32.2000 ;
	    RECT 138.8000 30.6000 143.0000 31.2000 ;
	    RECT 119.8000 27.8000 130.8000 28.4000 ;
	    RECT 120.2000 27.6000 121.0000 27.8000 ;
	    RECT 126.0000 27.6000 126.8000 27.8000 ;
	    RECT 129.2000 27.6000 130.8000 27.8000 ;
	    RECT 132.4000 28.2000 133.2000 28.4000 ;
	    RECT 132.4000 27.6000 134.0000 28.2000 ;
	    RECT 135.4000 27.6000 138.0000 28.4000 ;
	    RECT 113.2000 26.6000 117.0000 27.2000 ;
	    RECT 113.2000 22.2000 114.0000 26.6000 ;
	    RECT 116.2000 26.4000 117.0000 26.6000 ;
	    RECT 126.0000 25.6000 126.6000 27.6000 ;
	    RECT 133.2000 27.2000 134.0000 27.6000 ;
	    RECT 124.2000 25.4000 125.0000 25.6000 ;
	    RECT 118.0000 24.2000 118.8000 25.0000 ;
	    RECT 122.2000 24.8000 125.0000 25.4000 ;
	    RECT 126.0000 24.8000 126.8000 25.6000 ;
	    RECT 122.2000 24.2000 122.8000 24.8000 ;
	    RECT 127.6000 24.2000 128.4000 25.0000 ;
	    RECT 117.4000 23.6000 118.8000 24.2000 ;
	    RECT 117.4000 22.2000 118.6000 23.6000 ;
	    RECT 122.0000 22.2000 122.8000 24.2000 ;
	    RECT 126.4000 23.6000 128.4000 24.2000 ;
	    RECT 126.4000 22.2000 127.2000 23.6000 ;
	    RECT 130.8000 22.2000 131.6000 27.0000 ;
	    RECT 132.6000 26.2000 136.2000 26.6000 ;
	    RECT 137.2000 26.2000 137.8000 27.6000 ;
	    RECT 138.8000 27.2000 139.6000 30.6000 ;
	    RECT 142.2000 30.4000 143.0000 30.6000 ;
	    RECT 145.4000 30.4000 146.0000 31.6000 ;
	    RECT 147.4000 31.8000 148.0000 33.0000 ;
	    RECT 148.6000 33.0000 149.4000 33.2000 ;
	    RECT 153.2000 33.0000 154.0000 33.2000 ;
	    RECT 148.6000 32.4000 154.0000 33.0000 ;
	    RECT 147.4000 31.4000 152.2000 31.8000 ;
	    RECT 156.4000 31.4000 157.2000 39.8000 ;
	    RECT 160.2000 38.4000 161.0000 39.8000 ;
	    RECT 167.0000 38.4000 167.8000 39.8000 ;
	    RECT 160.2000 37.6000 162.0000 38.4000 ;
	    RECT 166.0000 37.6000 167.8000 38.4000 ;
	    RECT 158.8000 33.6000 159.6000 34.4000 ;
	    RECT 158.8000 32.4000 159.4000 33.6000 ;
	    RECT 160.2000 32.4000 161.0000 37.6000 ;
	    RECT 158.0000 31.8000 159.4000 32.4000 ;
	    RECT 160.0000 31.8000 161.0000 32.4000 ;
	    RECT 167.0000 32.4000 167.8000 37.6000 ;
	    RECT 168.4000 33.6000 169.2000 34.4000 ;
	    RECT 168.6000 32.4000 169.2000 33.6000 ;
	    RECT 167.0000 31.8000 168.0000 32.4000 ;
	    RECT 168.6000 31.8000 170.0000 32.4000 ;
	    RECT 158.0000 31.6000 158.8000 31.8000 ;
	    RECT 147.4000 31.2000 157.2000 31.4000 ;
	    RECT 151.4000 31.0000 157.2000 31.2000 ;
	    RECT 151.6000 30.8000 157.2000 31.0000 ;
	    RECT 140.6000 29.8000 141.4000 30.0000 ;
	    RECT 140.6000 29.2000 144.4000 29.8000 ;
	    RECT 145.2000 29.6000 146.0000 30.4000 ;
	    RECT 150.0000 30.2000 150.8000 30.4000 ;
	    RECT 150.0000 29.6000 155.0000 30.2000 ;
	    RECT 143.6000 29.0000 144.4000 29.2000 ;
	    RECT 145.4000 28.4000 146.0000 29.6000 ;
	    RECT 151.6000 29.4000 152.4000 29.6000 ;
	    RECT 154.2000 29.4000 155.0000 29.6000 ;
	    RECT 152.6000 28.4000 153.4000 28.6000 ;
	    RECT 160.0000 28.4000 160.6000 31.8000 ;
	    RECT 161.2000 30.3000 162.0000 30.4000 ;
	    RECT 166.0000 30.3000 166.8000 30.4000 ;
	    RECT 161.2000 29.7000 166.8000 30.3000 ;
	    RECT 161.2000 28.8000 162.0000 29.7000 ;
	    RECT 166.0000 28.8000 166.8000 29.7000 ;
	    RECT 167.4000 28.4000 168.0000 31.8000 ;
	    RECT 169.2000 31.6000 170.0000 31.8000 ;
	    RECT 170.8000 31.4000 171.6000 39.8000 ;
	    RECT 175.2000 36.4000 176.0000 39.8000 ;
	    RECT 174.0000 35.8000 176.0000 36.4000 ;
	    RECT 179.6000 35.8000 180.4000 39.8000 ;
	    RECT 183.8000 35.8000 185.0000 39.8000 ;
	    RECT 174.0000 35.0000 174.8000 35.8000 ;
	    RECT 179.6000 35.2000 180.2000 35.8000 ;
	    RECT 177.4000 34.6000 181.0000 35.2000 ;
	    RECT 183.6000 35.0000 184.4000 35.8000 ;
	    RECT 177.4000 34.4000 178.2000 34.6000 ;
	    RECT 180.2000 34.4000 181.0000 34.6000 ;
	    RECT 174.0000 33.0000 174.8000 33.2000 ;
	    RECT 178.6000 33.0000 179.4000 33.2000 ;
	    RECT 174.0000 32.4000 179.4000 33.0000 ;
	    RECT 180.0000 33.0000 182.2000 33.6000 ;
	    RECT 180.0000 31.8000 180.6000 33.0000 ;
	    RECT 181.4000 32.8000 182.2000 33.0000 ;
	    RECT 183.8000 33.2000 185.2000 34.0000 ;
	    RECT 183.8000 32.2000 184.4000 33.2000 ;
	    RECT 175.8000 31.4000 180.6000 31.8000 ;
	    RECT 170.8000 31.2000 180.6000 31.4000 ;
	    RECT 182.0000 31.6000 184.4000 32.2000 ;
	    RECT 170.8000 31.0000 176.6000 31.2000 ;
	    RECT 170.8000 30.8000 176.4000 31.0000 ;
	    RECT 177.2000 30.2000 178.0000 30.4000 ;
	    RECT 173.0000 29.6000 178.0000 30.2000 ;
	    RECT 173.0000 29.4000 173.8000 29.6000 ;
	    RECT 174.6000 28.4000 175.4000 28.6000 ;
	    RECT 182.0000 28.4000 182.6000 31.6000 ;
	    RECT 188.4000 31.2000 189.2000 39.8000 ;
	    RECT 193.8000 32.8000 194.6000 39.8000 ;
	    RECT 198.0000 35.0000 198.8000 39.0000 ;
	    RECT 193.0000 32.2000 194.6000 32.8000 ;
	    RECT 185.0000 30.6000 189.2000 31.2000 ;
	    RECT 185.0000 30.4000 185.8000 30.6000 ;
	    RECT 186.6000 29.8000 187.4000 30.0000 ;
	    RECT 183.6000 29.2000 187.4000 29.8000 ;
	    RECT 183.6000 29.0000 184.4000 29.2000 ;
	    RECT 145.4000 27.8000 156.4000 28.4000 ;
	    RECT 145.8000 27.6000 146.6000 27.8000 ;
	    RECT 138.8000 26.6000 142.6000 27.2000 ;
	    RECT 132.4000 26.0000 136.4000 26.2000 ;
	    RECT 132.4000 22.2000 133.2000 26.0000 ;
	    RECT 135.6000 22.2000 136.4000 26.0000 ;
	    RECT 137.2000 22.2000 138.0000 26.2000 ;
	    RECT 138.8000 22.2000 139.6000 26.6000 ;
	    RECT 141.8000 26.4000 142.6000 26.6000 ;
	    RECT 151.6000 25.6000 152.2000 27.8000 ;
	    RECT 154.8000 27.6000 156.4000 27.8000 ;
	    RECT 158.0000 27.6000 160.6000 28.4000 ;
	    RECT 162.8000 28.3000 163.6000 28.4000 ;
	    RECT 164.4000 28.3000 165.2000 28.4000 ;
	    RECT 162.8000 28.2000 165.2000 28.3000 ;
	    RECT 162.0000 27.7000 166.0000 28.2000 ;
	    RECT 162.0000 27.6000 163.6000 27.7000 ;
	    RECT 164.4000 27.6000 166.0000 27.7000 ;
	    RECT 167.4000 27.6000 170.0000 28.4000 ;
	    RECT 171.6000 27.8000 182.6000 28.4000 ;
	    RECT 171.6000 27.6000 173.2000 27.8000 ;
	    RECT 149.8000 25.4000 150.6000 25.6000 ;
	    RECT 143.6000 24.2000 144.4000 25.0000 ;
	    RECT 147.8000 24.8000 150.6000 25.4000 ;
	    RECT 151.6000 24.8000 152.4000 25.6000 ;
	    RECT 147.8000 24.2000 148.4000 24.8000 ;
	    RECT 153.2000 24.2000 154.0000 25.0000 ;
	    RECT 143.0000 23.6000 144.4000 24.2000 ;
	    RECT 143.0000 22.2000 144.2000 23.6000 ;
	    RECT 147.6000 22.2000 148.4000 24.2000 ;
	    RECT 152.0000 23.6000 154.0000 24.2000 ;
	    RECT 152.0000 22.2000 152.8000 23.6000 ;
	    RECT 156.4000 22.2000 157.2000 27.0000 ;
	    RECT 158.2000 26.2000 158.8000 27.6000 ;
	    RECT 162.0000 27.2000 162.8000 27.6000 ;
	    RECT 165.2000 27.2000 166.0000 27.6000 ;
	    RECT 159.8000 26.2000 163.4000 26.6000 ;
	    RECT 164.6000 26.2000 168.2000 26.6000 ;
	    RECT 169.2000 26.2000 169.8000 27.6000 ;
	    RECT 158.0000 22.2000 158.8000 26.2000 ;
	    RECT 159.6000 26.0000 163.6000 26.2000 ;
	    RECT 159.6000 22.2000 160.4000 26.0000 ;
	    RECT 162.8000 22.2000 163.6000 26.0000 ;
	    RECT 164.4000 26.0000 168.4000 26.2000 ;
	    RECT 164.4000 22.2000 165.2000 26.0000 ;
	    RECT 167.6000 22.2000 168.4000 26.0000 ;
	    RECT 169.2000 22.2000 170.0000 26.2000 ;
	    RECT 170.8000 22.2000 171.6000 27.0000 ;
	    RECT 175.8000 25.6000 176.4000 27.8000 ;
	    RECT 181.4000 27.6000 182.2000 27.8000 ;
	    RECT 188.4000 27.2000 189.2000 30.6000 ;
	    RECT 191.6000 29.6000 192.4000 31.2000 ;
	    RECT 193.0000 28.4000 193.6000 32.2000 ;
	    RECT 198.2000 31.6000 198.8000 35.0000 ;
	    RECT 203.4000 32.8000 204.2000 39.8000 ;
	    RECT 207.6000 35.0000 208.4000 39.0000 ;
	    RECT 195.0000 31.0000 198.8000 31.6000 ;
	    RECT 202.6000 32.2000 204.2000 32.8000 ;
	    RECT 195.0000 29.0000 195.6000 31.0000 ;
	    RECT 191.6000 27.6000 193.6000 28.4000 ;
	    RECT 194.2000 28.2000 195.6000 29.0000 ;
	    RECT 196.4000 28.8000 197.2000 30.4000 ;
	    RECT 198.0000 28.8000 198.8000 30.4000 ;
	    RECT 201.2000 29.6000 202.0000 31.2000 ;
	    RECT 202.6000 28.4000 203.2000 32.2000 ;
	    RECT 207.8000 31.6000 208.4000 35.0000 ;
	    RECT 209.2000 32.4000 210.0000 39.8000 ;
	    RECT 209.2000 31.8000 211.4000 32.4000 ;
	    RECT 212.4000 31.8000 213.2000 39.8000 ;
	    RECT 216.6000 31.8000 218.6000 39.8000 ;
	    RECT 222.8000 33.6000 223.6000 34.4000 ;
	    RECT 222.8000 32.4000 223.4000 33.6000 ;
	    RECT 224.2000 32.4000 225.0000 39.8000 ;
	    RECT 232.2000 38.4000 233.0000 39.8000 ;
	    RECT 231.6000 37.6000 233.0000 38.4000 ;
	    RECT 232.2000 32.8000 233.0000 37.6000 ;
	    RECT 236.4000 35.0000 237.2000 39.0000 ;
	    RECT 222.0000 31.8000 223.4000 32.4000 ;
	    RECT 224.0000 31.8000 225.0000 32.4000 ;
	    RECT 231.4000 32.2000 233.0000 32.8000 ;
	    RECT 204.6000 31.0000 208.4000 31.6000 ;
	    RECT 210.8000 31.2000 211.4000 31.8000 ;
	    RECT 204.6000 29.0000 205.2000 31.0000 ;
	    RECT 210.8000 30.4000 212.0000 31.2000 ;
	    RECT 185.2000 26.6000 189.2000 27.2000 ;
	    RECT 185.2000 26.4000 186.2000 26.6000 ;
	    RECT 185.2000 25.6000 186.0000 26.4000 ;
	    RECT 174.0000 24.2000 174.8000 25.0000 ;
	    RECT 175.6000 24.8000 176.4000 25.6000 ;
	    RECT 177.4000 25.4000 178.2000 25.6000 ;
	    RECT 177.4000 24.8000 180.2000 25.4000 ;
	    RECT 179.6000 24.2000 180.2000 24.8000 ;
	    RECT 183.6000 24.2000 184.4000 25.0000 ;
	    RECT 174.0000 23.6000 176.0000 24.2000 ;
	    RECT 175.2000 22.2000 176.0000 23.6000 ;
	    RECT 179.6000 22.2000 180.4000 24.2000 ;
	    RECT 183.6000 23.6000 185.0000 24.2000 ;
	    RECT 183.8000 22.2000 185.0000 23.6000 ;
	    RECT 188.4000 22.2000 189.2000 26.6000 ;
	    RECT 193.0000 27.0000 193.6000 27.6000 ;
	    RECT 194.6000 27.8000 195.6000 28.2000 ;
	    RECT 194.6000 27.2000 198.8000 27.8000 ;
	    RECT 201.2000 27.6000 203.2000 28.4000 ;
	    RECT 203.8000 28.2000 205.2000 29.0000 ;
	    RECT 206.0000 28.8000 206.8000 30.4000 ;
	    RECT 207.6000 28.8000 208.4000 30.4000 ;
	    RECT 193.0000 26.6000 193.8000 27.0000 ;
	    RECT 193.0000 26.4000 194.6000 26.6000 ;
	    RECT 193.0000 26.0000 195.6000 26.4000 ;
	    RECT 193.8000 25.6000 195.6000 26.0000 ;
	    RECT 193.8000 23.0000 194.6000 25.6000 ;
	    RECT 198.2000 25.0000 198.8000 27.2000 ;
	    RECT 202.6000 27.0000 203.2000 27.6000 ;
	    RECT 204.2000 27.8000 205.2000 28.2000 ;
	    RECT 204.2000 27.2000 208.4000 27.8000 ;
	    RECT 210.8000 27.4000 211.4000 30.4000 ;
	    RECT 212.6000 29.6000 213.2000 31.8000 ;
	    RECT 202.6000 26.6000 203.4000 27.0000 ;
	    RECT 202.6000 26.0000 204.2000 26.6000 ;
	    RECT 198.0000 23.0000 198.8000 25.0000 ;
	    RECT 203.4000 23.0000 204.2000 26.0000 ;
	    RECT 207.8000 25.0000 208.4000 27.2000 ;
	    RECT 207.6000 23.0000 208.4000 25.0000 ;
	    RECT 209.2000 26.8000 211.4000 27.4000 ;
	    RECT 212.4000 28.3000 213.2000 29.6000 ;
	    RECT 214.0000 28.3000 214.8000 30.4000 ;
	    RECT 215.6000 28.8000 216.4000 30.4000 ;
	    RECT 217.4000 28.4000 218.0000 31.8000 ;
	    RECT 222.0000 31.6000 222.8000 31.8000 ;
	    RECT 218.8000 28.8000 219.6000 30.4000 ;
	    RECT 224.0000 28.4000 224.6000 31.8000 ;
	    RECT 225.2000 28.8000 226.0000 30.4000 ;
	    RECT 230.0000 29.6000 230.8000 31.2000 ;
	    RECT 231.4000 28.4000 232.0000 32.2000 ;
	    RECT 236.6000 31.6000 237.2000 35.0000 ;
	    RECT 240.6000 32.6000 241.4000 39.8000 ;
	    RECT 246.6000 38.4000 247.4000 39.8000 ;
	    RECT 246.0000 37.6000 247.4000 38.4000 ;
	    RECT 246.6000 32.8000 247.4000 37.6000 ;
	    RECT 250.8000 35.0000 251.6000 39.0000 ;
	    RECT 261.4000 36.4000 263.4000 39.8000 ;
	    RECT 260.4000 35.6000 263.4000 36.4000 ;
	    RECT 239.6000 31.8000 241.4000 32.6000 ;
	    RECT 245.8000 32.2000 247.4000 32.8000 ;
	    RECT 233.4000 31.0000 237.2000 31.6000 ;
	    RECT 233.4000 29.0000 234.0000 31.0000 ;
	    RECT 212.4000 27.7000 214.8000 28.3000 ;
	    RECT 217.2000 28.2000 218.0000 28.4000 ;
	    RECT 220.4000 28.3000 221.2000 28.4000 ;
	    RECT 222.0000 28.3000 224.6000 28.4000 ;
	    RECT 220.4000 28.2000 224.6000 28.3000 ;
	    RECT 226.8000 28.2000 227.6000 28.4000 ;
	    RECT 209.2000 22.2000 210.0000 26.8000 ;
	    RECT 212.4000 22.2000 213.2000 27.7000 ;
	    RECT 214.0000 27.6000 214.8000 27.7000 ;
	    RECT 215.6000 27.6000 218.0000 28.2000 ;
	    RECT 219.6000 27.7000 224.6000 28.2000 ;
	    RECT 219.6000 27.6000 221.2000 27.7000 ;
	    RECT 222.0000 27.6000 224.6000 27.7000 ;
	    RECT 226.0000 27.6000 227.6000 28.2000 ;
	    RECT 230.0000 27.6000 232.0000 28.4000 ;
	    RECT 232.6000 28.2000 234.0000 29.0000 ;
	    RECT 234.8000 28.8000 235.6000 30.4000 ;
	    RECT 236.4000 28.8000 237.2000 30.4000 ;
	    RECT 239.8000 28.4000 240.4000 31.8000 ;
	    RECT 241.2000 30.3000 242.0000 31.2000 ;
	    RECT 242.8000 30.3000 243.6000 30.4000 ;
	    RECT 241.2000 29.7000 243.6000 30.3000 ;
	    RECT 241.2000 29.6000 242.0000 29.7000 ;
	    RECT 242.8000 29.6000 243.6000 29.7000 ;
	    RECT 244.4000 29.6000 245.2000 31.2000 ;
	    RECT 245.8000 28.4000 246.4000 32.2000 ;
	    RECT 251.0000 31.6000 251.6000 35.0000 ;
	    RECT 261.4000 31.8000 263.4000 35.6000 ;
	    RECT 267.4000 32.6000 268.2000 39.8000 ;
	    RECT 272.4000 33.6000 273.2000 34.4000 ;
	    RECT 267.4000 31.8000 269.2000 32.6000 ;
	    RECT 272.4000 32.4000 273.0000 33.6000 ;
	    RECT 273.8000 32.4000 274.6000 39.8000 ;
	    RECT 271.6000 31.8000 273.0000 32.4000 ;
	    RECT 273.6000 31.8000 274.6000 32.4000 ;
	    RECT 247.8000 31.0000 251.6000 31.6000 ;
	    RECT 247.8000 29.0000 248.4000 31.0000 ;
	    RECT 215.6000 26.2000 216.2000 27.6000 ;
	    RECT 219.6000 27.2000 220.4000 27.6000 ;
	    RECT 217.4000 26.2000 221.0000 26.6000 ;
	    RECT 222.2000 26.2000 222.8000 27.6000 ;
	    RECT 226.0000 27.2000 226.8000 27.6000 ;
	    RECT 231.4000 27.0000 232.0000 27.6000 ;
	    RECT 233.0000 27.8000 234.0000 28.2000 ;
	    RECT 233.0000 27.2000 237.2000 27.8000 ;
	    RECT 239.6000 27.6000 240.4000 28.4000 ;
	    RECT 244.4000 27.6000 246.4000 28.4000 ;
	    RECT 247.0000 28.2000 248.4000 29.0000 ;
	    RECT 249.2000 28.8000 250.0000 30.4000 ;
	    RECT 250.8000 28.8000 251.6000 30.4000 ;
	    RECT 231.4000 26.6000 232.2000 27.0000 ;
	    RECT 223.8000 26.2000 227.4000 26.6000 ;
	    RECT 214.0000 22.8000 214.8000 26.2000 ;
	    RECT 215.6000 23.4000 216.4000 26.2000 ;
	    RECT 217.2000 26.0000 221.2000 26.2000 ;
	    RECT 217.2000 22.8000 218.0000 26.0000 ;
	    RECT 214.0000 22.2000 218.0000 22.8000 ;
	    RECT 220.4000 22.2000 221.2000 26.0000 ;
	    RECT 222.0000 22.2000 222.8000 26.2000 ;
	    RECT 223.6000 26.0000 227.6000 26.2000 ;
	    RECT 231.4000 26.0000 233.0000 26.6000 ;
	    RECT 223.6000 22.2000 224.4000 26.0000 ;
	    RECT 226.8000 22.2000 227.6000 26.0000 ;
	    RECT 232.2000 23.0000 233.0000 26.0000 ;
	    RECT 236.6000 25.0000 237.2000 27.2000 ;
	    RECT 236.4000 23.0000 237.2000 25.0000 ;
	    RECT 238.0000 24.8000 238.8000 26.4000 ;
	    RECT 239.8000 24.4000 240.4000 27.6000 ;
	    RECT 245.8000 27.0000 246.4000 27.6000 ;
	    RECT 247.4000 27.8000 248.4000 28.2000 ;
	    RECT 257.2000 28.3000 258.0000 28.4000 ;
	    RECT 258.8000 28.3000 259.6000 29.2000 ;
	    RECT 260.4000 28.8000 261.2000 30.4000 ;
	    RECT 262.2000 28.4000 262.8000 31.8000 ;
	    RECT 263.6000 28.8000 264.4000 30.4000 ;
	    RECT 266.8000 29.6000 267.6000 31.2000 ;
	    RECT 268.4000 30.4000 269.0000 31.8000 ;
	    RECT 271.6000 31.6000 272.4000 31.8000 ;
	    RECT 268.4000 29.6000 269.2000 30.4000 ;
	    RECT 270.0000 30.3000 270.8000 30.4000 ;
	    RECT 273.6000 30.3000 274.2000 31.8000 ;
	    RECT 278.0000 31.2000 278.8000 39.8000 ;
	    RECT 282.2000 35.8000 283.4000 39.8000 ;
	    RECT 286.8000 35.8000 287.6000 39.8000 ;
	    RECT 291.2000 36.4000 292.0000 39.8000 ;
	    RECT 291.2000 35.8000 293.2000 36.4000 ;
	    RECT 282.8000 35.0000 283.6000 35.8000 ;
	    RECT 287.0000 35.2000 287.6000 35.8000 ;
	    RECT 286.2000 34.6000 289.8000 35.2000 ;
	    RECT 292.4000 35.0000 293.2000 35.8000 ;
	    RECT 286.2000 34.4000 287.0000 34.6000 ;
	    RECT 289.0000 34.4000 289.8000 34.6000 ;
	    RECT 282.0000 33.2000 283.4000 34.0000 ;
	    RECT 282.8000 32.2000 283.4000 33.2000 ;
	    RECT 285.0000 33.0000 287.2000 33.6000 ;
	    RECT 285.0000 32.8000 285.8000 33.0000 ;
	    RECT 282.8000 31.6000 285.2000 32.2000 ;
	    RECT 278.0000 30.6000 282.2000 31.2000 ;
	    RECT 270.0000 29.7000 274.2000 30.3000 ;
	    RECT 270.0000 29.6000 270.8000 29.7000 ;
	    RECT 268.4000 28.4000 269.0000 29.6000 ;
	    RECT 273.6000 28.4000 274.2000 29.7000 ;
	    RECT 274.8000 28.8000 275.6000 30.4000 ;
	    RECT 247.4000 27.2000 251.6000 27.8000 ;
	    RECT 257.2000 27.7000 259.6000 28.3000 ;
	    RECT 262.0000 28.2000 262.8000 28.4000 ;
	    RECT 265.2000 28.2000 266.0000 28.4000 ;
	    RECT 257.2000 27.6000 258.0000 27.7000 ;
	    RECT 258.8000 27.6000 259.6000 27.7000 ;
	    RECT 260.4000 27.6000 262.8000 28.2000 ;
	    RECT 264.4000 27.6000 266.0000 28.2000 ;
	    RECT 268.4000 27.6000 269.2000 28.4000 ;
	    RECT 271.6000 27.6000 274.2000 28.4000 ;
	    RECT 276.4000 28.2000 277.2000 28.4000 ;
	    RECT 275.6000 27.6000 277.2000 28.2000 ;
	    RECT 245.8000 26.6000 246.6000 27.0000 ;
	    RECT 245.8000 26.0000 247.4000 26.6000 ;
	    RECT 239.6000 22.2000 240.4000 24.4000 ;
	    RECT 246.6000 23.0000 247.4000 26.0000 ;
	    RECT 251.0000 25.0000 251.6000 27.2000 ;
	    RECT 260.4000 26.2000 261.0000 27.6000 ;
	    RECT 264.4000 27.2000 265.2000 27.6000 ;
	    RECT 262.2000 26.2000 265.8000 26.6000 ;
	    RECT 250.8000 23.0000 251.6000 25.0000 ;
	    RECT 258.8000 22.8000 259.6000 26.2000 ;
	    RECT 260.4000 23.4000 261.2000 26.2000 ;
	    RECT 262.0000 26.0000 266.0000 26.2000 ;
	    RECT 262.0000 22.8000 262.8000 26.0000 ;
	    RECT 258.8000 22.2000 262.8000 22.8000 ;
	    RECT 265.2000 22.2000 266.0000 26.0000 ;
	    RECT 268.4000 24.2000 269.0000 27.6000 ;
	    RECT 270.0000 24.8000 270.8000 26.4000 ;
	    RECT 271.8000 26.2000 272.4000 27.6000 ;
	    RECT 275.6000 27.2000 276.4000 27.6000 ;
	    RECT 278.0000 27.2000 278.8000 30.6000 ;
	    RECT 281.4000 30.4000 282.2000 30.6000 ;
	    RECT 279.8000 29.8000 280.6000 30.0000 ;
	    RECT 279.8000 29.2000 283.6000 29.8000 ;
	    RECT 282.8000 29.0000 283.6000 29.2000 ;
	    RECT 284.6000 28.4000 285.2000 31.6000 ;
	    RECT 286.6000 31.8000 287.2000 33.0000 ;
	    RECT 287.8000 33.0000 288.6000 33.2000 ;
	    RECT 292.4000 33.0000 293.2000 33.2000 ;
	    RECT 287.8000 32.4000 293.2000 33.0000 ;
	    RECT 286.6000 31.4000 291.4000 31.8000 ;
	    RECT 295.6000 31.4000 296.4000 39.8000 ;
	    RECT 299.8000 32.4000 300.6000 39.8000 ;
	    RECT 301.2000 33.6000 302.0000 34.4000 ;
	    RECT 301.4000 32.4000 302.0000 33.6000 ;
	    RECT 304.4000 33.6000 305.2000 34.4000 ;
	    RECT 304.4000 32.4000 305.0000 33.6000 ;
	    RECT 305.8000 32.4000 306.6000 39.8000 ;
	    RECT 313.8000 32.8000 314.6000 39.8000 ;
	    RECT 318.0000 35.0000 318.8000 39.0000 ;
	    RECT 299.8000 31.8000 300.8000 32.4000 ;
	    RECT 301.4000 31.8000 302.8000 32.4000 ;
	    RECT 286.6000 31.2000 296.4000 31.4000 ;
	    RECT 290.6000 31.0000 296.4000 31.2000 ;
	    RECT 290.8000 30.8000 296.4000 31.0000 ;
	    RECT 300.2000 30.4000 300.8000 31.8000 ;
	    RECT 302.0000 31.6000 302.8000 31.8000 ;
	    RECT 303.6000 31.8000 305.0000 32.4000 ;
	    RECT 305.6000 31.8000 306.6000 32.4000 ;
	    RECT 313.0000 32.2000 314.6000 32.8000 ;
	    RECT 303.6000 31.6000 304.4000 31.8000 ;
	    RECT 289.2000 30.2000 290.0000 30.4000 ;
	    RECT 289.2000 29.6000 294.2000 30.2000 ;
	    RECT 293.4000 29.4000 294.2000 29.6000 ;
	    RECT 298.8000 28.8000 299.6000 30.4000 ;
	    RECT 300.2000 29.6000 301.2000 30.4000 ;
	    RECT 302.1000 30.3000 302.7000 31.6000 ;
	    RECT 305.6000 30.3000 306.2000 31.8000 ;
	    RECT 302.1000 29.7000 306.2000 30.3000 ;
	    RECT 291.8000 28.4000 292.6000 28.6000 ;
	    RECT 300.2000 28.4000 300.8000 29.6000 ;
	    RECT 305.6000 28.4000 306.2000 29.7000 ;
	    RECT 306.8000 28.8000 307.6000 30.4000 ;
	    RECT 311.6000 29.6000 312.4000 31.2000 ;
	    RECT 313.0000 28.4000 313.6000 32.2000 ;
	    RECT 318.2000 31.6000 318.8000 35.0000 ;
	    RECT 322.2000 32.4000 323.0000 39.8000 ;
	    RECT 323.6000 33.6000 324.4000 34.4000 ;
	    RECT 323.8000 32.4000 324.4000 33.6000 ;
	    RECT 328.6000 32.4000 330.6000 39.8000 ;
	    RECT 322.2000 31.8000 323.2000 32.4000 ;
	    RECT 323.8000 31.8000 325.2000 32.4000 ;
	    RECT 315.0000 31.0000 318.8000 31.6000 ;
	    RECT 315.0000 29.0000 315.6000 31.0000 ;
	    RECT 284.6000 27.8000 295.6000 28.4000 ;
	    RECT 285.0000 27.6000 285.8000 27.8000 ;
	    RECT 290.8000 27.6000 291.6000 27.8000 ;
	    RECT 294.0000 27.6000 295.6000 27.8000 ;
	    RECT 297.2000 28.2000 298.0000 28.4000 ;
	    RECT 297.2000 27.6000 298.8000 28.2000 ;
	    RECT 300.2000 27.6000 302.8000 28.4000 ;
	    RECT 303.6000 27.6000 306.2000 28.4000 ;
	    RECT 308.4000 28.2000 309.2000 28.4000 ;
	    RECT 307.6000 27.6000 309.2000 28.2000 ;
	    RECT 310.0000 28.3000 310.8000 28.4000 ;
	    RECT 311.6000 28.3000 313.6000 28.4000 ;
	    RECT 310.0000 27.7000 313.6000 28.3000 ;
	    RECT 314.2000 28.2000 315.6000 29.0000 ;
	    RECT 316.4000 28.8000 317.2000 30.4000 ;
	    RECT 318.0000 28.8000 318.8000 30.4000 ;
	    RECT 321.2000 28.8000 322.0000 30.4000 ;
	    RECT 322.6000 28.4000 323.2000 31.8000 ;
	    RECT 324.4000 31.6000 325.2000 31.8000 ;
	    RECT 327.6000 31.8000 330.6000 32.4000 ;
	    RECT 334.0000 35.0000 334.8000 39.0000 ;
	    RECT 338.2000 38.4000 339.0000 39.8000 ;
	    RECT 337.2000 37.6000 339.0000 38.4000 ;
	    RECT 327.6000 31.6000 329.8000 31.8000 ;
	    RECT 326.0000 30.3000 326.8000 30.4000 ;
	    RECT 327.6000 30.3000 328.4000 30.4000 ;
	    RECT 326.0000 29.7000 328.4000 30.3000 ;
	    RECT 326.0000 29.6000 326.8000 29.7000 ;
	    RECT 327.6000 28.8000 328.4000 29.7000 ;
	    RECT 329.2000 28.4000 329.8000 31.6000 ;
	    RECT 334.0000 31.6000 334.6000 35.0000 ;
	    RECT 338.2000 32.8000 339.0000 37.6000 ;
	    RECT 338.2000 32.2000 339.8000 32.8000 ;
	    RECT 334.0000 31.0000 337.8000 31.6000 ;
	    RECT 330.8000 28.8000 331.6000 30.4000 ;
	    RECT 310.0000 27.6000 310.8000 27.7000 ;
	    RECT 311.6000 27.6000 313.6000 27.7000 ;
	    RECT 278.0000 26.6000 281.8000 27.2000 ;
	    RECT 273.4000 26.2000 277.0000 26.6000 ;
	    RECT 268.4000 22.2000 269.2000 24.2000 ;
	    RECT 271.6000 22.2000 272.4000 26.2000 ;
	    RECT 273.2000 26.0000 277.2000 26.2000 ;
	    RECT 273.2000 22.2000 274.0000 26.0000 ;
	    RECT 276.4000 22.2000 277.2000 26.0000 ;
	    RECT 278.0000 22.2000 278.8000 26.6000 ;
	    RECT 281.0000 26.4000 281.8000 26.6000 ;
	    RECT 290.8000 25.6000 291.4000 27.6000 ;
	    RECT 298.0000 27.2000 298.8000 27.6000 ;
	    RECT 289.0000 25.4000 289.8000 25.6000 ;
	    RECT 282.8000 24.2000 283.6000 25.0000 ;
	    RECT 287.0000 24.8000 289.8000 25.4000 ;
	    RECT 290.8000 24.8000 291.6000 25.6000 ;
	    RECT 287.0000 24.2000 287.6000 24.8000 ;
	    RECT 292.4000 24.2000 293.2000 25.0000 ;
	    RECT 282.2000 23.6000 283.6000 24.2000 ;
	    RECT 282.2000 22.2000 283.4000 23.6000 ;
	    RECT 286.8000 22.2000 287.6000 24.2000 ;
	    RECT 291.2000 23.6000 293.2000 24.2000 ;
	    RECT 291.2000 22.2000 292.0000 23.6000 ;
	    RECT 295.6000 22.2000 296.4000 27.0000 ;
	    RECT 297.4000 26.2000 301.0000 26.6000 ;
	    RECT 302.0000 26.2000 302.6000 27.6000 ;
	    RECT 303.8000 26.2000 304.4000 27.6000 ;
	    RECT 307.6000 27.2000 308.4000 27.6000 ;
	    RECT 313.0000 27.0000 313.6000 27.6000 ;
	    RECT 314.6000 27.8000 315.6000 28.2000 ;
	    RECT 319.6000 28.2000 320.4000 28.4000 ;
	    RECT 322.6000 28.3000 325.2000 28.4000 ;
	    RECT 326.0000 28.3000 326.8000 28.4000 ;
	    RECT 322.6000 28.2000 326.8000 28.3000 ;
	    RECT 329.2000 28.2000 330.0000 28.4000 ;
	    RECT 314.6000 27.2000 318.8000 27.8000 ;
	    RECT 319.6000 27.6000 321.2000 28.2000 ;
	    RECT 322.6000 27.7000 327.6000 28.2000 ;
	    RECT 322.6000 27.6000 325.2000 27.7000 ;
	    RECT 326.0000 27.6000 327.6000 27.7000 ;
	    RECT 329.2000 27.6000 331.6000 28.2000 ;
	    RECT 332.4000 27.6000 333.2000 29.2000 ;
	    RECT 334.0000 28.8000 334.8000 30.4000 ;
	    RECT 335.6000 28.8000 336.4000 30.4000 ;
	    RECT 337.2000 29.0000 337.8000 31.0000 ;
	    RECT 337.2000 28.2000 338.6000 29.0000 ;
	    RECT 339.2000 28.4000 339.8000 32.2000 ;
	    RECT 343.6000 31.2000 344.4000 39.8000 ;
	    RECT 347.8000 35.8000 349.0000 39.8000 ;
	    RECT 352.4000 35.8000 353.2000 39.8000 ;
	    RECT 356.8000 36.4000 357.6000 39.8000 ;
	    RECT 356.8000 35.8000 358.8000 36.4000 ;
	    RECT 348.4000 35.0000 349.2000 35.8000 ;
	    RECT 352.6000 35.2000 353.2000 35.8000 ;
	    RECT 351.8000 34.6000 355.4000 35.2000 ;
	    RECT 358.0000 35.0000 358.8000 35.8000 ;
	    RECT 351.8000 34.4000 352.6000 34.6000 ;
	    RECT 354.6000 34.4000 355.4000 34.6000 ;
	    RECT 346.8000 34.0000 348.2000 34.4000 ;
	    RECT 346.8000 33.6000 349.0000 34.0000 ;
	    RECT 347.6000 33.2000 349.0000 33.6000 ;
	    RECT 348.4000 32.2000 349.0000 33.2000 ;
	    RECT 350.6000 33.0000 352.8000 33.6000 ;
	    RECT 350.6000 32.8000 351.4000 33.0000 ;
	    RECT 348.4000 31.6000 350.8000 32.2000 ;
	    RECT 340.4000 30.3000 341.2000 31.2000 ;
	    RECT 343.6000 30.6000 347.8000 31.2000 ;
	    RECT 342.0000 30.3000 342.8000 30.4000 ;
	    RECT 340.4000 29.7000 342.8000 30.3000 ;
	    RECT 340.4000 29.6000 341.2000 29.7000 ;
	    RECT 342.0000 29.6000 342.8000 29.7000 ;
	    RECT 337.2000 27.8000 338.2000 28.2000 ;
	    RECT 320.4000 27.2000 321.2000 27.6000 ;
	    RECT 313.0000 26.6000 313.8000 27.0000 ;
	    RECT 305.4000 26.2000 309.0000 26.6000 ;
	    RECT 297.2000 26.0000 301.2000 26.2000 ;
	    RECT 297.2000 22.2000 298.0000 26.0000 ;
	    RECT 300.4000 22.2000 301.2000 26.0000 ;
	    RECT 302.0000 22.2000 302.8000 26.2000 ;
	    RECT 303.6000 22.2000 304.4000 26.2000 ;
	    RECT 305.2000 26.0000 309.2000 26.2000 ;
	    RECT 313.0000 26.0000 314.6000 26.6000 ;
	    RECT 305.2000 22.2000 306.0000 26.0000 ;
	    RECT 308.4000 22.2000 309.2000 26.0000 ;
	    RECT 313.8000 23.0000 314.6000 26.0000 ;
	    RECT 318.2000 25.0000 318.8000 27.2000 ;
	    RECT 319.8000 26.2000 323.4000 26.6000 ;
	    RECT 324.4000 26.2000 325.0000 27.6000 ;
	    RECT 326.8000 27.2000 327.6000 27.6000 ;
	    RECT 326.2000 26.2000 329.8000 26.6000 ;
	    RECT 331.0000 26.2000 331.6000 27.6000 ;
	    RECT 334.0000 27.2000 338.2000 27.8000 ;
	    RECT 339.2000 27.6000 341.2000 28.4000 ;
	    RECT 318.0000 23.0000 318.8000 25.0000 ;
	    RECT 319.6000 26.0000 323.6000 26.2000 ;
	    RECT 319.6000 22.2000 320.4000 26.0000 ;
	    RECT 322.8000 22.2000 323.6000 26.0000 ;
	    RECT 324.4000 22.2000 325.2000 26.2000 ;
	    RECT 326.0000 26.0000 330.0000 26.2000 ;
	    RECT 326.0000 22.2000 326.8000 26.0000 ;
	    RECT 329.2000 22.8000 330.0000 26.0000 ;
	    RECT 330.8000 23.4000 331.6000 26.2000 ;
	    RECT 332.4000 22.8000 333.2000 26.2000 ;
	    RECT 334.0000 25.0000 334.6000 27.2000 ;
	    RECT 339.2000 27.0000 339.8000 27.6000 ;
	    RECT 339.0000 26.6000 339.8000 27.0000 ;
	    RECT 338.2000 26.0000 339.8000 26.6000 ;
	    RECT 343.6000 27.2000 344.4000 30.6000 ;
	    RECT 347.0000 30.4000 347.8000 30.6000 ;
	    RECT 345.4000 29.8000 346.2000 30.0000 ;
	    RECT 345.4000 29.2000 349.2000 29.8000 ;
	    RECT 348.4000 29.0000 349.2000 29.2000 ;
	    RECT 350.2000 28.4000 350.8000 31.6000 ;
	    RECT 352.2000 31.8000 352.8000 33.0000 ;
	    RECT 353.4000 33.0000 354.2000 33.2000 ;
	    RECT 358.0000 33.0000 358.8000 33.2000 ;
	    RECT 353.4000 32.4000 358.8000 33.0000 ;
	    RECT 352.2000 31.4000 357.0000 31.8000 ;
	    RECT 361.2000 31.4000 362.0000 39.8000 ;
	    RECT 363.6000 33.6000 364.4000 34.4000 ;
	    RECT 363.6000 32.4000 364.2000 33.6000 ;
	    RECT 365.0000 32.4000 365.8000 39.8000 ;
	    RECT 362.8000 31.8000 364.2000 32.4000 ;
	    RECT 364.8000 31.8000 365.8000 32.4000 ;
	    RECT 371.8000 32.4000 372.6000 39.8000 ;
	    RECT 373.2000 33.6000 374.0000 34.4000 ;
	    RECT 373.4000 32.4000 374.0000 33.6000 ;
	    RECT 376.4000 33.6000 377.2000 34.4000 ;
	    RECT 376.4000 32.4000 377.0000 33.6000 ;
	    RECT 377.8000 32.4000 378.6000 39.8000 ;
	    RECT 371.8000 31.8000 372.8000 32.4000 ;
	    RECT 373.4000 31.8000 374.8000 32.4000 ;
	    RECT 362.8000 31.6000 363.6000 31.8000 ;
	    RECT 352.2000 31.2000 362.0000 31.4000 ;
	    RECT 356.2000 31.0000 362.0000 31.2000 ;
	    RECT 356.4000 30.8000 362.0000 31.0000 ;
	    RECT 364.8000 30.4000 365.4000 31.8000 ;
	    RECT 354.8000 30.2000 355.6000 30.4000 ;
	    RECT 354.8000 29.6000 359.8000 30.2000 ;
	    RECT 364.4000 29.6000 365.4000 30.4000 ;
	    RECT 356.4000 29.4000 357.2000 29.6000 ;
	    RECT 359.0000 29.4000 359.8000 29.6000 ;
	    RECT 357.4000 28.4000 358.2000 28.6000 ;
	    RECT 364.8000 28.4000 365.4000 29.6000 ;
	    RECT 366.0000 28.8000 366.8000 30.4000 ;
	    RECT 369.2000 30.3000 370.0000 30.4000 ;
	    RECT 370.8000 30.3000 371.6000 30.4000 ;
	    RECT 369.2000 29.7000 371.6000 30.3000 ;
	    RECT 369.2000 29.6000 370.0000 29.7000 ;
	    RECT 370.8000 28.8000 371.6000 29.7000 ;
	    RECT 372.2000 30.3000 372.8000 31.8000 ;
	    RECT 374.0000 31.6000 374.8000 31.8000 ;
	    RECT 375.6000 31.8000 377.0000 32.4000 ;
	    RECT 377.6000 31.8000 378.6000 32.4000 ;
	    RECT 375.6000 31.6000 376.4000 31.8000 ;
	    RECT 375.7000 30.3000 376.3000 31.6000 ;
	    RECT 372.2000 29.7000 376.3000 30.3000 ;
	    RECT 372.2000 28.4000 372.8000 29.7000 ;
	    RECT 377.6000 28.4000 378.2000 31.8000 ;
	    RECT 382.0000 31.2000 382.8000 39.8000 ;
	    RECT 386.2000 35.8000 387.4000 39.8000 ;
	    RECT 390.8000 35.8000 391.6000 39.8000 ;
	    RECT 395.2000 36.4000 396.0000 39.8000 ;
	    RECT 395.2000 35.8000 397.2000 36.4000 ;
	    RECT 386.8000 35.0000 387.6000 35.8000 ;
	    RECT 391.0000 35.2000 391.6000 35.8000 ;
	    RECT 390.2000 34.6000 393.8000 35.2000 ;
	    RECT 396.4000 35.0000 397.2000 35.8000 ;
	    RECT 390.2000 34.4000 391.0000 34.6000 ;
	    RECT 393.0000 34.4000 393.8000 34.6000 ;
	    RECT 385.2000 34.0000 386.6000 34.4000 ;
	    RECT 385.2000 33.6000 387.4000 34.0000 ;
	    RECT 386.0000 33.2000 387.4000 33.6000 ;
	    RECT 386.8000 32.2000 387.4000 33.2000 ;
	    RECT 389.0000 33.0000 391.2000 33.6000 ;
	    RECT 389.0000 32.8000 389.8000 33.0000 ;
	    RECT 386.8000 31.6000 389.2000 32.2000 ;
	    RECT 382.0000 30.6000 386.2000 31.2000 ;
	    RECT 378.8000 28.8000 379.6000 30.4000 ;
	    RECT 350.2000 27.8000 361.2000 28.4000 ;
	    RECT 350.6000 27.6000 351.4000 27.8000 ;
	    RECT 343.6000 26.6000 347.6000 27.2000 ;
	    RECT 334.0000 23.0000 334.8000 25.0000 ;
	    RECT 338.2000 23.0000 339.0000 26.0000 ;
	    RECT 329.2000 22.2000 333.2000 22.8000 ;
	    RECT 343.6000 22.2000 344.4000 26.6000 ;
	    RECT 346.6000 26.4000 347.6000 26.6000 ;
	    RECT 346.8000 26.3000 347.6000 26.4000 ;
	    RECT 350.0000 26.3000 350.8000 26.4000 ;
	    RECT 346.8000 25.7000 350.8000 26.3000 ;
	    RECT 350.0000 25.6000 350.8000 25.7000 ;
	    RECT 356.4000 25.6000 357.0000 27.8000 ;
	    RECT 359.6000 27.6000 361.2000 27.8000 ;
	    RECT 362.8000 27.6000 365.4000 28.4000 ;
	    RECT 367.6000 28.2000 368.4000 28.4000 ;
	    RECT 366.8000 27.6000 368.4000 28.2000 ;
	    RECT 369.2000 28.2000 370.0000 28.4000 ;
	    RECT 369.2000 27.6000 370.8000 28.2000 ;
	    RECT 372.2000 27.6000 374.8000 28.4000 ;
	    RECT 375.6000 27.6000 378.2000 28.4000 ;
	    RECT 380.4000 28.2000 381.2000 28.4000 ;
	    RECT 379.6000 27.6000 381.2000 28.2000 ;
	    RECT 354.6000 25.4000 355.4000 25.6000 ;
	    RECT 348.4000 24.2000 349.2000 25.0000 ;
	    RECT 352.6000 24.8000 355.4000 25.4000 ;
	    RECT 356.4000 24.8000 357.2000 25.6000 ;
	    RECT 352.6000 24.2000 353.2000 24.8000 ;
	    RECT 358.0000 24.2000 358.8000 25.0000 ;
	    RECT 347.8000 23.6000 349.2000 24.2000 ;
	    RECT 347.8000 22.2000 349.0000 23.6000 ;
	    RECT 352.4000 22.2000 353.2000 24.2000 ;
	    RECT 356.8000 23.6000 358.8000 24.2000 ;
	    RECT 356.8000 22.2000 357.6000 23.6000 ;
	    RECT 361.2000 22.2000 362.0000 27.0000 ;
	    RECT 363.0000 26.2000 363.6000 27.6000 ;
	    RECT 366.8000 27.2000 367.6000 27.6000 ;
	    RECT 370.0000 27.2000 370.8000 27.6000 ;
	    RECT 364.6000 26.2000 368.2000 26.6000 ;
	    RECT 369.4000 26.2000 373.0000 26.6000 ;
	    RECT 374.0000 26.2000 374.6000 27.6000 ;
	    RECT 375.8000 26.2000 376.4000 27.6000 ;
	    RECT 379.6000 27.2000 380.4000 27.6000 ;
	    RECT 382.0000 27.2000 382.8000 30.6000 ;
	    RECT 385.4000 30.4000 386.2000 30.6000 ;
	    RECT 383.8000 29.8000 384.6000 30.0000 ;
	    RECT 383.8000 29.2000 387.6000 29.8000 ;
	    RECT 386.8000 29.0000 387.6000 29.2000 ;
	    RECT 388.6000 28.4000 389.2000 31.6000 ;
	    RECT 390.6000 31.8000 391.2000 33.0000 ;
	    RECT 391.8000 33.0000 392.6000 33.2000 ;
	    RECT 396.4000 33.0000 397.2000 33.2000 ;
	    RECT 391.8000 32.4000 397.2000 33.0000 ;
	    RECT 390.6000 31.4000 395.4000 31.8000 ;
	    RECT 399.6000 31.4000 400.4000 39.8000 ;
	    RECT 390.6000 31.2000 400.4000 31.4000 ;
	    RECT 394.6000 31.0000 400.4000 31.2000 ;
	    RECT 394.8000 30.8000 400.4000 31.0000 ;
	    RECT 393.2000 30.2000 394.0000 30.4000 ;
	    RECT 402.8000 30.3000 403.6000 39.8000 ;
	    RECT 413.2000 33.6000 414.0000 34.4000 ;
	    RECT 404.4000 31.6000 405.2000 33.2000 ;
	    RECT 413.2000 32.4000 413.8000 33.6000 ;
	    RECT 414.6000 32.4000 415.4000 39.8000 ;
	    RECT 412.4000 31.8000 413.8000 32.4000 ;
	    RECT 414.4000 31.8000 415.4000 32.4000 ;
	    RECT 412.4000 31.6000 413.2000 31.8000 ;
	    RECT 412.5000 30.3000 413.1000 31.6000 ;
	    RECT 414.4000 30.4000 415.0000 31.8000 ;
	    RECT 418.8000 31.2000 419.6000 39.8000 ;
	    RECT 423.0000 35.8000 424.2000 39.8000 ;
	    RECT 427.6000 35.8000 428.4000 39.8000 ;
	    RECT 432.0000 36.4000 432.8000 39.8000 ;
	    RECT 432.0000 35.8000 434.0000 36.4000 ;
	    RECT 423.6000 35.0000 424.4000 35.8000 ;
	    RECT 427.8000 35.2000 428.4000 35.8000 ;
	    RECT 427.0000 34.6000 430.6000 35.2000 ;
	    RECT 433.2000 35.0000 434.0000 35.8000 ;
	    RECT 427.0000 34.4000 427.8000 34.6000 ;
	    RECT 429.8000 34.4000 430.6000 34.6000 ;
	    RECT 422.8000 33.2000 424.2000 34.0000 ;
	    RECT 423.6000 32.2000 424.2000 33.2000 ;
	    RECT 425.8000 33.0000 428.0000 33.6000 ;
	    RECT 425.8000 32.8000 426.6000 33.0000 ;
	    RECT 423.6000 31.6000 426.0000 32.2000 ;
	    RECT 418.8000 30.6000 423.0000 31.2000 ;
	    RECT 393.2000 29.6000 398.2000 30.2000 ;
	    RECT 394.8000 29.4000 395.6000 29.6000 ;
	    RECT 397.4000 29.4000 398.2000 29.6000 ;
	    RECT 402.8000 29.7000 413.1000 30.3000 ;
	    RECT 395.8000 28.4000 396.6000 28.6000 ;
	    RECT 388.6000 27.8000 399.6000 28.4000 ;
	    RECT 389.0000 27.6000 389.8000 27.8000 ;
	    RECT 382.0000 26.6000 385.8000 27.2000 ;
	    RECT 377.4000 26.2000 381.0000 26.6000 ;
	    RECT 362.8000 22.2000 363.6000 26.2000 ;
	    RECT 364.4000 26.0000 368.4000 26.2000 ;
	    RECT 364.4000 22.2000 365.2000 26.0000 ;
	    RECT 367.6000 22.2000 368.4000 26.0000 ;
	    RECT 369.2000 26.0000 373.2000 26.2000 ;
	    RECT 369.2000 22.2000 370.0000 26.0000 ;
	    RECT 372.4000 22.2000 373.2000 26.0000 ;
	    RECT 374.0000 22.2000 374.8000 26.2000 ;
	    RECT 375.6000 22.2000 376.4000 26.2000 ;
	    RECT 377.2000 26.0000 381.2000 26.2000 ;
	    RECT 377.2000 22.2000 378.0000 26.0000 ;
	    RECT 380.4000 22.2000 381.2000 26.0000 ;
	    RECT 382.0000 22.2000 382.8000 26.6000 ;
	    RECT 385.0000 26.4000 385.8000 26.6000 ;
	    RECT 394.8000 25.6000 395.4000 27.8000 ;
	    RECT 398.0000 27.6000 399.6000 27.8000 ;
	    RECT 393.0000 25.4000 393.8000 25.6000 ;
	    RECT 386.8000 24.2000 387.6000 25.0000 ;
	    RECT 391.0000 24.8000 393.8000 25.4000 ;
	    RECT 394.8000 24.8000 395.6000 25.6000 ;
	    RECT 391.0000 24.2000 391.6000 24.8000 ;
	    RECT 396.4000 24.2000 397.2000 25.0000 ;
	    RECT 386.2000 23.6000 387.6000 24.2000 ;
	    RECT 386.2000 22.2000 387.4000 23.6000 ;
	    RECT 390.8000 22.2000 391.6000 24.2000 ;
	    RECT 395.2000 23.6000 397.2000 24.2000 ;
	    RECT 395.2000 22.2000 396.0000 23.6000 ;
	    RECT 399.6000 22.2000 400.4000 27.0000 ;
	    RECT 401.2000 26.8000 402.0000 28.4000 ;
	    RECT 402.8000 26.2000 403.6000 29.7000 ;
	    RECT 414.0000 29.6000 415.0000 30.4000 ;
	    RECT 414.4000 28.4000 415.0000 29.6000 ;
	    RECT 415.6000 28.8000 416.4000 30.4000 ;
	    RECT 412.4000 27.6000 415.0000 28.4000 ;
	    RECT 417.2000 28.2000 418.0000 28.4000 ;
	    RECT 416.4000 27.6000 418.0000 28.2000 ;
	    RECT 412.6000 26.2000 413.2000 27.6000 ;
	    RECT 416.4000 27.2000 417.2000 27.6000 ;
	    RECT 418.8000 27.2000 419.6000 30.6000 ;
	    RECT 422.2000 30.4000 423.0000 30.6000 ;
	    RECT 425.4000 30.4000 426.0000 31.6000 ;
	    RECT 427.4000 31.8000 428.0000 33.0000 ;
	    RECT 428.6000 33.0000 429.4000 33.2000 ;
	    RECT 433.2000 33.0000 434.0000 33.2000 ;
	    RECT 428.6000 32.4000 434.0000 33.0000 ;
	    RECT 427.4000 31.4000 432.2000 31.8000 ;
	    RECT 436.4000 31.4000 437.2000 39.8000 ;
	    RECT 427.4000 31.2000 437.2000 31.4000 ;
	    RECT 431.4000 31.0000 437.2000 31.2000 ;
	    RECT 431.6000 30.8000 437.2000 31.0000 ;
	    RECT 438.0000 31.2000 438.8000 39.8000 ;
	    RECT 442.2000 35.8000 443.4000 39.8000 ;
	    RECT 446.8000 35.8000 447.6000 39.8000 ;
	    RECT 451.2000 36.4000 452.0000 39.8000 ;
	    RECT 451.2000 35.8000 453.2000 36.4000 ;
	    RECT 442.8000 35.0000 443.6000 35.8000 ;
	    RECT 447.0000 35.2000 447.6000 35.8000 ;
	    RECT 446.2000 34.6000 449.8000 35.2000 ;
	    RECT 452.4000 35.0000 453.2000 35.8000 ;
	    RECT 446.2000 34.4000 447.0000 34.6000 ;
	    RECT 449.0000 34.4000 449.8000 34.6000 ;
	    RECT 442.0000 33.2000 443.4000 34.0000 ;
	    RECT 442.8000 32.2000 443.4000 33.2000 ;
	    RECT 445.0000 33.0000 447.2000 33.6000 ;
	    RECT 445.0000 32.8000 445.8000 33.0000 ;
	    RECT 442.8000 31.6000 445.2000 32.2000 ;
	    RECT 438.0000 30.6000 442.2000 31.2000 ;
	    RECT 420.6000 29.8000 421.4000 30.0000 ;
	    RECT 420.6000 29.2000 424.4000 29.8000 ;
	    RECT 425.2000 29.6000 426.0000 30.4000 ;
	    RECT 426.8000 30.3000 427.6000 30.4000 ;
	    RECT 430.0000 30.3000 430.8000 30.4000 ;
	    RECT 426.8000 30.2000 430.8000 30.3000 ;
	    RECT 426.8000 29.7000 435.0000 30.2000 ;
	    RECT 426.8000 29.6000 427.6000 29.7000 ;
	    RECT 430.0000 29.6000 435.0000 29.7000 ;
	    RECT 423.6000 29.0000 424.4000 29.2000 ;
	    RECT 425.4000 28.4000 426.0000 29.6000 ;
	    RECT 434.2000 29.4000 435.0000 29.6000 ;
	    RECT 432.6000 28.4000 433.4000 28.6000 ;
	    RECT 425.4000 27.8000 436.4000 28.4000 ;
	    RECT 425.8000 27.6000 426.6000 27.8000 ;
	    RECT 418.8000 26.6000 422.6000 27.2000 ;
	    RECT 414.2000 26.2000 417.8000 26.6000 ;
	    RECT 402.8000 25.6000 404.6000 26.2000 ;
	    RECT 403.8000 22.2000 404.6000 25.6000 ;
	    RECT 412.4000 22.2000 413.2000 26.2000 ;
	    RECT 414.0000 26.0000 418.0000 26.2000 ;
	    RECT 414.0000 22.2000 414.8000 26.0000 ;
	    RECT 417.2000 22.2000 418.0000 26.0000 ;
	    RECT 418.8000 22.2000 419.6000 26.6000 ;
	    RECT 421.8000 26.4000 422.6000 26.6000 ;
	    RECT 431.6000 25.6000 432.2000 27.8000 ;
	    RECT 434.8000 27.6000 436.4000 27.8000 ;
	    RECT 438.0000 27.2000 438.8000 30.6000 ;
	    RECT 441.4000 30.4000 442.2000 30.6000 ;
	    RECT 439.8000 29.8000 440.6000 30.0000 ;
	    RECT 439.8000 29.2000 443.6000 29.8000 ;
	    RECT 442.8000 29.0000 443.6000 29.2000 ;
	    RECT 444.6000 28.4000 445.2000 31.6000 ;
	    RECT 446.6000 31.8000 447.2000 33.0000 ;
	    RECT 447.8000 33.0000 448.6000 33.2000 ;
	    RECT 452.4000 33.0000 453.2000 33.2000 ;
	    RECT 447.8000 32.4000 453.2000 33.0000 ;
	    RECT 446.6000 31.4000 451.4000 31.8000 ;
	    RECT 455.6000 31.4000 456.4000 39.8000 ;
	    RECT 457.2000 31.6000 458.0000 33.2000 ;
	    RECT 446.6000 31.2000 456.4000 31.4000 ;
	    RECT 450.6000 31.0000 456.4000 31.2000 ;
	    RECT 450.8000 30.8000 456.4000 31.0000 ;
	    RECT 449.2000 30.2000 450.0000 30.4000 ;
	    RECT 449.2000 29.6000 454.2000 30.2000 ;
	    RECT 453.4000 29.4000 454.2000 29.6000 ;
	    RECT 451.8000 28.4000 452.6000 28.6000 ;
	    RECT 444.6000 27.8000 455.6000 28.4000 ;
	    RECT 445.0000 27.6000 445.8000 27.8000 ;
	    RECT 450.8000 27.6000 451.6000 27.8000 ;
	    RECT 454.0000 27.6000 455.6000 27.8000 ;
	    RECT 429.8000 25.4000 430.6000 25.6000 ;
	    RECT 423.6000 24.2000 424.4000 25.0000 ;
	    RECT 427.8000 24.8000 430.6000 25.4000 ;
	    RECT 431.6000 24.8000 432.4000 25.6000 ;
	    RECT 427.8000 24.2000 428.4000 24.8000 ;
	    RECT 433.2000 24.2000 434.0000 25.0000 ;
	    RECT 423.0000 23.6000 424.4000 24.2000 ;
	    RECT 423.0000 22.2000 424.2000 23.6000 ;
	    RECT 427.6000 22.2000 428.4000 24.2000 ;
	    RECT 432.0000 23.6000 434.0000 24.2000 ;
	    RECT 432.0000 22.2000 432.8000 23.6000 ;
	    RECT 436.4000 22.2000 437.2000 27.0000 ;
	    RECT 438.0000 26.6000 441.8000 27.2000 ;
	    RECT 438.0000 22.2000 438.8000 26.6000 ;
	    RECT 441.0000 26.4000 441.8000 26.6000 ;
	    RECT 450.8000 25.6000 451.4000 27.6000 ;
	    RECT 449.0000 25.4000 449.8000 25.6000 ;
	    RECT 442.8000 24.2000 443.6000 25.0000 ;
	    RECT 447.0000 24.8000 449.8000 25.4000 ;
	    RECT 450.8000 24.8000 451.6000 25.6000 ;
	    RECT 447.0000 24.2000 447.6000 24.8000 ;
	    RECT 452.4000 24.2000 453.2000 25.0000 ;
	    RECT 442.2000 23.6000 443.6000 24.2000 ;
	    RECT 442.2000 22.2000 443.4000 23.6000 ;
	    RECT 446.8000 22.2000 447.6000 24.2000 ;
	    RECT 451.2000 23.6000 453.2000 24.2000 ;
	    RECT 451.2000 22.2000 452.0000 23.6000 ;
	    RECT 455.6000 22.2000 456.4000 27.0000 ;
	    RECT 458.8000 26.2000 459.6000 39.8000 ;
	    RECT 460.4000 26.8000 461.2000 28.4000 ;
	    RECT 463.6000 28.3000 464.4000 39.8000 ;
	    RECT 467.8000 32.4000 468.6000 39.8000 ;
	    RECT 469.2000 33.6000 470.0000 34.4000 ;
	    RECT 469.4000 32.4000 470.0000 33.6000 ;
	    RECT 466.8000 31.6000 468.8000 32.4000 ;
	    RECT 469.4000 31.8000 470.8000 32.4000 ;
	    RECT 470.0000 31.6000 470.8000 31.8000 ;
	    RECT 466.8000 28.8000 467.6000 30.4000 ;
	    RECT 468.2000 28.4000 468.8000 31.6000 ;
	    RECT 465.2000 28.3000 466.0000 28.4000 ;
	    RECT 463.6000 28.2000 466.0000 28.3000 ;
	    RECT 463.6000 27.7000 466.8000 28.2000 ;
	    RECT 457.8000 25.6000 459.6000 26.2000 ;
	    RECT 457.8000 24.4000 458.6000 25.6000 ;
	    RECT 462.0000 24.8000 462.8000 26.4000 ;
	    RECT 457.8000 23.6000 459.6000 24.4000 ;
	    RECT 457.8000 22.2000 458.6000 23.6000 ;
	    RECT 463.6000 22.2000 464.4000 27.7000 ;
	    RECT 465.2000 27.6000 466.8000 27.7000 ;
	    RECT 468.2000 27.6000 470.8000 28.4000 ;
	    RECT 473.2000 28.3000 474.0000 39.8000 ;
	    RECT 477.4000 32.4000 478.2000 39.8000 ;
	    RECT 478.8000 33.6000 479.6000 34.4000 ;
	    RECT 479.0000 32.4000 479.6000 33.6000 ;
	    RECT 477.4000 31.8000 478.4000 32.4000 ;
	    RECT 479.0000 31.8000 480.4000 32.4000 ;
	    RECT 476.4000 28.8000 477.2000 30.4000 ;
	    RECT 477.8000 28.4000 478.4000 31.8000 ;
	    RECT 479.6000 31.6000 480.4000 31.8000 ;
	    RECT 474.8000 28.3000 475.6000 28.4000 ;
	    RECT 473.2000 28.2000 475.6000 28.3000 ;
	    RECT 473.2000 27.7000 476.4000 28.2000 ;
	    RECT 466.0000 27.2000 466.8000 27.6000 ;
	    RECT 465.4000 26.2000 469.0000 26.6000 ;
	    RECT 470.0000 26.2000 470.6000 27.6000 ;
	    RECT 465.2000 26.0000 469.2000 26.2000 ;
	    RECT 465.2000 22.2000 466.0000 26.0000 ;
	    RECT 468.4000 22.2000 469.2000 26.0000 ;
	    RECT 470.0000 22.2000 470.8000 26.2000 ;
	    RECT 471.6000 24.8000 472.4000 26.4000 ;
	    RECT 473.2000 22.2000 474.0000 27.7000 ;
	    RECT 474.8000 27.6000 476.4000 27.7000 ;
	    RECT 477.8000 27.6000 480.4000 28.4000 ;
	    RECT 482.8000 28.3000 483.6000 39.8000 ;
	    RECT 487.0000 32.4000 487.8000 39.8000 ;
	    RECT 488.4000 33.6000 489.2000 34.4000 ;
	    RECT 488.6000 32.4000 489.2000 33.6000 ;
	    RECT 487.0000 31.8000 488.0000 32.4000 ;
	    RECT 488.6000 31.8000 490.0000 32.4000 ;
	    RECT 486.0000 28.8000 486.8000 30.4000 ;
	    RECT 487.4000 30.3000 488.0000 31.8000 ;
	    RECT 489.2000 31.6000 490.0000 31.8000 ;
	    RECT 490.8000 31.2000 491.6000 39.8000 ;
	    RECT 495.0000 35.8000 496.2000 39.8000 ;
	    RECT 499.6000 35.8000 500.4000 39.8000 ;
	    RECT 504.0000 36.4000 504.8000 39.8000 ;
	    RECT 504.0000 35.8000 506.0000 36.4000 ;
	    RECT 495.6000 35.0000 496.4000 35.8000 ;
	    RECT 499.8000 35.2000 500.4000 35.8000 ;
	    RECT 499.0000 34.6000 502.6000 35.2000 ;
	    RECT 505.2000 35.0000 506.0000 35.8000 ;
	    RECT 499.0000 34.4000 499.8000 34.6000 ;
	    RECT 501.8000 34.4000 502.6000 34.6000 ;
	    RECT 494.8000 33.2000 496.2000 34.0000 ;
	    RECT 495.6000 32.2000 496.2000 33.2000 ;
	    RECT 497.8000 33.0000 500.0000 33.6000 ;
	    RECT 497.8000 32.8000 498.6000 33.0000 ;
	    RECT 495.6000 31.6000 498.0000 32.2000 ;
	    RECT 490.8000 30.6000 495.0000 31.2000 ;
	    RECT 489.2000 30.3000 490.0000 30.4000 ;
	    RECT 487.4000 29.7000 490.0000 30.3000 ;
	    RECT 487.4000 28.4000 488.0000 29.7000 ;
	    RECT 489.2000 29.6000 490.0000 29.7000 ;
	    RECT 484.4000 28.3000 485.2000 28.4000 ;
	    RECT 482.8000 28.2000 485.2000 28.3000 ;
	    RECT 482.8000 27.7000 486.0000 28.2000 ;
	    RECT 475.6000 27.2000 476.4000 27.6000 ;
	    RECT 475.0000 26.2000 478.6000 26.6000 ;
	    RECT 479.6000 26.2000 480.2000 27.6000 ;
	    RECT 474.8000 26.0000 478.8000 26.2000 ;
	    RECT 474.8000 22.2000 475.6000 26.0000 ;
	    RECT 478.0000 22.2000 478.8000 26.0000 ;
	    RECT 479.6000 22.2000 480.4000 26.2000 ;
	    RECT 481.2000 24.8000 482.0000 26.4000 ;
	    RECT 482.8000 22.2000 483.6000 27.7000 ;
	    RECT 484.4000 27.6000 486.0000 27.7000 ;
	    RECT 487.4000 27.6000 490.0000 28.4000 ;
	    RECT 485.2000 27.2000 486.0000 27.6000 ;
	    RECT 484.6000 26.2000 488.2000 26.6000 ;
	    RECT 489.2000 26.2000 489.8000 27.6000 ;
	    RECT 490.8000 27.2000 491.6000 30.6000 ;
	    RECT 494.2000 30.4000 495.0000 30.6000 ;
	    RECT 492.6000 29.8000 493.4000 30.0000 ;
	    RECT 492.6000 29.2000 496.4000 29.8000 ;
	    RECT 495.6000 29.0000 496.4000 29.2000 ;
	    RECT 497.4000 28.4000 498.0000 31.6000 ;
	    RECT 499.4000 31.8000 500.0000 33.0000 ;
	    RECT 500.6000 33.0000 501.4000 33.2000 ;
	    RECT 505.2000 33.0000 506.0000 33.2000 ;
	    RECT 500.6000 32.4000 506.0000 33.0000 ;
	    RECT 499.4000 31.4000 504.2000 31.8000 ;
	    RECT 508.4000 31.4000 509.2000 39.8000 ;
	    RECT 499.4000 31.2000 509.2000 31.4000 ;
	    RECT 503.4000 31.0000 509.2000 31.2000 ;
	    RECT 503.6000 30.8000 509.2000 31.0000 ;
	    RECT 500.4000 30.3000 501.2000 30.4000 ;
	    RECT 502.0000 30.3000 502.8000 30.4000 ;
	    RECT 500.4000 30.2000 502.8000 30.3000 ;
	    RECT 500.4000 29.7000 507.0000 30.2000 ;
	    RECT 500.4000 29.6000 501.2000 29.7000 ;
	    RECT 502.0000 29.6000 507.0000 29.7000 ;
	    RECT 506.2000 29.4000 507.0000 29.6000 ;
	    RECT 504.6000 28.4000 505.4000 28.6000 ;
	    RECT 497.2000 27.8000 508.4000 28.4000 ;
	    RECT 497.2000 27.6000 498.6000 27.8000 ;
	    RECT 502.0000 27.6000 502.8000 27.8000 ;
	    RECT 490.8000 26.6000 494.6000 27.2000 ;
	    RECT 484.4000 26.0000 488.4000 26.2000 ;
	    RECT 484.4000 22.2000 485.2000 26.0000 ;
	    RECT 487.6000 22.2000 488.4000 26.0000 ;
	    RECT 489.2000 22.2000 490.0000 26.2000 ;
	    RECT 490.8000 22.2000 491.6000 26.6000 ;
	    RECT 493.8000 26.4000 494.6000 26.6000 ;
	    RECT 503.6000 25.6000 504.2000 27.8000 ;
	    RECT 506.8000 27.6000 508.4000 27.8000 ;
	    RECT 501.8000 25.4000 502.6000 25.6000 ;
	    RECT 495.6000 24.2000 496.4000 25.0000 ;
	    RECT 499.8000 24.8000 502.6000 25.4000 ;
	    RECT 503.6000 24.8000 504.4000 25.6000 ;
	    RECT 499.8000 24.2000 500.4000 24.8000 ;
	    RECT 505.2000 24.2000 506.0000 25.0000 ;
	    RECT 495.0000 23.6000 496.4000 24.2000 ;
	    RECT 495.0000 22.2000 496.2000 23.6000 ;
	    RECT 499.6000 22.2000 500.4000 24.2000 ;
	    RECT 504.0000 23.6000 506.0000 24.2000 ;
	    RECT 504.0000 22.2000 504.8000 23.6000 ;
	    RECT 508.4000 22.2000 509.2000 27.0000 ;
	    RECT 4.4000 15.2000 5.2000 19.8000 ;
	    RECT 9.2000 15.2000 10.0000 19.8000 ;
	    RECT 3.0000 14.6000 5.2000 15.2000 ;
	    RECT 7.8000 14.6000 10.0000 15.2000 ;
	    RECT 10.8000 15.4000 11.6000 19.8000 ;
	    RECT 15.0000 18.4000 16.2000 19.8000 ;
	    RECT 15.0000 17.8000 16.4000 18.4000 ;
	    RECT 19.6000 17.8000 20.4000 19.8000 ;
	    RECT 24.0000 18.4000 24.8000 19.8000 ;
	    RECT 24.0000 17.8000 26.0000 18.4000 ;
	    RECT 15.6000 17.0000 16.4000 17.8000 ;
	    RECT 19.8000 17.2000 20.4000 17.8000 ;
	    RECT 19.8000 16.6000 22.6000 17.2000 ;
	    RECT 21.8000 16.4000 22.6000 16.6000 ;
	    RECT 23.6000 16.4000 24.4000 17.2000 ;
	    RECT 25.2000 17.0000 26.0000 17.8000 ;
	    RECT 13.8000 15.4000 14.6000 15.6000 ;
	    RECT 10.8000 14.8000 14.6000 15.4000 ;
	    RECT 3.0000 11.6000 3.6000 14.6000 ;
	    RECT 4.4000 11.6000 5.2000 13.2000 ;
	    RECT 7.8000 11.6000 8.4000 14.6000 ;
	    RECT 9.2000 11.6000 10.0000 13.2000 ;
	    RECT 2.4000 10.8000 3.6000 11.6000 ;
	    RECT 7.2000 10.8000 8.4000 11.6000 ;
	    RECT 3.0000 10.2000 3.6000 10.8000 ;
	    RECT 7.8000 10.2000 8.4000 10.8000 ;
	    RECT 10.8000 11.4000 11.6000 14.8000 ;
	    RECT 17.8000 14.2000 18.6000 14.4000 ;
	    RECT 22.0000 14.2000 22.8000 14.4000 ;
	    RECT 23.6000 14.2000 24.2000 16.4000 ;
	    RECT 28.4000 15.0000 29.2000 19.8000 ;
	    RECT 30.0000 15.8000 30.8000 19.8000 ;
	    RECT 31.6000 16.0000 32.4000 19.8000 ;
	    RECT 34.8000 16.0000 35.6000 19.8000 ;
	    RECT 31.6000 15.8000 35.6000 16.0000 ;
	    RECT 30.2000 14.4000 30.8000 15.8000 ;
	    RECT 31.8000 15.4000 35.4000 15.8000 ;
	    RECT 39.6000 15.2000 40.4000 19.8000 ;
	    RECT 41.2000 15.8000 42.0000 19.8000 ;
	    RECT 42.8000 16.0000 43.6000 19.8000 ;
	    RECT 46.0000 16.0000 46.8000 19.8000 ;
	    RECT 42.8000 15.8000 46.8000 16.0000 ;
	    RECT 34.0000 14.4000 34.8000 14.8000 ;
	    RECT 38.2000 14.6000 40.4000 15.2000 ;
	    RECT 26.8000 14.2000 28.4000 14.4000 ;
	    RECT 17.4000 13.6000 28.4000 14.2000 ;
	    RECT 30.0000 13.6000 32.6000 14.4000 ;
	    RECT 34.0000 13.8000 35.6000 14.4000 ;
	    RECT 34.8000 13.6000 35.6000 13.8000 ;
	    RECT 15.6000 12.8000 16.4000 13.0000 ;
	    RECT 12.6000 12.2000 16.4000 12.8000 ;
	    RECT 17.4000 12.4000 18.0000 13.6000 ;
	    RECT 24.6000 13.4000 25.4000 13.6000 ;
	    RECT 23.6000 12.4000 24.4000 12.6000 ;
	    RECT 26.2000 12.4000 27.0000 12.6000 ;
	    RECT 12.6000 12.0000 13.4000 12.2000 ;
	    RECT 17.2000 11.6000 18.0000 12.4000 ;
	    RECT 22.0000 11.8000 27.0000 12.4000 ;
	    RECT 22.0000 11.6000 22.8000 11.8000 ;
	    RECT 14.2000 11.4000 15.0000 11.6000 ;
	    RECT 10.8000 10.8000 15.0000 11.4000 ;
	    RECT 3.0000 9.6000 5.2000 10.2000 ;
	    RECT 7.8000 9.6000 10.0000 10.2000 ;
	    RECT 4.4000 2.2000 5.2000 9.6000 ;
	    RECT 9.2000 2.2000 10.0000 9.6000 ;
	    RECT 10.8000 2.2000 11.6000 10.8000 ;
	    RECT 17.4000 10.4000 18.0000 11.6000 ;
	    RECT 23.6000 11.0000 29.2000 11.2000 ;
	    RECT 23.4000 10.8000 29.2000 11.0000 ;
	    RECT 15.6000 9.8000 18.0000 10.4000 ;
	    RECT 19.4000 10.6000 29.2000 10.8000 ;
	    RECT 19.4000 10.2000 24.2000 10.6000 ;
	    RECT 15.6000 8.8000 16.2000 9.8000 ;
	    RECT 14.8000 8.0000 16.2000 8.8000 ;
	    RECT 17.8000 9.0000 18.6000 9.2000 ;
	    RECT 19.4000 9.0000 20.0000 10.2000 ;
	    RECT 17.8000 8.4000 20.0000 9.0000 ;
	    RECT 20.6000 9.0000 26.0000 9.6000 ;
	    RECT 20.6000 8.8000 21.4000 9.0000 ;
	    RECT 25.2000 8.8000 26.0000 9.0000 ;
	    RECT 19.0000 7.4000 19.8000 7.6000 ;
	    RECT 21.8000 7.4000 22.6000 7.6000 ;
	    RECT 15.6000 6.2000 16.4000 7.0000 ;
	    RECT 19.0000 6.8000 22.6000 7.4000 ;
	    RECT 19.8000 6.2000 20.4000 6.8000 ;
	    RECT 25.2000 6.2000 26.0000 7.0000 ;
	    RECT 15.0000 2.2000 16.2000 6.2000 ;
	    RECT 19.6000 2.2000 20.4000 6.2000 ;
	    RECT 24.0000 5.6000 26.0000 6.2000 ;
	    RECT 24.0000 2.2000 24.8000 5.6000 ;
	    RECT 28.4000 2.2000 29.2000 10.6000 ;
	    RECT 32.0000 10.4000 32.6000 13.6000 ;
	    RECT 33.2000 11.6000 34.0000 13.2000 ;
	    RECT 38.2000 11.6000 38.8000 14.6000 ;
	    RECT 41.4000 14.4000 42.0000 15.8000 ;
	    RECT 43.0000 15.4000 46.6000 15.8000 ;
	    RECT 50.8000 15.2000 51.6000 19.8000 ;
	    RECT 45.2000 14.4000 46.0000 14.8000 ;
	    RECT 49.4000 14.6000 51.6000 15.2000 ;
	    RECT 52.4000 15.4000 53.2000 19.8000 ;
	    RECT 56.6000 18.4000 57.8000 19.8000 ;
	    RECT 56.6000 17.8000 58.0000 18.4000 ;
	    RECT 61.2000 17.8000 62.0000 19.8000 ;
	    RECT 65.6000 18.4000 66.4000 19.8000 ;
	    RECT 65.6000 17.8000 67.6000 18.4000 ;
	    RECT 57.2000 17.0000 58.0000 17.8000 ;
	    RECT 61.4000 17.2000 62.0000 17.8000 ;
	    RECT 61.4000 16.6000 64.2000 17.2000 ;
	    RECT 63.4000 16.4000 64.2000 16.6000 ;
	    RECT 65.2000 16.4000 66.0000 17.2000 ;
	    RECT 66.8000 17.0000 67.6000 17.8000 ;
	    RECT 55.6000 15.6000 56.4000 16.4000 ;
	    RECT 55.4000 15.4000 56.4000 15.6000 ;
	    RECT 52.4000 14.8000 56.4000 15.4000 ;
	    RECT 41.2000 13.6000 43.8000 14.4000 ;
	    RECT 45.2000 13.8000 46.8000 14.4000 ;
	    RECT 46.0000 13.6000 46.8000 13.8000 ;
	    RECT 39.6000 11.6000 40.4000 13.2000 ;
	    RECT 41.2000 12.3000 42.0000 12.4000 ;
	    RECT 43.2000 12.3000 43.8000 13.6000 ;
	    RECT 41.2000 11.7000 43.8000 12.3000 ;
	    RECT 41.2000 11.6000 42.0000 11.7000 ;
	    RECT 37.6000 10.8000 38.8000 11.6000 ;
	    RECT 30.0000 10.2000 30.8000 10.4000 ;
	    RECT 30.0000 9.6000 31.4000 10.2000 ;
	    RECT 32.0000 9.6000 34.0000 10.4000 ;
	    RECT 38.2000 10.2000 38.8000 10.8000 ;
	    RECT 41.2000 10.2000 42.0000 10.4000 ;
	    RECT 43.2000 10.2000 43.8000 11.7000 ;
	    RECT 44.4000 11.6000 45.2000 13.2000 ;
	    RECT 49.4000 11.6000 50.0000 14.6000 ;
	    RECT 50.8000 11.6000 51.6000 13.2000 ;
	    RECT 48.8000 10.8000 50.0000 11.6000 ;
	    RECT 49.4000 10.2000 50.0000 10.8000 ;
	    RECT 52.4000 11.4000 53.2000 14.8000 ;
	    RECT 59.4000 14.2000 60.2000 14.4000 ;
	    RECT 65.2000 14.2000 65.8000 16.4000 ;
	    RECT 70.0000 15.0000 70.8000 19.8000 ;
	    RECT 71.6000 16.0000 72.4000 19.8000 ;
	    RECT 74.8000 16.0000 75.6000 19.8000 ;
	    RECT 71.6000 15.8000 75.6000 16.0000 ;
	    RECT 76.4000 15.8000 77.2000 19.8000 ;
	    RECT 71.8000 15.4000 75.4000 15.8000 ;
	    RECT 72.4000 14.4000 73.2000 14.8000 ;
	    RECT 76.4000 14.4000 77.0000 15.8000 ;
	    RECT 81.2000 15.2000 82.0000 19.8000 ;
	    RECT 79.8000 14.6000 82.0000 15.2000 ;
	    RECT 82.8000 15.0000 83.6000 19.8000 ;
	    RECT 87.2000 18.4000 88.0000 19.8000 ;
	    RECT 86.0000 17.8000 88.0000 18.4000 ;
	    RECT 91.6000 17.8000 92.4000 19.8000 ;
	    RECT 95.8000 18.4000 97.0000 19.8000 ;
	    RECT 95.6000 17.8000 97.0000 18.4000 ;
	    RECT 86.0000 17.0000 86.8000 17.8000 ;
	    RECT 91.6000 17.2000 92.2000 17.8000 ;
	    RECT 87.6000 16.4000 88.4000 17.2000 ;
	    RECT 89.4000 16.6000 92.2000 17.2000 ;
	    RECT 95.6000 17.0000 96.4000 17.8000 ;
	    RECT 89.4000 16.4000 90.2000 16.6000 ;
	    RECT 68.4000 14.2000 70.0000 14.4000 ;
	    RECT 59.0000 13.6000 70.0000 14.2000 ;
	    RECT 71.6000 13.8000 73.2000 14.4000 ;
	    RECT 71.6000 13.6000 72.4000 13.8000 ;
	    RECT 74.6000 13.6000 77.2000 14.4000 ;
	    RECT 57.2000 12.8000 58.0000 13.0000 ;
	    RECT 54.2000 12.2000 58.0000 12.8000 ;
	    RECT 59.0000 12.4000 59.6000 13.6000 ;
	    RECT 66.2000 13.4000 67.0000 13.6000 ;
	    RECT 67.8000 12.4000 68.6000 12.6000 ;
	    RECT 54.2000 12.0000 55.0000 12.2000 ;
	    RECT 58.8000 11.6000 59.6000 12.4000 ;
	    RECT 60.4000 12.3000 61.2000 12.4000 ;
	    RECT 63.6000 12.3000 68.6000 12.4000 ;
	    RECT 60.4000 11.8000 68.6000 12.3000 ;
	    RECT 60.4000 11.7000 64.4000 11.8000 ;
	    RECT 60.4000 11.6000 61.2000 11.7000 ;
	    RECT 63.6000 11.6000 64.4000 11.7000 ;
	    RECT 73.2000 11.6000 74.0000 13.2000 ;
	    RECT 74.6000 12.3000 75.2000 13.6000 ;
	    RECT 76.4000 12.3000 77.2000 12.4000 ;
	    RECT 74.6000 11.7000 77.2000 12.3000 ;
	    RECT 55.8000 11.4000 56.6000 11.6000 ;
	    RECT 52.4000 10.8000 56.6000 11.4000 ;
	    RECT 38.2000 9.6000 40.4000 10.2000 ;
	    RECT 41.2000 9.6000 42.6000 10.2000 ;
	    RECT 43.2000 9.6000 44.2000 10.2000 ;
	    RECT 49.4000 9.6000 51.6000 10.2000 ;
	    RECT 30.8000 8.4000 31.4000 9.6000 ;
	    RECT 30.8000 7.6000 31.6000 8.4000 ;
	    RECT 32.2000 2.2000 33.0000 9.6000 ;
	    RECT 39.6000 2.2000 40.4000 9.6000 ;
	    RECT 42.0000 8.4000 42.6000 9.6000 ;
	    RECT 42.0000 7.6000 42.8000 8.4000 ;
	    RECT 43.4000 2.2000 44.2000 9.6000 ;
	    RECT 50.8000 2.2000 51.6000 9.6000 ;
	    RECT 52.4000 2.2000 53.2000 10.8000 ;
	    RECT 59.0000 10.4000 59.6000 11.6000 ;
	    RECT 65.2000 11.0000 70.8000 11.2000 ;
	    RECT 65.0000 10.8000 70.8000 11.0000 ;
	    RECT 57.2000 9.8000 59.6000 10.4000 ;
	    RECT 61.0000 10.6000 70.8000 10.8000 ;
	    RECT 61.0000 10.2000 65.8000 10.6000 ;
	    RECT 57.2000 8.8000 57.8000 9.8000 ;
	    RECT 56.4000 8.0000 57.8000 8.8000 ;
	    RECT 59.4000 9.0000 60.2000 9.2000 ;
	    RECT 61.0000 9.0000 61.6000 10.2000 ;
	    RECT 59.4000 8.4000 61.6000 9.0000 ;
	    RECT 62.2000 9.0000 67.6000 9.6000 ;
	    RECT 62.2000 8.8000 63.0000 9.0000 ;
	    RECT 66.8000 8.8000 67.6000 9.0000 ;
	    RECT 60.6000 7.4000 61.4000 7.6000 ;
	    RECT 63.4000 7.4000 64.2000 7.6000 ;
	    RECT 57.2000 6.2000 58.0000 7.0000 ;
	    RECT 60.6000 6.8000 64.2000 7.4000 ;
	    RECT 61.4000 6.2000 62.0000 6.8000 ;
	    RECT 66.8000 6.2000 67.6000 7.0000 ;
	    RECT 56.6000 2.2000 57.8000 6.2000 ;
	    RECT 61.2000 2.2000 62.0000 6.2000 ;
	    RECT 65.6000 5.6000 67.6000 6.2000 ;
	    RECT 65.6000 2.2000 66.4000 5.6000 ;
	    RECT 70.0000 2.2000 70.8000 10.6000 ;
	    RECT 74.6000 10.2000 75.2000 11.7000 ;
	    RECT 76.4000 11.6000 77.2000 11.7000 ;
	    RECT 79.8000 11.6000 80.4000 14.6000 ;
	    RECT 83.6000 14.2000 85.2000 14.4000 ;
	    RECT 87.8000 14.2000 88.4000 16.4000 ;
	    RECT 97.4000 15.4000 98.2000 15.6000 ;
	    RECT 100.4000 15.4000 101.2000 19.8000 ;
	    RECT 97.4000 14.8000 101.2000 15.4000 ;
	    RECT 93.4000 14.2000 94.2000 14.4000 ;
	    RECT 83.6000 13.6000 94.6000 14.2000 ;
	    RECT 86.6000 13.4000 87.4000 13.6000 ;
	    RECT 81.2000 11.6000 82.0000 13.2000 ;
	    RECT 85.0000 12.4000 85.8000 12.6000 ;
	    RECT 85.0000 12.3000 90.0000 12.4000 ;
	    RECT 92.4000 12.3000 93.2000 12.4000 ;
	    RECT 85.0000 11.8000 93.2000 12.3000 ;
	    RECT 89.2000 11.7000 93.2000 11.8000 ;
	    RECT 89.2000 11.6000 90.0000 11.7000 ;
	    RECT 92.4000 11.6000 93.2000 11.7000 ;
	    RECT 79.2000 10.8000 80.4000 11.6000 ;
	    RECT 76.4000 10.2000 77.2000 10.4000 ;
	    RECT 74.2000 9.6000 75.2000 10.2000 ;
	    RECT 75.8000 9.6000 77.2000 10.2000 ;
	    RECT 79.8000 10.2000 80.4000 10.8000 ;
	    RECT 82.8000 11.0000 88.4000 11.2000 ;
	    RECT 82.8000 10.8000 88.6000 11.0000 ;
	    RECT 82.8000 10.6000 92.6000 10.8000 ;
	    RECT 79.8000 9.6000 82.0000 10.2000 ;
	    RECT 74.2000 2.2000 75.0000 9.6000 ;
	    RECT 75.8000 8.4000 76.4000 9.6000 ;
	    RECT 75.6000 7.6000 76.4000 8.4000 ;
	    RECT 81.2000 2.2000 82.0000 9.6000 ;
	    RECT 82.8000 2.2000 83.6000 10.6000 ;
	    RECT 87.8000 10.2000 92.6000 10.6000 ;
	    RECT 86.0000 9.0000 91.4000 9.6000 ;
	    RECT 86.0000 8.8000 86.8000 9.0000 ;
	    RECT 90.6000 8.8000 91.4000 9.0000 ;
	    RECT 92.0000 9.0000 92.6000 10.2000 ;
	    RECT 94.0000 10.4000 94.6000 13.6000 ;
	    RECT 95.6000 12.8000 96.4000 13.0000 ;
	    RECT 95.6000 12.2000 99.4000 12.8000 ;
	    RECT 98.6000 12.0000 99.4000 12.2000 ;
	    RECT 97.0000 11.4000 97.8000 11.6000 ;
	    RECT 100.4000 11.4000 101.2000 14.8000 ;
	    RECT 102.0000 15.2000 102.8000 19.8000 ;
	    RECT 113.2000 15.8000 114.0000 19.8000 ;
	    RECT 114.8000 16.0000 115.6000 19.8000 ;
	    RECT 118.0000 16.0000 118.8000 19.8000 ;
	    RECT 114.8000 15.8000 118.8000 16.0000 ;
	    RECT 119.6000 15.8000 120.4000 19.8000 ;
	    RECT 121.2000 16.0000 122.0000 19.8000 ;
	    RECT 124.4000 16.0000 125.2000 19.8000 ;
	    RECT 121.2000 15.8000 125.2000 16.0000 ;
	    RECT 126.0000 15.8000 126.8000 19.8000 ;
	    RECT 127.6000 16.0000 128.4000 19.8000 ;
	    RECT 130.8000 16.0000 131.6000 19.8000 ;
	    RECT 127.6000 15.8000 131.6000 16.0000 ;
	    RECT 102.0000 14.6000 104.2000 15.2000 ;
	    RECT 102.0000 11.6000 102.8000 13.2000 ;
	    RECT 103.6000 11.6000 104.2000 14.6000 ;
	    RECT 113.4000 14.4000 114.0000 15.8000 ;
	    RECT 115.0000 15.4000 118.6000 15.8000 ;
	    RECT 117.2000 14.4000 118.0000 14.8000 ;
	    RECT 119.8000 14.4000 120.4000 15.8000 ;
	    RECT 121.4000 15.4000 125.0000 15.8000 ;
	    RECT 123.6000 14.4000 124.4000 14.8000 ;
	    RECT 126.2000 14.4000 126.8000 15.8000 ;
	    RECT 127.8000 15.4000 131.4000 15.8000 ;
	    RECT 135.6000 15.2000 136.4000 19.8000 ;
	    RECT 140.4000 15.2000 141.2000 19.8000 ;
	    RECT 130.0000 14.4000 130.8000 14.8000 ;
	    RECT 134.2000 14.6000 136.4000 15.2000 ;
	    RECT 139.0000 14.6000 141.2000 15.2000 ;
	    RECT 142.0000 15.4000 142.8000 19.8000 ;
	    RECT 146.2000 18.4000 147.4000 19.8000 ;
	    RECT 146.2000 17.8000 147.6000 18.4000 ;
	    RECT 150.8000 17.8000 151.6000 19.8000 ;
	    RECT 155.2000 18.4000 156.0000 19.8000 ;
	    RECT 155.2000 17.8000 157.2000 18.4000 ;
	    RECT 146.8000 17.0000 147.6000 17.8000 ;
	    RECT 151.0000 17.2000 151.6000 17.8000 ;
	    RECT 151.0000 16.6000 153.8000 17.2000 ;
	    RECT 153.0000 16.4000 153.8000 16.6000 ;
	    RECT 154.8000 15.6000 155.6000 17.2000 ;
	    RECT 156.4000 17.0000 157.2000 17.8000 ;
	    RECT 145.0000 15.4000 145.8000 15.6000 ;
	    RECT 142.0000 14.8000 145.8000 15.4000 ;
	    RECT 113.2000 13.6000 115.8000 14.4000 ;
	    RECT 117.2000 13.8000 118.8000 14.4000 ;
	    RECT 118.0000 13.6000 118.8000 13.8000 ;
	    RECT 119.6000 13.6000 122.2000 14.4000 ;
	    RECT 123.6000 13.8000 125.2000 14.4000 ;
	    RECT 124.4000 13.6000 125.2000 13.8000 ;
	    RECT 126.0000 13.6000 128.6000 14.4000 ;
	    RECT 130.0000 13.8000 131.6000 14.4000 ;
	    RECT 130.8000 13.6000 131.6000 13.8000 ;
	    RECT 97.0000 10.8000 101.2000 11.4000 ;
	    RECT 94.0000 9.8000 96.4000 10.4000 ;
	    RECT 93.4000 9.0000 94.2000 9.2000 ;
	    RECT 92.0000 8.4000 94.2000 9.0000 ;
	    RECT 95.8000 8.8000 96.4000 9.8000 ;
	    RECT 95.8000 8.0000 97.2000 8.8000 ;
	    RECT 89.4000 7.4000 90.2000 7.6000 ;
	    RECT 92.2000 7.4000 93.0000 7.6000 ;
	    RECT 86.0000 6.2000 86.8000 7.0000 ;
	    RECT 89.4000 6.8000 93.0000 7.4000 ;
	    RECT 91.6000 6.2000 92.2000 6.8000 ;
	    RECT 95.6000 6.2000 96.4000 7.0000 ;
	    RECT 86.0000 5.6000 88.0000 6.2000 ;
	    RECT 87.2000 2.2000 88.0000 5.6000 ;
	    RECT 91.6000 2.2000 92.4000 6.2000 ;
	    RECT 95.8000 2.2000 97.0000 6.2000 ;
	    RECT 100.4000 2.2000 101.2000 10.8000 ;
	    RECT 103.6000 10.8000 104.8000 11.6000 ;
	    RECT 103.6000 10.2000 104.2000 10.8000 ;
	    RECT 102.0000 9.6000 104.2000 10.2000 ;
	    RECT 113.2000 10.2000 114.0000 10.4000 ;
	    RECT 115.2000 10.2000 115.8000 13.6000 ;
	    RECT 116.4000 12.3000 117.2000 13.2000 ;
	    RECT 121.6000 12.3000 122.2000 13.6000 ;
	    RECT 116.4000 11.7000 122.2000 12.3000 ;
	    RECT 116.4000 11.6000 117.2000 11.7000 ;
	    RECT 119.6000 10.2000 120.4000 10.4000 ;
	    RECT 121.6000 10.2000 122.2000 11.7000 ;
	    RECT 122.8000 12.3000 123.6000 13.2000 ;
	    RECT 124.4000 12.3000 125.2000 12.4000 ;
	    RECT 122.8000 11.7000 125.2000 12.3000 ;
	    RECT 122.8000 11.6000 123.6000 11.7000 ;
	    RECT 124.4000 11.6000 125.2000 11.7000 ;
	    RECT 126.0000 10.2000 126.8000 10.4000 ;
	    RECT 128.0000 10.2000 128.6000 13.6000 ;
	    RECT 129.2000 11.6000 130.0000 13.2000 ;
	    RECT 134.2000 11.6000 134.8000 14.6000 ;
	    RECT 135.6000 11.6000 136.4000 13.2000 ;
	    RECT 139.0000 11.6000 139.6000 14.6000 ;
	    RECT 140.4000 11.6000 141.2000 13.2000 ;
	    RECT 133.6000 10.8000 134.8000 11.6000 ;
	    RECT 138.4000 10.8000 139.6000 11.6000 ;
	    RECT 134.2000 10.2000 134.8000 10.8000 ;
	    RECT 139.0000 10.2000 139.6000 10.8000 ;
	    RECT 142.0000 11.4000 142.8000 14.8000 ;
	    RECT 149.0000 14.2000 149.8000 14.4000 ;
	    RECT 154.8000 14.2000 155.4000 15.6000 ;
	    RECT 159.6000 15.0000 160.4000 19.8000 ;
	    RECT 164.4000 15.2000 165.2000 19.8000 ;
	    RECT 163.0000 14.6000 165.2000 15.2000 ;
	    RECT 166.0000 15.4000 166.8000 19.8000 ;
	    RECT 170.2000 18.4000 171.4000 19.8000 ;
	    RECT 170.2000 17.8000 171.6000 18.4000 ;
	    RECT 174.8000 17.8000 175.6000 19.8000 ;
	    RECT 179.2000 18.4000 180.0000 19.8000 ;
	    RECT 179.2000 17.8000 181.2000 18.4000 ;
	    RECT 170.8000 17.0000 171.6000 17.8000 ;
	    RECT 175.0000 17.2000 175.6000 17.8000 ;
	    RECT 175.0000 16.6000 177.8000 17.2000 ;
	    RECT 177.0000 16.4000 177.8000 16.6000 ;
	    RECT 178.8000 16.4000 179.6000 17.2000 ;
	    RECT 180.4000 17.0000 181.2000 17.8000 ;
	    RECT 169.0000 15.4000 169.8000 15.6000 ;
	    RECT 166.0000 14.8000 169.8000 15.4000 ;
	    RECT 158.0000 14.2000 159.6000 14.4000 ;
	    RECT 148.6000 13.6000 159.6000 14.2000 ;
	    RECT 146.8000 12.8000 147.6000 13.0000 ;
	    RECT 143.8000 12.2000 147.6000 12.8000 ;
	    RECT 143.8000 12.0000 144.6000 12.2000 ;
	    RECT 145.4000 11.4000 146.2000 11.6000 ;
	    RECT 142.0000 10.8000 146.2000 11.4000 ;
	    RECT 113.2000 9.6000 114.6000 10.2000 ;
	    RECT 115.2000 9.6000 116.2000 10.2000 ;
	    RECT 119.6000 9.6000 121.0000 10.2000 ;
	    RECT 121.6000 9.6000 122.6000 10.2000 ;
	    RECT 126.0000 9.6000 127.4000 10.2000 ;
	    RECT 128.0000 9.6000 129.0000 10.2000 ;
	    RECT 134.2000 9.6000 136.4000 10.2000 ;
	    RECT 139.0000 9.6000 141.2000 10.2000 ;
	    RECT 102.0000 2.2000 102.8000 9.6000 ;
	    RECT 114.0000 8.4000 114.6000 9.6000 ;
	    RECT 114.0000 7.6000 114.8000 8.4000 ;
	    RECT 115.4000 2.2000 116.2000 9.6000 ;
	    RECT 120.4000 8.4000 121.0000 9.6000 ;
	    RECT 120.4000 7.6000 121.2000 8.4000 ;
	    RECT 121.8000 2.2000 122.6000 9.6000 ;
	    RECT 126.8000 8.4000 127.4000 9.6000 ;
	    RECT 126.8000 7.6000 127.6000 8.4000 ;
	    RECT 128.2000 2.2000 129.0000 9.6000 ;
	    RECT 135.6000 2.2000 136.4000 9.6000 ;
	    RECT 140.4000 2.2000 141.2000 9.6000 ;
	    RECT 142.0000 2.2000 142.8000 10.8000 ;
	    RECT 148.6000 10.4000 149.2000 13.6000 ;
	    RECT 155.8000 13.4000 156.6000 13.6000 ;
	    RECT 154.8000 12.4000 155.6000 12.6000 ;
	    RECT 157.4000 12.4000 158.2000 12.6000 ;
	    RECT 153.2000 11.8000 158.2000 12.4000 ;
	    RECT 153.2000 11.6000 154.0000 11.8000 ;
	    RECT 163.0000 11.6000 163.6000 14.6000 ;
	    RECT 164.4000 12.3000 165.2000 13.2000 ;
	    RECT 166.0000 12.3000 166.8000 14.8000 ;
	    RECT 173.0000 14.2000 173.8000 14.4000 ;
	    RECT 178.8000 14.2000 179.4000 16.4000 ;
	    RECT 183.6000 15.0000 184.4000 19.8000 ;
	    RECT 185.2000 15.2000 186.0000 19.8000 ;
	    RECT 190.0000 15.4000 190.8000 19.8000 ;
	    RECT 194.2000 18.4000 195.4000 19.8000 ;
	    RECT 194.2000 17.8000 195.6000 18.4000 ;
	    RECT 198.8000 17.8000 199.6000 19.8000 ;
	    RECT 203.2000 18.4000 204.0000 19.8000 ;
	    RECT 203.2000 17.8000 205.2000 18.4000 ;
	    RECT 194.8000 17.0000 195.6000 17.8000 ;
	    RECT 199.0000 17.2000 199.6000 17.8000 ;
	    RECT 199.0000 16.6000 201.8000 17.2000 ;
	    RECT 201.0000 16.4000 201.8000 16.6000 ;
	    RECT 202.8000 15.6000 203.6000 17.2000 ;
	    RECT 204.4000 17.0000 205.2000 17.8000 ;
	    RECT 193.0000 15.4000 193.8000 15.6000 ;
	    RECT 185.2000 14.6000 187.4000 15.2000 ;
	    RECT 182.0000 14.2000 183.6000 14.4000 ;
	    RECT 172.6000 13.6000 183.6000 14.2000 ;
	    RECT 170.8000 12.8000 171.6000 13.0000 ;
	    RECT 164.4000 11.7000 166.8000 12.3000 ;
	    RECT 167.8000 12.2000 171.6000 12.8000 ;
	    RECT 172.6000 12.4000 173.2000 13.6000 ;
	    RECT 179.8000 13.4000 180.6000 13.6000 ;
	    RECT 178.8000 12.4000 179.6000 12.6000 ;
	    RECT 181.4000 12.4000 182.2000 12.6000 ;
	    RECT 167.8000 12.0000 168.6000 12.2000 ;
	    RECT 164.4000 11.6000 165.2000 11.7000 ;
	    RECT 154.8000 11.0000 160.4000 11.2000 ;
	    RECT 154.6000 10.8000 160.4000 11.0000 ;
	    RECT 162.4000 10.8000 163.6000 11.6000 ;
	    RECT 146.8000 9.8000 149.2000 10.4000 ;
	    RECT 150.6000 10.6000 160.4000 10.8000 ;
	    RECT 150.6000 10.2000 155.4000 10.6000 ;
	    RECT 146.8000 8.8000 147.4000 9.8000 ;
	    RECT 146.0000 8.0000 147.4000 8.8000 ;
	    RECT 149.0000 9.0000 149.8000 9.2000 ;
	    RECT 150.6000 9.0000 151.2000 10.2000 ;
	    RECT 149.0000 8.4000 151.2000 9.0000 ;
	    RECT 151.8000 9.0000 157.2000 9.6000 ;
	    RECT 151.8000 8.8000 152.6000 9.0000 ;
	    RECT 156.4000 8.8000 157.2000 9.0000 ;
	    RECT 150.2000 7.4000 151.0000 7.6000 ;
	    RECT 153.0000 7.4000 153.8000 7.6000 ;
	    RECT 146.8000 6.2000 147.6000 7.0000 ;
	    RECT 150.2000 6.8000 153.8000 7.4000 ;
	    RECT 151.0000 6.2000 151.6000 6.8000 ;
	    RECT 156.4000 6.2000 157.2000 7.0000 ;
	    RECT 146.2000 2.2000 147.4000 6.2000 ;
	    RECT 150.8000 2.2000 151.6000 6.2000 ;
	    RECT 155.2000 5.6000 157.2000 6.2000 ;
	    RECT 155.2000 2.2000 156.0000 5.6000 ;
	    RECT 159.6000 2.2000 160.4000 10.6000 ;
	    RECT 163.0000 10.2000 163.6000 10.8000 ;
	    RECT 166.0000 11.4000 166.8000 11.7000 ;
	    RECT 172.4000 11.6000 173.2000 12.4000 ;
	    RECT 177.2000 11.8000 182.2000 12.4000 ;
	    RECT 177.2000 11.6000 178.0000 11.8000 ;
	    RECT 185.2000 11.6000 186.0000 13.2000 ;
	    RECT 186.8000 11.6000 187.4000 14.6000 ;
	    RECT 190.0000 14.8000 193.8000 15.4000 ;
	    RECT 169.4000 11.4000 170.2000 11.6000 ;
	    RECT 166.0000 10.8000 170.2000 11.4000 ;
	    RECT 163.0000 9.6000 165.2000 10.2000 ;
	    RECT 164.4000 2.2000 165.2000 9.6000 ;
	    RECT 166.0000 2.2000 166.8000 10.8000 ;
	    RECT 172.6000 10.4000 173.2000 11.6000 ;
	    RECT 178.8000 11.0000 184.4000 11.2000 ;
	    RECT 178.6000 10.8000 184.4000 11.0000 ;
	    RECT 170.8000 9.8000 173.2000 10.4000 ;
	    RECT 174.6000 10.6000 184.4000 10.8000 ;
	    RECT 174.6000 10.2000 179.4000 10.6000 ;
	    RECT 170.8000 8.8000 171.4000 9.8000 ;
	    RECT 170.0000 8.0000 171.4000 8.8000 ;
	    RECT 173.0000 9.0000 173.8000 9.2000 ;
	    RECT 174.6000 9.0000 175.2000 10.2000 ;
	    RECT 173.0000 8.4000 175.2000 9.0000 ;
	    RECT 175.8000 9.0000 181.2000 9.6000 ;
	    RECT 175.8000 8.8000 176.6000 9.0000 ;
	    RECT 180.4000 8.8000 181.2000 9.0000 ;
	    RECT 174.2000 7.4000 175.0000 7.6000 ;
	    RECT 177.0000 7.4000 177.8000 7.6000 ;
	    RECT 170.8000 6.2000 171.6000 7.0000 ;
	    RECT 174.2000 6.8000 177.8000 7.4000 ;
	    RECT 175.0000 6.2000 175.6000 6.8000 ;
	    RECT 180.4000 6.2000 181.2000 7.0000 ;
	    RECT 170.2000 2.2000 171.4000 6.2000 ;
	    RECT 174.8000 2.2000 175.6000 6.2000 ;
	    RECT 179.2000 5.6000 181.2000 6.2000 ;
	    RECT 179.2000 2.2000 180.0000 5.6000 ;
	    RECT 183.6000 2.2000 184.4000 10.6000 ;
	    RECT 186.8000 10.8000 188.0000 11.6000 ;
	    RECT 190.0000 11.4000 190.8000 14.8000 ;
	    RECT 197.0000 14.2000 197.8000 14.4000 ;
	    RECT 202.8000 14.2000 203.4000 15.6000 ;
	    RECT 207.6000 15.0000 208.4000 19.8000 ;
	    RECT 211.8000 16.4000 212.6000 19.8000 ;
	    RECT 210.8000 15.8000 212.6000 16.4000 ;
	    RECT 214.0000 15.8000 214.8000 19.8000 ;
	    RECT 215.6000 16.0000 216.4000 19.8000 ;
	    RECT 218.8000 16.0000 219.6000 19.8000 ;
	    RECT 215.6000 15.8000 219.6000 16.0000 ;
	    RECT 220.4000 19.2000 224.4000 19.8000 ;
	    RECT 220.4000 15.8000 221.2000 19.2000 ;
	    RECT 206.0000 14.2000 207.6000 14.4000 ;
	    RECT 196.6000 13.6000 207.6000 14.2000 ;
	    RECT 209.2000 13.6000 210.0000 15.2000 ;
	    RECT 194.8000 12.8000 195.6000 13.0000 ;
	    RECT 191.8000 12.2000 195.6000 12.8000 ;
	    RECT 196.6000 12.4000 197.2000 13.6000 ;
	    RECT 203.8000 13.4000 204.6000 13.6000 ;
	    RECT 202.8000 12.4000 203.6000 12.6000 ;
	    RECT 205.4000 12.4000 206.2000 12.6000 ;
	    RECT 191.8000 12.0000 192.6000 12.2000 ;
	    RECT 196.4000 11.6000 197.2000 12.4000 ;
	    RECT 201.2000 11.8000 206.2000 12.4000 ;
	    RECT 210.8000 12.3000 211.6000 15.8000 ;
	    RECT 214.2000 14.4000 214.8000 15.8000 ;
	    RECT 215.8000 15.4000 219.4000 15.8000 ;
	    RECT 222.0000 15.6000 222.8000 18.6000 ;
	    RECT 223.6000 16.0000 224.4000 19.2000 ;
	    RECT 226.8000 16.0000 227.6000 19.8000 ;
	    RECT 223.6000 15.8000 227.6000 16.0000 ;
	    RECT 228.4000 15.8000 229.2000 19.8000 ;
	    RECT 230.0000 16.0000 230.8000 19.8000 ;
	    RECT 233.2000 16.0000 234.0000 19.8000 ;
	    RECT 230.0000 15.8000 234.0000 16.0000 ;
	    RECT 236.4000 17.8000 237.2000 19.8000 ;
	    RECT 218.0000 14.4000 218.8000 14.8000 ;
	    RECT 222.0000 14.4000 222.6000 15.6000 ;
	    RECT 223.8000 15.4000 227.4000 15.8000 ;
	    RECT 226.0000 14.4000 226.8000 14.8000 ;
	    RECT 228.6000 14.4000 229.2000 15.8000 ;
	    RECT 230.2000 15.4000 233.8000 15.8000 ;
	    RECT 232.4000 14.4000 233.2000 14.8000 ;
	    RECT 236.4000 14.4000 237.0000 17.8000 ;
	    RECT 238.0000 15.6000 238.8000 17.2000 ;
	    RECT 239.6000 15.0000 240.4000 19.8000 ;
	    RECT 244.0000 18.4000 244.8000 19.8000 ;
	    RECT 242.8000 17.8000 244.8000 18.4000 ;
	    RECT 248.4000 17.8000 249.2000 19.8000 ;
	    RECT 252.6000 18.4000 253.8000 19.8000 ;
	    RECT 252.4000 17.8000 253.8000 18.4000 ;
	    RECT 257.2000 18.3000 258.0000 19.8000 ;
	    RECT 262.0000 18.3000 262.8000 18.4000 ;
	    RECT 242.8000 17.0000 243.6000 17.8000 ;
	    RECT 248.4000 17.2000 249.0000 17.8000 ;
	    RECT 244.4000 16.4000 245.2000 17.2000 ;
	    RECT 246.2000 16.6000 249.0000 17.2000 ;
	    RECT 252.4000 17.0000 253.2000 17.8000 ;
	    RECT 257.2000 17.7000 262.8000 18.3000 ;
	    RECT 246.2000 16.4000 247.0000 16.6000 ;
	    RECT 214.0000 13.6000 216.6000 14.4000 ;
	    RECT 218.0000 13.8000 219.6000 14.4000 ;
	    RECT 218.8000 13.6000 219.6000 13.8000 ;
	    RECT 201.2000 11.6000 202.0000 11.8000 ;
	    RECT 210.8000 11.7000 214.7000 12.3000 ;
	    RECT 193.4000 11.4000 194.2000 11.6000 ;
	    RECT 190.0000 10.8000 194.2000 11.4000 ;
	    RECT 186.8000 10.2000 187.4000 10.8000 ;
	    RECT 185.2000 9.6000 187.4000 10.2000 ;
	    RECT 185.2000 2.2000 186.0000 9.6000 ;
	    RECT 190.0000 2.2000 190.8000 10.8000 ;
	    RECT 196.6000 10.4000 197.2000 11.6000 ;
	    RECT 202.8000 11.0000 208.4000 11.2000 ;
	    RECT 202.6000 10.8000 208.4000 11.0000 ;
	    RECT 194.8000 9.8000 197.2000 10.4000 ;
	    RECT 198.6000 10.6000 208.4000 10.8000 ;
	    RECT 198.6000 10.2000 203.4000 10.6000 ;
	    RECT 194.8000 8.8000 195.4000 9.8000 ;
	    RECT 194.0000 8.0000 195.4000 8.8000 ;
	    RECT 197.0000 9.0000 197.8000 9.2000 ;
	    RECT 198.6000 9.0000 199.2000 10.2000 ;
	    RECT 197.0000 8.4000 199.2000 9.0000 ;
	    RECT 199.8000 9.0000 205.2000 9.6000 ;
	    RECT 199.8000 8.8000 200.6000 9.0000 ;
	    RECT 204.4000 8.8000 205.2000 9.0000 ;
	    RECT 198.2000 7.4000 199.0000 7.6000 ;
	    RECT 201.0000 7.4000 201.8000 7.6000 ;
	    RECT 194.8000 6.2000 195.6000 7.0000 ;
	    RECT 198.2000 6.8000 201.8000 7.4000 ;
	    RECT 199.0000 6.2000 199.6000 6.8000 ;
	    RECT 204.4000 6.2000 205.2000 7.0000 ;
	    RECT 194.2000 2.2000 195.4000 6.2000 ;
	    RECT 198.8000 2.2000 199.6000 6.2000 ;
	    RECT 203.2000 5.6000 205.2000 6.2000 ;
	    RECT 203.2000 2.2000 204.0000 5.6000 ;
	    RECT 207.6000 2.2000 208.4000 10.6000 ;
	    RECT 210.8000 2.2000 211.6000 11.7000 ;
	    RECT 214.1000 10.4000 214.7000 11.7000 ;
	    RECT 212.4000 8.8000 213.2000 10.4000 ;
	    RECT 214.0000 10.2000 214.8000 10.4000 ;
	    RECT 216.0000 10.2000 216.6000 13.6000 ;
	    RECT 217.2000 11.6000 218.0000 13.2000 ;
	    RECT 220.4000 12.8000 221.2000 14.4000 ;
	    RECT 222.0000 13.8000 224.4000 14.4000 ;
	    RECT 226.0000 14.3000 227.6000 14.4000 ;
	    RECT 228.4000 14.3000 231.0000 14.4000 ;
	    RECT 226.0000 13.8000 231.0000 14.3000 ;
	    RECT 232.4000 14.3000 234.0000 14.4000 ;
	    RECT 234.8000 14.3000 235.6000 14.4000 ;
	    RECT 232.4000 13.8000 235.6000 14.3000 ;
	    RECT 223.6000 13.6000 224.4000 13.8000 ;
	    RECT 226.8000 13.7000 231.0000 13.8000 ;
	    RECT 226.8000 13.6000 227.6000 13.7000 ;
	    RECT 228.4000 13.6000 231.0000 13.7000 ;
	    RECT 233.2000 13.7000 235.6000 13.8000 ;
	    RECT 233.2000 13.6000 234.0000 13.7000 ;
	    RECT 234.8000 13.6000 235.6000 13.7000 ;
	    RECT 236.4000 13.6000 237.2000 14.4000 ;
	    RECT 240.4000 14.2000 242.0000 14.4000 ;
	    RECT 244.6000 14.2000 245.2000 16.4000 ;
	    RECT 254.2000 15.4000 255.0000 15.6000 ;
	    RECT 257.2000 15.4000 258.0000 17.7000 ;
	    RECT 262.0000 17.6000 262.8000 17.7000 ;
	    RECT 263.6000 18.3000 264.4000 18.4000 ;
	    RECT 265.2000 18.3000 266.0000 19.8000 ;
	    RECT 263.6000 17.7000 266.0000 18.3000 ;
	    RECT 263.6000 17.6000 264.4000 17.7000 ;
	    RECT 254.2000 14.8000 258.0000 15.4000 ;
	    RECT 250.2000 14.2000 251.0000 14.4000 ;
	    RECT 240.4000 13.6000 251.4000 14.2000 ;
	    RECT 222.0000 11.6000 222.8000 13.2000 ;
	    RECT 223.8000 10.2000 224.4000 13.6000 ;
	    RECT 225.2000 11.6000 226.0000 13.2000 ;
	    RECT 228.4000 10.2000 229.2000 10.4000 ;
	    RECT 230.4000 10.2000 231.0000 13.6000 ;
	    RECT 231.6000 11.6000 232.4000 13.2000 ;
	    RECT 233.2000 12.3000 234.0000 12.4000 ;
	    RECT 234.8000 12.3000 235.6000 12.4000 ;
	    RECT 233.2000 11.7000 235.6000 12.3000 ;
	    RECT 233.2000 11.6000 234.0000 11.7000 ;
	    RECT 234.8000 10.8000 235.6000 11.7000 ;
	    RECT 236.4000 10.2000 237.0000 13.6000 ;
	    RECT 243.4000 13.4000 244.2000 13.6000 ;
	    RECT 241.8000 12.4000 242.6000 12.6000 ;
	    RECT 241.8000 12.3000 246.8000 12.4000 ;
	    RECT 247.6000 12.3000 248.4000 12.4000 ;
	    RECT 241.8000 11.8000 248.4000 12.3000 ;
	    RECT 246.0000 11.7000 248.4000 11.8000 ;
	    RECT 246.0000 11.6000 246.8000 11.7000 ;
	    RECT 247.6000 11.6000 248.4000 11.7000 ;
	    RECT 239.6000 11.0000 245.2000 11.2000 ;
	    RECT 239.6000 10.8000 245.4000 11.0000 ;
	    RECT 239.6000 10.6000 249.4000 10.8000 ;
	    RECT 214.0000 9.6000 215.4000 10.2000 ;
	    RECT 216.0000 9.6000 217.0000 10.2000 ;
	    RECT 214.8000 8.4000 215.4000 9.6000 ;
	    RECT 214.8000 7.6000 215.6000 8.4000 ;
	    RECT 216.2000 2.2000 217.0000 9.6000 ;
	    RECT 223.0000 2.2000 225.0000 10.2000 ;
	    RECT 228.4000 9.6000 229.8000 10.2000 ;
	    RECT 230.4000 9.6000 231.4000 10.2000 ;
	    RECT 229.2000 8.4000 229.8000 9.6000 ;
	    RECT 229.2000 7.6000 230.0000 8.4000 ;
	    RECT 230.6000 2.2000 231.4000 9.6000 ;
	    RECT 235.4000 9.4000 237.2000 10.2000 ;
	    RECT 235.4000 8.4000 236.2000 9.4000 ;
	    RECT 234.8000 7.6000 236.2000 8.4000 ;
	    RECT 235.4000 2.2000 236.2000 7.6000 ;
	    RECT 239.6000 2.2000 240.4000 10.6000 ;
	    RECT 244.6000 10.2000 249.4000 10.6000 ;
	    RECT 242.8000 9.0000 248.2000 9.6000 ;
	    RECT 242.8000 8.8000 243.6000 9.0000 ;
	    RECT 247.4000 8.8000 248.2000 9.0000 ;
	    RECT 248.8000 9.0000 249.4000 10.2000 ;
	    RECT 250.8000 10.4000 251.4000 13.6000 ;
	    RECT 252.4000 12.8000 253.2000 13.0000 ;
	    RECT 252.4000 12.2000 256.2000 12.8000 ;
	    RECT 255.4000 12.0000 256.2000 12.2000 ;
	    RECT 253.8000 11.4000 254.6000 11.6000 ;
	    RECT 257.2000 11.4000 258.0000 14.8000 ;
	    RECT 253.8000 10.8000 258.0000 11.4000 ;
	    RECT 250.8000 9.8000 253.2000 10.4000 ;
	    RECT 250.2000 9.0000 251.0000 9.2000 ;
	    RECT 248.8000 8.4000 251.0000 9.0000 ;
	    RECT 252.6000 8.8000 253.2000 9.8000 ;
	    RECT 252.6000 8.0000 254.0000 8.8000 ;
	    RECT 246.2000 7.4000 247.0000 7.6000 ;
	    RECT 249.0000 7.4000 249.8000 7.6000 ;
	    RECT 242.8000 6.2000 243.6000 7.0000 ;
	    RECT 246.2000 6.8000 249.8000 7.4000 ;
	    RECT 248.4000 6.2000 249.0000 6.8000 ;
	    RECT 252.4000 6.2000 253.2000 7.0000 ;
	    RECT 242.8000 5.6000 244.8000 6.2000 ;
	    RECT 244.0000 2.2000 244.8000 5.6000 ;
	    RECT 248.4000 2.2000 249.2000 6.2000 ;
	    RECT 252.6000 2.2000 253.8000 6.2000 ;
	    RECT 257.2000 2.2000 258.0000 10.8000 ;
	    RECT 265.2000 12.4000 266.0000 17.7000 ;
	    RECT 268.4000 15.2000 269.2000 19.8000 ;
	    RECT 267.0000 14.6000 269.2000 15.2000 ;
	    RECT 270.0000 15.4000 270.8000 19.8000 ;
	    RECT 274.2000 18.4000 275.4000 19.8000 ;
	    RECT 274.2000 17.8000 275.6000 18.4000 ;
	    RECT 278.8000 17.8000 279.6000 19.8000 ;
	    RECT 283.2000 18.4000 284.0000 19.8000 ;
	    RECT 283.2000 17.8000 285.2000 18.4000 ;
	    RECT 274.8000 17.0000 275.6000 17.8000 ;
	    RECT 279.0000 17.2000 279.6000 17.8000 ;
	    RECT 279.0000 16.6000 281.8000 17.2000 ;
	    RECT 281.0000 16.4000 281.8000 16.6000 ;
	    RECT 282.8000 16.4000 283.6000 17.2000 ;
	    RECT 284.4000 17.0000 285.2000 17.8000 ;
	    RECT 273.0000 15.4000 273.8000 15.6000 ;
	    RECT 270.0000 14.8000 273.8000 15.4000 ;
	    RECT 265.2000 10.2000 265.8000 12.4000 ;
	    RECT 267.0000 11.6000 267.6000 14.6000 ;
	    RECT 266.4000 10.8000 267.6000 11.6000 ;
	    RECT 267.0000 10.2000 267.6000 10.8000 ;
	    RECT 270.0000 11.4000 270.8000 14.8000 ;
	    RECT 277.0000 14.2000 277.8000 14.4000 ;
	    RECT 282.8000 14.2000 283.4000 16.4000 ;
	    RECT 287.6000 15.0000 288.4000 19.8000 ;
	    RECT 291.8000 16.4000 292.6000 19.8000 ;
	    RECT 290.8000 15.8000 292.6000 16.4000 ;
	    RECT 294.0000 15.8000 294.8000 19.8000 ;
	    RECT 295.6000 16.0000 296.4000 19.8000 ;
	    RECT 298.8000 16.0000 299.6000 19.8000 ;
	    RECT 295.6000 15.8000 299.6000 16.0000 ;
	    RECT 286.0000 14.2000 287.6000 14.4000 ;
	    RECT 276.6000 13.6000 287.6000 14.2000 ;
	    RECT 289.2000 13.6000 290.0000 15.2000 ;
	    RECT 274.8000 12.8000 275.6000 13.0000 ;
	    RECT 271.8000 12.2000 275.6000 12.8000 ;
	    RECT 276.6000 12.3000 277.2000 13.6000 ;
	    RECT 283.8000 13.4000 284.6000 13.6000 ;
	    RECT 282.8000 12.4000 283.6000 12.6000 ;
	    RECT 285.4000 12.4000 286.2000 12.6000 ;
	    RECT 278.0000 12.3000 278.8000 12.4000 ;
	    RECT 271.8000 12.0000 272.6000 12.2000 ;
	    RECT 276.5000 11.7000 278.8000 12.3000 ;
	    RECT 273.4000 11.4000 274.2000 11.6000 ;
	    RECT 270.0000 10.8000 274.2000 11.4000 ;
	    RECT 265.2000 2.2000 266.0000 10.2000 ;
	    RECT 267.0000 9.6000 269.2000 10.2000 ;
	    RECT 268.4000 2.2000 269.2000 9.6000 ;
	    RECT 270.0000 2.2000 270.8000 10.8000 ;
	    RECT 276.6000 10.4000 277.2000 11.7000 ;
	    RECT 278.0000 11.6000 278.8000 11.7000 ;
	    RECT 281.2000 11.8000 286.2000 12.4000 ;
	    RECT 290.8000 12.3000 291.6000 15.8000 ;
	    RECT 294.2000 14.4000 294.8000 15.8000 ;
	    RECT 295.8000 15.4000 299.4000 15.8000 ;
	    RECT 300.4000 15.4000 301.2000 19.8000 ;
	    RECT 304.6000 18.4000 305.8000 19.8000 ;
	    RECT 304.6000 17.8000 306.0000 18.4000 ;
	    RECT 309.2000 17.8000 310.0000 19.8000 ;
	    RECT 313.6000 18.4000 314.4000 19.8000 ;
	    RECT 313.6000 17.8000 315.6000 18.4000 ;
	    RECT 305.2000 17.0000 306.0000 17.8000 ;
	    RECT 309.4000 17.2000 310.0000 17.8000 ;
	    RECT 309.4000 16.6000 312.2000 17.2000 ;
	    RECT 311.4000 16.4000 312.2000 16.6000 ;
	    RECT 313.2000 15.6000 314.0000 17.2000 ;
	    RECT 314.8000 17.0000 315.6000 17.8000 ;
	    RECT 303.4000 15.4000 304.2000 15.6000 ;
	    RECT 300.4000 14.8000 304.2000 15.4000 ;
	    RECT 298.0000 14.4000 298.8000 14.8000 ;
	    RECT 294.0000 13.6000 296.6000 14.4000 ;
	    RECT 298.0000 13.8000 299.6000 14.4000 ;
	    RECT 298.8000 13.6000 299.6000 13.8000 ;
	    RECT 281.2000 11.6000 282.0000 11.8000 ;
	    RECT 290.8000 11.7000 294.7000 12.3000 ;
	    RECT 282.8000 11.0000 288.4000 11.2000 ;
	    RECT 282.6000 10.8000 288.4000 11.0000 ;
	    RECT 274.8000 9.8000 277.2000 10.4000 ;
	    RECT 278.6000 10.6000 288.4000 10.8000 ;
	    RECT 278.6000 10.2000 283.4000 10.6000 ;
	    RECT 274.8000 8.8000 275.4000 9.8000 ;
	    RECT 274.0000 8.0000 275.4000 8.8000 ;
	    RECT 277.0000 9.0000 277.8000 9.2000 ;
	    RECT 278.6000 9.0000 279.2000 10.2000 ;
	    RECT 277.0000 8.4000 279.2000 9.0000 ;
	    RECT 279.8000 9.0000 285.2000 9.6000 ;
	    RECT 279.8000 8.8000 280.6000 9.0000 ;
	    RECT 284.4000 8.8000 285.2000 9.0000 ;
	    RECT 278.2000 7.4000 279.0000 7.6000 ;
	    RECT 281.0000 7.4000 281.8000 7.6000 ;
	    RECT 274.8000 6.2000 275.6000 7.0000 ;
	    RECT 278.2000 6.8000 281.8000 7.4000 ;
	    RECT 279.0000 6.2000 279.6000 6.8000 ;
	    RECT 284.4000 6.2000 285.2000 7.0000 ;
	    RECT 274.2000 2.2000 275.4000 6.2000 ;
	    RECT 278.8000 2.2000 279.6000 6.2000 ;
	    RECT 283.2000 5.6000 285.2000 6.2000 ;
	    RECT 283.2000 2.2000 284.0000 5.6000 ;
	    RECT 287.6000 2.2000 288.4000 10.6000 ;
	    RECT 290.8000 2.2000 291.6000 11.7000 ;
	    RECT 294.1000 10.4000 294.7000 11.7000 ;
	    RECT 292.4000 8.8000 293.2000 10.4000 ;
	    RECT 294.0000 10.2000 294.8000 10.4000 ;
	    RECT 296.0000 10.2000 296.6000 13.6000 ;
	    RECT 297.2000 11.6000 298.0000 13.2000 ;
	    RECT 300.4000 11.4000 301.2000 14.8000 ;
	    RECT 307.4000 14.2000 308.2000 14.4000 ;
	    RECT 313.2000 14.2000 313.8000 15.6000 ;
	    RECT 318.0000 15.0000 318.8000 19.8000 ;
	    RECT 322.2000 16.4000 323.0000 19.8000 ;
	    RECT 321.2000 15.8000 323.0000 16.4000 ;
	    RECT 324.4000 15.8000 325.2000 19.8000 ;
	    RECT 326.0000 16.0000 326.8000 19.8000 ;
	    RECT 329.2000 16.0000 330.0000 19.8000 ;
	    RECT 326.0000 15.8000 330.0000 16.0000 ;
	    RECT 330.8000 16.0000 331.6000 19.8000 ;
	    RECT 334.0000 16.0000 334.8000 19.8000 ;
	    RECT 330.8000 15.8000 334.8000 16.0000 ;
	    RECT 335.6000 15.8000 336.4000 19.8000 ;
	    RECT 337.2000 19.2000 341.2000 19.8000 ;
	    RECT 337.2000 15.8000 338.0000 19.2000 ;
	    RECT 338.8000 15.8000 339.6000 18.6000 ;
	    RECT 340.4000 16.0000 341.2000 19.2000 ;
	    RECT 343.6000 16.0000 344.4000 19.8000 ;
	    RECT 346.8000 17.8000 347.6000 19.8000 ;
	    RECT 353.8000 18.4000 354.6000 19.0000 ;
	    RECT 340.4000 15.8000 344.4000 16.0000 ;
	    RECT 345.2000 16.3000 346.0000 16.4000 ;
	    RECT 346.8000 16.3000 347.4000 17.8000 ;
	    RECT 353.2000 17.6000 354.6000 18.4000 ;
	    RECT 316.4000 14.2000 318.0000 14.4000 ;
	    RECT 307.0000 13.6000 318.0000 14.2000 ;
	    RECT 319.6000 13.6000 320.4000 15.2000 ;
	    RECT 305.2000 12.8000 306.0000 13.0000 ;
	    RECT 302.2000 12.2000 306.0000 12.8000 ;
	    RECT 302.2000 12.0000 303.0000 12.2000 ;
	    RECT 303.8000 11.4000 304.6000 11.6000 ;
	    RECT 300.4000 10.8000 304.6000 11.4000 ;
	    RECT 294.0000 9.6000 295.4000 10.2000 ;
	    RECT 296.0000 9.6000 297.0000 10.2000 ;
	    RECT 294.8000 8.4000 295.4000 9.6000 ;
	    RECT 294.8000 7.6000 295.6000 8.4000 ;
	    RECT 296.2000 2.2000 297.0000 9.6000 ;
	    RECT 300.4000 2.2000 301.2000 10.8000 ;
	    RECT 307.0000 10.4000 307.6000 13.6000 ;
	    RECT 314.2000 13.4000 315.0000 13.6000 ;
	    RECT 313.2000 12.4000 314.0000 12.6000 ;
	    RECT 315.8000 12.4000 316.6000 12.6000 ;
	    RECT 311.6000 11.8000 316.6000 12.4000 ;
	    RECT 321.2000 12.3000 322.0000 15.8000 ;
	    RECT 324.6000 14.4000 325.2000 15.8000 ;
	    RECT 326.2000 15.4000 329.8000 15.8000 ;
	    RECT 331.0000 15.4000 334.6000 15.8000 ;
	    RECT 328.4000 14.4000 329.2000 14.8000 ;
	    RECT 331.6000 14.4000 332.4000 14.8000 ;
	    RECT 335.6000 14.4000 336.2000 15.8000 ;
	    RECT 338.8000 14.4000 339.4000 15.8000 ;
	    RECT 340.6000 15.4000 344.2000 15.8000 ;
	    RECT 345.2000 15.7000 347.5000 16.3000 ;
	    RECT 345.2000 15.6000 346.0000 15.7000 ;
	    RECT 342.8000 14.4000 343.6000 14.8000 ;
	    RECT 346.8000 14.4000 347.4000 15.7000 ;
	    RECT 348.4000 15.6000 349.2000 17.2000 ;
	    RECT 353.8000 16.0000 354.6000 17.6000 ;
	    RECT 358.0000 17.0000 358.8000 19.0000 ;
	    RECT 353.0000 15.4000 354.6000 16.0000 ;
	    RECT 353.0000 15.0000 353.8000 15.4000 ;
	    RECT 353.0000 14.4000 353.6000 15.0000 ;
	    RECT 358.2000 14.8000 358.8000 17.0000 ;
	    RECT 324.4000 13.6000 327.0000 14.4000 ;
	    RECT 328.4000 13.8000 330.0000 14.4000 ;
	    RECT 329.2000 13.6000 330.0000 13.8000 ;
	    RECT 330.8000 13.8000 332.4000 14.4000 ;
	    RECT 330.8000 13.6000 331.6000 13.8000 ;
	    RECT 333.8000 13.6000 336.4000 14.4000 ;
	    RECT 311.6000 11.6000 312.4000 11.8000 ;
	    RECT 321.2000 11.7000 325.1000 12.3000 ;
	    RECT 313.2000 11.0000 318.8000 11.2000 ;
	    RECT 313.0000 10.8000 318.8000 11.0000 ;
	    RECT 305.2000 9.8000 307.6000 10.4000 ;
	    RECT 309.0000 10.6000 318.8000 10.8000 ;
	    RECT 309.0000 10.2000 313.8000 10.6000 ;
	    RECT 305.2000 8.8000 305.8000 9.8000 ;
	    RECT 304.4000 8.0000 305.8000 8.8000 ;
	    RECT 307.4000 9.0000 308.2000 9.2000 ;
	    RECT 309.0000 9.0000 309.6000 10.2000 ;
	    RECT 307.4000 8.4000 309.6000 9.0000 ;
	    RECT 310.2000 9.0000 315.6000 9.6000 ;
	    RECT 310.2000 8.8000 311.0000 9.0000 ;
	    RECT 314.8000 8.8000 315.6000 9.0000 ;
	    RECT 308.6000 7.4000 309.4000 7.6000 ;
	    RECT 311.4000 7.4000 312.2000 7.6000 ;
	    RECT 305.2000 6.2000 306.0000 7.0000 ;
	    RECT 308.6000 6.8000 312.2000 7.4000 ;
	    RECT 309.4000 6.2000 310.0000 6.8000 ;
	    RECT 314.8000 6.2000 315.6000 7.0000 ;
	    RECT 304.6000 2.2000 305.8000 6.2000 ;
	    RECT 309.2000 2.2000 310.0000 6.2000 ;
	    RECT 313.6000 5.6000 315.6000 6.2000 ;
	    RECT 313.6000 2.2000 314.4000 5.6000 ;
	    RECT 318.0000 2.2000 318.8000 10.6000 ;
	    RECT 321.2000 2.2000 322.0000 11.7000 ;
	    RECT 324.5000 10.4000 325.1000 11.7000 ;
	    RECT 322.8000 8.8000 323.6000 10.4000 ;
	    RECT 324.4000 10.2000 325.2000 10.4000 ;
	    RECT 326.4000 10.2000 327.0000 13.6000 ;
	    RECT 327.6000 11.6000 328.4000 13.2000 ;
	    RECT 332.4000 11.6000 333.2000 13.2000 ;
	    RECT 333.8000 10.2000 334.4000 13.6000 ;
	    RECT 337.2000 12.3000 338.0000 14.4000 ;
	    RECT 338.8000 13.8000 341.2000 14.4000 ;
	    RECT 342.8000 14.3000 344.4000 14.4000 ;
	    RECT 345.2000 14.3000 346.0000 14.4000 ;
	    RECT 342.8000 13.8000 346.0000 14.3000 ;
	    RECT 340.4000 13.6000 341.2000 13.8000 ;
	    RECT 343.6000 13.7000 346.0000 13.8000 ;
	    RECT 343.6000 13.6000 344.4000 13.7000 ;
	    RECT 345.2000 13.6000 346.0000 13.7000 ;
	    RECT 346.8000 13.6000 347.6000 14.4000 ;
	    RECT 351.6000 13.6000 353.6000 14.4000 ;
	    RECT 354.6000 14.2000 358.8000 14.8000 ;
	    RECT 359.6000 17.0000 360.4000 19.0000 ;
	    RECT 359.6000 14.8000 360.2000 17.0000 ;
	    RECT 363.8000 16.0000 364.6000 19.0000 ;
	    RECT 363.8000 15.4000 365.4000 16.0000 ;
	    RECT 364.6000 15.0000 365.4000 15.4000 ;
	    RECT 359.6000 14.2000 363.8000 14.8000 ;
	    RECT 354.6000 13.8000 355.6000 14.2000 ;
	    RECT 335.7000 11.7000 338.0000 12.3000 ;
	    RECT 335.7000 10.4000 336.3000 11.7000 ;
	    RECT 338.8000 11.6000 339.6000 13.2000 ;
	    RECT 335.6000 10.2000 336.4000 10.4000 ;
	    RECT 340.6000 10.2000 341.2000 13.6000 ;
	    RECT 342.0000 11.6000 342.8000 13.2000 ;
	    RECT 343.6000 12.3000 344.4000 12.4000 ;
	    RECT 345.2000 12.3000 346.0000 12.4000 ;
	    RECT 343.6000 11.7000 346.0000 12.3000 ;
	    RECT 343.6000 11.6000 344.4000 11.7000 ;
	    RECT 345.2000 10.8000 346.0000 11.7000 ;
	    RECT 346.8000 10.2000 347.4000 13.6000 ;
	    RECT 350.0000 12.3000 350.8000 12.4000 ;
	    RECT 351.6000 12.3000 352.4000 12.4000 ;
	    RECT 350.0000 11.7000 352.4000 12.3000 ;
	    RECT 350.0000 11.6000 350.8000 11.7000 ;
	    RECT 351.6000 10.8000 352.4000 11.7000 ;
	    RECT 324.4000 9.6000 325.8000 10.2000 ;
	    RECT 326.4000 9.6000 327.4000 10.2000 ;
	    RECT 325.2000 8.4000 325.8000 9.6000 ;
	    RECT 325.2000 7.6000 326.0000 8.4000 ;
	    RECT 326.6000 2.2000 327.4000 9.6000 ;
	    RECT 333.4000 9.6000 334.4000 10.2000 ;
	    RECT 335.0000 9.6000 336.4000 10.2000 ;
	    RECT 333.4000 2.2000 334.2000 9.6000 ;
	    RECT 335.0000 8.4000 335.6000 9.6000 ;
	    RECT 334.8000 7.6000 335.6000 8.4000 ;
	    RECT 339.8000 4.4000 341.8000 10.2000 ;
	    RECT 338.8000 3.6000 341.8000 4.4000 ;
	    RECT 339.8000 2.2000 341.8000 3.6000 ;
	    RECT 345.8000 9.4000 347.6000 10.2000 ;
	    RECT 353.0000 9.8000 353.6000 13.6000 ;
	    RECT 354.2000 13.0000 355.6000 13.8000 ;
	    RECT 362.8000 13.8000 363.8000 14.2000 ;
	    RECT 364.8000 14.4000 365.4000 15.0000 ;
	    RECT 369.2000 15.4000 370.0000 19.8000 ;
	    RECT 373.4000 18.4000 374.6000 19.8000 ;
	    RECT 373.4000 17.8000 374.8000 18.4000 ;
	    RECT 378.0000 17.8000 378.8000 19.8000 ;
	    RECT 382.4000 18.4000 383.2000 19.8000 ;
	    RECT 382.4000 17.8000 384.4000 18.4000 ;
	    RECT 374.0000 17.0000 374.8000 17.8000 ;
	    RECT 378.2000 17.2000 378.8000 17.8000 ;
	    RECT 378.2000 16.6000 381.0000 17.2000 ;
	    RECT 380.2000 16.4000 381.0000 16.6000 ;
	    RECT 382.0000 16.4000 382.8000 17.2000 ;
	    RECT 383.6000 17.0000 384.4000 17.8000 ;
	    RECT 372.2000 15.4000 373.0000 15.6000 ;
	    RECT 369.2000 14.8000 373.0000 15.4000 ;
	    RECT 355.0000 11.0000 355.6000 13.0000 ;
	    RECT 356.4000 11.6000 357.2000 13.2000 ;
	    RECT 358.0000 12.3000 358.8000 13.2000 ;
	    RECT 359.6000 12.3000 360.4000 13.2000 ;
	    RECT 358.0000 11.7000 360.4000 12.3000 ;
	    RECT 358.0000 11.6000 358.8000 11.7000 ;
	    RECT 359.6000 11.6000 360.4000 11.7000 ;
	    RECT 361.2000 11.6000 362.0000 13.2000 ;
	    RECT 362.8000 13.0000 364.2000 13.8000 ;
	    RECT 364.8000 13.6000 366.8000 14.4000 ;
	    RECT 362.8000 11.0000 363.4000 13.0000 ;
	    RECT 355.0000 10.4000 358.8000 11.0000 ;
	    RECT 345.8000 2.2000 346.6000 9.4000 ;
	    RECT 353.0000 9.2000 354.6000 9.8000 ;
	    RECT 353.8000 2.2000 354.6000 9.2000 ;
	    RECT 358.2000 7.0000 358.8000 10.4000 ;
	    RECT 358.0000 3.0000 358.8000 7.0000 ;
	    RECT 359.6000 10.4000 363.4000 11.0000 ;
	    RECT 359.6000 7.0000 360.2000 10.4000 ;
	    RECT 364.8000 9.8000 365.4000 13.6000 ;
	    RECT 366.0000 10.8000 366.8000 12.4000 ;
	    RECT 369.2000 11.4000 370.0000 14.8000 ;
	    RECT 376.2000 14.2000 377.0000 14.4000 ;
	    RECT 382.0000 14.2000 382.6000 16.4000 ;
	    RECT 386.8000 15.0000 387.6000 19.8000 ;
	    RECT 388.4000 15.4000 389.2000 19.8000 ;
	    RECT 392.6000 18.4000 393.8000 19.8000 ;
	    RECT 392.6000 17.8000 394.0000 18.4000 ;
	    RECT 397.2000 17.8000 398.0000 19.8000 ;
	    RECT 401.6000 18.4000 402.4000 19.8000 ;
	    RECT 401.6000 17.8000 403.6000 18.4000 ;
	    RECT 393.2000 17.0000 394.0000 17.8000 ;
	    RECT 397.4000 17.2000 398.0000 17.8000 ;
	    RECT 397.4000 16.6000 400.2000 17.2000 ;
	    RECT 399.4000 16.4000 400.2000 16.6000 ;
	    RECT 401.2000 16.4000 402.0000 17.2000 ;
	    RECT 402.8000 17.0000 403.6000 17.8000 ;
	    RECT 391.4000 15.4000 392.2000 15.6000 ;
	    RECT 388.4000 14.8000 392.2000 15.4000 ;
	    RECT 385.2000 14.2000 386.8000 14.4000 ;
	    RECT 375.8000 13.6000 386.8000 14.2000 ;
	    RECT 374.0000 12.8000 374.8000 13.0000 ;
	    RECT 371.0000 12.2000 374.8000 12.8000 ;
	    RECT 371.0000 12.0000 371.8000 12.2000 ;
	    RECT 372.6000 11.4000 373.4000 11.6000 ;
	    RECT 369.2000 10.8000 373.4000 11.4000 ;
	    RECT 363.8000 9.2000 365.4000 9.8000 ;
	    RECT 359.6000 3.0000 360.4000 7.0000 ;
	    RECT 363.8000 6.4000 364.6000 9.2000 ;
	    RECT 362.8000 5.6000 364.6000 6.4000 ;
	    RECT 363.8000 2.2000 364.6000 5.6000 ;
	    RECT 369.2000 2.2000 370.0000 10.8000 ;
	    RECT 375.8000 10.4000 376.4000 13.6000 ;
	    RECT 383.0000 13.4000 383.8000 13.6000 ;
	    RECT 384.6000 12.4000 385.4000 12.6000 ;
	    RECT 377.2000 12.3000 378.0000 12.4000 ;
	    RECT 380.4000 12.3000 385.4000 12.4000 ;
	    RECT 377.2000 11.8000 385.4000 12.3000 ;
	    RECT 377.2000 11.7000 381.2000 11.8000 ;
	    RECT 377.2000 11.6000 378.0000 11.7000 ;
	    RECT 380.4000 11.6000 381.2000 11.7000 ;
	    RECT 388.4000 11.4000 389.2000 14.8000 ;
	    RECT 395.4000 14.2000 396.2000 14.4000 ;
	    RECT 398.0000 14.2000 398.8000 14.4000 ;
	    RECT 401.2000 14.2000 401.8000 16.4000 ;
	    RECT 406.0000 15.0000 406.8000 19.8000 ;
	    RECT 416.6000 16.4000 417.4000 19.8000 ;
	    RECT 415.6000 15.8000 417.4000 16.4000 ;
	    RECT 404.4000 14.2000 406.0000 14.4000 ;
	    RECT 395.0000 13.6000 406.0000 14.2000 ;
	    RECT 414.0000 13.6000 414.8000 15.2000 ;
	    RECT 393.2000 12.8000 394.0000 13.0000 ;
	    RECT 390.2000 12.2000 394.0000 12.8000 ;
	    RECT 390.2000 12.0000 391.0000 12.2000 ;
	    RECT 391.8000 11.4000 392.6000 11.6000 ;
	    RECT 382.0000 11.0000 387.6000 11.2000 ;
	    RECT 381.8000 10.8000 387.6000 11.0000 ;
	    RECT 374.0000 9.8000 376.4000 10.4000 ;
	    RECT 377.8000 10.6000 387.6000 10.8000 ;
	    RECT 377.8000 10.2000 382.6000 10.6000 ;
	    RECT 374.0000 8.8000 374.6000 9.8000 ;
	    RECT 373.2000 8.0000 374.6000 8.8000 ;
	    RECT 376.2000 9.0000 377.0000 9.2000 ;
	    RECT 377.8000 9.0000 378.4000 10.2000 ;
	    RECT 376.2000 8.4000 378.4000 9.0000 ;
	    RECT 379.0000 9.0000 384.4000 9.6000 ;
	    RECT 379.0000 8.8000 379.8000 9.0000 ;
	    RECT 383.6000 8.8000 384.4000 9.0000 ;
	    RECT 377.4000 7.4000 378.2000 7.6000 ;
	    RECT 380.2000 7.4000 381.0000 7.6000 ;
	    RECT 374.0000 6.2000 374.8000 7.0000 ;
	    RECT 377.4000 6.8000 381.0000 7.4000 ;
	    RECT 378.2000 6.2000 378.8000 6.8000 ;
	    RECT 383.6000 6.2000 384.4000 7.0000 ;
	    RECT 373.4000 2.2000 374.6000 6.2000 ;
	    RECT 378.0000 2.2000 378.8000 6.2000 ;
	    RECT 382.4000 5.6000 384.4000 6.2000 ;
	    RECT 382.4000 2.2000 383.2000 5.6000 ;
	    RECT 386.8000 2.2000 387.6000 10.6000 ;
	    RECT 388.4000 10.8000 392.6000 11.4000 ;
	    RECT 388.4000 2.2000 389.2000 10.8000 ;
	    RECT 395.0000 10.4000 395.6000 13.6000 ;
	    RECT 402.2000 13.4000 403.0000 13.6000 ;
	    RECT 401.2000 12.4000 402.0000 12.6000 ;
	    RECT 403.8000 12.4000 404.6000 12.6000 ;
	    RECT 399.6000 11.8000 404.6000 12.4000 ;
	    RECT 415.6000 12.3000 416.4000 15.8000 ;
	    RECT 418.8000 15.6000 419.6000 19.8000 ;
	    RECT 420.4000 16.0000 421.2000 19.8000 ;
	    RECT 423.6000 16.0000 424.4000 19.8000 ;
	    RECT 420.4000 15.8000 424.4000 16.0000 ;
	    RECT 419.0000 14.4000 419.6000 15.6000 ;
	    RECT 420.6000 15.4000 424.2000 15.8000 ;
	    RECT 425.2000 15.4000 426.0000 19.8000 ;
	    RECT 429.4000 18.4000 430.6000 19.8000 ;
	    RECT 429.4000 17.8000 430.8000 18.4000 ;
	    RECT 434.0000 17.8000 434.8000 19.8000 ;
	    RECT 438.4000 18.4000 439.2000 19.8000 ;
	    RECT 438.4000 17.8000 440.4000 18.4000 ;
	    RECT 430.0000 17.0000 430.8000 17.8000 ;
	    RECT 434.2000 17.2000 434.8000 17.8000 ;
	    RECT 434.2000 16.6000 437.0000 17.2000 ;
	    RECT 436.2000 16.4000 437.0000 16.6000 ;
	    RECT 438.0000 16.4000 438.8000 17.2000 ;
	    RECT 439.6000 17.0000 440.4000 17.8000 ;
	    RECT 428.2000 15.4000 429.0000 15.6000 ;
	    RECT 425.2000 14.8000 429.0000 15.4000 ;
	    RECT 422.8000 14.4000 423.6000 14.8000 ;
	    RECT 418.8000 13.6000 421.4000 14.4000 ;
	    RECT 422.8000 13.8000 424.4000 14.4000 ;
	    RECT 423.6000 13.6000 424.4000 13.8000 ;
	    RECT 399.6000 11.6000 400.4000 11.8000 ;
	    RECT 415.6000 11.7000 419.5000 12.3000 ;
	    RECT 401.2000 11.0000 406.8000 11.2000 ;
	    RECT 401.0000 10.8000 406.8000 11.0000 ;
	    RECT 393.2000 9.8000 395.6000 10.4000 ;
	    RECT 397.0000 10.6000 406.8000 10.8000 ;
	    RECT 397.0000 10.2000 401.8000 10.6000 ;
	    RECT 393.2000 8.8000 393.8000 9.8000 ;
	    RECT 392.4000 8.0000 393.8000 8.8000 ;
	    RECT 395.4000 9.0000 396.2000 9.2000 ;
	    RECT 397.0000 9.0000 397.6000 10.2000 ;
	    RECT 395.4000 8.4000 397.6000 9.0000 ;
	    RECT 398.2000 9.0000 403.6000 9.6000 ;
	    RECT 398.2000 8.8000 399.0000 9.0000 ;
	    RECT 402.8000 8.8000 403.6000 9.0000 ;
	    RECT 396.6000 7.4000 397.4000 7.6000 ;
	    RECT 399.4000 7.4000 400.2000 7.6000 ;
	    RECT 393.2000 6.2000 394.0000 7.0000 ;
	    RECT 396.6000 6.8000 400.2000 7.4000 ;
	    RECT 397.4000 6.2000 398.0000 6.8000 ;
	    RECT 402.8000 6.2000 403.6000 7.0000 ;
	    RECT 392.6000 2.2000 393.8000 6.2000 ;
	    RECT 397.2000 2.2000 398.0000 6.2000 ;
	    RECT 401.6000 5.6000 403.6000 6.2000 ;
	    RECT 401.6000 2.2000 402.4000 5.6000 ;
	    RECT 406.0000 2.2000 406.8000 10.6000 ;
	    RECT 415.6000 2.2000 416.4000 11.7000 ;
	    RECT 418.9000 10.4000 419.5000 11.7000 ;
	    RECT 417.2000 8.8000 418.0000 10.4000 ;
	    RECT 418.8000 10.2000 419.6000 10.4000 ;
	    RECT 420.8000 10.2000 421.4000 13.6000 ;
	    RECT 422.0000 11.6000 422.8000 13.2000 ;
	    RECT 425.2000 11.4000 426.0000 14.8000 ;
	    RECT 432.2000 14.2000 433.0000 14.4000 ;
	    RECT 434.8000 14.2000 435.6000 14.4000 ;
	    RECT 438.0000 14.2000 438.6000 16.4000 ;
	    RECT 442.8000 15.0000 443.6000 19.8000 ;
	    RECT 444.4000 16.0000 445.2000 19.8000 ;
	    RECT 447.6000 16.0000 448.4000 19.8000 ;
	    RECT 444.4000 15.8000 448.4000 16.0000 ;
	    RECT 449.2000 15.8000 450.0000 19.8000 ;
	    RECT 451.4000 16.4000 452.2000 19.8000 ;
	    RECT 451.4000 15.8000 453.2000 16.4000 ;
	    RECT 455.6000 16.0000 456.4000 19.8000 ;
	    RECT 458.8000 16.0000 459.6000 19.8000 ;
	    RECT 455.6000 15.8000 459.6000 16.0000 ;
	    RECT 460.4000 15.8000 461.2000 19.8000 ;
	    RECT 444.6000 15.4000 448.2000 15.8000 ;
	    RECT 445.2000 14.4000 446.0000 14.8000 ;
	    RECT 449.2000 14.4000 449.8000 15.8000 ;
	    RECT 441.2000 14.2000 442.8000 14.4000 ;
	    RECT 431.8000 13.6000 442.8000 14.2000 ;
	    RECT 444.4000 13.8000 446.0000 14.4000 ;
	    RECT 444.4000 13.6000 445.2000 13.8000 ;
	    RECT 447.4000 13.6000 450.0000 14.4000 ;
	    RECT 430.0000 12.8000 430.8000 13.0000 ;
	    RECT 427.0000 12.2000 430.8000 12.8000 ;
	    RECT 427.0000 12.0000 427.8000 12.2000 ;
	    RECT 428.6000 11.4000 429.4000 11.6000 ;
	    RECT 425.2000 10.8000 429.4000 11.4000 ;
	    RECT 418.8000 9.6000 420.2000 10.2000 ;
	    RECT 420.8000 9.6000 421.8000 10.2000 ;
	    RECT 419.6000 8.4000 420.2000 9.6000 ;
	    RECT 419.6000 7.6000 420.4000 8.4000 ;
	    RECT 421.0000 2.2000 421.8000 9.6000 ;
	    RECT 425.2000 2.2000 426.0000 10.8000 ;
	    RECT 431.8000 10.4000 432.4000 13.6000 ;
	    RECT 439.0000 13.4000 439.8000 13.6000 ;
	    RECT 438.0000 12.4000 438.8000 12.6000 ;
	    RECT 440.6000 12.4000 441.4000 12.6000 ;
	    RECT 436.4000 11.8000 441.4000 12.4000 ;
	    RECT 436.4000 11.6000 437.2000 11.8000 ;
	    RECT 446.0000 11.6000 446.8000 13.2000 ;
	    RECT 447.4000 12.4000 448.0000 13.6000 ;
	    RECT 447.4000 11.6000 448.4000 12.4000 ;
	    RECT 452.4000 12.3000 453.2000 15.8000 ;
	    RECT 455.8000 15.4000 459.4000 15.8000 ;
	    RECT 454.0000 13.6000 454.8000 15.2000 ;
	    RECT 456.4000 14.4000 457.2000 14.8000 ;
	    RECT 460.4000 14.4000 461.0000 15.8000 ;
	    RECT 462.0000 15.4000 462.8000 19.8000 ;
	    RECT 466.2000 18.4000 467.4000 19.8000 ;
	    RECT 466.2000 17.8000 467.6000 18.4000 ;
	    RECT 470.8000 17.8000 471.6000 19.8000 ;
	    RECT 475.2000 18.4000 476.0000 19.8000 ;
	    RECT 475.2000 17.8000 477.2000 18.4000 ;
	    RECT 466.8000 17.0000 467.6000 17.8000 ;
	    RECT 471.0000 17.2000 471.6000 17.8000 ;
	    RECT 471.0000 16.6000 473.8000 17.2000 ;
	    RECT 473.0000 16.4000 473.8000 16.6000 ;
	    RECT 474.8000 16.4000 475.6000 17.2000 ;
	    RECT 476.4000 17.0000 477.2000 17.8000 ;
	    RECT 465.0000 15.4000 465.8000 15.6000 ;
	    RECT 462.0000 14.8000 465.8000 15.4000 ;
	    RECT 455.6000 13.8000 457.2000 14.4000 ;
	    RECT 455.6000 13.6000 456.4000 13.8000 ;
	    RECT 458.6000 13.6000 461.2000 14.4000 ;
	    RECT 449.3000 11.7000 453.2000 12.3000 ;
	    RECT 438.0000 11.0000 443.6000 11.2000 ;
	    RECT 437.8000 10.8000 443.6000 11.0000 ;
	    RECT 430.0000 9.8000 432.4000 10.4000 ;
	    RECT 433.8000 10.6000 443.6000 10.8000 ;
	    RECT 433.8000 10.2000 438.6000 10.6000 ;
	    RECT 430.0000 8.8000 430.6000 9.8000 ;
	    RECT 429.2000 8.0000 430.6000 8.8000 ;
	    RECT 432.2000 9.0000 433.0000 9.2000 ;
	    RECT 433.8000 9.0000 434.4000 10.2000 ;
	    RECT 432.2000 8.4000 434.4000 9.0000 ;
	    RECT 435.0000 9.0000 440.4000 9.6000 ;
	    RECT 435.0000 8.8000 435.8000 9.0000 ;
	    RECT 439.6000 8.8000 440.4000 9.0000 ;
	    RECT 433.4000 7.4000 434.2000 7.6000 ;
	    RECT 436.2000 7.4000 437.0000 7.6000 ;
	    RECT 430.0000 6.2000 430.8000 7.0000 ;
	    RECT 433.4000 6.8000 437.0000 7.4000 ;
	    RECT 434.2000 6.2000 434.8000 6.8000 ;
	    RECT 439.6000 6.2000 440.4000 7.0000 ;
	    RECT 429.4000 2.2000 430.6000 6.2000 ;
	    RECT 434.0000 2.2000 434.8000 6.2000 ;
	    RECT 438.4000 5.6000 440.4000 6.2000 ;
	    RECT 438.4000 2.2000 439.2000 5.6000 ;
	    RECT 442.8000 2.2000 443.6000 10.6000 ;
	    RECT 447.4000 10.2000 448.0000 11.6000 ;
	    RECT 449.3000 10.4000 449.9000 11.7000 ;
	    RECT 449.2000 10.2000 450.0000 10.4000 ;
	    RECT 447.0000 9.6000 448.0000 10.2000 ;
	    RECT 448.6000 9.6000 450.0000 10.2000 ;
	    RECT 447.0000 2.2000 447.8000 9.6000 ;
	    RECT 448.6000 8.4000 449.2000 9.6000 ;
	    RECT 450.8000 8.8000 451.6000 10.4000 ;
	    RECT 448.4000 7.6000 449.2000 8.4000 ;
	    RECT 452.4000 2.2000 453.2000 11.7000 ;
	    RECT 457.2000 11.6000 458.0000 13.2000 ;
	    RECT 458.6000 10.2000 459.2000 13.6000 ;
	    RECT 462.0000 11.4000 462.8000 14.8000 ;
	    RECT 468.4000 14.2000 469.8000 14.4000 ;
	    RECT 474.8000 14.2000 475.4000 16.4000 ;
	    RECT 479.6000 15.0000 480.4000 19.8000 ;
	    RECT 481.2000 15.4000 482.0000 19.8000 ;
	    RECT 485.4000 18.4000 486.6000 19.8000 ;
	    RECT 485.4000 17.8000 486.8000 18.4000 ;
	    RECT 490.0000 17.8000 490.8000 19.8000 ;
	    RECT 494.4000 18.4000 495.2000 19.8000 ;
	    RECT 494.4000 17.8000 496.4000 18.4000 ;
	    RECT 486.0000 17.0000 486.8000 17.8000 ;
	    RECT 490.2000 17.2000 490.8000 17.8000 ;
	    RECT 490.2000 16.6000 493.0000 17.2000 ;
	    RECT 492.2000 16.4000 493.0000 16.6000 ;
	    RECT 494.0000 16.4000 494.8000 17.2000 ;
	    RECT 495.6000 17.0000 496.4000 17.8000 ;
	    RECT 484.2000 15.4000 485.0000 15.6000 ;
	    RECT 481.2000 14.8000 485.0000 15.4000 ;
	    RECT 478.0000 14.2000 479.6000 14.4000 ;
	    RECT 468.4000 13.6000 479.6000 14.2000 ;
	    RECT 466.8000 12.8000 467.6000 13.0000 ;
	    RECT 463.8000 12.2000 467.6000 12.8000 ;
	    RECT 463.8000 12.0000 464.6000 12.2000 ;
	    RECT 465.4000 11.4000 466.2000 11.6000 ;
	    RECT 462.0000 10.8000 466.2000 11.4000 ;
	    RECT 460.4000 10.2000 461.2000 10.4000 ;
	    RECT 458.2000 9.6000 459.2000 10.2000 ;
	    RECT 459.8000 9.6000 461.2000 10.2000 ;
	    RECT 458.2000 2.2000 459.0000 9.6000 ;
	    RECT 459.8000 8.4000 460.4000 9.6000 ;
	    RECT 459.6000 7.6000 460.4000 8.4000 ;
	    RECT 462.0000 2.2000 462.8000 10.8000 ;
	    RECT 468.6000 10.4000 469.2000 13.6000 ;
	    RECT 475.8000 13.4000 476.6000 13.6000 ;
	    RECT 477.4000 12.4000 478.2000 12.6000 ;
	    RECT 470.0000 12.3000 470.8000 12.4000 ;
	    RECT 473.2000 12.3000 478.2000 12.4000 ;
	    RECT 470.0000 11.8000 478.2000 12.3000 ;
	    RECT 470.0000 11.7000 474.0000 11.8000 ;
	    RECT 470.0000 11.6000 470.8000 11.7000 ;
	    RECT 473.2000 11.6000 474.0000 11.7000 ;
	    RECT 481.2000 11.4000 482.0000 14.8000 ;
	    RECT 487.6000 14.2000 489.0000 14.4000 ;
	    RECT 494.0000 14.2000 494.6000 16.4000 ;
	    RECT 498.8000 15.0000 499.6000 19.8000 ;
	    RECT 502.0000 15.2000 502.8000 19.8000 ;
	    RECT 505.2000 15.2000 506.0000 19.8000 ;
	    RECT 508.4000 15.2000 509.2000 19.8000 ;
	    RECT 511.6000 15.2000 512.4000 19.8000 ;
	    RECT 500.4000 14.4000 502.8000 15.2000 ;
	    RECT 503.8000 14.4000 506.0000 15.2000 ;
	    RECT 507.0000 14.4000 509.2000 15.2000 ;
	    RECT 510.6000 14.4000 512.4000 15.2000 ;
	    RECT 497.2000 14.2000 498.8000 14.4000 ;
	    RECT 487.6000 13.6000 498.8000 14.2000 ;
	    RECT 486.0000 12.8000 486.8000 13.0000 ;
	    RECT 483.0000 12.2000 486.8000 12.8000 ;
	    RECT 483.0000 12.0000 483.8000 12.2000 ;
	    RECT 484.6000 11.4000 485.4000 11.6000 ;
	    RECT 474.8000 11.0000 480.4000 11.2000 ;
	    RECT 474.6000 10.8000 480.4000 11.0000 ;
	    RECT 466.8000 9.8000 469.2000 10.4000 ;
	    RECT 470.6000 10.6000 480.4000 10.8000 ;
	    RECT 470.6000 10.2000 475.4000 10.6000 ;
	    RECT 466.8000 8.8000 467.4000 9.8000 ;
	    RECT 466.0000 8.0000 467.4000 8.8000 ;
	    RECT 469.0000 9.0000 469.8000 9.2000 ;
	    RECT 470.6000 9.0000 471.2000 10.2000 ;
	    RECT 469.0000 8.4000 471.2000 9.0000 ;
	    RECT 471.8000 9.0000 477.2000 9.6000 ;
	    RECT 471.8000 8.8000 472.6000 9.0000 ;
	    RECT 476.4000 8.8000 477.2000 9.0000 ;
	    RECT 470.2000 7.4000 471.0000 7.6000 ;
	    RECT 473.0000 7.4000 473.8000 7.6000 ;
	    RECT 466.8000 6.2000 467.6000 7.0000 ;
	    RECT 470.2000 6.8000 473.8000 7.4000 ;
	    RECT 471.0000 6.2000 471.6000 6.8000 ;
	    RECT 476.4000 6.2000 477.2000 7.0000 ;
	    RECT 466.2000 2.2000 467.4000 6.2000 ;
	    RECT 470.8000 2.2000 471.6000 6.2000 ;
	    RECT 475.2000 5.6000 477.2000 6.2000 ;
	    RECT 475.2000 2.2000 476.0000 5.6000 ;
	    RECT 479.6000 2.2000 480.4000 10.6000 ;
	    RECT 481.2000 10.8000 485.4000 11.4000 ;
	    RECT 481.2000 2.2000 482.0000 10.8000 ;
	    RECT 487.8000 10.4000 488.4000 13.6000 ;
	    RECT 495.0000 13.4000 495.8000 13.6000 ;
	    RECT 496.6000 12.4000 497.4000 12.6000 ;
	    RECT 492.4000 11.8000 497.4000 12.4000 ;
	    RECT 492.4000 11.6000 493.2000 11.8000 ;
	    RECT 500.4000 11.6000 501.2000 14.4000 ;
	    RECT 503.8000 13.8000 504.6000 14.4000 ;
	    RECT 507.0000 13.8000 507.8000 14.4000 ;
	    RECT 510.6000 13.8000 511.4000 14.4000 ;
	    RECT 502.0000 13.0000 504.6000 13.8000 ;
	    RECT 505.4000 13.0000 507.8000 13.8000 ;
	    RECT 508.8000 13.0000 511.4000 13.8000 ;
	    RECT 503.8000 11.6000 504.6000 13.0000 ;
	    RECT 507.0000 11.6000 507.8000 13.0000 ;
	    RECT 510.6000 11.6000 511.4000 13.0000 ;
	    RECT 494.0000 11.0000 499.6000 11.2000 ;
	    RECT 493.8000 10.8000 499.6000 11.0000 ;
	    RECT 500.4000 10.8000 502.8000 11.6000 ;
	    RECT 503.8000 10.8000 506.0000 11.6000 ;
	    RECT 507.0000 10.8000 509.2000 11.6000 ;
	    RECT 510.6000 10.8000 512.4000 11.6000 ;
	    RECT 486.0000 9.8000 488.4000 10.4000 ;
	    RECT 489.8000 10.6000 499.6000 10.8000 ;
	    RECT 489.8000 10.2000 494.6000 10.6000 ;
	    RECT 486.0000 8.8000 486.6000 9.8000 ;
	    RECT 485.2000 8.0000 486.6000 8.8000 ;
	    RECT 488.2000 9.0000 489.0000 9.2000 ;
	    RECT 489.8000 9.0000 490.4000 10.2000 ;
	    RECT 488.2000 8.4000 490.4000 9.0000 ;
	    RECT 491.0000 9.0000 496.4000 9.6000 ;
	    RECT 491.0000 8.8000 491.8000 9.0000 ;
	    RECT 495.6000 8.8000 496.4000 9.0000 ;
	    RECT 489.4000 7.4000 490.2000 7.6000 ;
	    RECT 492.2000 7.4000 493.0000 7.6000 ;
	    RECT 486.0000 6.2000 486.8000 7.0000 ;
	    RECT 489.4000 6.8000 493.0000 7.4000 ;
	    RECT 490.2000 6.2000 490.8000 6.8000 ;
	    RECT 495.6000 6.2000 496.4000 7.0000 ;
	    RECT 485.4000 2.2000 486.6000 6.2000 ;
	    RECT 490.0000 2.2000 490.8000 6.2000 ;
	    RECT 494.4000 5.6000 496.4000 6.2000 ;
	    RECT 494.4000 2.2000 495.2000 5.6000 ;
	    RECT 498.8000 2.2000 499.6000 10.6000 ;
	    RECT 502.0000 2.2000 502.8000 10.8000 ;
	    RECT 505.2000 2.2000 506.0000 10.8000 ;
	    RECT 508.4000 2.2000 509.2000 10.8000 ;
	    RECT 511.6000 2.2000 512.4000 10.8000 ;
         LAYER metal2 ;
	    RECT 1.2000 331.6000 2.0000 332.4000 ;
	    RECT 1.3000 328.4000 1.9000 331.6000 ;
	    RECT 1.2000 327.6000 2.0000 328.4000 ;
	    RECT 6.0000 326.2000 6.8000 337.8000 ;
	    RECT 14.0000 335.6000 14.8000 336.4000 ;
	    RECT 12.4000 333.6000 13.2000 334.4000 ;
	    RECT 12.5000 318.4000 13.1000 333.6000 ;
	    RECT 14.1000 332.6000 14.7000 335.6000 ;
	    RECT 14.0000 331.8000 14.8000 332.6000 ;
	    RECT 15.6000 326.2000 16.4000 337.8000 ;
	    RECT 18.8000 330.2000 19.6000 335.8000 ;
	    RECT 36.4000 335.6000 37.2000 336.4000 ;
	    RECT 34.8000 333.6000 35.6000 334.4000 ;
	    RECT 41.2000 333.6000 42.0000 334.4000 ;
	    RECT 47.6000 333.6000 48.4000 334.4000 ;
	    RECT 23.6000 331.6000 24.4000 332.4000 ;
	    RECT 25.2000 331.6000 26.0000 332.4000 ;
	    RECT 30.0000 331.6000 30.8000 332.4000 ;
	    RECT 34.8000 331.6000 35.6000 332.4000 ;
	    RECT 39.6000 331.6000 40.4000 332.4000 ;
	    RECT 12.4000 317.6000 13.2000 318.4000 ;
	    RECT 25.3000 316.3000 25.9000 331.6000 ;
	    RECT 30.1000 330.4000 30.7000 331.6000 ;
	    RECT 30.0000 329.6000 30.8000 330.4000 ;
	    RECT 33.2000 329.6000 34.0000 330.4000 ;
	    RECT 25.3000 315.7000 27.5000 316.3000 ;
	    RECT 9.2000 313.6000 10.0000 314.4000 ;
	    RECT 25.2000 313.6000 26.0000 314.4000 ;
	    RECT 9.3000 310.4000 9.9000 313.6000 ;
	    RECT 4.4000 309.6000 5.2000 310.4000 ;
	    RECT 9.2000 309.6000 10.0000 310.4000 ;
	    RECT 4.5000 300.4000 5.1000 309.6000 ;
	    RECT 12.4000 303.6000 13.2000 304.4000 ;
	    RECT 1.2000 299.6000 2.0000 300.4000 ;
	    RECT 4.4000 299.6000 5.2000 300.4000 ;
	    RECT 1.3000 298.4000 1.9000 299.6000 ;
	    RECT 1.2000 297.6000 2.0000 298.4000 ;
	    RECT 4.5000 274.3000 5.1000 299.6000 ;
	    RECT 6.0000 286.2000 6.8000 297.8000 ;
	    RECT 12.5000 294.4000 13.1000 303.6000 ;
	    RECT 26.9000 298.4000 27.5000 315.7000 ;
	    RECT 30.0000 304.2000 30.8000 315.8000 ;
	    RECT 34.9000 310.4000 35.5000 331.6000 ;
	    RECT 36.4000 329.6000 37.2000 330.4000 ;
	    RECT 39.7000 328.4000 40.3000 331.6000 ;
	    RECT 39.6000 327.6000 40.4000 328.4000 ;
	    RECT 36.4000 325.6000 37.2000 326.4000 ;
	    RECT 34.8000 309.6000 35.6000 310.4000 ;
	    RECT 36.5000 308.4000 37.1000 325.6000 ;
	    RECT 41.3000 324.4000 41.9000 333.6000 ;
	    RECT 46.0000 331.6000 46.8000 332.4000 ;
	    RECT 46.1000 330.4000 46.7000 331.6000 ;
	    RECT 46.0000 329.6000 46.8000 330.4000 ;
	    RECT 47.7000 330.3000 48.3000 333.6000 ;
	    RECT 49.2000 331.6000 50.0000 332.4000 ;
	    RECT 52.4000 331.6000 53.2000 332.4000 ;
	    RECT 47.7000 329.7000 49.9000 330.3000 ;
	    RECT 41.2000 323.6000 42.0000 324.4000 ;
	    RECT 38.0000 315.6000 38.8000 316.4000 ;
	    RECT 38.1000 310.2000 38.7000 315.6000 ;
	    RECT 38.0000 309.4000 38.8000 310.2000 ;
	    RECT 36.4000 307.6000 37.2000 308.4000 ;
	    RECT 12.4000 293.6000 13.2000 294.4000 ;
	    RECT 12.5000 292.4000 13.1000 293.6000 ;
	    RECT 12.4000 291.6000 13.2000 292.4000 ;
	    RECT 14.0000 291.8000 14.8000 292.6000 ;
	    RECT 14.1000 274.4000 14.7000 291.8000 ;
	    RECT 15.6000 286.2000 16.4000 297.8000 ;
	    RECT 18.8000 290.2000 19.6000 295.8000 ;
	    RECT 25.2000 286.2000 26.0000 297.8000 ;
	    RECT 26.8000 297.6000 27.6000 298.4000 ;
	    RECT 26.8000 291.6000 27.6000 292.4000 ;
	    RECT 33.2000 291.8000 34.0000 292.6000 ;
	    RECT 20.4000 283.6000 21.2000 284.4000 ;
	    RECT 20.5000 278.4000 21.1000 283.6000 ;
	    RECT 20.4000 277.6000 21.2000 278.4000 ;
	    RECT 4.5000 273.7000 6.7000 274.3000 ;
	    RECT 6.1000 272.4000 6.7000 273.7000 ;
	    RECT 14.0000 273.6000 14.8000 274.4000 ;
	    RECT 4.4000 271.6000 5.2000 272.4000 ;
	    RECT 6.0000 271.6000 6.8000 272.4000 ;
	    RECT 17.2000 271.6000 18.0000 272.4000 ;
	    RECT 4.5000 270.4000 5.1000 271.6000 ;
	    RECT 4.4000 269.6000 5.2000 270.4000 ;
	    RECT 14.0000 269.6000 14.8000 270.4000 ;
	    RECT 17.2000 269.6000 18.0000 270.4000 ;
	    RECT 4.4000 267.6000 5.2000 268.4000 ;
	    RECT 10.8000 268.3000 11.6000 268.4000 ;
	    RECT 9.3000 267.7000 11.6000 268.3000 ;
	    RECT 4.5000 252.4000 5.1000 267.6000 ;
	    RECT 6.0000 263.6000 6.8000 264.4000 ;
	    RECT 4.4000 251.6000 5.2000 252.4000 ;
	    RECT 4.4000 231.6000 5.2000 232.4000 ;
	    RECT 4.5000 230.4000 5.1000 231.6000 ;
	    RECT 4.4000 229.6000 5.2000 230.4000 ;
	    RECT 9.3000 218.4000 9.9000 267.7000 ;
	    RECT 10.8000 267.6000 11.6000 267.7000 ;
	    RECT 10.9000 266.4000 11.5000 267.6000 ;
	    RECT 10.8000 265.6000 11.6000 266.4000 ;
	    RECT 12.4000 245.6000 13.2000 246.4000 ;
	    RECT 10.8000 243.6000 11.6000 244.4000 ;
	    RECT 12.5000 238.4000 13.1000 245.6000 ;
	    RECT 12.4000 237.6000 13.2000 238.4000 ;
	    RECT 10.8000 235.6000 11.6000 236.4000 ;
	    RECT 10.9000 230.4000 11.5000 235.6000 ;
	    RECT 14.1000 230.4000 14.7000 269.6000 ;
	    RECT 20.5000 268.4000 21.1000 277.6000 ;
	    RECT 20.4000 267.6000 21.2000 268.4000 ;
	    RECT 23.6000 264.2000 24.4000 275.8000 ;
	    RECT 26.9000 270.4000 27.5000 291.6000 ;
	    RECT 33.3000 282.4000 33.9000 291.8000 ;
	    RECT 34.8000 286.2000 35.6000 297.8000 ;
	    RECT 36.5000 294.4000 37.1000 307.6000 ;
	    RECT 39.6000 304.2000 40.4000 315.8000 ;
	    RECT 44.4000 313.6000 45.2000 314.4000 ;
	    RECT 42.8000 306.2000 43.6000 311.8000 ;
	    RECT 47.6000 311.6000 48.4000 312.4000 ;
	    RECT 47.6000 309.6000 48.4000 310.4000 ;
	    RECT 39.6000 297.6000 40.4000 298.4000 ;
	    RECT 36.4000 293.6000 37.2000 294.4000 ;
	    RECT 38.0000 290.2000 38.8000 295.8000 ;
	    RECT 42.8000 289.6000 43.6000 290.4000 ;
	    RECT 33.2000 281.6000 34.0000 282.4000 ;
	    RECT 26.8000 269.6000 27.6000 270.4000 ;
	    RECT 31.6000 269.4000 32.4000 270.2000 ;
	    RECT 31.7000 268.4000 32.3000 269.4000 ;
	    RECT 31.6000 267.6000 32.4000 268.4000 ;
	    RECT 33.2000 264.2000 34.0000 275.8000 ;
	    RECT 36.4000 266.2000 37.2000 271.8000 ;
	    RECT 38.0000 271.6000 38.8000 272.4000 ;
	    RECT 42.9000 272.3000 43.5000 289.6000 ;
	    RECT 44.4000 286.2000 45.2000 297.8000 ;
	    RECT 46.0000 291.6000 46.8000 292.4000 ;
	    RECT 47.7000 282.3000 48.3000 309.6000 ;
	    RECT 49.3000 308.4000 49.9000 329.7000 ;
	    RECT 52.4000 329.6000 53.2000 330.4000 ;
	    RECT 58.8000 326.2000 59.6000 337.8000 ;
	    RECT 66.8000 333.6000 67.6000 334.4000 ;
	    RECT 66.9000 332.6000 67.5000 333.6000 ;
	    RECT 60.4000 331.6000 61.2000 332.4000 ;
	    RECT 66.8000 331.8000 67.6000 332.6000 ;
	    RECT 60.5000 326.4000 61.1000 331.6000 ;
	    RECT 65.2000 327.6000 66.0000 328.4000 ;
	    RECT 60.4000 325.6000 61.2000 326.4000 ;
	    RECT 58.8000 323.6000 59.6000 324.4000 ;
	    RECT 58.9000 318.4000 59.5000 323.6000 ;
	    RECT 65.3000 318.4000 65.9000 327.6000 ;
	    RECT 68.4000 326.2000 69.2000 337.8000 ;
	    RECT 71.6000 330.2000 72.4000 335.8000 ;
	    RECT 73.2000 333.6000 74.0000 334.4000 ;
	    RECT 78.0000 333.6000 78.8000 334.4000 ;
	    RECT 73.2000 331.6000 74.0000 332.4000 ;
	    RECT 76.4000 332.3000 77.2000 332.4000 ;
	    RECT 74.9000 331.7000 77.2000 332.3000 ;
	    RECT 73.3000 330.4000 73.9000 331.6000 ;
	    RECT 73.2000 329.6000 74.0000 330.4000 ;
	    RECT 71.6000 323.6000 72.4000 324.4000 ;
	    RECT 58.8000 317.6000 59.6000 318.4000 ;
	    RECT 65.2000 317.6000 66.0000 318.4000 ;
	    RECT 54.0000 315.6000 54.8000 316.4000 ;
	    RECT 66.8000 315.6000 67.6000 316.4000 ;
	    RECT 55.6000 313.6000 56.4000 314.4000 ;
	    RECT 50.8000 311.6000 51.6000 312.4000 ;
	    RECT 54.0000 309.6000 54.8000 310.4000 ;
	    RECT 55.7000 308.4000 56.3000 313.6000 ;
	    RECT 62.0000 312.3000 62.8000 312.4000 ;
	    RECT 63.6000 312.3000 64.4000 312.4000 ;
	    RECT 62.0000 311.7000 64.4000 312.3000 ;
	    RECT 62.0000 311.6000 62.8000 311.7000 ;
	    RECT 63.6000 311.6000 64.4000 311.7000 ;
	    RECT 60.4000 309.6000 61.2000 310.4000 ;
	    RECT 49.2000 307.6000 50.0000 308.4000 ;
	    RECT 55.6000 307.6000 56.4000 308.4000 ;
	    RECT 46.1000 281.7000 48.3000 282.3000 ;
	    RECT 46.1000 274.3000 46.7000 281.7000 ;
	    RECT 47.6000 275.6000 48.4000 276.4000 ;
	    RECT 46.1000 273.7000 48.3000 274.3000 ;
	    RECT 44.4000 272.3000 45.2000 272.4000 ;
	    RECT 42.9000 271.7000 45.2000 272.3000 ;
	    RECT 44.4000 271.6000 45.2000 271.7000 ;
	    RECT 38.1000 270.4000 38.7000 271.6000 ;
	    RECT 47.7000 270.4000 48.3000 273.7000 ;
	    RECT 38.0000 269.6000 38.8000 270.4000 ;
	    RECT 41.2000 269.6000 42.0000 270.4000 ;
	    RECT 47.6000 269.6000 48.4000 270.4000 ;
	    RECT 38.0000 267.6000 38.8000 268.4000 ;
	    RECT 41.3000 262.4000 41.9000 269.6000 ;
	    RECT 42.8000 267.6000 43.6000 268.4000 ;
	    RECT 41.2000 261.6000 42.0000 262.4000 ;
	    RECT 47.7000 260.4000 48.3000 269.6000 ;
	    RECT 49.3000 268.4000 49.9000 307.6000 ;
	    RECT 57.2000 306.3000 58.0000 306.4000 ;
	    RECT 57.2000 305.7000 59.5000 306.3000 ;
	    RECT 57.2000 305.6000 58.0000 305.7000 ;
	    RECT 52.4000 291.8000 53.2000 292.6000 ;
	    RECT 52.5000 270.4000 53.1000 291.8000 ;
	    RECT 54.0000 286.2000 54.8000 297.8000 ;
	    RECT 58.9000 296.4000 59.5000 305.7000 ;
	    RECT 60.5000 302.4000 61.1000 309.6000 ;
	    RECT 60.4000 301.6000 61.2000 302.4000 ;
	    RECT 57.2000 290.2000 58.0000 295.8000 ;
	    RECT 58.8000 295.6000 59.6000 296.4000 ;
	    RECT 58.9000 294.4000 59.5000 295.6000 ;
	    RECT 58.8000 293.6000 59.6000 294.4000 ;
	    RECT 62.0000 293.6000 62.8000 294.4000 ;
	    RECT 63.7000 290.4000 64.3000 311.6000 ;
	    RECT 66.9000 310.4000 67.5000 315.6000 ;
	    RECT 65.2000 309.6000 66.0000 310.4000 ;
	    RECT 66.8000 309.6000 67.6000 310.4000 ;
	    RECT 65.3000 294.4000 65.9000 309.6000 ;
	    RECT 68.4000 303.6000 69.2000 304.4000 ;
	    RECT 70.0000 303.6000 70.8000 304.4000 ;
	    RECT 68.5000 294.4000 69.1000 303.6000 ;
	    RECT 70.1000 296.4000 70.7000 303.6000 ;
	    RECT 71.7000 298.4000 72.3000 323.6000 ;
	    RECT 74.9000 318.4000 75.5000 331.7000 ;
	    RECT 76.4000 331.6000 77.2000 331.7000 ;
	    RECT 78.1000 324.4000 78.7000 333.6000 ;
	    RECT 86.0000 325.6000 86.8000 326.4000 ;
	    RECT 98.8000 326.2000 99.6000 337.8000 ;
	    RECT 106.8000 333.6000 107.6000 334.4000 ;
	    RECT 106.9000 332.6000 107.5000 333.6000 ;
	    RECT 100.4000 331.6000 101.2000 332.4000 ;
	    RECT 106.8000 331.8000 107.6000 332.6000 ;
	    RECT 106.9000 331.7000 107.5000 331.8000 ;
	    RECT 100.5000 330.4000 101.1000 331.6000 ;
	    RECT 100.4000 329.6000 101.2000 330.4000 ;
	    RECT 100.5000 326.4000 101.1000 329.6000 ;
	    RECT 100.4000 325.6000 101.2000 326.4000 ;
	    RECT 108.4000 326.2000 109.2000 337.8000 ;
	    RECT 130.8000 337.6000 131.6000 338.4000 ;
	    RECT 111.6000 330.2000 112.4000 335.8000 ;
	    RECT 116.4000 333.6000 117.2000 334.4000 ;
	    RECT 122.8000 333.6000 123.6000 334.4000 ;
	    RECT 129.2000 333.6000 130.0000 334.4000 ;
	    RECT 78.0000 323.6000 78.8000 324.4000 ;
	    RECT 81.2000 323.6000 82.0000 324.4000 ;
	    RECT 81.3000 318.4000 81.9000 323.6000 ;
	    RECT 74.8000 317.6000 75.6000 318.4000 ;
	    RECT 81.2000 317.6000 82.0000 318.4000 ;
	    RECT 82.8000 317.6000 83.6000 318.4000 ;
	    RECT 81.2000 313.6000 82.0000 314.4000 ;
	    RECT 78.0000 311.6000 78.8000 312.4000 ;
	    RECT 82.9000 310.4000 83.5000 317.6000 ;
	    RECT 74.8000 309.6000 75.6000 310.4000 ;
	    RECT 82.8000 309.6000 83.6000 310.4000 ;
	    RECT 73.2000 307.6000 74.0000 308.4000 ;
	    RECT 71.6000 297.6000 72.4000 298.4000 ;
	    RECT 70.0000 295.6000 70.8000 296.4000 ;
	    RECT 71.6000 295.6000 72.4000 296.4000 ;
	    RECT 65.2000 293.6000 66.0000 294.4000 ;
	    RECT 68.4000 293.6000 69.2000 294.4000 ;
	    RECT 70.0000 292.3000 70.8000 292.4000 ;
	    RECT 71.7000 292.3000 72.3000 295.6000 ;
	    RECT 73.3000 294.4000 73.9000 307.6000 ;
	    RECT 74.9000 306.4000 75.5000 309.6000 ;
	    RECT 74.8000 305.6000 75.6000 306.4000 ;
	    RECT 79.6000 305.6000 80.4000 306.4000 ;
	    RECT 84.4000 306.2000 85.2000 311.8000 ;
	    RECT 86.1000 308.4000 86.7000 325.6000 ;
	    RECT 116.5000 324.4000 117.1000 333.6000 ;
	    RECT 122.8000 331.6000 123.6000 332.4000 ;
	    RECT 127.6000 331.6000 128.4000 332.4000 ;
	    RECT 122.9000 330.4000 123.5000 331.6000 ;
	    RECT 122.8000 329.6000 123.6000 330.4000 ;
	    RECT 129.3000 328.4000 129.9000 333.6000 ;
	    RECT 134.0000 329.6000 134.8000 330.4000 ;
	    RECT 119.6000 327.6000 120.4000 328.4000 ;
	    RECT 129.2000 327.6000 130.0000 328.4000 ;
	    RECT 118.0000 325.6000 118.8000 326.4000 ;
	    RECT 94.0000 323.6000 94.8000 324.4000 ;
	    RECT 116.4000 323.6000 117.2000 324.4000 ;
	    RECT 86.0000 307.6000 86.8000 308.4000 ;
	    RECT 79.7000 304.4000 80.3000 305.6000 ;
	    RECT 79.6000 303.6000 80.4000 304.4000 ;
	    RECT 87.6000 304.2000 88.4000 315.8000 ;
	    RECT 90.8000 311.6000 91.6000 312.4000 ;
	    RECT 90.9000 310.4000 91.5000 311.6000 ;
	    RECT 90.8000 309.6000 91.6000 310.4000 ;
	    RECT 89.2000 305.6000 90.0000 306.4000 ;
	    RECT 84.4000 299.6000 85.2000 300.4000 ;
	    RECT 84.5000 294.4000 85.1000 299.6000 ;
	    RECT 73.2000 293.6000 74.0000 294.4000 ;
	    RECT 74.8000 293.6000 75.6000 294.4000 ;
	    RECT 84.4000 293.6000 85.2000 294.4000 ;
	    RECT 86.0000 293.6000 86.8000 294.4000 ;
	    RECT 70.0000 291.7000 72.3000 292.3000 ;
	    RECT 70.0000 291.6000 70.8000 291.7000 ;
	    RECT 73.2000 291.6000 74.0000 292.4000 ;
	    RECT 78.0000 291.6000 78.8000 292.4000 ;
	    RECT 81.2000 291.6000 82.0000 292.4000 ;
	    RECT 82.8000 291.6000 83.6000 292.4000 ;
	    RECT 86.0000 291.6000 86.8000 292.4000 ;
	    RECT 63.6000 289.6000 64.4000 290.4000 ;
	    RECT 63.7000 288.4000 64.3000 289.6000 ;
	    RECT 63.6000 287.6000 64.4000 288.4000 ;
	    RECT 73.3000 284.4000 73.9000 291.6000 ;
	    RECT 78.1000 290.4000 78.7000 291.6000 ;
	    RECT 78.0000 289.6000 78.8000 290.4000 ;
	    RECT 76.4000 287.6000 77.2000 288.4000 ;
	    RECT 73.2000 283.6000 74.0000 284.4000 ;
	    RECT 65.2000 281.6000 66.0000 282.4000 ;
	    RECT 55.6000 277.6000 56.4000 278.4000 ;
	    RECT 55.7000 272.4000 56.3000 277.6000 ;
	    RECT 58.8000 273.6000 59.6000 274.4000 ;
	    RECT 54.0000 271.6000 54.8000 272.4000 ;
	    RECT 55.6000 271.6000 56.4000 272.4000 ;
	    RECT 57.2000 271.6000 58.0000 272.4000 ;
	    RECT 54.1000 270.4000 54.7000 271.6000 ;
	    RECT 52.4000 269.6000 53.2000 270.4000 ;
	    RECT 54.0000 269.6000 54.8000 270.4000 ;
	    RECT 49.2000 267.6000 50.0000 268.4000 ;
	    RECT 49.3000 266.4000 49.9000 267.6000 ;
	    RECT 49.2000 265.6000 50.0000 266.4000 ;
	    RECT 57.3000 264.4000 57.9000 271.6000 ;
	    RECT 58.9000 270.4000 59.5000 273.6000 ;
	    RECT 63.6000 271.6000 64.4000 272.4000 ;
	    RECT 65.3000 270.4000 65.9000 281.6000 ;
	    RECT 70.0000 275.6000 70.8000 276.4000 ;
	    RECT 73.2000 275.6000 74.0000 276.4000 ;
	    RECT 66.8000 273.6000 67.6000 274.4000 ;
	    RECT 66.9000 270.4000 67.5000 273.6000 ;
	    RECT 70.1000 272.4000 70.7000 275.6000 ;
	    RECT 70.0000 271.6000 70.8000 272.4000 ;
	    RECT 73.3000 270.4000 73.9000 275.6000 ;
	    RECT 76.5000 272.4000 77.1000 287.6000 ;
	    RECT 79.6000 273.6000 80.4000 274.4000 ;
	    RECT 76.4000 271.6000 77.2000 272.4000 ;
	    RECT 58.8000 269.6000 59.6000 270.4000 ;
	    RECT 60.4000 269.6000 61.2000 270.4000 ;
	    RECT 65.2000 269.6000 66.0000 270.4000 ;
	    RECT 66.8000 269.6000 67.6000 270.4000 ;
	    RECT 71.6000 269.6000 72.4000 270.4000 ;
	    RECT 73.2000 269.6000 74.0000 270.4000 ;
	    RECT 74.8000 269.6000 75.6000 270.4000 ;
	    RECT 60.5000 268.4000 61.1000 269.6000 ;
	    RECT 74.9000 268.4000 75.5000 269.6000 ;
	    RECT 60.4000 267.6000 61.2000 268.4000 ;
	    RECT 62.0000 267.6000 62.8000 268.4000 ;
	    RECT 68.4000 267.6000 69.2000 268.4000 ;
	    RECT 74.8000 267.6000 75.6000 268.4000 ;
	    RECT 57.2000 263.6000 58.0000 264.4000 ;
	    RECT 57.2000 261.6000 58.0000 262.4000 ;
	    RECT 60.4000 261.6000 61.2000 262.4000 ;
	    RECT 44.4000 259.6000 45.2000 260.4000 ;
	    RECT 47.6000 259.6000 48.4000 260.4000 ;
	    RECT 15.6000 246.2000 16.4000 257.8000 ;
	    RECT 23.6000 251.6000 24.4000 252.6000 ;
	    RECT 25.2000 246.2000 26.0000 257.8000 ;
	    RECT 26.8000 253.6000 27.6000 254.4000 ;
	    RECT 28.4000 250.2000 29.2000 255.8000 ;
	    RECT 33.2000 255.6000 34.0000 256.4000 ;
	    RECT 31.6000 253.6000 32.4000 254.4000 ;
	    RECT 30.0000 251.6000 30.8000 252.4000 ;
	    RECT 30.0000 249.6000 30.8000 250.4000 ;
	    RECT 30.1000 246.4000 30.7000 249.6000 ;
	    RECT 30.0000 245.6000 30.8000 246.4000 ;
	    RECT 15.6000 243.6000 16.4000 244.4000 ;
	    RECT 15.7000 234.4000 16.3000 243.6000 ;
	    RECT 15.6000 233.6000 16.4000 234.4000 ;
	    RECT 18.8000 233.6000 19.6000 234.4000 ;
	    RECT 22.0000 231.6000 22.8000 232.4000 ;
	    RECT 10.8000 229.6000 11.6000 230.4000 ;
	    RECT 12.4000 229.6000 13.2000 230.4000 ;
	    RECT 14.0000 229.6000 14.8000 230.4000 ;
	    RECT 18.8000 229.6000 19.6000 230.4000 ;
	    RECT 10.8000 227.6000 11.6000 228.4000 ;
	    RECT 9.2000 217.6000 10.0000 218.4000 ;
	    RECT 10.9000 214.4000 11.5000 227.6000 ;
	    RECT 10.8000 213.6000 11.6000 214.4000 ;
	    RECT 12.5000 212.4000 13.1000 229.6000 ;
	    RECT 17.2000 227.6000 18.0000 228.4000 ;
	    RECT 4.4000 211.6000 5.2000 212.4000 ;
	    RECT 12.4000 211.6000 13.2000 212.4000 ;
	    RECT 14.0000 211.6000 14.8000 212.4000 ;
	    RECT 15.6000 211.6000 16.4000 212.4000 ;
	    RECT 4.4000 191.6000 5.2000 192.4000 ;
	    RECT 4.5000 190.4000 5.1000 191.6000 ;
	    RECT 12.5000 190.4000 13.1000 211.6000 ;
	    RECT 14.1000 210.4000 14.7000 211.6000 ;
	    RECT 15.7000 210.4000 16.3000 211.6000 ;
	    RECT 14.0000 209.6000 14.8000 210.4000 ;
	    RECT 15.6000 209.6000 16.4000 210.4000 ;
	    RECT 17.3000 204.4000 17.9000 227.6000 ;
	    RECT 28.4000 224.2000 29.2000 235.8000 ;
	    RECT 31.7000 230.4000 32.3000 253.6000 ;
	    RECT 33.3000 252.4000 33.9000 255.6000 ;
	    RECT 34.8000 253.6000 35.6000 254.4000 ;
	    RECT 36.4000 253.6000 37.2000 254.4000 ;
	    RECT 34.9000 252.4000 35.5000 253.6000 ;
	    RECT 33.2000 251.6000 34.0000 252.4000 ;
	    RECT 34.8000 251.6000 35.6000 252.4000 ;
	    RECT 36.4000 231.6000 37.2000 232.4000 ;
	    RECT 31.6000 229.6000 32.4000 230.4000 ;
	    RECT 36.5000 230.2000 37.1000 231.6000 ;
	    RECT 36.4000 229.4000 37.2000 230.2000 ;
	    RECT 30.0000 227.6000 30.8000 228.4000 ;
	    RECT 22.0000 206.2000 22.8000 217.8000 ;
	    RECT 30.1000 216.4000 30.7000 227.6000 ;
	    RECT 38.0000 224.2000 38.8000 235.8000 ;
	    RECT 41.2000 226.2000 42.0000 231.8000 ;
	    RECT 44.5000 230.4000 45.1000 259.6000 ;
	    RECT 57.3000 258.4000 57.9000 261.6000 ;
	    RECT 58.8000 259.6000 59.6000 260.4000 ;
	    RECT 57.2000 257.6000 58.0000 258.4000 ;
	    RECT 50.8000 253.6000 51.6000 254.4000 ;
	    RECT 55.6000 253.6000 56.4000 254.4000 ;
	    RECT 54.0000 251.6000 54.8000 252.4000 ;
	    RECT 50.8000 249.6000 51.6000 250.4000 ;
	    RECT 54.1000 248.4000 54.7000 251.6000 ;
	    RECT 55.6000 250.3000 56.4000 250.4000 ;
	    RECT 57.2000 250.3000 58.0000 250.4000 ;
	    RECT 55.6000 249.7000 58.0000 250.3000 ;
	    RECT 55.6000 249.6000 56.4000 249.7000 ;
	    RECT 57.2000 249.6000 58.0000 249.7000 ;
	    RECT 54.0000 247.6000 54.8000 248.4000 ;
	    RECT 47.6000 235.6000 48.4000 236.4000 ;
	    RECT 47.7000 232.4000 48.3000 235.6000 ;
	    RECT 49.2000 233.6000 50.0000 234.4000 ;
	    RECT 49.3000 232.4000 49.9000 233.6000 ;
	    RECT 55.7000 232.4000 56.3000 249.6000 ;
	    RECT 46.0000 231.6000 46.8000 232.4000 ;
	    RECT 47.6000 231.6000 48.4000 232.4000 ;
	    RECT 49.2000 231.6000 50.0000 232.4000 ;
	    RECT 55.6000 231.6000 56.4000 232.4000 ;
	    RECT 44.4000 229.6000 45.2000 230.4000 ;
	    RECT 46.1000 230.3000 46.7000 231.6000 ;
	    RECT 47.6000 230.3000 48.4000 230.4000 ;
	    RECT 46.1000 229.7000 48.4000 230.3000 ;
	    RECT 47.6000 229.6000 48.4000 229.7000 ;
	    RECT 42.8000 227.6000 43.6000 228.4000 ;
	    RECT 30.0000 215.6000 30.8000 216.4000 ;
	    RECT 30.0000 211.6000 30.8000 212.6000 ;
	    RECT 31.6000 206.2000 32.4000 217.8000 ;
	    RECT 33.2000 213.6000 34.0000 214.4000 ;
	    RECT 14.0000 203.6000 14.8000 204.4000 ;
	    RECT 17.2000 203.6000 18.0000 204.4000 ;
	    RECT 14.1000 198.4000 14.7000 203.6000 ;
	    RECT 14.0000 197.6000 14.8000 198.4000 ;
	    RECT 20.4000 191.6000 21.2000 192.4000 ;
	    RECT 4.4000 189.6000 5.2000 190.4000 ;
	    RECT 6.0000 189.6000 6.8000 190.4000 ;
	    RECT 9.2000 189.6000 10.0000 190.4000 ;
	    RECT 12.4000 189.6000 13.2000 190.4000 ;
	    RECT 17.2000 189.6000 18.0000 190.4000 ;
	    RECT 6.1000 186.4000 6.7000 189.6000 ;
	    RECT 9.3000 188.4000 9.9000 189.6000 ;
	    RECT 9.2000 187.6000 10.0000 188.4000 ;
	    RECT 20.4000 187.6000 21.2000 188.4000 ;
	    RECT 6.0000 185.6000 6.8000 186.4000 ;
	    RECT 6.1000 178.4000 6.7000 185.6000 ;
	    RECT 14.0000 183.6000 14.8000 184.4000 ;
	    RECT 26.8000 184.2000 27.6000 195.8000 ;
	    RECT 28.4000 193.6000 29.2000 194.4000 ;
	    RECT 6.0000 177.6000 6.8000 178.4000 ;
	    RECT 14.1000 174.4000 14.7000 183.6000 ;
	    RECT 22.0000 181.6000 22.8000 182.4000 ;
	    RECT 22.1000 178.4000 22.7000 181.6000 ;
	    RECT 28.5000 178.4000 29.1000 193.6000 ;
	    RECT 33.3000 188.4000 33.9000 213.6000 ;
	    RECT 34.8000 210.2000 35.6000 215.8000 ;
	    RECT 39.6000 215.6000 40.4000 216.4000 ;
	    RECT 39.7000 212.4000 40.3000 215.6000 ;
	    RECT 41.2000 213.6000 42.0000 214.4000 ;
	    RECT 36.4000 211.6000 37.2000 212.4000 ;
	    RECT 39.6000 211.6000 40.4000 212.4000 ;
	    RECT 41.2000 211.6000 42.0000 212.4000 ;
	    RECT 36.4000 209.6000 37.2000 210.4000 ;
	    RECT 34.8000 189.4000 35.6000 190.4000 ;
	    RECT 33.2000 187.6000 34.0000 188.4000 ;
	    RECT 36.4000 184.2000 37.2000 195.8000 ;
	    RECT 41.3000 192.4000 41.9000 211.6000 ;
	    RECT 44.5000 198.4000 45.1000 229.6000 ;
	    RECT 47.6000 227.6000 48.4000 228.4000 ;
	    RECT 54.0000 227.6000 54.8000 228.4000 ;
	    RECT 54.1000 216.4000 54.7000 227.6000 ;
	    RECT 47.6000 215.6000 48.4000 216.4000 ;
	    RECT 52.4000 215.6000 53.2000 216.4000 ;
	    RECT 54.0000 215.6000 54.8000 216.4000 ;
	    RECT 52.5000 214.4000 53.1000 215.6000 ;
	    RECT 52.4000 213.6000 53.2000 214.4000 ;
	    RECT 50.8000 211.6000 51.6000 212.4000 ;
	    RECT 54.0000 211.6000 54.8000 212.4000 ;
	    RECT 50.9000 208.4000 51.5000 211.6000 ;
	    RECT 50.8000 207.6000 51.6000 208.4000 ;
	    RECT 46.0000 203.6000 46.8000 204.4000 ;
	    RECT 44.4000 197.6000 45.2000 198.4000 ;
	    RECT 46.1000 196.4000 46.7000 203.6000 ;
	    RECT 54.1000 198.4000 54.7000 211.6000 ;
	    RECT 54.0000 197.6000 54.8000 198.4000 ;
	    RECT 55.7000 196.4000 56.3000 231.6000 ;
	    RECT 58.9000 216.4000 59.5000 259.6000 ;
	    RECT 60.5000 252.4000 61.1000 261.6000 ;
	    RECT 62.1000 258.4000 62.7000 267.6000 ;
	    RECT 68.5000 264.4000 69.1000 267.6000 ;
	    RECT 68.4000 263.6000 69.2000 264.4000 ;
	    RECT 63.6000 259.6000 64.4000 260.4000 ;
	    RECT 62.0000 257.6000 62.8000 258.4000 ;
	    RECT 63.7000 256.4000 64.3000 259.6000 ;
	    RECT 63.6000 255.6000 64.4000 256.4000 ;
	    RECT 63.6000 253.6000 64.4000 254.4000 ;
	    RECT 60.4000 251.6000 61.2000 252.4000 ;
	    RECT 62.0000 251.6000 62.8000 252.4000 ;
	    RECT 62.0000 235.6000 62.8000 236.4000 ;
	    RECT 60.4000 233.6000 61.2000 234.4000 ;
	    RECT 60.5000 230.4000 61.1000 233.6000 ;
	    RECT 60.4000 229.6000 61.2000 230.4000 ;
	    RECT 60.4000 227.6000 61.2000 228.4000 ;
	    RECT 60.5000 226.3000 61.1000 227.6000 ;
	    RECT 60.5000 225.7000 62.7000 226.3000 ;
	    RECT 62.1000 216.4000 62.7000 225.7000 ;
	    RECT 63.7000 218.4000 64.3000 253.6000 ;
	    RECT 66.8000 251.6000 67.6000 252.4000 ;
	    RECT 66.9000 250.4000 67.5000 251.6000 ;
	    RECT 66.8000 249.6000 67.6000 250.4000 ;
	    RECT 68.4000 250.2000 69.2000 255.8000 ;
	    RECT 71.6000 246.2000 72.4000 257.8000 ;
	    RECT 76.5000 256.4000 77.1000 271.6000 ;
	    RECT 81.3000 270.4000 81.9000 291.6000 ;
	    RECT 86.1000 290.4000 86.7000 291.6000 ;
	    RECT 86.0000 289.6000 86.8000 290.4000 ;
	    RECT 89.3000 282.4000 89.9000 305.6000 ;
	    RECT 97.2000 304.2000 98.0000 315.8000 ;
	    RECT 113.2000 311.6000 114.0000 312.4000 ;
	    RECT 114.8000 311.6000 115.6000 312.4000 ;
	    RECT 113.3000 310.4000 113.9000 311.6000 ;
	    RECT 113.2000 309.6000 114.0000 310.4000 ;
	    RECT 114.9000 308.4000 115.5000 311.6000 ;
	    RECT 103.6000 307.6000 104.4000 308.4000 ;
	    RECT 114.8000 307.6000 115.6000 308.4000 ;
	    RECT 100.4000 305.6000 101.2000 306.4000 ;
	    RECT 94.0000 295.6000 94.8000 296.4000 ;
	    RECT 94.1000 292.4000 94.7000 295.6000 ;
	    RECT 95.6000 293.6000 96.4000 294.4000 ;
	    RECT 97.2000 293.6000 98.0000 294.4000 ;
	    RECT 98.8000 293.6000 99.6000 294.4000 ;
	    RECT 97.3000 292.4000 97.9000 293.6000 ;
	    RECT 98.9000 292.4000 99.5000 293.6000 ;
	    RECT 100.5000 292.4000 101.1000 305.6000 ;
	    RECT 103.7000 304.4000 104.3000 307.6000 ;
	    RECT 103.6000 303.6000 104.4000 304.4000 ;
	    RECT 103.6000 295.6000 104.4000 296.4000 ;
	    RECT 103.7000 294.4000 104.3000 295.6000 ;
	    RECT 103.6000 293.6000 104.4000 294.4000 ;
	    RECT 116.5000 292.4000 117.1000 323.6000 ;
	    RECT 118.1000 310.4000 118.7000 325.6000 ;
	    RECT 118.0000 309.6000 118.8000 310.4000 ;
	    RECT 119.7000 308.4000 120.3000 327.6000 ;
	    RECT 122.8000 317.6000 123.6000 318.4000 ;
	    RECT 130.8000 315.6000 131.6000 316.4000 ;
	    RECT 129.2000 311.6000 130.0000 312.4000 ;
	    RECT 122.8000 309.6000 123.6000 310.4000 ;
	    RECT 126.0000 309.6000 126.8000 310.4000 ;
	    RECT 119.6000 307.6000 120.4000 308.4000 ;
	    RECT 121.2000 307.6000 122.0000 308.4000 ;
	    RECT 118.0000 299.6000 118.8000 300.4000 ;
	    RECT 118.1000 292.4000 118.7000 299.6000 ;
	    RECT 119.7000 298.4000 120.3000 307.6000 ;
	    RECT 119.6000 297.6000 120.4000 298.4000 ;
	    RECT 90.8000 291.6000 91.6000 292.4000 ;
	    RECT 94.0000 291.6000 94.8000 292.4000 ;
	    RECT 97.2000 291.6000 98.0000 292.4000 ;
	    RECT 98.8000 291.6000 99.6000 292.4000 ;
	    RECT 100.4000 291.6000 101.2000 292.4000 ;
	    RECT 102.0000 291.6000 102.8000 292.4000 ;
	    RECT 116.4000 291.6000 117.2000 292.4000 ;
	    RECT 118.0000 291.6000 118.8000 292.4000 ;
	    RECT 90.9000 290.4000 91.5000 291.6000 ;
	    RECT 100.5000 290.4000 101.1000 291.6000 ;
	    RECT 90.8000 289.6000 91.6000 290.4000 ;
	    RECT 97.2000 289.6000 98.0000 290.4000 ;
	    RECT 100.4000 289.6000 101.2000 290.4000 ;
	    RECT 89.2000 281.6000 90.0000 282.4000 ;
	    RECT 86.0000 277.6000 86.8000 278.4000 ;
	    RECT 84.4000 275.6000 85.2000 276.4000 ;
	    RECT 82.8000 271.6000 83.6000 272.4000 ;
	    RECT 78.0000 269.6000 78.8000 270.4000 ;
	    RECT 81.2000 269.6000 82.0000 270.4000 ;
	    RECT 82.8000 270.3000 83.6000 270.4000 ;
	    RECT 84.5000 270.3000 85.1000 275.6000 ;
	    RECT 86.1000 270.4000 86.7000 277.6000 ;
	    RECT 90.9000 274.4000 91.5000 289.6000 ;
	    RECT 92.4000 279.6000 93.2000 280.4000 ;
	    RECT 87.6000 273.6000 88.4000 274.4000 ;
	    RECT 90.8000 273.6000 91.6000 274.4000 ;
	    RECT 87.7000 270.4000 88.3000 273.6000 ;
	    RECT 89.2000 271.6000 90.0000 272.4000 ;
	    RECT 90.8000 271.6000 91.6000 272.4000 ;
	    RECT 82.8000 269.7000 85.1000 270.3000 ;
	    RECT 82.8000 269.6000 83.6000 269.7000 ;
	    RECT 86.0000 269.6000 86.8000 270.4000 ;
	    RECT 87.6000 269.6000 88.4000 270.4000 ;
	    RECT 78.1000 264.3000 78.7000 269.6000 ;
	    RECT 79.6000 267.6000 80.4000 268.4000 ;
	    RECT 81.2000 267.6000 82.0000 268.4000 ;
	    RECT 87.6000 267.6000 88.4000 268.4000 ;
	    RECT 79.7000 266.3000 80.3000 267.6000 ;
	    RECT 82.8000 266.3000 83.6000 266.4000 ;
	    RECT 79.7000 265.7000 83.6000 266.3000 ;
	    RECT 82.8000 265.6000 83.6000 265.7000 ;
	    RECT 90.9000 264.3000 91.5000 271.6000 ;
	    RECT 92.5000 270.4000 93.1000 279.6000 ;
	    RECT 92.4000 269.6000 93.2000 270.4000 ;
	    RECT 92.4000 268.3000 93.2000 268.4000 ;
	    RECT 94.0000 268.3000 94.8000 268.4000 ;
	    RECT 92.4000 267.7000 94.8000 268.3000 ;
	    RECT 92.4000 267.6000 93.2000 267.7000 ;
	    RECT 94.0000 267.6000 94.8000 267.7000 ;
	    RECT 78.1000 263.7000 91.5000 264.3000 ;
	    RECT 73.2000 255.6000 74.0000 256.4000 ;
	    RECT 76.4000 255.6000 77.2000 256.4000 ;
	    RECT 76.4000 253.6000 77.2000 254.4000 ;
	    RECT 76.5000 252.4000 77.1000 253.6000 ;
	    RECT 76.4000 251.6000 77.2000 252.4000 ;
	    RECT 78.0000 251.6000 78.8000 252.4000 ;
	    RECT 66.8000 224.2000 67.6000 235.8000 ;
	    RECT 68.4000 229.6000 69.2000 230.4000 ;
	    RECT 74.8000 229.4000 75.6000 230.4000 ;
	    RECT 68.4000 225.6000 69.2000 226.4000 ;
	    RECT 68.5000 218.4000 69.1000 225.6000 ;
	    RECT 76.4000 224.2000 77.2000 235.8000 ;
	    RECT 63.6000 217.6000 64.4000 218.4000 ;
	    RECT 68.4000 217.6000 69.2000 218.4000 ;
	    RECT 58.8000 215.6000 59.6000 216.4000 ;
	    RECT 62.0000 215.6000 62.8000 216.4000 ;
	    RECT 57.2000 213.6000 58.0000 214.4000 ;
	    RECT 58.9000 200.4000 59.5000 215.6000 ;
	    RECT 62.0000 213.6000 62.8000 214.4000 ;
	    RECT 62.1000 212.4000 62.7000 213.6000 ;
	    RECT 62.0000 211.6000 62.8000 212.4000 ;
	    RECT 71.6000 211.6000 72.4000 212.4000 ;
	    RECT 73.2000 210.2000 74.0000 215.8000 ;
	    RECT 62.0000 205.6000 62.8000 206.4000 ;
	    RECT 76.4000 206.2000 77.2000 217.8000 ;
	    RECT 78.1000 216.4000 78.7000 251.6000 ;
	    RECT 81.2000 246.2000 82.0000 257.8000 ;
	    RECT 86.0000 257.6000 86.8000 258.4000 ;
	    RECT 86.1000 256.3000 86.7000 257.6000 ;
	    RECT 87.6000 256.3000 88.4000 256.4000 ;
	    RECT 86.1000 255.7000 88.4000 256.3000 ;
	    RECT 87.6000 255.6000 88.4000 255.7000 ;
	    RECT 87.7000 254.4000 88.3000 255.6000 ;
	    RECT 87.6000 253.6000 88.4000 254.4000 ;
	    RECT 90.8000 253.6000 91.6000 254.4000 ;
	    RECT 90.8000 251.6000 91.6000 252.4000 ;
	    RECT 90.9000 250.4000 91.5000 251.6000 ;
	    RECT 90.8000 249.6000 91.6000 250.4000 ;
	    RECT 86.0000 243.6000 86.8000 244.4000 ;
	    RECT 79.6000 226.2000 80.4000 231.8000 ;
	    RECT 81.2000 231.6000 82.0000 232.4000 ;
	    RECT 81.3000 228.4000 81.9000 231.6000 ;
	    RECT 82.8000 229.6000 83.6000 230.4000 ;
	    RECT 86.1000 228.4000 86.7000 243.6000 ;
	    RECT 87.6000 231.6000 88.4000 232.4000 ;
	    RECT 90.8000 231.6000 91.6000 232.4000 ;
	    RECT 81.2000 227.6000 82.0000 228.4000 ;
	    RECT 86.0000 227.6000 86.8000 228.4000 ;
	    RECT 87.7000 226.4000 88.3000 231.6000 ;
	    RECT 90.9000 230.4000 91.5000 231.6000 ;
	    RECT 90.8000 229.6000 91.6000 230.4000 ;
	    RECT 92.5000 228.4000 93.1000 267.6000 ;
	    RECT 95.6000 266.2000 96.4000 271.8000 ;
	    RECT 97.3000 256.3000 97.9000 289.6000 ;
	    RECT 113.2000 285.6000 114.0000 286.4000 ;
	    RECT 114.8000 285.6000 115.6000 286.4000 ;
	    RECT 102.0000 281.6000 102.8000 282.4000 ;
	    RECT 98.8000 264.2000 99.6000 275.8000 ;
	    RECT 100.4000 269.4000 101.2000 270.4000 ;
	    RECT 102.1000 268.4000 102.7000 281.6000 ;
	    RECT 111.6000 279.6000 112.4000 280.4000 ;
	    RECT 103.6000 269.6000 104.4000 270.4000 ;
	    RECT 102.0000 267.6000 102.8000 268.4000 ;
	    RECT 103.7000 266.4000 104.3000 269.6000 ;
	    RECT 103.6000 265.6000 104.4000 266.4000 ;
	    RECT 108.4000 264.2000 109.2000 275.8000 ;
	    RECT 111.7000 268.4000 112.3000 279.6000 ;
	    RECT 113.3000 278.4000 113.9000 285.6000 ;
	    RECT 114.9000 278.4000 115.5000 285.6000 ;
	    RECT 119.6000 283.6000 120.4000 284.4000 ;
	    RECT 113.2000 277.6000 114.0000 278.4000 ;
	    RECT 114.8000 277.6000 115.6000 278.4000 ;
	    RECT 114.8000 273.6000 115.6000 274.4000 ;
	    RECT 111.6000 267.6000 112.4000 268.4000 ;
	    RECT 97.3000 255.7000 99.5000 256.3000 ;
	    RECT 97.2000 253.6000 98.0000 254.4000 ;
	    RECT 95.6000 251.6000 96.4000 252.4000 ;
	    RECT 97.3000 238.3000 97.9000 253.6000 ;
	    RECT 98.9000 252.4000 99.5000 255.7000 ;
	    RECT 100.4000 255.6000 101.2000 256.4000 ;
	    RECT 100.5000 252.4000 101.1000 255.6000 ;
	    RECT 114.9000 254.4000 115.5000 273.6000 ;
	    RECT 119.7000 266.4000 120.3000 283.6000 ;
	    RECT 121.3000 274.4000 121.9000 307.6000 ;
	    RECT 122.9000 298.4000 123.5000 309.6000 ;
	    RECT 129.3000 308.4000 129.9000 311.6000 ;
	    RECT 129.2000 307.6000 130.0000 308.4000 ;
	    RECT 122.8000 297.6000 123.6000 298.4000 ;
	    RECT 130.9000 296.4000 131.5000 315.6000 ;
	    RECT 132.4000 309.6000 133.2000 310.4000 ;
	    RECT 132.5000 306.4000 133.1000 309.6000 ;
	    RECT 134.1000 308.4000 134.7000 329.6000 ;
	    RECT 135.6000 326.2000 136.4000 337.8000 ;
	    RECT 137.2000 331.6000 138.0000 332.4000 ;
	    RECT 143.6000 331.6000 144.4000 332.6000 ;
	    RECT 137.3000 330.4000 137.9000 331.6000 ;
	    RECT 137.2000 329.6000 138.0000 330.4000 ;
	    RECT 145.2000 326.2000 146.0000 337.8000 ;
	    RECT 150.0000 337.6000 150.8000 338.4000 ;
	    RECT 148.4000 330.2000 149.2000 335.8000 ;
	    RECT 150.1000 334.4000 150.7000 337.6000 ;
	    RECT 150.0000 333.6000 150.8000 334.4000 ;
	    RECT 153.2000 333.6000 154.0000 334.4000 ;
	    RECT 159.6000 333.6000 160.4000 334.4000 ;
	    RECT 153.3000 332.4000 153.9000 333.6000 ;
	    RECT 153.2000 331.6000 154.0000 332.4000 ;
	    RECT 158.0000 331.6000 158.8000 332.4000 ;
	    RECT 153.2000 329.6000 154.0000 330.4000 ;
	    RECT 156.4000 329.6000 157.2000 330.4000 ;
	    RECT 153.3000 322.4000 153.9000 329.6000 ;
	    RECT 153.2000 321.6000 154.0000 322.4000 ;
	    RECT 137.2000 309.6000 138.0000 310.4000 ;
	    RECT 142.0000 309.6000 142.8000 310.4000 ;
	    RECT 143.6000 309.6000 144.4000 310.4000 ;
	    RECT 146.8000 309.6000 147.6000 310.4000 ;
	    RECT 134.0000 307.6000 134.8000 308.4000 ;
	    RECT 132.4000 305.6000 133.2000 306.4000 ;
	    RECT 124.4000 295.6000 125.2000 296.4000 ;
	    RECT 130.8000 295.6000 131.6000 296.4000 ;
	    RECT 124.5000 292.4000 125.1000 295.6000 ;
	    RECT 126.0000 293.6000 126.8000 294.4000 ;
	    RECT 122.8000 291.6000 123.6000 292.4000 ;
	    RECT 124.4000 291.6000 125.2000 292.4000 ;
	    RECT 126.0000 291.6000 126.8000 292.4000 ;
	    RECT 121.2000 273.6000 122.0000 274.4000 ;
	    RECT 124.5000 268.4000 125.1000 291.6000 ;
	    RECT 132.5000 280.4000 133.1000 305.6000 ;
	    RECT 137.3000 304.4000 137.9000 309.6000 ;
	    RECT 142.1000 306.4000 142.7000 309.6000 ;
	    RECT 142.0000 305.6000 142.8000 306.4000 ;
	    RECT 137.2000 303.6000 138.0000 304.4000 ;
	    RECT 138.8000 303.6000 139.6000 304.4000 ;
	    RECT 135.6000 295.6000 136.4000 296.4000 ;
	    RECT 134.0000 293.6000 134.8000 294.4000 ;
	    RECT 134.1000 292.4000 134.7000 293.6000 ;
	    RECT 135.7000 292.4000 136.3000 295.6000 ;
	    RECT 137.3000 292.4000 137.9000 303.6000 ;
	    RECT 138.9000 298.4000 139.5000 303.6000 ;
	    RECT 138.8000 297.6000 139.6000 298.4000 ;
	    RECT 140.4000 297.6000 141.2000 298.4000 ;
	    RECT 142.1000 292.4000 142.7000 305.6000 ;
	    RECT 143.7000 292.4000 144.3000 309.6000 ;
	    RECT 148.4000 307.6000 149.2000 308.4000 ;
	    RECT 148.5000 306.4000 149.1000 307.6000 ;
	    RECT 148.4000 305.6000 149.2000 306.4000 ;
	    RECT 150.0000 303.6000 150.8000 304.4000 ;
	    RECT 154.8000 304.2000 155.6000 315.8000 ;
	    RECT 156.5000 310.4000 157.1000 329.6000 ;
	    RECT 158.1000 322.4000 158.7000 331.6000 ;
	    RECT 161.2000 328.3000 162.0000 328.4000 ;
	    RECT 159.7000 327.7000 162.0000 328.3000 ;
	    RECT 158.0000 321.6000 158.8000 322.4000 ;
	    RECT 156.4000 309.6000 157.2000 310.4000 ;
	    RECT 150.1000 300.4000 150.7000 303.6000 ;
	    RECT 150.0000 299.6000 150.8000 300.4000 ;
	    RECT 146.8000 297.6000 147.6000 298.4000 ;
	    RECT 151.6000 297.6000 152.4000 298.4000 ;
	    RECT 145.2000 293.6000 146.0000 294.4000 ;
	    RECT 134.0000 291.6000 134.8000 292.4000 ;
	    RECT 135.6000 291.6000 136.4000 292.4000 ;
	    RECT 137.2000 291.6000 138.0000 292.4000 ;
	    RECT 142.0000 291.6000 142.8000 292.4000 ;
	    RECT 143.6000 291.6000 144.4000 292.4000 ;
	    RECT 134.0000 283.6000 134.8000 284.4000 ;
	    RECT 138.8000 283.6000 139.6000 284.4000 ;
	    RECT 129.2000 279.6000 130.0000 280.4000 ;
	    RECT 132.4000 279.6000 133.2000 280.4000 ;
	    RECT 129.3000 278.4000 129.9000 279.6000 ;
	    RECT 126.0000 277.6000 126.8000 278.4000 ;
	    RECT 127.6000 277.6000 128.4000 278.4000 ;
	    RECT 129.2000 277.6000 130.0000 278.4000 ;
	    RECT 126.1000 272.4000 126.7000 277.6000 ;
	    RECT 126.0000 271.6000 126.8000 272.4000 ;
	    RECT 127.7000 268.4000 128.3000 277.6000 ;
	    RECT 134.1000 270.4000 134.7000 283.6000 ;
	    RECT 138.9000 270.4000 139.5000 283.6000 ;
	    RECT 145.3000 278.4000 145.9000 293.6000 ;
	    RECT 146.9000 292.4000 147.5000 297.6000 ;
	    RECT 151.7000 294.4000 152.3000 297.6000 ;
	    RECT 153.2000 295.6000 154.0000 296.4000 ;
	    RECT 153.3000 294.4000 153.9000 295.6000 ;
	    RECT 151.6000 293.6000 152.4000 294.4000 ;
	    RECT 153.2000 293.6000 154.0000 294.4000 ;
	    RECT 146.8000 291.6000 147.6000 292.4000 ;
	    RECT 150.0000 291.6000 150.8000 292.4000 ;
	    RECT 154.8000 291.6000 155.6000 292.4000 ;
	    RECT 150.1000 290.4000 150.7000 291.6000 ;
	    RECT 150.0000 289.6000 150.8000 290.4000 ;
	    RECT 146.8000 283.6000 147.6000 284.4000 ;
	    RECT 145.2000 277.6000 146.0000 278.4000 ;
	    RECT 145.2000 273.6000 146.0000 274.4000 ;
	    RECT 142.0000 271.6000 142.8000 272.4000 ;
	    RECT 143.6000 271.6000 144.4000 272.4000 ;
	    RECT 143.7000 270.4000 144.3000 271.6000 ;
	    RECT 129.2000 269.6000 130.0000 270.4000 ;
	    RECT 134.0000 269.6000 134.8000 270.4000 ;
	    RECT 138.8000 269.6000 139.6000 270.4000 ;
	    RECT 143.6000 269.6000 144.4000 270.4000 ;
	    RECT 121.2000 267.6000 122.0000 268.4000 ;
	    RECT 122.8000 267.6000 123.6000 268.4000 ;
	    RECT 124.4000 267.6000 125.2000 268.4000 ;
	    RECT 127.6000 267.6000 128.4000 268.4000 ;
	    RECT 119.6000 265.6000 120.4000 266.4000 ;
	    RECT 122.9000 254.4000 123.5000 267.6000 ;
	    RECT 129.3000 266.4000 129.9000 269.6000 ;
	    RECT 134.0000 267.6000 134.8000 268.4000 ;
	    RECT 145.3000 268.3000 145.9000 273.6000 ;
	    RECT 146.9000 272.4000 147.5000 283.6000 ;
	    RECT 150.0000 279.6000 150.8000 280.4000 ;
	    RECT 150.1000 278.4000 150.7000 279.6000 ;
	    RECT 150.0000 277.6000 150.8000 278.4000 ;
	    RECT 150.0000 275.6000 150.8000 276.4000 ;
	    RECT 146.8000 271.6000 147.6000 272.4000 ;
	    RECT 148.4000 271.6000 149.2000 272.4000 ;
	    RECT 148.5000 270.4000 149.1000 271.6000 ;
	    RECT 146.8000 269.6000 147.6000 270.4000 ;
	    RECT 148.4000 269.6000 149.2000 270.4000 ;
	    RECT 150.1000 268.4000 150.7000 275.6000 ;
	    RECT 143.7000 267.7000 145.9000 268.3000 ;
	    RECT 134.1000 266.4000 134.7000 267.6000 ;
	    RECT 129.2000 265.6000 130.0000 266.4000 ;
	    RECT 130.8000 265.6000 131.6000 266.4000 ;
	    RECT 134.0000 265.6000 134.8000 266.4000 ;
	    RECT 135.6000 265.6000 136.4000 266.4000 ;
	    RECT 140.4000 265.6000 141.2000 266.4000 ;
	    RECT 126.0000 264.3000 126.8000 264.4000 ;
	    RECT 130.9000 264.3000 131.5000 265.6000 ;
	    RECT 126.0000 263.7000 131.5000 264.3000 ;
	    RECT 126.0000 263.6000 126.8000 263.7000 ;
	    RECT 137.2000 263.6000 138.0000 264.4000 ;
	    RECT 126.0000 261.6000 126.8000 262.4000 ;
	    RECT 135.6000 261.6000 136.4000 262.4000 ;
	    RECT 126.1000 258.4000 126.7000 261.6000 ;
	    RECT 132.4000 259.6000 133.2000 260.4000 ;
	    RECT 124.4000 257.6000 125.2000 258.4000 ;
	    RECT 126.0000 257.6000 126.8000 258.4000 ;
	    RECT 113.2000 253.6000 114.0000 254.4000 ;
	    RECT 114.8000 253.6000 115.6000 254.4000 ;
	    RECT 116.4000 253.6000 117.2000 254.4000 ;
	    RECT 121.2000 253.6000 122.0000 254.4000 ;
	    RECT 122.8000 253.6000 123.6000 254.4000 ;
	    RECT 116.5000 252.4000 117.1000 253.6000 ;
	    RECT 98.8000 251.6000 99.6000 252.4000 ;
	    RECT 100.4000 251.6000 101.2000 252.4000 ;
	    RECT 113.2000 251.6000 114.0000 252.4000 ;
	    RECT 116.4000 251.6000 117.2000 252.4000 ;
	    RECT 119.6000 251.6000 120.4000 252.4000 ;
	    RECT 119.7000 250.4000 120.3000 251.6000 ;
	    RECT 111.6000 249.6000 112.4000 250.4000 ;
	    RECT 119.6000 249.6000 120.4000 250.4000 ;
	    RECT 111.7000 240.4000 112.3000 249.6000 ;
	    RECT 121.3000 248.4000 121.9000 253.6000 ;
	    RECT 122.9000 252.4000 123.5000 253.6000 ;
	    RECT 124.5000 252.4000 125.1000 257.6000 ;
	    RECT 132.5000 256.4000 133.1000 259.6000 ;
	    RECT 132.4000 255.6000 133.2000 256.4000 ;
	    RECT 135.7000 252.4000 136.3000 261.6000 ;
	    RECT 140.4000 259.6000 141.2000 260.4000 ;
	    RECT 140.5000 256.4000 141.1000 259.6000 ;
	    RECT 140.4000 255.6000 141.2000 256.4000 ;
	    RECT 138.8000 253.6000 139.6000 254.4000 ;
	    RECT 122.8000 251.6000 123.6000 252.4000 ;
	    RECT 124.4000 251.6000 125.2000 252.4000 ;
	    RECT 129.2000 251.6000 130.0000 252.4000 ;
	    RECT 135.6000 251.6000 136.4000 252.4000 ;
	    RECT 137.2000 251.6000 138.0000 252.4000 ;
	    RECT 134.0000 249.6000 134.8000 250.4000 ;
	    RECT 137.3000 248.4000 137.9000 251.6000 ;
	    RECT 116.4000 247.6000 117.2000 248.4000 ;
	    RECT 121.2000 247.6000 122.0000 248.4000 ;
	    RECT 137.2000 247.6000 138.0000 248.4000 ;
	    RECT 113.2000 245.6000 114.0000 246.4000 ;
	    RECT 111.6000 239.6000 112.4000 240.4000 ;
	    RECT 98.8000 238.3000 99.6000 238.4000 ;
	    RECT 97.3000 237.7000 99.6000 238.3000 ;
	    RECT 98.8000 237.6000 99.6000 237.7000 ;
	    RECT 94.0000 231.6000 94.8000 232.4000 ;
	    RECT 92.4000 227.6000 93.2000 228.4000 ;
	    RECT 87.6000 225.6000 88.4000 226.4000 ;
	    RECT 92.4000 225.6000 93.2000 226.4000 ;
	    RECT 78.0000 215.6000 78.8000 216.4000 ;
	    RECT 79.6000 213.6000 80.4000 214.4000 ;
	    RECT 81.2000 213.6000 82.0000 214.4000 ;
	    RECT 58.8000 199.6000 59.6000 200.4000 ;
	    RECT 46.0000 195.6000 46.8000 196.4000 ;
	    RECT 52.4000 195.6000 53.2000 196.4000 ;
	    RECT 55.6000 195.6000 56.4000 196.4000 ;
	    RECT 58.8000 195.6000 59.6000 196.4000 ;
	    RECT 52.5000 192.4000 53.1000 195.6000 ;
	    RECT 58.9000 192.4000 59.5000 195.6000 ;
	    RECT 38.0000 187.6000 38.8000 188.4000 ;
	    RECT 22.0000 177.6000 22.8000 178.4000 ;
	    RECT 28.4000 177.6000 29.2000 178.4000 ;
	    RECT 34.8000 177.6000 35.6000 178.4000 ;
	    RECT 34.9000 174.4000 35.5000 177.6000 ;
	    RECT 14.0000 173.6000 14.8000 174.4000 ;
	    RECT 34.8000 173.6000 35.6000 174.4000 ;
	    RECT 12.4000 171.6000 13.2000 172.4000 ;
	    RECT 20.4000 171.6000 21.2000 172.4000 ;
	    RECT 31.6000 171.6000 32.4000 172.4000 ;
	    RECT 33.2000 171.6000 34.0000 172.4000 ;
	    RECT 17.2000 169.6000 18.0000 170.4000 ;
	    RECT 28.4000 169.6000 29.2000 170.4000 ;
	    RECT 30.0000 169.6000 30.8000 170.4000 ;
	    RECT 6.0000 163.6000 6.8000 164.4000 ;
	    RECT 4.4000 151.6000 5.2000 152.4000 ;
	    RECT 4.5000 150.4000 5.1000 151.6000 ;
	    RECT 6.1000 150.4000 6.7000 163.6000 ;
	    RECT 17.3000 158.4000 17.9000 169.6000 ;
	    RECT 28.5000 168.4000 29.1000 169.6000 ;
	    RECT 18.8000 167.6000 19.6000 168.4000 ;
	    RECT 28.4000 167.6000 29.2000 168.4000 ;
	    RECT 17.2000 157.6000 18.0000 158.4000 ;
	    RECT 20.4000 151.6000 21.2000 152.4000 ;
	    RECT 4.4000 149.6000 5.2000 150.4000 ;
	    RECT 6.0000 149.6000 6.8000 150.4000 ;
	    RECT 9.2000 149.6000 10.0000 150.4000 ;
	    RECT 17.2000 149.6000 18.0000 150.4000 ;
	    RECT 9.3000 148.4000 9.9000 149.6000 ;
	    RECT 9.2000 147.6000 10.0000 148.4000 ;
	    RECT 14.0000 143.6000 14.8000 144.4000 ;
	    RECT 26.8000 144.2000 27.6000 155.8000 ;
	    RECT 31.7000 150.4000 32.3000 171.6000 ;
	    RECT 36.4000 170.2000 37.2000 175.8000 ;
	    RECT 38.1000 174.4000 38.7000 187.6000 ;
	    RECT 39.6000 186.2000 40.4000 191.8000 ;
	    RECT 41.2000 191.6000 42.0000 192.4000 ;
	    RECT 46.0000 191.6000 46.8000 192.4000 ;
	    RECT 52.4000 191.6000 53.2000 192.4000 ;
	    RECT 58.8000 191.6000 59.6000 192.4000 ;
	    RECT 41.2000 189.6000 42.0000 190.4000 ;
	    RECT 41.3000 186.4000 41.9000 189.6000 ;
	    RECT 46.1000 188.4000 46.7000 191.6000 ;
	    RECT 62.1000 190.4000 62.7000 205.6000 ;
	    RECT 68.4000 195.6000 69.2000 196.4000 ;
	    RECT 68.5000 190.4000 69.1000 195.6000 ;
	    RECT 47.6000 189.6000 48.4000 190.4000 ;
	    RECT 50.8000 189.6000 51.6000 190.4000 ;
	    RECT 55.6000 189.6000 56.4000 190.4000 ;
	    RECT 62.0000 189.6000 62.8000 190.4000 ;
	    RECT 63.6000 189.6000 64.4000 190.4000 ;
	    RECT 68.4000 189.6000 69.2000 190.4000 ;
	    RECT 50.9000 188.4000 51.5000 189.6000 ;
	    RECT 46.0000 187.6000 46.8000 188.4000 ;
	    RECT 50.8000 187.6000 51.6000 188.4000 ;
	    RECT 55.7000 186.4000 56.3000 189.6000 ;
	    RECT 57.2000 187.6000 58.0000 188.4000 ;
	    RECT 63.6000 187.6000 64.4000 188.4000 ;
	    RECT 68.4000 187.6000 69.2000 188.4000 ;
	    RECT 41.2000 185.6000 42.0000 186.4000 ;
	    RECT 46.0000 185.6000 46.8000 186.4000 ;
	    RECT 55.6000 185.6000 56.4000 186.4000 ;
	    RECT 65.2000 185.6000 66.0000 186.4000 ;
	    RECT 38.0000 173.6000 38.8000 174.4000 ;
	    RECT 31.6000 149.6000 32.4000 150.4000 ;
	    RECT 33.2000 149.6000 34.0000 150.4000 ;
	    RECT 28.4000 147.6000 29.2000 148.4000 ;
	    RECT 4.4000 137.6000 5.2000 138.4000 ;
	    RECT 10.8000 137.6000 11.6000 138.4000 ;
	    RECT 4.5000 132.4000 5.1000 137.6000 ;
	    RECT 14.1000 134.4000 14.7000 143.6000 ;
	    RECT 28.5000 138.3000 29.1000 147.6000 ;
	    RECT 14.0000 133.6000 14.8000 134.4000 ;
	    RECT 4.4000 131.6000 5.2000 132.4000 ;
	    RECT 9.2000 131.6000 10.0000 132.4000 ;
	    RECT 9.3000 130.4000 9.9000 131.6000 ;
	    RECT 9.2000 129.6000 10.0000 130.4000 ;
	    RECT 15.6000 126.2000 16.4000 137.8000 ;
	    RECT 23.6000 135.6000 24.4000 136.4000 ;
	    RECT 18.8000 133.6000 19.6000 134.4000 ;
	    RECT 4.4000 111.6000 5.2000 112.4000 ;
	    RECT 4.5000 110.4000 5.1000 111.6000 ;
	    RECT 4.4000 109.6000 5.2000 110.4000 ;
	    RECT 6.0000 104.3000 6.8000 104.4000 ;
	    RECT 4.5000 103.7000 6.8000 104.3000 ;
	    RECT 10.8000 104.2000 11.6000 115.8000 ;
	    RECT 17.2000 109.6000 18.0000 110.4000 ;
	    RECT 4.5000 92.4000 5.1000 103.7000 ;
	    RECT 6.0000 103.6000 6.8000 103.7000 ;
	    RECT 17.3000 98.4000 17.9000 109.6000 ;
	    RECT 18.9000 108.4000 19.5000 133.6000 ;
	    RECT 23.7000 132.6000 24.3000 135.6000 ;
	    RECT 23.6000 131.8000 24.4000 132.6000 ;
	    RECT 25.2000 126.2000 26.0000 137.8000 ;
	    RECT 26.9000 137.7000 29.1000 138.3000 ;
	    RECT 26.9000 134.4000 27.5000 137.7000 ;
	    RECT 30.0000 137.6000 30.8000 138.4000 ;
	    RECT 26.8000 133.6000 27.6000 134.4000 ;
	    RECT 28.4000 130.2000 29.2000 135.8000 ;
	    RECT 30.1000 130.4000 30.7000 137.6000 ;
	    RECT 33.3000 132.4000 33.9000 149.6000 ;
	    RECT 36.4000 144.2000 37.2000 155.8000 ;
	    RECT 38.1000 148.4000 38.7000 173.6000 ;
	    RECT 39.6000 166.2000 40.4000 177.8000 ;
	    RECT 42.8000 171.6000 43.6000 172.4000 ;
	    RECT 42.9000 152.4000 43.5000 171.6000 ;
	    RECT 38.0000 147.6000 38.8000 148.4000 ;
	    RECT 39.6000 146.2000 40.4000 151.8000 ;
	    RECT 41.2000 146.2000 42.0000 151.8000 ;
	    RECT 42.8000 151.6000 43.6000 152.4000 ;
	    RECT 44.4000 144.2000 45.2000 155.8000 ;
	    RECT 34.8000 133.6000 35.6000 134.4000 ;
	    RECT 33.2000 131.6000 34.0000 132.4000 ;
	    RECT 30.0000 129.6000 30.8000 130.4000 ;
	    RECT 33.3000 130.3000 33.9000 131.6000 ;
	    RECT 31.7000 129.7000 33.9000 130.3000 ;
	    RECT 18.8000 107.6000 19.6000 108.4000 ;
	    RECT 20.4000 104.2000 21.2000 115.8000 ;
	    RECT 22.0000 115.6000 22.8000 116.4000 ;
	    RECT 17.2000 97.6000 18.0000 98.4000 ;
	    RECT 22.1000 94.4000 22.7000 115.6000 ;
	    RECT 26.8000 113.6000 27.6000 114.4000 ;
	    RECT 23.6000 106.2000 24.4000 111.8000 ;
	    RECT 30.0000 111.6000 30.8000 112.4000 ;
	    RECT 31.7000 110.4000 32.3000 129.7000 ;
	    RECT 33.2000 127.6000 34.0000 128.4000 ;
	    RECT 33.2000 125.6000 34.0000 126.4000 ;
	    RECT 33.3000 118.4000 33.9000 125.6000 ;
	    RECT 33.2000 117.6000 34.0000 118.4000 ;
	    RECT 26.8000 109.6000 27.6000 110.4000 ;
	    RECT 31.6000 109.6000 32.4000 110.4000 ;
	    RECT 25.2000 107.6000 26.0000 108.4000 ;
	    RECT 15.6000 93.6000 16.4000 94.4000 ;
	    RECT 22.0000 93.6000 22.8000 94.4000 ;
	    RECT 23.6000 94.3000 24.4000 94.4000 ;
	    RECT 25.3000 94.3000 25.9000 107.6000 ;
	    RECT 23.6000 93.7000 25.9000 94.3000 ;
	    RECT 23.6000 93.6000 24.4000 93.7000 ;
	    RECT 4.4000 91.6000 5.2000 92.4000 ;
	    RECT 9.2000 91.6000 10.0000 92.4000 ;
	    RECT 10.8000 91.6000 11.6000 92.4000 ;
	    RECT 14.0000 91.6000 14.8000 92.4000 ;
	    RECT 22.0000 91.6000 22.8000 92.4000 ;
	    RECT 25.2000 92.3000 26.0000 92.4000 ;
	    RECT 26.9000 92.3000 27.5000 109.6000 ;
	    RECT 34.9000 108.4000 35.5000 133.6000 ;
	    RECT 41.2000 131.6000 42.0000 132.4000 ;
	    RECT 41.2000 129.6000 42.0000 130.4000 ;
	    RECT 36.4000 113.6000 37.2000 114.4000 ;
	    RECT 36.5000 112.4000 37.1000 113.6000 ;
	    RECT 36.4000 111.6000 37.2000 112.4000 ;
	    RECT 34.8000 107.6000 35.6000 108.4000 ;
	    RECT 34.9000 106.4000 35.5000 107.6000 ;
	    RECT 34.8000 105.6000 35.6000 106.4000 ;
	    RECT 33.2000 103.6000 34.0000 104.4000 ;
	    RECT 41.2000 104.2000 42.0000 115.8000 ;
	    RECT 25.2000 91.7000 27.5000 92.3000 ;
	    RECT 25.2000 91.6000 26.0000 91.7000 ;
	    RECT 28.4000 91.6000 29.2000 92.4000 ;
	    RECT 9.3000 90.4000 9.9000 91.6000 ;
	    RECT 10.9000 90.4000 11.5000 91.6000 ;
	    RECT 9.2000 89.6000 10.0000 90.4000 ;
	    RECT 10.8000 89.6000 11.6000 90.4000 ;
	    RECT 17.2000 89.6000 18.0000 90.4000 ;
	    RECT 17.3000 88.4000 17.9000 89.6000 ;
	    RECT 14.0000 87.6000 14.8000 88.4000 ;
	    RECT 17.2000 87.6000 18.0000 88.4000 ;
	    RECT 22.1000 76.4000 22.7000 91.6000 ;
	    RECT 28.4000 89.6000 29.2000 90.4000 ;
	    RECT 33.3000 84.4000 33.9000 103.6000 ;
	    RECT 34.8000 86.2000 35.6000 97.8000 ;
	    RECT 42.8000 93.6000 43.6000 94.4000 ;
	    RECT 42.9000 92.6000 43.5000 93.6000 ;
	    RECT 36.4000 91.6000 37.2000 92.4000 ;
	    RECT 42.8000 91.8000 43.6000 92.6000 ;
	    RECT 33.2000 83.6000 34.0000 84.4000 ;
	    RECT 4.4000 73.6000 5.2000 74.4000 ;
	    RECT 15.6000 73.6000 16.4000 74.4000 ;
	    RECT 4.5000 70.4000 5.1000 73.6000 ;
	    RECT 4.4000 69.6000 5.2000 70.4000 ;
	    RECT 9.2000 63.6000 10.0000 64.4000 ;
	    RECT 14.0000 63.6000 14.8000 64.4000 ;
	    RECT 20.4000 64.2000 21.2000 75.8000 ;
	    RECT 22.0000 75.6000 22.8000 76.4000 ;
	    RECT 28.4000 69.4000 29.2000 70.4000 ;
	    RECT 26.8000 67.6000 27.6000 68.4000 ;
	    RECT 14.1000 62.4000 14.7000 63.6000 ;
	    RECT 14.0000 61.6000 14.8000 62.4000 ;
	    RECT 4.4000 51.6000 5.2000 52.4000 ;
	    RECT 4.5000 48.4000 5.1000 51.6000 ;
	    RECT 4.4000 47.6000 5.2000 48.4000 ;
	    RECT 20.4000 47.6000 21.2000 48.4000 ;
	    RECT 25.2000 46.2000 26.0000 57.8000 ;
	    RECT 26.9000 52.4000 27.5000 67.6000 ;
	    RECT 30.0000 64.2000 30.8000 75.8000 ;
	    RECT 33.2000 66.2000 34.0000 71.8000 ;
	    RECT 34.8000 71.6000 35.6000 72.4000 ;
	    RECT 34.9000 70.4000 35.5000 71.6000 ;
	    RECT 34.8000 69.6000 35.6000 70.4000 ;
	    RECT 33.2000 55.6000 34.0000 56.4000 ;
	    RECT 33.3000 52.6000 33.9000 55.6000 ;
	    RECT 26.8000 51.6000 27.6000 52.4000 ;
	    RECT 28.4000 51.6000 29.2000 52.4000 ;
	    RECT 33.2000 51.8000 34.0000 52.6000 ;
	    RECT 17.2000 43.6000 18.0000 44.4000 ;
	    RECT 1.2000 33.6000 2.0000 34.4000 ;
	    RECT 4.4000 25.6000 5.2000 26.4000 ;
	    RECT 4.5000 12.4000 5.1000 25.6000 ;
	    RECT 6.0000 24.2000 6.8000 35.8000 ;
	    RECT 14.0000 35.6000 14.8000 36.4000 ;
	    RECT 14.1000 30.2000 14.7000 35.6000 ;
	    RECT 14.0000 29.4000 14.8000 30.2000 ;
	    RECT 15.6000 24.2000 16.4000 35.8000 ;
	    RECT 17.3000 28.4000 17.9000 43.6000 ;
	    RECT 17.2000 27.6000 18.0000 28.4000 ;
	    RECT 4.4000 11.6000 5.2000 12.4000 ;
	    RECT 9.2000 11.6000 10.0000 12.4000 ;
	    RECT 9.3000 8.3000 9.9000 11.6000 ;
	    RECT 10.8000 9.6000 11.6000 10.4000 ;
	    RECT 10.9000 8.4000 11.5000 9.6000 ;
	    RECT 10.8000 8.3000 11.6000 8.4000 ;
	    RECT 9.3000 7.7000 11.6000 8.3000 ;
	    RECT 10.8000 7.6000 11.6000 7.7000 ;
	    RECT 15.6000 6.2000 16.4000 17.8000 ;
	    RECT 17.3000 12.4000 17.9000 27.6000 ;
	    RECT 18.8000 26.2000 19.6000 31.8000 ;
	    RECT 20.4000 26.2000 21.2000 31.8000 ;
	    RECT 22.0000 27.6000 22.8000 28.4000 ;
	    RECT 22.1000 14.4000 22.7000 27.6000 ;
	    RECT 23.6000 24.2000 24.4000 35.8000 ;
	    RECT 26.9000 28.4000 27.5000 51.6000 ;
	    RECT 28.5000 30.4000 29.1000 51.6000 ;
	    RECT 34.8000 46.2000 35.6000 57.8000 ;
	    RECT 36.5000 54.4000 37.1000 91.6000 ;
	    RECT 44.4000 86.2000 45.2000 97.8000 ;
	    RECT 39.6000 73.6000 40.4000 74.4000 ;
	    RECT 42.8000 73.6000 43.6000 74.4000 ;
	    RECT 39.7000 72.4000 40.3000 73.6000 ;
	    RECT 46.1000 72.4000 46.7000 185.6000 ;
	    RECT 55.6000 183.6000 56.4000 184.4000 ;
	    RECT 58.8000 183.6000 59.6000 184.4000 ;
	    RECT 55.7000 178.4000 56.3000 183.6000 ;
	    RECT 49.2000 166.2000 50.0000 177.8000 ;
	    RECT 55.6000 177.6000 56.4000 178.4000 ;
	    RECT 58.9000 172.4000 59.5000 183.6000 ;
	    RECT 58.8000 171.6000 59.6000 172.4000 ;
	    RECT 60.4000 166.2000 61.2000 177.8000 ;
	    RECT 65.3000 164.4000 65.9000 185.6000 ;
	    RECT 66.8000 171.6000 67.6000 172.4000 ;
	    RECT 54.0000 163.6000 54.8000 164.4000 ;
	    RECT 65.2000 163.6000 66.0000 164.4000 ;
	    RECT 54.1000 162.4000 54.7000 163.6000 ;
	    RECT 54.0000 161.6000 54.8000 162.4000 ;
	    RECT 58.8000 157.6000 59.6000 158.4000 ;
	    RECT 47.6000 155.6000 48.4000 156.4000 ;
	    RECT 47.7000 150.4000 48.3000 155.6000 ;
	    RECT 47.6000 149.6000 48.4000 150.4000 ;
	    RECT 52.4000 147.6000 53.2000 148.4000 ;
	    RECT 47.6000 126.2000 48.4000 137.8000 ;
	    RECT 52.5000 134.4000 53.1000 147.6000 ;
	    RECT 54.0000 144.2000 54.8000 155.8000 ;
	    RECT 60.4000 146.2000 61.2000 151.8000 ;
	    RECT 62.0000 147.6000 62.8000 148.4000 ;
	    RECT 63.6000 144.2000 64.4000 155.8000 ;
	    RECT 65.3000 148.4000 65.9000 163.6000 ;
	    RECT 65.2000 147.6000 66.0000 148.4000 ;
	    RECT 66.8000 143.6000 67.6000 144.4000 ;
	    RECT 65.2000 139.6000 66.0000 140.4000 ;
	    RECT 52.4000 133.6000 53.2000 134.4000 ;
	    RECT 49.2000 109.4000 50.0000 110.4000 ;
	    RECT 50.8000 104.2000 51.6000 115.8000 ;
	    RECT 52.5000 108.4000 53.1000 133.6000 ;
	    RECT 55.6000 131.8000 56.4000 132.6000 ;
	    RECT 55.7000 128.4000 56.3000 131.8000 ;
	    RECT 55.6000 127.6000 56.4000 128.4000 ;
	    RECT 57.2000 126.2000 58.0000 137.8000 ;
	    RECT 60.4000 130.2000 61.2000 135.8000 ;
	    RECT 62.0000 135.6000 62.8000 136.4000 ;
	    RECT 65.3000 132.4000 65.9000 139.6000 ;
	    RECT 66.9000 134.4000 67.5000 143.6000 ;
	    RECT 68.5000 142.4000 69.1000 187.6000 ;
	    RECT 70.0000 186.2000 70.8000 191.8000 ;
	    RECT 71.6000 187.6000 72.4000 188.4000 ;
	    RECT 70.0000 166.2000 70.8000 177.8000 ;
	    RECT 71.7000 174.4000 72.3000 187.6000 ;
	    RECT 73.2000 184.2000 74.0000 195.8000 ;
	    RECT 79.7000 190.4000 80.3000 213.6000 ;
	    RECT 81.3000 212.4000 81.9000 213.6000 ;
	    RECT 81.2000 211.6000 82.0000 212.4000 ;
	    RECT 86.0000 206.2000 86.8000 217.8000 ;
	    RECT 90.8000 217.6000 91.6000 218.4000 ;
	    RECT 92.5000 214.4000 93.1000 225.6000 ;
	    RECT 94.1000 218.4000 94.7000 231.6000 ;
	    RECT 95.6000 229.6000 96.4000 230.4000 ;
	    RECT 97.2000 229.6000 98.0000 230.4000 ;
	    RECT 97.3000 222.4000 97.9000 229.6000 ;
	    RECT 98.9000 228.4000 99.5000 237.6000 ;
	    RECT 98.8000 227.6000 99.6000 228.4000 ;
	    RECT 106.8000 226.2000 107.6000 231.8000 ;
	    RECT 110.0000 224.2000 110.8000 235.8000 ;
	    RECT 111.6000 229.4000 112.4000 230.4000 ;
	    RECT 111.6000 225.6000 112.4000 226.4000 ;
	    RECT 97.2000 222.3000 98.0000 222.4000 ;
	    RECT 95.7000 221.7000 98.0000 222.3000 ;
	    RECT 94.0000 217.6000 94.8000 218.4000 ;
	    RECT 92.4000 213.6000 93.2000 214.4000 ;
	    RECT 92.4000 211.6000 93.2000 212.4000 ;
	    RECT 81.2000 199.6000 82.0000 200.4000 ;
	    RECT 78.0000 189.6000 78.8000 190.4000 ;
	    RECT 79.6000 189.6000 80.4000 190.4000 ;
	    RECT 74.8000 183.6000 75.6000 184.4000 ;
	    RECT 71.6000 173.6000 72.4000 174.4000 ;
	    RECT 73.2000 170.2000 74.0000 175.8000 ;
	    RECT 74.9000 174.4000 75.5000 183.6000 ;
	    RECT 74.8000 173.6000 75.6000 174.4000 ;
	    RECT 79.6000 173.6000 80.4000 174.4000 ;
	    RECT 79.7000 172.4000 80.3000 173.6000 ;
	    RECT 79.6000 171.6000 80.4000 172.4000 ;
	    RECT 81.3000 170.4000 81.9000 199.6000 ;
	    RECT 92.5000 198.4000 93.1000 211.6000 ;
	    RECT 95.7000 210.4000 96.3000 221.7000 ;
	    RECT 97.2000 221.6000 98.0000 221.7000 ;
	    RECT 97.2000 217.6000 98.0000 218.4000 ;
	    RECT 97.3000 214.4000 97.9000 217.6000 ;
	    RECT 105.2000 215.6000 106.0000 216.4000 ;
	    RECT 97.2000 213.6000 98.0000 214.4000 ;
	    RECT 100.4000 213.6000 101.2000 214.4000 ;
	    RECT 105.3000 212.4000 105.9000 215.6000 ;
	    RECT 111.7000 214.4000 112.3000 225.6000 ;
	    RECT 106.8000 213.6000 107.6000 214.4000 ;
	    RECT 111.6000 213.6000 112.4000 214.4000 ;
	    RECT 105.2000 211.6000 106.0000 212.4000 ;
	    RECT 105.3000 210.4000 105.9000 211.6000 ;
	    RECT 95.6000 209.6000 96.4000 210.4000 ;
	    RECT 100.4000 209.6000 101.2000 210.4000 ;
	    RECT 105.2000 209.6000 106.0000 210.4000 ;
	    RECT 106.9000 204.4000 107.5000 213.6000 ;
	    RECT 94.0000 203.6000 94.8000 204.4000 ;
	    RECT 106.8000 203.6000 107.6000 204.4000 ;
	    RECT 92.4000 197.6000 93.2000 198.4000 ;
	    RECT 82.8000 184.2000 83.6000 195.8000 ;
	    RECT 87.6000 193.6000 88.4000 194.4000 ;
	    RECT 87.7000 192.4000 88.3000 193.6000 ;
	    RECT 87.6000 191.6000 88.4000 192.4000 ;
	    RECT 94.1000 188.4000 94.7000 203.6000 ;
	    RECT 100.4000 191.6000 101.2000 192.4000 ;
	    RECT 105.2000 191.6000 106.0000 192.4000 ;
	    RECT 105.3000 190.4000 105.9000 191.6000 ;
	    RECT 95.6000 189.6000 96.4000 190.4000 ;
	    RECT 97.2000 189.6000 98.0000 190.4000 ;
	    RECT 103.6000 189.6000 104.4000 190.4000 ;
	    RECT 105.2000 189.6000 106.0000 190.4000 ;
	    RECT 94.0000 187.6000 94.8000 188.4000 ;
	    RECT 84.4000 175.6000 85.2000 176.4000 ;
	    RECT 84.5000 174.4000 85.1000 175.6000 ;
	    RECT 84.4000 173.6000 85.2000 174.4000 ;
	    RECT 82.8000 171.6000 83.6000 172.4000 ;
	    RECT 78.0000 169.6000 78.8000 170.4000 ;
	    RECT 81.2000 169.6000 82.0000 170.4000 ;
	    RECT 78.1000 168.4000 78.7000 169.6000 ;
	    RECT 78.0000 167.6000 78.8000 168.4000 ;
	    RECT 70.0000 153.6000 70.8000 154.4000 ;
	    RECT 70.1000 150.4000 70.7000 153.6000 ;
	    RECT 70.0000 149.6000 70.8000 150.4000 ;
	    RECT 70.0000 147.6000 70.8000 148.4000 ;
	    RECT 68.4000 141.6000 69.2000 142.4000 ;
	    RECT 68.5000 134.4000 69.1000 141.6000 ;
	    RECT 70.1000 138.4000 70.7000 147.6000 ;
	    RECT 73.2000 144.2000 74.0000 155.8000 ;
	    RECT 78.0000 143.6000 78.8000 144.4000 ;
	    RECT 79.6000 143.6000 80.4000 144.4000 ;
	    RECT 78.1000 138.4000 78.7000 143.6000 ;
	    RECT 79.7000 142.4000 80.3000 143.6000 ;
	    RECT 79.6000 141.6000 80.4000 142.4000 ;
	    RECT 81.3000 140.3000 81.9000 169.6000 ;
	    RECT 82.9000 168.4000 83.5000 171.6000 ;
	    RECT 86.0000 170.2000 86.8000 175.8000 ;
	    RECT 87.6000 173.6000 88.4000 174.4000 ;
	    RECT 82.8000 167.6000 83.6000 168.4000 ;
	    RECT 86.0000 167.6000 86.8000 168.4000 ;
	    RECT 84.4000 147.6000 85.2000 148.4000 ;
	    RECT 79.7000 139.7000 81.9000 140.3000 ;
	    RECT 70.0000 137.6000 70.8000 138.4000 ;
	    RECT 78.0000 137.6000 78.8000 138.4000 ;
	    RECT 79.7000 136.4000 80.3000 139.7000 ;
	    RECT 82.8000 139.6000 83.6000 140.4000 ;
	    RECT 82.9000 136.4000 83.5000 139.6000 ;
	    RECT 84.5000 138.4000 85.1000 147.6000 ;
	    RECT 84.4000 137.6000 85.2000 138.4000 ;
	    RECT 79.6000 135.6000 80.4000 136.4000 ;
	    RECT 81.2000 135.6000 82.0000 136.4000 ;
	    RECT 82.8000 135.6000 83.6000 136.4000 ;
	    RECT 66.8000 133.6000 67.6000 134.4000 ;
	    RECT 68.4000 133.6000 69.2000 134.4000 ;
	    RECT 78.0000 133.6000 78.8000 134.4000 ;
	    RECT 65.2000 131.6000 66.0000 132.4000 ;
	    RECT 66.8000 131.6000 67.6000 132.4000 ;
	    RECT 71.6000 131.6000 72.4000 132.4000 ;
	    RECT 79.6000 132.3000 80.4000 132.4000 ;
	    RECT 81.3000 132.3000 81.9000 135.6000 ;
	    RECT 79.6000 131.7000 81.9000 132.3000 ;
	    RECT 79.6000 131.6000 80.4000 131.7000 ;
	    RECT 82.8000 131.6000 83.6000 132.4000 ;
	    RECT 62.0000 129.6000 62.8000 130.4000 ;
	    RECT 55.6000 113.6000 56.4000 114.4000 ;
	    RECT 58.8000 113.6000 59.6000 114.4000 ;
	    RECT 55.7000 112.4000 56.3000 113.6000 ;
	    RECT 52.4000 107.6000 53.2000 108.4000 ;
	    RECT 54.0000 106.2000 54.8000 111.8000 ;
	    RECT 55.6000 111.6000 56.4000 112.4000 ;
	    RECT 58.9000 110.4000 59.5000 113.6000 ;
	    RECT 55.6000 109.6000 56.4000 110.4000 ;
	    RECT 58.8000 109.6000 59.6000 110.4000 ;
	    RECT 55.7000 108.4000 56.3000 109.6000 ;
	    RECT 55.6000 107.6000 56.4000 108.4000 ;
	    RECT 60.4000 107.6000 61.2000 108.4000 ;
	    RECT 62.0000 106.2000 62.8000 111.8000 ;
	    RECT 63.6000 107.6000 64.4000 108.4000 ;
	    RECT 55.6000 101.6000 56.4000 102.4000 ;
	    RECT 60.4000 101.6000 61.2000 102.4000 ;
	    RECT 55.7000 96.4000 56.3000 101.6000 ;
	    RECT 60.5000 96.4000 61.1000 101.6000 ;
	    RECT 47.6000 90.2000 48.4000 95.8000 ;
	    RECT 55.6000 95.6000 56.4000 96.4000 ;
	    RECT 58.8000 95.6000 59.6000 96.4000 ;
	    RECT 60.4000 95.6000 61.2000 96.4000 ;
	    RECT 49.2000 93.6000 50.0000 94.4000 ;
	    RECT 52.4000 93.6000 53.2000 94.4000 ;
	    RECT 52.5000 92.4000 53.1000 93.6000 ;
	    RECT 58.9000 92.4000 59.5000 95.6000 ;
	    RECT 63.7000 94.4000 64.3000 107.6000 ;
	    RECT 65.2000 104.2000 66.0000 115.8000 ;
	    RECT 65.2000 96.3000 66.0000 96.4000 ;
	    RECT 66.9000 96.3000 67.5000 131.6000 ;
	    RECT 71.7000 114.4000 72.3000 131.6000 ;
	    RECT 73.2000 129.6000 74.0000 130.4000 ;
	    RECT 71.6000 113.6000 72.4000 114.4000 ;
	    RECT 71.6000 111.6000 72.4000 112.4000 ;
	    RECT 71.7000 110.4000 72.3000 111.6000 ;
	    RECT 71.6000 109.6000 72.4000 110.4000 ;
	    RECT 68.4000 107.6000 69.2000 108.4000 ;
	    RECT 68.5000 98.4000 69.1000 107.6000 ;
	    RECT 70.0000 101.6000 70.8000 102.4000 ;
	    RECT 73.3000 102.3000 73.9000 129.6000 ;
	    RECT 82.9000 126.4000 83.5000 131.6000 ;
	    RECT 84.4000 129.6000 85.2000 130.4000 ;
	    RECT 82.8000 125.6000 83.6000 126.4000 ;
	    RECT 81.2000 123.6000 82.0000 124.4000 ;
	    RECT 81.3000 116.4000 81.9000 123.6000 ;
	    RECT 74.8000 104.2000 75.6000 115.8000 ;
	    RECT 81.2000 115.6000 82.0000 116.4000 ;
	    RECT 86.1000 116.3000 86.7000 167.6000 ;
	    RECT 89.2000 166.2000 90.0000 177.8000 ;
	    RECT 94.1000 176.4000 94.7000 187.6000 ;
	    RECT 94.0000 175.6000 94.8000 176.4000 ;
	    RECT 94.0000 171.6000 94.8000 172.4000 ;
	    RECT 90.8000 153.6000 91.6000 154.4000 ;
	    RECT 94.0000 153.6000 94.8000 154.4000 ;
	    RECT 87.6000 151.6000 88.4000 152.4000 ;
	    RECT 87.7000 150.4000 88.3000 151.6000 ;
	    RECT 90.9000 150.4000 91.5000 153.6000 ;
	    RECT 87.6000 149.6000 88.4000 150.4000 ;
	    RECT 90.8000 149.6000 91.6000 150.4000 ;
	    RECT 92.4000 149.6000 93.2000 150.4000 ;
	    RECT 89.2000 133.6000 90.0000 134.4000 ;
	    RECT 87.6000 131.6000 88.4000 132.4000 ;
	    RECT 90.8000 131.6000 91.6000 132.4000 ;
	    RECT 87.7000 116.4000 88.3000 131.6000 ;
	    RECT 90.9000 130.4000 91.5000 131.6000 ;
	    RECT 90.8000 129.6000 91.6000 130.4000 ;
	    RECT 92.5000 118.4000 93.1000 149.6000 ;
	    RECT 94.1000 148.4000 94.7000 153.6000 ;
	    RECT 95.7000 150.3000 96.3000 189.6000 ;
	    RECT 103.7000 188.4000 104.3000 189.6000 ;
	    RECT 100.4000 187.6000 101.2000 188.4000 ;
	    RECT 103.6000 187.6000 104.4000 188.4000 ;
	    RECT 105.2000 187.6000 106.0000 188.4000 ;
	    RECT 98.8000 166.2000 99.6000 177.8000 ;
	    RECT 98.8000 151.6000 99.6000 152.4000 ;
	    RECT 98.9000 150.4000 99.5000 151.6000 ;
	    RECT 97.2000 150.3000 98.0000 150.4000 ;
	    RECT 95.7000 149.7000 98.0000 150.3000 ;
	    RECT 97.2000 149.6000 98.0000 149.7000 ;
	    RECT 98.8000 149.6000 99.6000 150.4000 ;
	    RECT 97.3000 148.4000 97.9000 149.6000 ;
	    RECT 94.0000 147.6000 94.8000 148.4000 ;
	    RECT 97.2000 147.6000 98.0000 148.4000 ;
	    RECT 100.5000 146.4000 101.1000 187.6000 ;
	    RECT 103.6000 177.6000 104.4000 178.4000 ;
	    RECT 111.7000 174.4000 112.3000 213.6000 ;
	    RECT 113.3000 188.4000 113.9000 245.6000 ;
	    RECT 127.6000 243.6000 128.4000 244.4000 ;
	    RECT 137.2000 243.6000 138.0000 244.4000 ;
	    RECT 114.8000 227.6000 115.6000 228.4000 ;
	    RECT 114.9000 214.4000 115.5000 227.6000 ;
	    RECT 119.6000 224.2000 120.4000 235.8000 ;
	    RECT 124.4000 233.6000 125.2000 234.4000 ;
	    RECT 124.5000 232.4000 125.1000 233.6000 ;
	    RECT 122.8000 231.6000 123.6000 232.4000 ;
	    RECT 124.4000 231.6000 125.2000 232.4000 ;
	    RECT 122.9000 224.3000 123.5000 231.6000 ;
	    RECT 124.5000 226.4000 125.1000 231.6000 ;
	    RECT 127.7000 230.4000 128.3000 243.6000 ;
	    RECT 137.3000 242.4000 137.9000 243.6000 ;
	    RECT 130.8000 241.6000 131.6000 242.4000 ;
	    RECT 137.2000 241.6000 138.0000 242.4000 ;
	    RECT 130.9000 230.4000 131.5000 241.6000 ;
	    RECT 135.6000 235.6000 136.4000 236.4000 ;
	    RECT 134.0000 231.6000 134.8000 232.4000 ;
	    RECT 134.1000 230.4000 134.7000 231.6000 ;
	    RECT 126.0000 229.6000 126.8000 230.4000 ;
	    RECT 127.6000 229.6000 128.4000 230.4000 ;
	    RECT 130.8000 229.6000 131.6000 230.4000 ;
	    RECT 134.0000 229.6000 134.8000 230.4000 ;
	    RECT 126.1000 228.4000 126.7000 229.6000 ;
	    RECT 126.0000 227.6000 126.8000 228.4000 ;
	    RECT 124.4000 225.6000 125.2000 226.4000 ;
	    RECT 127.6000 224.3000 128.4000 224.4000 ;
	    RECT 122.9000 223.7000 128.4000 224.3000 ;
	    RECT 127.6000 223.6000 128.4000 223.7000 ;
	    RECT 119.6000 219.6000 120.4000 220.4000 ;
	    RECT 114.8000 213.6000 115.6000 214.4000 ;
	    RECT 114.9000 210.4000 115.5000 213.6000 ;
	    RECT 119.7000 212.4000 120.3000 219.6000 ;
	    RECT 127.6000 213.6000 128.4000 214.4000 ;
	    RECT 116.4000 211.6000 117.2000 212.4000 ;
	    RECT 119.6000 211.6000 120.4000 212.4000 ;
	    RECT 121.2000 211.6000 122.0000 212.4000 ;
	    RECT 126.0000 211.6000 126.8000 212.4000 ;
	    RECT 114.8000 209.6000 115.6000 210.4000 ;
	    RECT 116.5000 198.4000 117.1000 211.6000 ;
	    RECT 118.0000 207.6000 118.8000 208.4000 ;
	    RECT 116.4000 197.6000 117.2000 198.4000 ;
	    RECT 121.3000 190.4000 121.9000 211.6000 ;
	    RECT 122.8000 209.6000 123.6000 210.4000 ;
	    RECT 119.6000 189.6000 120.4000 190.4000 ;
	    RECT 121.2000 189.6000 122.0000 190.4000 ;
	    RECT 122.8000 189.6000 123.6000 190.4000 ;
	    RECT 124.4000 189.6000 125.2000 190.4000 ;
	    RECT 119.7000 188.4000 120.3000 189.6000 ;
	    RECT 124.5000 188.4000 125.1000 189.6000 ;
	    RECT 127.7000 188.4000 128.3000 213.6000 ;
	    RECT 129.2000 210.2000 130.0000 215.8000 ;
	    RECT 130.8000 213.6000 131.6000 214.4000 ;
	    RECT 132.4000 206.2000 133.2000 217.8000 ;
	    RECT 134.1000 204.3000 134.7000 229.6000 ;
	    RECT 135.7000 212.4000 136.3000 235.6000 ;
	    RECT 137.2000 231.6000 138.0000 232.4000 ;
	    RECT 137.3000 230.4000 137.9000 231.6000 ;
	    RECT 137.2000 229.6000 138.0000 230.4000 ;
	    RECT 138.9000 228.4000 139.5000 253.6000 ;
	    RECT 142.0000 251.6000 142.8000 252.4000 ;
	    RECT 140.4000 249.6000 141.2000 250.4000 ;
	    RECT 140.5000 246.3000 141.1000 249.6000 ;
	    RECT 142.1000 248.4000 142.7000 251.6000 ;
	    RECT 142.0000 247.6000 142.8000 248.4000 ;
	    RECT 140.5000 245.7000 142.7000 246.3000 ;
	    RECT 142.1000 238.4000 142.7000 245.7000 ;
	    RECT 142.0000 237.6000 142.8000 238.4000 ;
	    RECT 143.7000 232.3000 144.3000 267.7000 ;
	    RECT 150.0000 267.6000 150.8000 268.4000 ;
	    RECT 145.2000 265.6000 146.0000 266.4000 ;
	    RECT 154.8000 266.2000 155.6000 271.8000 ;
	    RECT 156.5000 268.4000 157.1000 309.6000 ;
	    RECT 159.7000 308.4000 160.3000 327.7000 ;
	    RECT 161.2000 327.6000 162.0000 327.7000 ;
	    RECT 166.0000 326.2000 166.8000 337.8000 ;
	    RECT 170.8000 333.6000 171.6000 334.4000 ;
	    RECT 162.9000 310.2000 163.5000 310.3000 ;
	    RECT 162.8000 309.4000 163.6000 310.2000 ;
	    RECT 159.6000 307.6000 160.4000 308.4000 ;
	    RECT 158.0000 297.6000 158.8000 298.4000 ;
	    RECT 159.7000 296.4000 160.3000 307.6000 ;
	    RECT 162.9000 298.4000 163.5000 309.4000 ;
	    RECT 164.4000 304.2000 165.2000 315.8000 ;
	    RECT 167.6000 306.2000 168.4000 311.8000 ;
	    RECT 170.9000 310.4000 171.5000 333.6000 ;
	    RECT 174.0000 331.6000 174.8000 332.6000 ;
	    RECT 175.6000 326.2000 176.4000 337.8000 ;
	    RECT 178.8000 330.2000 179.6000 335.8000 ;
	    RECT 193.2000 335.6000 194.0000 336.4000 ;
	    RECT 183.6000 333.6000 184.4000 334.4000 ;
	    RECT 185.2000 333.6000 186.0000 334.4000 ;
	    RECT 186.8000 333.6000 187.6000 334.4000 ;
	    RECT 183.7000 332.4000 184.3000 333.6000 ;
	    RECT 183.6000 331.6000 184.4000 332.4000 ;
	    RECT 183.6000 329.6000 184.4000 330.4000 ;
	    RECT 180.4000 327.6000 181.2000 328.4000 ;
	    RECT 185.3000 324.4000 185.9000 333.6000 ;
	    RECT 186.9000 332.4000 187.5000 333.6000 ;
	    RECT 186.8000 331.6000 187.6000 332.4000 ;
	    RECT 190.0000 331.6000 190.8000 332.4000 ;
	    RECT 186.8000 329.6000 187.6000 330.4000 ;
	    RECT 196.4000 330.2000 197.2000 335.8000 ;
	    RECT 199.6000 326.2000 200.4000 337.8000 ;
	    RECT 202.8000 331.6000 203.6000 332.4000 ;
	    RECT 207.6000 331.6000 208.4000 332.4000 ;
	    RECT 202.9000 328.4000 203.5000 331.6000 ;
	    RECT 207.7000 330.4000 208.3000 331.6000 ;
	    RECT 207.6000 329.6000 208.4000 330.4000 ;
	    RECT 202.8000 327.6000 203.6000 328.4000 ;
	    RECT 209.2000 326.2000 210.0000 337.8000 ;
	    RECT 242.8000 337.6000 243.6000 338.4000 ;
	    RECT 242.9000 336.4000 243.5000 337.6000 ;
	    RECT 242.8000 335.6000 243.6000 336.4000 ;
	    RECT 215.6000 333.6000 216.4000 334.4000 ;
	    RECT 217.2000 333.6000 218.0000 334.4000 ;
	    RECT 222.0000 333.6000 222.8000 334.4000 ;
	    RECT 226.8000 333.6000 227.6000 334.4000 ;
	    RECT 214.0000 327.6000 214.8000 328.4000 ;
	    RECT 215.7000 324.4000 216.3000 333.6000 ;
	    RECT 217.3000 332.4000 217.9000 333.6000 ;
	    RECT 217.2000 331.6000 218.0000 332.4000 ;
	    RECT 225.2000 331.6000 226.0000 332.4000 ;
	    RECT 185.2000 323.6000 186.0000 324.4000 ;
	    RECT 215.6000 323.6000 216.4000 324.4000 ;
	    RECT 194.8000 321.6000 195.6000 322.4000 ;
	    RECT 201.2000 321.6000 202.0000 322.4000 ;
	    RECT 210.8000 321.6000 211.6000 322.4000 ;
	    RECT 180.4000 319.6000 181.2000 320.4000 ;
	    RECT 172.4000 313.6000 173.2000 314.4000 ;
	    RECT 170.8000 309.6000 171.6000 310.4000 ;
	    RECT 169.2000 305.6000 170.0000 306.4000 ;
	    RECT 169.3000 304.4000 169.9000 305.6000 ;
	    RECT 169.2000 303.6000 170.0000 304.4000 ;
	    RECT 172.5000 300.4000 173.1000 313.6000 ;
	    RECT 174.0000 304.2000 174.8000 315.8000 ;
	    RECT 175.6000 309.6000 176.4000 310.4000 ;
	    RECT 170.8000 299.6000 171.6000 300.4000 ;
	    RECT 172.4000 299.6000 173.2000 300.4000 ;
	    RECT 162.8000 297.6000 163.6000 298.4000 ;
	    RECT 169.2000 297.6000 170.0000 298.4000 ;
	    RECT 159.6000 295.6000 160.4000 296.4000 ;
	    RECT 162.8000 293.6000 163.6000 294.4000 ;
	    RECT 164.4000 293.6000 165.2000 294.4000 ;
	    RECT 169.2000 293.6000 170.0000 294.4000 ;
	    RECT 162.9000 292.4000 163.5000 293.6000 ;
	    RECT 162.8000 291.6000 163.6000 292.4000 ;
	    RECT 164.4000 291.6000 165.2000 292.4000 ;
	    RECT 162.9000 290.4000 163.5000 291.6000 ;
	    RECT 158.0000 289.6000 158.8000 290.4000 ;
	    RECT 161.2000 289.6000 162.0000 290.4000 ;
	    RECT 162.8000 289.6000 163.6000 290.4000 ;
	    RECT 158.1000 278.4000 158.7000 289.6000 ;
	    RECT 164.5000 288.3000 165.1000 291.6000 ;
	    RECT 166.0000 289.6000 166.8000 290.4000 ;
	    RECT 162.9000 287.7000 165.1000 288.3000 ;
	    RECT 158.0000 277.6000 158.8000 278.4000 ;
	    RECT 156.4000 267.6000 157.2000 268.4000 ;
	    RECT 145.3000 242.4000 145.9000 265.6000 ;
	    RECT 150.0000 263.6000 150.8000 264.4000 ;
	    RECT 158.0000 264.2000 158.8000 275.8000 ;
	    RECT 161.2000 269.6000 162.0000 270.4000 ;
	    RECT 148.4000 261.6000 149.2000 262.4000 ;
	    RECT 146.8000 246.2000 147.6000 257.8000 ;
	    RECT 145.2000 241.6000 146.0000 242.4000 ;
	    RECT 145.2000 232.3000 146.0000 232.4000 ;
	    RECT 143.7000 231.7000 146.0000 232.3000 ;
	    RECT 145.2000 231.6000 146.0000 231.7000 ;
	    RECT 142.0000 229.6000 142.8000 230.4000 ;
	    RECT 146.8000 230.3000 147.6000 230.4000 ;
	    RECT 148.5000 230.3000 149.1000 261.6000 ;
	    RECT 150.1000 250.4000 150.7000 263.6000 ;
	    RECT 154.8000 251.6000 155.6000 252.6000 ;
	    RECT 150.0000 249.6000 150.8000 250.4000 ;
	    RECT 150.0000 247.6000 150.8000 248.4000 ;
	    RECT 146.8000 229.7000 149.1000 230.3000 ;
	    RECT 146.8000 229.6000 147.6000 229.7000 ;
	    RECT 138.8000 227.6000 139.6000 228.4000 ;
	    RECT 150.1000 228.3000 150.7000 247.6000 ;
	    RECT 156.4000 246.2000 157.2000 257.8000 ;
	    RECT 158.0000 255.6000 158.8000 256.4000 ;
	    RECT 158.1000 254.4000 158.7000 255.6000 ;
	    RECT 158.0000 253.6000 158.8000 254.4000 ;
	    RECT 153.2000 243.6000 154.0000 244.4000 ;
	    RECT 158.1000 244.3000 158.7000 253.6000 ;
	    RECT 159.6000 250.2000 160.4000 255.8000 ;
	    RECT 161.2000 253.6000 162.0000 254.4000 ;
	    RECT 156.5000 243.7000 158.7000 244.3000 ;
	    RECT 153.3000 238.4000 153.9000 243.6000 ;
	    RECT 153.2000 237.6000 154.0000 238.4000 ;
	    RECT 151.6000 233.6000 152.4000 234.4000 ;
	    RECT 151.7000 228.4000 152.3000 233.6000 ;
	    RECT 154.8000 229.6000 155.6000 230.4000 ;
	    RECT 148.5000 227.7000 150.7000 228.3000 ;
	    RECT 135.6000 211.6000 136.4000 212.4000 ;
	    RECT 137.2000 209.6000 138.0000 210.4000 ;
	    RECT 132.5000 203.7000 134.7000 204.3000 ;
	    RECT 129.2000 191.6000 130.0000 192.4000 ;
	    RECT 130.8000 191.6000 131.6000 192.4000 ;
	    RECT 129.3000 190.4000 129.9000 191.6000 ;
	    RECT 129.2000 189.6000 130.0000 190.4000 ;
	    RECT 130.9000 188.4000 131.5000 191.6000 ;
	    RECT 132.5000 188.4000 133.1000 203.7000 ;
	    RECT 134.0000 191.6000 134.8000 192.4000 ;
	    RECT 134.1000 190.4000 134.7000 191.6000 ;
	    RECT 137.3000 190.4000 137.9000 209.6000 ;
	    RECT 138.9000 190.4000 139.5000 227.6000 ;
	    RECT 146.8000 225.6000 147.6000 226.4000 ;
	    RECT 146.9000 220.4000 147.5000 225.6000 ;
	    RECT 146.8000 219.6000 147.6000 220.4000 ;
	    RECT 142.0000 206.2000 142.8000 217.8000 ;
	    RECT 148.5000 212.4000 149.1000 227.7000 ;
	    RECT 151.6000 227.6000 152.4000 228.4000 ;
	    RECT 150.0000 225.6000 150.8000 226.4000 ;
	    RECT 151.6000 225.6000 152.4000 226.4000 ;
	    RECT 150.1000 216.3000 150.7000 225.6000 ;
	    RECT 151.7000 220.4000 152.3000 225.6000 ;
	    RECT 151.6000 219.6000 152.4000 220.4000 ;
	    RECT 154.9000 216.4000 155.5000 229.6000 ;
	    RECT 151.6000 216.3000 152.4000 216.4000 ;
	    RECT 150.1000 215.7000 152.4000 216.3000 ;
	    RECT 151.6000 215.6000 152.4000 215.7000 ;
	    RECT 154.8000 215.6000 155.6000 216.4000 ;
	    RECT 156.5000 214.4000 157.1000 243.7000 ;
	    RECT 158.0000 241.6000 158.8000 242.4000 ;
	    RECT 158.1000 230.4000 158.7000 241.6000 ;
	    RECT 161.3000 238.4000 161.9000 253.6000 ;
	    RECT 162.9000 252.4000 163.5000 287.7000 ;
	    RECT 166.1000 286.4000 166.7000 289.6000 ;
	    RECT 166.0000 285.6000 166.8000 286.4000 ;
	    RECT 167.6000 264.2000 168.4000 275.8000 ;
	    RECT 164.4000 257.6000 165.2000 258.4000 ;
	    RECT 162.8000 251.6000 163.6000 252.4000 ;
	    RECT 162.9000 250.4000 163.5000 251.6000 ;
	    RECT 164.5000 250.4000 165.1000 257.6000 ;
	    RECT 166.0000 253.6000 166.8000 254.4000 ;
	    RECT 167.6000 253.6000 168.4000 254.4000 ;
	    RECT 166.1000 252.4000 166.7000 253.6000 ;
	    RECT 166.0000 251.6000 166.8000 252.4000 ;
	    RECT 167.7000 250.4000 168.3000 253.6000 ;
	    RECT 162.8000 249.6000 163.6000 250.4000 ;
	    RECT 164.4000 249.6000 165.2000 250.4000 ;
	    RECT 167.6000 249.6000 168.4000 250.4000 ;
	    RECT 169.3000 246.4000 169.9000 293.6000 ;
	    RECT 170.9000 290.4000 171.5000 299.6000 ;
	    RECT 180.5000 298.3000 181.1000 319.6000 ;
	    RECT 191.6000 317.6000 192.4000 318.4000 ;
	    RECT 182.0000 313.6000 182.8000 314.4000 ;
	    RECT 182.1000 310.2000 182.7000 313.6000 ;
	    RECT 182.0000 309.4000 182.8000 310.2000 ;
	    RECT 183.6000 304.2000 184.4000 315.8000 ;
	    RECT 186.8000 306.2000 187.6000 311.8000 ;
	    RECT 191.7000 308.4000 192.3000 317.6000 ;
	    RECT 194.9000 312.4000 195.5000 321.6000 ;
	    RECT 194.8000 311.6000 195.6000 312.4000 ;
	    RECT 198.0000 311.6000 198.8000 312.4000 ;
	    RECT 199.6000 311.6000 200.4000 312.4000 ;
	    RECT 194.9000 310.4000 195.5000 311.6000 ;
	    RECT 194.8000 309.6000 195.6000 310.4000 ;
	    RECT 191.6000 307.6000 192.4000 308.4000 ;
	    RECT 198.1000 308.3000 198.7000 311.6000 ;
	    RECT 199.6000 309.6000 200.4000 310.4000 ;
	    RECT 201.3000 308.4000 201.9000 321.6000 ;
	    RECT 204.4000 317.6000 205.2000 318.4000 ;
	    RECT 198.1000 307.7000 200.3000 308.3000 ;
	    RECT 188.4000 305.6000 189.2000 306.4000 ;
	    RECT 190.0000 305.6000 190.8000 306.4000 ;
	    RECT 199.7000 306.3000 200.3000 307.7000 ;
	    RECT 201.2000 307.6000 202.0000 308.4000 ;
	    RECT 199.7000 305.7000 201.9000 306.3000 ;
	    RECT 202.8000 306.2000 203.6000 311.8000 ;
	    RECT 204.5000 310.4000 205.1000 317.6000 ;
	    RECT 204.4000 309.6000 205.2000 310.4000 ;
	    RECT 204.4000 307.6000 205.2000 308.4000 ;
	    RECT 201.3000 304.3000 201.9000 305.7000 ;
	    RECT 201.3000 303.7000 205.1000 304.3000 ;
	    RECT 206.0000 304.2000 206.8000 315.8000 ;
	    RECT 207.6000 311.6000 208.4000 312.4000 ;
	    RECT 207.7000 310.2000 208.3000 311.6000 ;
	    RECT 207.6000 309.4000 208.4000 310.2000 ;
	    RECT 209.2000 307.6000 210.0000 308.4000 ;
	    RECT 204.5000 302.3000 205.1000 303.7000 ;
	    RECT 204.5000 301.7000 208.3000 302.3000 ;
	    RECT 207.7000 298.4000 208.3000 301.7000 ;
	    RECT 182.0000 298.3000 182.8000 298.4000 ;
	    RECT 180.5000 297.7000 182.8000 298.3000 ;
	    RECT 198.0000 298.3000 198.8000 298.4000 ;
	    RECT 182.0000 297.6000 182.8000 297.7000 ;
	    RECT 177.2000 295.6000 178.0000 296.4000 ;
	    RECT 175.6000 293.6000 176.4000 294.4000 ;
	    RECT 174.0000 291.6000 174.8000 292.4000 ;
	    RECT 170.8000 289.6000 171.6000 290.4000 ;
	    RECT 174.1000 286.4000 174.7000 291.6000 ;
	    RECT 170.8000 285.6000 171.6000 286.4000 ;
	    RECT 174.0000 285.6000 174.8000 286.4000 ;
	    RECT 186.8000 286.2000 187.6000 297.8000 ;
	    RECT 194.8000 295.6000 195.6000 296.4000 ;
	    RECT 194.9000 292.6000 195.5000 295.6000 ;
	    RECT 194.8000 291.8000 195.6000 292.6000 ;
	    RECT 194.9000 291.7000 195.5000 291.8000 ;
	    RECT 196.4000 286.2000 197.2000 297.8000 ;
	    RECT 198.0000 297.7000 205.1000 298.3000 ;
	    RECT 198.0000 297.6000 198.8000 297.7000 ;
	    RECT 198.0000 293.6000 198.8000 294.4000 ;
	    RECT 199.6000 290.2000 200.4000 295.8000 ;
	    RECT 201.2000 295.6000 202.0000 296.4000 ;
	    RECT 201.3000 294.4000 201.9000 295.6000 ;
	    RECT 204.5000 294.4000 205.1000 297.7000 ;
	    RECT 206.0000 297.6000 206.8000 298.4000 ;
	    RECT 207.6000 297.6000 208.4000 298.4000 ;
	    RECT 209.3000 294.4000 209.9000 307.6000 ;
	    RECT 210.9000 296.4000 211.5000 321.6000 ;
	    RECT 214.0000 311.6000 214.8000 312.4000 ;
	    RECT 214.1000 310.4000 214.7000 311.6000 ;
	    RECT 214.0000 309.6000 214.8000 310.4000 ;
	    RECT 215.6000 304.2000 216.4000 315.8000 ;
	    RECT 217.3000 302.3000 217.9000 331.6000 ;
	    RECT 220.4000 327.6000 221.2000 328.4000 ;
	    RECT 218.8000 323.6000 219.6000 324.4000 ;
	    RECT 214.1000 301.7000 217.9000 302.3000 ;
	    RECT 210.8000 295.6000 211.6000 296.4000 ;
	    RECT 201.2000 293.6000 202.0000 294.4000 ;
	    RECT 204.4000 293.6000 205.2000 294.4000 ;
	    RECT 209.2000 293.6000 210.0000 294.4000 ;
	    RECT 210.8000 293.6000 211.6000 294.4000 ;
	    RECT 212.4000 293.6000 213.2000 294.4000 ;
	    RECT 170.9000 256.4000 171.5000 285.6000 ;
	    RECT 196.5000 283.7000 200.3000 284.3000 ;
	    RECT 196.5000 278.3000 197.1000 283.7000 ;
	    RECT 199.7000 282.4000 200.3000 283.7000 ;
	    RECT 198.0000 281.6000 198.8000 282.4000 ;
	    RECT 199.6000 281.6000 200.4000 282.4000 ;
	    RECT 182.1000 277.7000 197.1000 278.3000 ;
	    RECT 182.1000 276.4000 182.7000 277.7000 ;
	    RECT 182.0000 275.6000 182.8000 276.4000 ;
	    RECT 183.7000 275.7000 195.5000 276.3000 ;
	    RECT 180.4000 271.6000 181.2000 272.4000 ;
	    RECT 183.7000 270.4000 184.3000 275.7000 ;
	    RECT 185.2000 273.6000 186.0000 274.4000 ;
	    RECT 186.8000 273.6000 187.6000 274.4000 ;
	    RECT 174.0000 270.3000 174.8000 270.4000 ;
	    RECT 174.0000 269.7000 176.3000 270.3000 ;
	    RECT 174.0000 269.6000 174.8000 269.7000 ;
	    RECT 172.4000 263.6000 173.2000 264.4000 ;
	    RECT 172.5000 258.4000 173.1000 263.6000 ;
	    RECT 175.7000 262.4000 176.3000 269.7000 ;
	    RECT 183.6000 269.6000 184.4000 270.4000 ;
	    RECT 185.3000 268.4000 185.9000 273.6000 ;
	    RECT 186.9000 270.4000 187.5000 273.6000 ;
	    RECT 194.9000 272.4000 195.5000 275.7000 ;
	    RECT 198.1000 274.4000 198.7000 281.6000 ;
	    RECT 196.4000 273.6000 197.2000 274.4000 ;
	    RECT 198.0000 273.6000 198.8000 274.4000 ;
	    RECT 193.2000 271.6000 194.0000 272.4000 ;
	    RECT 194.8000 271.6000 195.6000 272.4000 ;
	    RECT 201.3000 272.3000 201.9000 293.6000 ;
	    RECT 202.8000 291.6000 203.6000 292.4000 ;
	    RECT 202.9000 288.4000 203.5000 291.6000 ;
	    RECT 207.6000 289.6000 208.4000 290.4000 ;
	    RECT 212.5000 290.3000 213.1000 293.6000 ;
	    RECT 214.1000 292.4000 214.7000 301.7000 ;
	    RECT 217.2000 297.6000 218.0000 298.4000 ;
	    RECT 215.6000 293.6000 216.4000 294.4000 ;
	    RECT 214.0000 291.6000 214.8000 292.4000 ;
	    RECT 210.9000 289.7000 213.1000 290.3000 ;
	    RECT 207.7000 288.4000 208.3000 289.6000 ;
	    RECT 202.8000 287.6000 203.6000 288.4000 ;
	    RECT 207.6000 287.6000 208.4000 288.4000 ;
	    RECT 209.2000 287.6000 210.0000 288.4000 ;
	    RECT 209.3000 286.3000 209.9000 287.6000 ;
	    RECT 206.1000 285.7000 209.9000 286.3000 ;
	    RECT 206.1000 284.4000 206.7000 285.7000 ;
	    RECT 206.0000 283.6000 206.8000 284.4000 ;
	    RECT 207.6000 283.6000 208.4000 284.4000 ;
	    RECT 206.0000 281.6000 206.8000 282.4000 ;
	    RECT 206.1000 278.4000 206.7000 281.6000 ;
	    RECT 206.0000 277.6000 206.8000 278.4000 ;
	    RECT 199.7000 271.7000 201.9000 272.3000 ;
	    RECT 186.8000 269.6000 187.6000 270.4000 ;
	    RECT 190.0000 269.6000 190.8000 270.4000 ;
	    RECT 196.4000 269.6000 197.2000 270.4000 ;
	    RECT 198.0000 269.6000 198.8000 270.4000 ;
	    RECT 178.8000 268.3000 179.6000 268.4000 ;
	    RECT 178.8000 267.7000 184.3000 268.3000 ;
	    RECT 178.8000 267.6000 179.6000 267.7000 ;
	    RECT 177.2000 265.6000 178.0000 266.4000 ;
	    RECT 182.0000 265.6000 182.8000 266.4000 ;
	    RECT 175.6000 261.6000 176.4000 262.4000 ;
	    RECT 177.3000 258.4000 177.9000 265.6000 ;
	    RECT 182.1000 258.4000 182.7000 265.6000 ;
	    RECT 183.7000 264.3000 184.3000 267.7000 ;
	    RECT 185.2000 267.6000 186.0000 268.4000 ;
	    RECT 185.3000 266.4000 185.9000 267.6000 ;
	    RECT 185.2000 265.6000 186.0000 266.4000 ;
	    RECT 188.4000 265.6000 189.2000 266.4000 ;
	    RECT 186.8000 264.3000 187.6000 264.4000 ;
	    RECT 183.7000 263.7000 187.6000 264.3000 ;
	    RECT 186.8000 263.6000 187.6000 263.7000 ;
	    RECT 188.5000 258.4000 189.1000 265.6000 ;
	    RECT 172.4000 257.6000 173.2000 258.4000 ;
	    RECT 177.2000 257.6000 178.0000 258.4000 ;
	    RECT 182.0000 257.6000 182.8000 258.4000 ;
	    RECT 188.4000 257.6000 189.2000 258.4000 ;
	    RECT 170.8000 255.6000 171.6000 256.4000 ;
	    RECT 183.6000 255.6000 184.4000 256.4000 ;
	    RECT 170.9000 252.4000 171.5000 255.6000 ;
	    RECT 190.1000 254.4000 190.7000 269.6000 ;
	    RECT 191.6000 267.6000 192.4000 268.4000 ;
	    RECT 191.7000 266.4000 192.3000 267.6000 ;
	    RECT 198.1000 266.4000 198.7000 269.6000 ;
	    RECT 199.7000 268.4000 200.3000 271.7000 ;
	    RECT 207.7000 270.4000 208.3000 283.6000 ;
	    RECT 210.9000 278.4000 211.5000 289.7000 ;
	    RECT 214.1000 286.4000 214.7000 291.6000 ;
	    RECT 214.0000 285.6000 214.8000 286.4000 ;
	    RECT 214.1000 282.4000 214.7000 285.6000 ;
	    RECT 214.0000 281.6000 214.8000 282.4000 ;
	    RECT 210.8000 277.6000 211.6000 278.4000 ;
	    RECT 209.2000 275.6000 210.0000 276.4000 ;
	    RECT 209.3000 272.4000 209.9000 275.6000 ;
	    RECT 209.2000 271.6000 210.0000 272.4000 ;
	    RECT 210.9000 271.7000 214.7000 272.3000 ;
	    RECT 202.8000 270.3000 203.6000 270.4000 ;
	    RECT 201.3000 269.7000 203.6000 270.3000 ;
	    RECT 199.6000 267.6000 200.4000 268.4000 ;
	    RECT 191.6000 265.6000 192.4000 266.4000 ;
	    RECT 198.0000 265.6000 198.8000 266.4000 ;
	    RECT 199.6000 265.6000 200.4000 266.4000 ;
	    RECT 194.8000 261.6000 195.6000 262.4000 ;
	    RECT 193.2000 257.6000 194.0000 258.4000 ;
	    RECT 172.4000 253.6000 173.2000 254.4000 ;
	    RECT 182.0000 253.6000 182.8000 254.4000 ;
	    RECT 190.0000 253.6000 190.8000 254.4000 ;
	    RECT 170.8000 251.6000 171.6000 252.4000 ;
	    RECT 172.5000 246.4000 173.1000 253.6000 ;
	    RECT 169.2000 245.6000 170.0000 246.4000 ;
	    RECT 172.4000 245.6000 173.2000 246.4000 ;
	    RECT 182.1000 244.4000 182.7000 253.6000 ;
	    RECT 186.8000 251.6000 187.6000 252.4000 ;
	    RECT 164.4000 243.6000 165.2000 244.4000 ;
	    RECT 177.2000 243.6000 178.0000 244.4000 ;
	    RECT 182.0000 243.6000 182.8000 244.4000 ;
	    RECT 161.2000 237.6000 162.0000 238.4000 ;
	    RECT 164.5000 230.4000 165.1000 243.6000 ;
	    RECT 177.3000 233.7000 181.1000 234.3000 ;
	    RECT 177.3000 232.3000 177.9000 233.7000 ;
	    RECT 175.7000 231.7000 177.9000 232.3000 ;
	    RECT 158.0000 229.6000 158.8000 230.4000 ;
	    RECT 159.6000 229.6000 160.4000 230.4000 ;
	    RECT 162.8000 229.6000 163.6000 230.4000 ;
	    RECT 164.4000 229.6000 165.2000 230.4000 ;
	    RECT 167.6000 229.6000 168.4000 230.4000 ;
	    RECT 175.7000 230.3000 176.3000 231.7000 ;
	    RECT 178.8000 231.6000 179.6000 232.4000 ;
	    RECT 178.9000 230.4000 179.5000 231.6000 ;
	    RECT 180.5000 230.4000 181.1000 233.7000 ;
	    RECT 182.1000 230.4000 182.7000 243.6000 ;
	    RECT 174.1000 229.7000 176.3000 230.3000 ;
	    RECT 156.4000 213.6000 157.2000 214.4000 ;
	    RECT 158.1000 212.4000 158.7000 229.6000 ;
	    RECT 162.9000 218.4000 163.5000 229.6000 ;
	    RECT 174.1000 228.4000 174.7000 229.7000 ;
	    RECT 177.2000 229.6000 178.0000 230.4000 ;
	    RECT 178.8000 229.6000 179.6000 230.4000 ;
	    RECT 180.4000 229.6000 181.2000 230.4000 ;
	    RECT 182.0000 229.6000 182.8000 230.4000 ;
	    RECT 166.0000 227.6000 166.8000 228.4000 ;
	    RECT 174.0000 227.6000 174.8000 228.4000 ;
	    RECT 175.6000 227.6000 176.4000 228.4000 ;
	    RECT 177.2000 227.6000 178.0000 228.4000 ;
	    RECT 166.1000 226.4000 166.7000 227.6000 ;
	    RECT 166.0000 225.6000 166.8000 226.4000 ;
	    RECT 174.0000 226.3000 174.8000 226.4000 ;
	    RECT 172.5000 225.7000 174.8000 226.3000 ;
	    RECT 167.6000 223.6000 168.4000 224.4000 ;
	    RECT 159.6000 217.6000 160.4000 218.4000 ;
	    RECT 162.8000 217.6000 163.6000 218.4000 ;
	    RECT 159.7000 212.4000 160.3000 217.6000 ;
	    RECT 148.4000 211.6000 149.2000 212.4000 ;
	    RECT 154.8000 211.6000 155.6000 212.4000 ;
	    RECT 158.0000 211.6000 158.8000 212.4000 ;
	    RECT 159.6000 211.6000 160.4000 212.4000 ;
	    RECT 161.2000 211.6000 162.0000 212.4000 ;
	    RECT 148.4000 209.6000 149.2000 210.4000 ;
	    RECT 154.8000 209.6000 155.6000 210.4000 ;
	    RECT 161.3000 210.3000 161.9000 211.6000 ;
	    RECT 159.7000 209.7000 161.9000 210.3000 ;
	    RECT 148.5000 208.4000 149.1000 209.6000 ;
	    RECT 146.8000 207.6000 147.6000 208.4000 ;
	    RECT 148.4000 207.6000 149.2000 208.4000 ;
	    RECT 153.2000 203.6000 154.0000 204.4000 ;
	    RECT 148.4000 201.6000 149.2000 202.4000 ;
	    RECT 142.0000 192.3000 142.8000 192.4000 ;
	    RECT 140.5000 191.7000 142.8000 192.3000 ;
	    RECT 134.0000 189.6000 134.8000 190.4000 ;
	    RECT 137.2000 189.6000 138.0000 190.4000 ;
	    RECT 138.8000 189.6000 139.6000 190.4000 ;
	    RECT 113.2000 187.6000 114.0000 188.4000 ;
	    RECT 119.6000 187.6000 120.4000 188.4000 ;
	    RECT 124.4000 187.6000 125.2000 188.4000 ;
	    RECT 127.6000 187.6000 128.4000 188.4000 ;
	    RECT 130.8000 187.6000 131.6000 188.4000 ;
	    RECT 132.4000 187.6000 133.2000 188.4000 ;
	    RECT 138.8000 188.3000 139.6000 188.4000 ;
	    RECT 140.5000 188.3000 141.1000 191.7000 ;
	    RECT 142.0000 191.6000 142.8000 191.7000 ;
	    RECT 145.2000 191.6000 146.0000 192.4000 ;
	    RECT 146.8000 191.6000 147.6000 192.4000 ;
	    RECT 142.0000 189.6000 142.8000 190.4000 ;
	    RECT 142.1000 188.4000 142.7000 189.6000 ;
	    RECT 146.9000 188.4000 147.5000 191.6000 ;
	    RECT 148.5000 190.4000 149.1000 201.6000 ;
	    RECT 150.0000 195.6000 150.8000 196.4000 ;
	    RECT 148.4000 189.6000 149.2000 190.4000 ;
	    RECT 151.6000 189.6000 152.4000 190.4000 ;
	    RECT 138.8000 187.7000 141.1000 188.3000 ;
	    RECT 138.8000 187.6000 139.6000 187.7000 ;
	    RECT 142.0000 187.6000 142.8000 188.4000 ;
	    RECT 146.8000 187.6000 147.6000 188.4000 ;
	    RECT 119.7000 184.4000 120.3000 187.6000 ;
	    RECT 119.6000 183.6000 120.4000 184.4000 ;
	    RECT 127.7000 180.4000 128.3000 187.6000 ;
	    RECT 129.2000 185.6000 130.0000 186.4000 ;
	    RECT 122.8000 179.6000 123.6000 180.4000 ;
	    RECT 127.6000 179.6000 128.4000 180.4000 ;
	    RECT 122.9000 178.4000 123.5000 179.6000 ;
	    RECT 121.2000 177.6000 122.0000 178.4000 ;
	    RECT 122.8000 177.6000 123.6000 178.4000 ;
	    RECT 121.3000 174.4000 121.9000 177.6000 ;
	    RECT 111.6000 173.6000 112.4000 174.4000 ;
	    RECT 121.2000 173.6000 122.0000 174.4000 ;
	    RECT 111.6000 171.6000 112.4000 172.4000 ;
	    RECT 113.2000 171.6000 114.0000 172.4000 ;
	    RECT 114.8000 171.6000 115.6000 172.4000 ;
	    RECT 102.0000 161.6000 102.8000 162.4000 ;
	    RECT 102.1000 152.4000 102.7000 161.6000 ;
	    RECT 111.7000 154.4000 112.3000 171.6000 ;
	    RECT 113.3000 168.4000 113.9000 171.6000 ;
	    RECT 118.0000 169.6000 118.8000 170.4000 ;
	    RECT 118.1000 168.4000 118.7000 169.6000 ;
	    RECT 113.2000 167.6000 114.0000 168.4000 ;
	    RECT 118.0000 167.6000 118.8000 168.4000 ;
	    RECT 111.6000 153.6000 112.4000 154.4000 ;
	    RECT 102.0000 151.6000 102.8000 152.4000 ;
	    RECT 108.4000 151.6000 109.2000 152.4000 ;
	    RECT 100.4000 145.6000 101.2000 146.4000 ;
	    RECT 102.1000 144.4000 102.7000 151.6000 ;
	    RECT 105.2000 149.6000 106.0000 150.4000 ;
	    RECT 103.6000 147.6000 104.4000 148.4000 ;
	    RECT 102.0000 143.6000 102.8000 144.4000 ;
	    RECT 95.6000 141.6000 96.4000 142.4000 ;
	    RECT 95.7000 134.4000 96.3000 141.6000 ;
	    RECT 95.6000 133.6000 96.4000 134.4000 ;
	    RECT 97.2000 133.6000 98.0000 134.4000 ;
	    RECT 94.0000 131.6000 94.8000 132.4000 ;
	    RECT 94.0000 127.6000 94.8000 128.4000 ;
	    RECT 92.4000 117.6000 93.2000 118.4000 ;
	    RECT 84.5000 115.7000 86.7000 116.3000 ;
	    RECT 79.6000 113.6000 80.4000 114.4000 ;
	    RECT 84.5000 112.4000 85.1000 115.7000 ;
	    RECT 87.6000 115.6000 88.4000 116.4000 ;
	    RECT 84.4000 111.6000 85.2000 112.4000 ;
	    RECT 86.0000 111.6000 86.8000 112.4000 ;
	    RECT 84.5000 110.4000 85.1000 111.6000 ;
	    RECT 84.4000 109.6000 85.2000 110.4000 ;
	    RECT 86.1000 108.4000 86.7000 111.6000 ;
	    RECT 89.2000 109.6000 90.0000 110.4000 ;
	    RECT 94.0000 109.6000 94.8000 110.4000 ;
	    RECT 95.6000 109.6000 96.4000 110.4000 ;
	    RECT 78.0000 107.6000 78.8000 108.4000 ;
	    RECT 86.0000 107.6000 86.8000 108.4000 ;
	    RECT 90.8000 107.6000 91.6000 108.4000 ;
	    RECT 73.3000 101.7000 75.5000 102.3000 ;
	    RECT 68.4000 97.6000 69.2000 98.4000 ;
	    RECT 70.1000 96.4000 70.7000 101.6000 ;
	    RECT 65.2000 95.7000 67.5000 96.3000 ;
	    RECT 65.2000 95.6000 66.0000 95.7000 ;
	    RECT 70.0000 95.6000 70.8000 96.4000 ;
	    RECT 63.6000 93.6000 64.4000 94.4000 ;
	    RECT 73.2000 93.6000 74.0000 94.4000 ;
	    RECT 49.2000 91.6000 50.0000 92.4000 ;
	    RECT 52.4000 91.6000 53.2000 92.4000 ;
	    RECT 58.8000 91.6000 59.6000 92.4000 ;
	    RECT 63.6000 91.6000 64.4000 92.4000 ;
	    RECT 68.4000 91.6000 69.2000 92.4000 ;
	    RECT 73.2000 91.6000 74.0000 92.4000 ;
	    RECT 49.3000 90.4000 49.9000 91.6000 ;
	    RECT 49.2000 89.6000 50.0000 90.4000 ;
	    RECT 55.6000 87.6000 56.4000 88.4000 ;
	    RECT 50.8000 73.6000 51.6000 74.4000 ;
	    RECT 50.9000 72.4000 51.5000 73.6000 ;
	    RECT 39.6000 71.6000 40.4000 72.4000 ;
	    RECT 46.0000 71.6000 46.8000 72.4000 ;
	    RECT 50.8000 71.6000 51.6000 72.4000 ;
	    RECT 46.1000 70.4000 46.7000 71.6000 ;
	    RECT 42.8000 69.6000 43.6000 70.4000 ;
	    RECT 46.0000 69.6000 46.8000 70.4000 ;
	    RECT 52.4000 69.6000 53.2000 70.4000 ;
	    RECT 42.9000 66.4000 43.5000 69.6000 ;
	    RECT 55.7000 68.4000 56.3000 87.6000 ;
	    RECT 62.0000 83.6000 62.8000 84.4000 ;
	    RECT 65.2000 83.6000 66.0000 84.4000 ;
	    RECT 57.2000 70.3000 58.0000 70.4000 ;
	    RECT 57.2000 69.7000 59.5000 70.3000 ;
	    RECT 57.2000 69.6000 58.0000 69.7000 ;
	    RECT 44.4000 67.6000 45.2000 68.4000 ;
	    RECT 55.6000 67.6000 56.4000 68.4000 ;
	    RECT 38.0000 65.6000 38.8000 66.4000 ;
	    RECT 42.8000 65.6000 43.6000 66.4000 ;
	    RECT 36.4000 53.6000 37.2000 54.4000 ;
	    RECT 38.0000 50.2000 38.8000 55.8000 ;
	    RECT 42.9000 52.4000 43.5000 65.6000 ;
	    RECT 44.5000 64.4000 45.1000 67.6000 ;
	    RECT 54.0000 65.6000 54.8000 66.4000 ;
	    RECT 44.4000 63.6000 45.2000 64.4000 ;
	    RECT 49.2000 63.6000 50.0000 64.4000 ;
	    RECT 44.5000 54.4000 45.1000 63.6000 ;
	    RECT 44.4000 53.6000 45.2000 54.4000 ;
	    RECT 42.8000 51.6000 43.6000 52.4000 ;
	    RECT 42.8000 49.6000 43.6000 50.4000 ;
	    RECT 39.6000 47.6000 40.4000 48.4000 ;
	    RECT 42.8000 47.6000 43.6000 48.4000 ;
	    RECT 42.9000 38.4000 43.5000 47.6000 ;
	    RECT 42.8000 37.6000 43.6000 38.4000 ;
	    RECT 28.4000 29.6000 29.2000 30.4000 ;
	    RECT 26.8000 27.6000 27.6000 28.4000 ;
	    RECT 33.2000 24.2000 34.0000 35.8000 ;
	    RECT 39.6000 31.6000 40.4000 32.4000 ;
	    RECT 34.8000 27.6000 35.6000 28.4000 ;
	    RECT 33.2000 19.6000 34.0000 20.4000 ;
	    RECT 22.0000 13.6000 22.8000 14.4000 ;
	    RECT 17.2000 11.6000 18.0000 12.4000 ;
	    RECT 23.6000 11.6000 24.4000 12.6000 ;
	    RECT 25.2000 6.2000 26.0000 17.8000 ;
	    RECT 28.4000 10.2000 29.2000 15.8000 ;
	    RECT 33.3000 12.4000 33.9000 19.6000 ;
	    RECT 34.9000 14.4000 35.5000 27.6000 ;
	    RECT 34.8000 13.6000 35.6000 14.4000 ;
	    RECT 39.7000 12.4000 40.3000 31.6000 ;
	    RECT 42.8000 29.6000 43.6000 30.4000 ;
	    RECT 42.9000 20.4000 43.5000 29.6000 ;
	    RECT 44.5000 28.4000 45.1000 53.6000 ;
	    RECT 46.0000 51.6000 46.8000 52.4000 ;
	    RECT 46.0000 49.6000 46.8000 50.4000 ;
	    RECT 46.1000 48.4000 46.7000 49.6000 ;
	    RECT 46.0000 47.6000 46.8000 48.4000 ;
	    RECT 47.6000 45.6000 48.4000 46.4000 ;
	    RECT 46.0000 33.6000 46.8000 34.4000 ;
	    RECT 47.7000 30.4000 48.3000 45.6000 ;
	    RECT 49.3000 38.4000 49.9000 63.6000 ;
	    RECT 52.4000 55.6000 53.2000 56.4000 ;
	    RECT 50.8000 53.6000 51.6000 54.4000 ;
	    RECT 50.8000 51.6000 51.6000 52.4000 ;
	    RECT 52.4000 49.6000 53.2000 50.4000 ;
	    RECT 49.2000 37.6000 50.0000 38.4000 ;
	    RECT 49.3000 30.4000 49.9000 37.6000 ;
	    RECT 54.1000 30.4000 54.7000 65.6000 ;
	    RECT 58.9000 64.4000 59.5000 69.7000 ;
	    RECT 58.8000 63.6000 59.6000 64.4000 ;
	    RECT 55.6000 57.6000 56.4000 58.4000 ;
	    RECT 55.7000 52.4000 56.3000 57.6000 ;
	    RECT 62.1000 54.4000 62.7000 83.6000 ;
	    RECT 63.6000 73.6000 64.4000 74.4000 ;
	    RECT 63.7000 54.4000 64.3000 73.6000 ;
	    RECT 65.3000 54.4000 65.9000 83.6000 ;
	    RECT 68.5000 80.4000 69.1000 91.6000 ;
	    RECT 74.9000 90.4000 75.5000 101.7000 ;
	    RECT 78.1000 92.4000 78.7000 107.6000 ;
	    RECT 79.6000 105.6000 80.4000 106.4000 ;
	    RECT 79.7000 94.4000 80.3000 105.6000 ;
	    RECT 79.6000 93.6000 80.4000 94.4000 ;
	    RECT 78.0000 91.6000 78.8000 92.4000 ;
	    RECT 74.8000 89.6000 75.6000 90.4000 ;
	    RECT 74.9000 86.3000 75.5000 89.6000 ;
	    RECT 79.7000 88.3000 80.3000 93.6000 ;
	    RECT 81.2000 90.2000 82.0000 95.8000 ;
	    RECT 82.8000 91.6000 83.6000 92.4000 ;
	    RECT 82.9000 88.4000 83.5000 91.6000 ;
	    RECT 79.7000 87.7000 81.9000 88.3000 ;
	    RECT 73.3000 85.7000 75.5000 86.3000 ;
	    RECT 71.6000 83.6000 72.4000 84.4000 ;
	    RECT 68.4000 79.6000 69.2000 80.4000 ;
	    RECT 71.7000 74.4000 72.3000 83.6000 ;
	    RECT 71.6000 73.6000 72.4000 74.4000 ;
	    RECT 71.6000 71.6000 72.4000 72.4000 ;
	    RECT 68.4000 63.6000 69.2000 64.4000 ;
	    RECT 57.2000 53.6000 58.0000 54.4000 ;
	    RECT 58.8000 53.6000 59.6000 54.4000 ;
	    RECT 62.0000 53.6000 62.8000 54.4000 ;
	    RECT 63.6000 53.6000 64.4000 54.4000 ;
	    RECT 65.2000 53.6000 66.0000 54.4000 ;
	    RECT 55.6000 51.6000 56.4000 52.4000 ;
	    RECT 58.9000 52.3000 59.5000 53.6000 ;
	    RECT 68.5000 52.4000 69.1000 63.6000 ;
	    RECT 57.3000 51.7000 59.5000 52.3000 ;
	    RECT 57.3000 36.4000 57.9000 51.7000 ;
	    RECT 62.0000 51.6000 62.8000 52.4000 ;
	    RECT 68.4000 51.6000 69.2000 52.4000 ;
	    RECT 58.8000 49.6000 59.6000 50.4000 ;
	    RECT 58.9000 46.4000 59.5000 49.6000 ;
	    RECT 62.1000 48.4000 62.7000 51.6000 ;
	    RECT 62.0000 47.6000 62.8000 48.4000 ;
	    RECT 58.8000 45.6000 59.6000 46.4000 ;
	    RECT 70.0000 46.2000 70.8000 57.8000 ;
	    RECT 71.7000 56.4000 72.3000 71.6000 ;
	    RECT 73.3000 56.4000 73.9000 85.7000 ;
	    RECT 74.8000 83.6000 75.6000 84.4000 ;
	    RECT 74.9000 78.4000 75.5000 83.6000 ;
	    RECT 78.0000 81.6000 78.8000 82.4000 ;
	    RECT 74.8000 77.6000 75.6000 78.4000 ;
	    RECT 74.8000 69.6000 75.6000 70.4000 ;
	    RECT 74.9000 66.4000 75.5000 69.6000 ;
	    RECT 76.4000 67.6000 77.2000 68.4000 ;
	    RECT 74.8000 65.6000 75.6000 66.4000 ;
	    RECT 76.5000 62.4000 77.1000 67.6000 ;
	    RECT 76.4000 61.6000 77.2000 62.4000 ;
	    RECT 71.6000 55.6000 72.4000 56.4000 ;
	    RECT 73.2000 55.6000 74.0000 56.4000 ;
	    RECT 65.2000 43.6000 66.0000 44.4000 ;
	    RECT 57.2000 35.6000 58.0000 36.4000 ;
	    RECT 62.0000 33.6000 62.8000 34.4000 ;
	    RECT 57.2000 31.6000 58.0000 32.4000 ;
	    RECT 47.6000 29.6000 48.4000 30.4000 ;
	    RECT 49.2000 29.6000 50.0000 30.4000 ;
	    RECT 54.0000 29.6000 54.8000 30.4000 ;
	    RECT 44.4000 27.6000 45.2000 28.4000 ;
	    RECT 50.8000 27.6000 51.6000 28.4000 ;
	    RECT 42.8000 19.6000 43.6000 20.4000 ;
	    RECT 44.4000 17.6000 45.2000 18.4000 ;
	    RECT 44.5000 12.4000 45.1000 17.6000 ;
	    RECT 46.0000 15.6000 46.8000 16.4000 ;
	    RECT 46.1000 14.4000 46.7000 15.6000 ;
	    RECT 46.0000 13.6000 46.8000 14.4000 ;
	    RECT 54.1000 12.4000 54.7000 29.6000 ;
	    RECT 57.3000 28.3000 57.9000 31.6000 ;
	    RECT 62.1000 30.4000 62.7000 33.6000 ;
	    RECT 65.3000 30.4000 65.9000 43.6000 ;
	    RECT 62.0000 29.6000 62.8000 30.4000 ;
	    RECT 63.6000 29.6000 64.4000 30.4000 ;
	    RECT 65.2000 29.6000 66.0000 30.4000 ;
	    RECT 63.7000 28.4000 64.3000 29.6000 ;
	    RECT 55.7000 27.7000 57.9000 28.3000 ;
	    RECT 55.7000 16.4000 56.3000 27.7000 ;
	    RECT 60.4000 27.6000 61.2000 28.4000 ;
	    RECT 63.6000 27.6000 64.4000 28.4000 ;
	    RECT 71.6000 27.6000 72.4000 28.4000 ;
	    RECT 55.6000 15.6000 56.4000 16.4000 ;
	    RECT 33.2000 11.6000 34.0000 12.4000 ;
	    RECT 39.6000 11.6000 40.4000 12.4000 ;
	    RECT 41.2000 11.6000 42.0000 12.4000 ;
	    RECT 44.4000 11.6000 45.2000 12.4000 ;
	    RECT 50.8000 11.6000 51.6000 12.4000 ;
	    RECT 54.0000 11.6000 54.8000 12.4000 ;
	    RECT 30.0000 9.6000 30.8000 10.4000 ;
	    RECT 33.2000 9.6000 34.0000 10.4000 ;
	    RECT 41.2000 9.6000 42.0000 10.4000 ;
	    RECT 50.9000 8.3000 51.5000 11.6000 ;
	    RECT 52.4000 8.3000 53.2000 8.4000 ;
	    RECT 50.9000 7.7000 53.2000 8.3000 ;
	    RECT 52.4000 7.6000 53.2000 7.7000 ;
	    RECT 57.2000 6.2000 58.0000 17.8000 ;
	    RECT 58.8000 13.6000 59.6000 14.4000 ;
	    RECT 58.9000 12.4000 59.5000 13.6000 ;
	    RECT 60.5000 12.4000 61.1000 27.6000 ;
	    RECT 70.0000 23.6000 70.8000 24.4000 ;
	    RECT 58.8000 11.6000 59.6000 12.4000 ;
	    RECT 60.4000 11.6000 61.2000 12.4000 ;
	    RECT 66.8000 6.2000 67.6000 17.8000 ;
	    RECT 70.0000 10.2000 70.8000 15.8000 ;
	    RECT 71.7000 14.4000 72.3000 27.6000 ;
	    RECT 74.8000 24.2000 75.6000 35.8000 ;
	    RECT 76.5000 28.4000 77.1000 61.6000 ;
	    RECT 78.1000 52.6000 78.7000 81.6000 ;
	    RECT 81.3000 78.4000 81.9000 87.7000 ;
	    RECT 82.8000 87.6000 83.6000 88.4000 ;
	    RECT 84.4000 86.2000 85.2000 97.8000 ;
	    RECT 87.6000 97.6000 88.4000 98.4000 ;
	    RECT 87.7000 94.4000 88.3000 97.6000 ;
	    RECT 87.6000 93.6000 88.4000 94.4000 ;
	    RECT 89.2000 93.6000 90.0000 94.4000 ;
	    RECT 81.2000 77.6000 82.0000 78.4000 ;
	    RECT 81.3000 72.4000 81.9000 77.6000 ;
	    RECT 81.2000 71.6000 82.0000 72.4000 ;
	    RECT 81.2000 65.6000 82.0000 66.4000 ;
	    RECT 82.8000 66.2000 83.6000 71.8000 ;
	    RECT 84.4000 67.6000 85.2000 68.4000 ;
	    RECT 84.5000 66.4000 85.1000 67.6000 ;
	    RECT 84.4000 65.6000 85.2000 66.4000 ;
	    RECT 78.0000 51.8000 78.8000 52.6000 ;
	    RECT 78.1000 51.7000 78.7000 51.8000 ;
	    RECT 79.6000 46.2000 80.4000 57.8000 ;
	    RECT 81.3000 54.4000 81.9000 65.6000 ;
	    RECT 86.0000 64.2000 86.8000 75.8000 ;
	    RECT 87.7000 68.4000 88.3000 93.6000 ;
	    RECT 89.3000 92.4000 89.9000 93.6000 ;
	    RECT 89.2000 91.6000 90.0000 92.4000 ;
	    RECT 90.9000 86.4000 91.5000 107.6000 ;
	    RECT 94.1000 102.4000 94.7000 109.6000 ;
	    RECT 97.3000 106.4000 97.9000 133.6000 ;
	    RECT 98.8000 131.6000 99.6000 132.4000 ;
	    RECT 100.4000 131.6000 101.2000 132.4000 ;
	    RECT 98.9000 128.4000 99.5000 131.6000 ;
	    RECT 102.0000 129.6000 102.8000 130.4000 ;
	    RECT 98.8000 127.6000 99.6000 128.4000 ;
	    RECT 103.7000 124.3000 104.3000 147.6000 ;
	    RECT 105.3000 146.4000 105.9000 149.6000 ;
	    RECT 106.8000 147.6000 107.6000 148.4000 ;
	    RECT 105.2000 145.6000 106.0000 146.4000 ;
	    RECT 106.9000 124.4000 107.5000 147.6000 ;
	    RECT 108.5000 142.4000 109.1000 151.6000 ;
	    RECT 111.6000 149.6000 112.4000 150.4000 ;
	    RECT 116.4000 149.6000 117.2000 150.4000 ;
	    RECT 108.4000 141.6000 109.2000 142.4000 ;
	    RECT 110.0000 141.6000 110.8000 142.4000 ;
	    RECT 110.1000 136.4000 110.7000 141.6000 ;
	    RECT 110.0000 135.6000 110.8000 136.4000 ;
	    RECT 111.7000 132.4000 112.3000 149.6000 ;
	    RECT 116.5000 144.4000 117.1000 149.6000 ;
	    RECT 118.1000 144.4000 118.7000 167.6000 ;
	    RECT 121.3000 150.4000 121.9000 173.6000 ;
	    RECT 127.6000 166.2000 128.4000 177.8000 ;
	    RECT 129.3000 170.4000 129.9000 185.6000 ;
	    RECT 132.5000 180.4000 133.1000 187.6000 ;
	    RECT 134.0000 183.6000 134.8000 184.4000 ;
	    RECT 132.4000 179.6000 133.2000 180.4000 ;
	    RECT 132.4000 173.6000 133.2000 174.4000 ;
	    RECT 135.6000 171.6000 136.4000 172.6000 ;
	    RECT 129.2000 169.6000 130.0000 170.4000 ;
	    RECT 124.4000 163.6000 125.2000 164.4000 ;
	    RECT 121.2000 149.6000 122.0000 150.4000 ;
	    RECT 122.8000 149.6000 123.6000 150.4000 ;
	    RECT 124.5000 146.4000 125.1000 163.6000 ;
	    RECT 127.6000 159.6000 128.4000 160.4000 ;
	    RECT 127.7000 150.4000 128.3000 159.6000 ;
	    RECT 127.6000 149.6000 128.4000 150.4000 ;
	    RECT 129.3000 146.4000 129.9000 169.6000 ;
	    RECT 137.2000 166.2000 138.0000 177.8000 ;
	    RECT 140.4000 170.2000 141.2000 175.8000 ;
	    RECT 142.1000 174.4000 142.7000 187.6000 ;
	    RECT 146.9000 180.4000 147.5000 187.6000 ;
	    RECT 151.7000 184.4000 152.3000 189.6000 ;
	    RECT 151.6000 183.6000 152.4000 184.4000 ;
	    RECT 153.3000 182.3000 153.9000 203.6000 ;
	    RECT 154.9000 192.4000 155.5000 209.6000 ;
	    RECT 158.0000 207.6000 158.8000 208.4000 ;
	    RECT 156.4000 203.6000 157.2000 204.4000 ;
	    RECT 156.5000 202.4000 157.1000 203.6000 ;
	    RECT 156.4000 201.6000 157.2000 202.4000 ;
	    RECT 156.4000 193.6000 157.2000 194.4000 ;
	    RECT 154.8000 191.6000 155.6000 192.4000 ;
	    RECT 154.8000 185.6000 155.6000 186.4000 ;
	    RECT 151.7000 181.7000 153.9000 182.3000 ;
	    RECT 146.8000 180.3000 147.6000 180.4000 ;
	    RECT 146.8000 179.7000 149.1000 180.3000 ;
	    RECT 146.8000 179.6000 147.6000 179.7000 ;
	    RECT 142.0000 173.6000 142.8000 174.4000 ;
	    RECT 146.8000 173.6000 147.6000 174.4000 ;
	    RECT 146.9000 172.4000 147.5000 173.6000 ;
	    RECT 146.8000 171.6000 147.6000 172.4000 ;
	    RECT 145.2000 170.3000 146.0000 170.4000 ;
	    RECT 145.2000 169.7000 147.5000 170.3000 ;
	    RECT 145.2000 169.6000 146.0000 169.7000 ;
	    RECT 140.4000 167.6000 141.2000 168.4000 ;
	    RECT 135.6000 155.6000 136.4000 156.4000 ;
	    RECT 135.6000 153.6000 136.4000 154.4000 ;
	    RECT 130.8000 151.6000 131.6000 152.4000 ;
	    RECT 134.0000 151.6000 134.8000 152.4000 ;
	    RECT 134.1000 150.4000 134.7000 151.6000 ;
	    RECT 132.4000 149.6000 133.2000 150.4000 ;
	    RECT 134.0000 149.6000 134.8000 150.4000 ;
	    RECT 124.4000 145.6000 125.2000 146.4000 ;
	    RECT 129.2000 145.6000 130.0000 146.4000 ;
	    RECT 132.5000 146.3000 133.1000 149.6000 ;
	    RECT 134.0000 148.3000 134.8000 148.4000 ;
	    RECT 135.7000 148.3000 136.3000 153.6000 ;
	    RECT 140.5000 152.4000 141.1000 167.6000 ;
	    RECT 143.6000 155.6000 144.4000 156.4000 ;
	    RECT 140.4000 151.6000 141.2000 152.4000 ;
	    RECT 142.0000 151.6000 142.8000 152.4000 ;
	    RECT 134.0000 147.7000 136.3000 148.3000 ;
	    RECT 134.0000 147.6000 134.8000 147.7000 ;
	    RECT 132.5000 145.7000 134.7000 146.3000 ;
	    RECT 116.4000 143.6000 117.2000 144.4000 ;
	    RECT 118.0000 143.6000 118.8000 144.4000 ;
	    RECT 119.6000 143.6000 120.4000 144.4000 ;
	    RECT 126.0000 143.6000 126.8000 144.4000 ;
	    RECT 113.2000 135.6000 114.0000 136.4000 ;
	    RECT 110.0000 131.6000 110.8000 132.4000 ;
	    RECT 111.6000 131.6000 112.4000 132.4000 ;
	    RECT 102.1000 123.7000 104.3000 124.3000 ;
	    RECT 98.8000 113.6000 99.6000 114.4000 ;
	    RECT 98.9000 110.4000 99.5000 113.6000 ;
	    RECT 98.8000 109.6000 99.6000 110.4000 ;
	    RECT 100.4000 109.6000 101.2000 110.4000 ;
	    RECT 97.2000 105.6000 98.0000 106.4000 ;
	    RECT 100.5000 102.4000 101.1000 109.6000 ;
	    RECT 94.0000 101.6000 94.8000 102.4000 ;
	    RECT 98.8000 101.6000 99.6000 102.4000 ;
	    RECT 100.4000 101.6000 101.2000 102.4000 ;
	    RECT 98.9000 98.4000 99.5000 101.6000 ;
	    RECT 90.8000 85.6000 91.6000 86.4000 ;
	    RECT 94.0000 86.2000 94.8000 97.8000 ;
	    RECT 98.8000 97.6000 99.6000 98.4000 ;
	    RECT 98.9000 92.4000 99.5000 97.6000 ;
	    RECT 100.4000 93.6000 101.2000 94.4000 ;
	    RECT 98.8000 91.6000 99.6000 92.4000 ;
	    RECT 100.5000 86.4000 101.1000 93.6000 ;
	    RECT 102.1000 92.4000 102.7000 123.7000 ;
	    RECT 106.8000 123.6000 107.6000 124.4000 ;
	    RECT 111.6000 119.6000 112.4000 120.4000 ;
	    RECT 113.3000 120.3000 113.9000 135.6000 ;
	    RECT 114.8000 133.6000 115.6000 134.4000 ;
	    RECT 114.9000 132.4000 115.5000 133.6000 ;
	    RECT 116.5000 132.4000 117.1000 143.6000 ;
	    RECT 118.0000 133.6000 118.8000 134.4000 ;
	    RECT 114.8000 131.6000 115.6000 132.4000 ;
	    RECT 116.4000 131.6000 117.2000 132.4000 ;
	    RECT 118.1000 130.4000 118.7000 133.6000 ;
	    RECT 118.0000 129.6000 118.8000 130.4000 ;
	    RECT 113.3000 119.7000 115.5000 120.3000 ;
	    RECT 111.7000 116.4000 112.3000 119.6000 ;
	    RECT 113.2000 117.6000 114.0000 118.4000 ;
	    RECT 111.6000 115.6000 112.4000 116.4000 ;
	    RECT 110.0000 109.6000 110.8000 110.4000 ;
	    RECT 108.4000 107.6000 109.2000 108.4000 ;
	    RECT 110.0000 105.6000 110.8000 106.4000 ;
	    RECT 111.6000 105.6000 112.4000 106.4000 ;
	    RECT 103.6000 93.6000 104.4000 94.4000 ;
	    RECT 111.7000 92.4000 112.3000 105.6000 ;
	    RECT 102.0000 91.6000 102.8000 92.4000 ;
	    RECT 111.6000 91.6000 112.4000 92.4000 ;
	    RECT 111.7000 90.4000 112.3000 91.6000 ;
	    RECT 111.6000 89.6000 112.4000 90.4000 ;
	    RECT 100.4000 85.6000 101.2000 86.4000 ;
	    RECT 102.0000 79.6000 102.8000 80.4000 ;
	    RECT 100.4000 77.6000 101.2000 78.4000 ;
	    RECT 102.1000 78.3000 102.7000 79.6000 ;
	    RECT 102.1000 77.7000 104.3000 78.3000 ;
	    RECT 103.7000 76.3000 104.3000 77.7000 ;
	    RECT 92.4000 73.6000 93.2000 74.4000 ;
	    RECT 92.5000 70.4000 93.1000 73.6000 ;
	    RECT 94.0000 71.6000 94.8000 72.4000 ;
	    RECT 92.4000 69.6000 93.2000 70.4000 ;
	    RECT 87.6000 67.6000 88.4000 68.4000 ;
	    RECT 89.2000 57.6000 90.0000 58.4000 ;
	    RECT 81.2000 53.6000 82.0000 54.4000 ;
	    RECT 81.3000 28.4000 81.9000 53.6000 ;
	    RECT 82.8000 50.2000 83.6000 55.8000 ;
	    RECT 84.4000 55.6000 85.2000 56.4000 ;
	    RECT 89.2000 55.6000 90.0000 56.4000 ;
	    RECT 90.8000 55.6000 91.6000 56.4000 ;
	    RECT 87.6000 53.6000 88.4000 54.4000 ;
	    RECT 87.7000 52.4000 88.3000 53.6000 ;
	    RECT 87.6000 51.6000 88.4000 52.4000 ;
	    RECT 89.3000 50.4000 89.9000 55.6000 ;
	    RECT 90.9000 50.4000 91.5000 55.6000 ;
	    RECT 94.1000 54.4000 94.7000 71.6000 ;
	    RECT 95.6000 64.2000 96.4000 75.8000 ;
	    RECT 103.7000 75.7000 107.5000 76.3000 ;
	    RECT 106.9000 74.4000 107.5000 75.7000 ;
	    RECT 105.2000 73.6000 106.0000 74.4000 ;
	    RECT 106.8000 73.6000 107.6000 74.4000 ;
	    RECT 103.6000 71.6000 104.4000 72.4000 ;
	    RECT 103.7000 70.4000 104.3000 71.6000 ;
	    RECT 105.3000 70.4000 105.9000 73.6000 ;
	    RECT 113.3000 72.4000 113.9000 117.6000 ;
	    RECT 114.9000 110.4000 115.5000 119.7000 ;
	    RECT 116.4000 111.6000 117.2000 112.4000 ;
	    RECT 114.8000 109.6000 115.6000 110.4000 ;
	    RECT 116.5000 108.4000 117.1000 111.6000 ;
	    RECT 118.1000 108.4000 118.7000 129.6000 ;
	    RECT 119.7000 116.4000 120.3000 143.6000 ;
	    RECT 121.2000 133.6000 122.0000 134.4000 ;
	    RECT 121.3000 132.4000 121.9000 133.6000 ;
	    RECT 121.2000 131.6000 122.0000 132.4000 ;
	    RECT 121.2000 127.6000 122.0000 128.4000 ;
	    RECT 119.6000 115.6000 120.4000 116.4000 ;
	    RECT 124.4000 113.6000 125.2000 114.4000 ;
	    RECT 121.2000 111.6000 122.0000 112.4000 ;
	    RECT 119.6000 109.6000 120.4000 110.4000 ;
	    RECT 116.4000 107.6000 117.2000 108.4000 ;
	    RECT 118.0000 107.6000 118.8000 108.4000 ;
	    RECT 119.7000 102.4000 120.3000 109.6000 ;
	    RECT 121.3000 108.4000 121.9000 111.6000 ;
	    RECT 124.5000 110.4000 125.1000 113.6000 ;
	    RECT 122.8000 109.6000 123.6000 110.4000 ;
	    RECT 124.4000 109.6000 125.2000 110.4000 ;
	    RECT 121.2000 107.6000 122.0000 108.4000 ;
	    RECT 119.6000 101.6000 120.4000 102.4000 ;
	    RECT 119.6000 97.6000 120.4000 98.4000 ;
	    RECT 118.0000 93.6000 118.8000 94.4000 ;
	    RECT 121.3000 92.4000 121.9000 107.6000 ;
	    RECT 122.8000 101.6000 123.6000 102.4000 ;
	    RECT 116.4000 91.6000 117.2000 92.4000 ;
	    RECT 118.0000 91.6000 118.8000 92.4000 ;
	    RECT 121.2000 91.6000 122.0000 92.4000 ;
	    RECT 114.8000 79.6000 115.6000 80.4000 ;
	    RECT 113.2000 71.6000 114.0000 72.4000 ;
	    RECT 103.6000 69.6000 104.4000 70.4000 ;
	    RECT 105.2000 69.6000 106.0000 70.4000 ;
	    RECT 102.0000 67.6000 102.8000 68.4000 ;
	    RECT 100.4000 57.6000 101.2000 58.4000 ;
	    RECT 100.5000 54.4000 101.1000 57.6000 ;
	    RECT 94.0000 53.6000 94.8000 54.4000 ;
	    RECT 100.4000 53.6000 101.2000 54.4000 ;
	    RECT 105.2000 53.6000 106.0000 54.4000 ;
	    RECT 105.3000 52.4000 105.9000 53.6000 ;
	    RECT 94.0000 51.6000 94.8000 52.4000 ;
	    RECT 97.2000 51.6000 98.0000 52.4000 ;
	    RECT 98.8000 51.6000 99.6000 52.4000 ;
	    RECT 105.2000 51.6000 106.0000 52.4000 ;
	    RECT 106.8000 51.6000 107.6000 52.4000 ;
	    RECT 89.2000 49.6000 90.0000 50.4000 ;
	    RECT 90.8000 49.6000 91.6000 50.4000 ;
	    RECT 92.4000 49.6000 93.2000 50.4000 ;
	    RECT 82.8000 45.6000 83.6000 46.4000 ;
	    RECT 82.9000 30.2000 83.5000 45.6000 ;
	    RECT 92.5000 38.4000 93.1000 49.6000 ;
	    RECT 94.1000 42.3000 94.7000 51.6000 ;
	    RECT 95.6000 49.6000 96.4000 50.4000 ;
	    RECT 97.3000 46.4000 97.9000 51.6000 ;
	    RECT 98.9000 50.4000 99.5000 51.6000 ;
	    RECT 106.9000 50.4000 107.5000 51.6000 ;
	    RECT 98.8000 49.6000 99.6000 50.4000 ;
	    RECT 106.8000 49.6000 107.6000 50.4000 ;
	    RECT 113.2000 49.6000 114.0000 50.4000 ;
	    RECT 113.3000 46.4000 113.9000 49.6000 ;
	    RECT 97.2000 45.6000 98.0000 46.4000 ;
	    RECT 102.0000 45.6000 102.8000 46.4000 ;
	    RECT 113.2000 45.6000 114.0000 46.4000 ;
	    RECT 94.1000 41.7000 96.3000 42.3000 ;
	    RECT 95.7000 38.4000 96.3000 41.7000 ;
	    RECT 92.4000 37.6000 93.2000 38.4000 ;
	    RECT 94.0000 37.6000 94.8000 38.4000 ;
	    RECT 95.6000 37.6000 96.4000 38.4000 ;
	    RECT 82.8000 29.4000 83.6000 30.2000 ;
	    RECT 76.4000 27.6000 77.2000 28.4000 ;
	    RECT 81.2000 27.6000 82.0000 28.4000 ;
	    RECT 79.6000 23.6000 80.4000 24.4000 ;
	    RECT 71.6000 13.6000 72.4000 14.4000 ;
	    RECT 73.2000 11.6000 74.0000 12.4000 ;
	    RECT 76.4000 11.6000 77.2000 12.4000 ;
	    RECT 79.7000 12.3000 80.3000 23.6000 ;
	    RECT 81.3000 14.4000 81.9000 27.6000 ;
	    RECT 84.4000 24.2000 85.2000 35.8000 ;
	    RECT 94.1000 32.4000 94.7000 37.6000 ;
	    RECT 102.1000 36.4000 102.7000 45.6000 ;
	    RECT 111.6000 43.6000 112.4000 44.4000 ;
	    RECT 95.6000 35.6000 96.4000 36.4000 ;
	    RECT 102.0000 35.6000 102.8000 36.4000 ;
	    RECT 95.7000 32.4000 96.3000 35.6000 ;
	    RECT 111.7000 34.4000 112.3000 43.6000 ;
	    RECT 98.8000 33.6000 99.6000 34.4000 ;
	    RECT 111.6000 33.6000 112.4000 34.4000 ;
	    RECT 87.6000 26.2000 88.4000 31.8000 ;
	    RECT 89.2000 31.6000 90.0000 32.4000 ;
	    RECT 94.0000 31.6000 94.8000 32.4000 ;
	    RECT 95.6000 31.6000 96.4000 32.4000 ;
	    RECT 89.3000 24.4000 89.9000 31.6000 ;
	    RECT 94.1000 30.4000 94.7000 31.6000 ;
	    RECT 111.7000 30.4000 112.3000 33.6000 ;
	    RECT 94.0000 29.6000 94.8000 30.4000 ;
	    RECT 98.8000 29.6000 99.6000 30.4000 ;
	    RECT 111.6000 29.6000 112.4000 30.4000 ;
	    RECT 94.0000 27.6000 94.8000 28.4000 ;
	    RECT 89.2000 23.6000 90.0000 24.4000 ;
	    RECT 98.9000 22.4000 99.5000 29.6000 ;
	    RECT 100.4000 27.6000 101.2000 28.4000 ;
	    RECT 100.5000 24.4000 101.1000 27.6000 ;
	    RECT 100.4000 23.6000 101.2000 24.4000 ;
	    RECT 98.8000 21.6000 99.6000 22.4000 ;
	    RECT 113.3000 20.4000 113.9000 45.6000 ;
	    RECT 113.2000 19.6000 114.0000 20.4000 ;
	    RECT 81.2000 13.6000 82.0000 14.4000 ;
	    RECT 81.2000 12.3000 82.0000 12.4000 ;
	    RECT 79.7000 11.7000 82.0000 12.3000 ;
	    RECT 81.2000 11.6000 82.0000 11.7000 ;
	    RECT 76.4000 9.6000 77.2000 10.4000 ;
	    RECT 82.8000 10.2000 83.6000 15.8000 ;
	    RECT 84.4000 13.6000 85.2000 14.4000 ;
	    RECT 86.0000 6.2000 86.8000 17.8000 ;
	    RECT 92.4000 13.6000 93.2000 14.4000 ;
	    RECT 92.5000 12.4000 93.1000 13.6000 ;
	    RECT 92.4000 11.6000 93.2000 12.4000 ;
	    RECT 95.6000 6.2000 96.4000 17.8000 ;
	    RECT 114.9000 16.4000 115.5000 79.6000 ;
	    RECT 118.1000 78.4000 118.7000 91.6000 ;
	    RECT 119.6000 89.6000 120.4000 90.4000 ;
	    RECT 119.7000 84.4000 120.3000 89.6000 ;
	    RECT 119.6000 83.6000 120.4000 84.4000 ;
	    RECT 121.2000 83.6000 122.0000 84.4000 ;
	    RECT 118.0000 77.6000 118.8000 78.4000 ;
	    RECT 118.1000 68.4000 118.7000 77.6000 ;
	    RECT 118.0000 67.6000 118.8000 68.4000 ;
	    RECT 116.4000 59.6000 117.2000 60.4000 ;
	    RECT 116.5000 52.4000 117.1000 59.6000 ;
	    RECT 116.4000 51.6000 117.2000 52.4000 ;
	    RECT 119.6000 43.6000 120.4000 44.4000 ;
	    RECT 118.0000 24.2000 118.8000 35.8000 ;
	    RECT 119.7000 24.4000 120.3000 43.6000 ;
	    RECT 119.6000 23.6000 120.4000 24.4000 ;
	    RECT 119.6000 19.6000 120.4000 20.4000 ;
	    RECT 114.8000 15.6000 115.6000 16.4000 ;
	    RECT 113.2000 13.6000 114.0000 14.4000 ;
	    RECT 118.0000 13.6000 118.8000 14.4000 ;
	    RECT 102.0000 11.6000 102.8000 12.4000 ;
	    RECT 113.2000 11.6000 114.0000 12.4000 ;
	    RECT 100.4000 9.6000 101.2000 10.4000 ;
	    RECT 100.5000 8.4000 101.1000 9.6000 ;
	    RECT 100.4000 8.3000 101.2000 8.4000 ;
	    RECT 102.1000 8.3000 102.7000 11.6000 ;
	    RECT 113.3000 10.4000 113.9000 11.6000 ;
	    RECT 119.7000 10.4000 120.3000 19.6000 ;
	    RECT 121.3000 14.4000 121.9000 83.6000 ;
	    RECT 122.9000 70.3000 123.5000 101.6000 ;
	    RECT 124.4000 94.3000 125.2000 94.4000 ;
	    RECT 126.1000 94.3000 126.7000 143.6000 ;
	    RECT 134.1000 142.4000 134.7000 145.7000 ;
	    RECT 142.1000 142.4000 142.7000 151.6000 ;
	    RECT 143.7000 150.4000 144.3000 155.6000 ;
	    RECT 143.6000 149.6000 144.4000 150.4000 ;
	    RECT 145.2000 149.6000 146.0000 150.4000 ;
	    RECT 145.3000 148.4000 145.9000 149.6000 ;
	    RECT 145.2000 147.6000 146.0000 148.4000 ;
	    RECT 132.4000 141.6000 133.2000 142.4000 ;
	    RECT 134.0000 141.6000 134.8000 142.4000 ;
	    RECT 142.0000 141.6000 142.8000 142.4000 ;
	    RECT 132.5000 140.3000 133.1000 141.6000 ;
	    RECT 132.5000 139.7000 136.3000 140.3000 ;
	    RECT 135.7000 138.4000 136.3000 139.7000 ;
	    RECT 132.4000 137.6000 133.2000 138.4000 ;
	    RECT 135.6000 137.6000 136.4000 138.4000 ;
	    RECT 132.5000 134.4000 133.1000 137.6000 ;
	    RECT 145.3000 136.4000 145.9000 147.6000 ;
	    RECT 143.6000 136.3000 144.4000 136.4000 ;
	    RECT 138.9000 135.7000 144.4000 136.3000 ;
	    RECT 132.4000 133.6000 133.2000 134.4000 ;
	    RECT 134.0000 133.6000 134.8000 134.4000 ;
	    RECT 138.9000 134.3000 139.5000 135.7000 ;
	    RECT 143.6000 135.6000 144.4000 135.7000 ;
	    RECT 145.2000 135.6000 146.0000 136.4000 ;
	    RECT 137.3000 133.7000 139.5000 134.3000 ;
	    RECT 127.6000 132.3000 128.4000 132.4000 ;
	    RECT 127.6000 131.7000 129.9000 132.3000 ;
	    RECT 127.6000 131.6000 128.4000 131.7000 ;
	    RECT 129.3000 130.4000 129.9000 131.7000 ;
	    RECT 130.8000 131.6000 131.6000 132.4000 ;
	    RECT 135.6000 131.6000 136.4000 132.4000 ;
	    RECT 127.6000 129.6000 128.4000 130.4000 ;
	    RECT 129.2000 129.6000 130.0000 130.4000 ;
	    RECT 127.6000 127.6000 128.4000 128.4000 ;
	    RECT 127.7000 118.4000 128.3000 127.6000 ;
	    RECT 127.6000 117.6000 128.4000 118.4000 ;
	    RECT 129.2000 109.6000 130.0000 110.4000 ;
	    RECT 129.3000 106.4000 129.9000 109.6000 ;
	    RECT 129.2000 105.6000 130.0000 106.4000 ;
	    RECT 130.9000 102.4000 131.5000 131.6000 ;
	    RECT 135.7000 128.4000 136.3000 131.6000 ;
	    RECT 135.6000 127.6000 136.4000 128.4000 ;
	    RECT 134.0000 121.6000 134.8000 122.4000 ;
	    RECT 134.1000 118.4000 134.7000 121.6000 ;
	    RECT 134.0000 117.6000 134.8000 118.4000 ;
	    RECT 137.3000 116.3000 137.9000 133.7000 ;
	    RECT 140.4000 133.6000 141.2000 134.4000 ;
	    RECT 142.0000 133.6000 142.8000 134.4000 ;
	    RECT 138.8000 131.6000 139.6000 132.4000 ;
	    RECT 140.5000 122.4000 141.1000 133.6000 ;
	    RECT 140.4000 121.6000 141.2000 122.4000 ;
	    RECT 135.7000 115.7000 137.9000 116.3000 ;
	    RECT 134.0000 111.6000 134.8000 112.4000 ;
	    RECT 134.1000 110.4000 134.7000 111.6000 ;
	    RECT 132.4000 109.6000 133.2000 110.4000 ;
	    RECT 134.0000 109.6000 134.8000 110.4000 ;
	    RECT 132.5000 108.4000 133.1000 109.6000 ;
	    RECT 132.4000 107.6000 133.2000 108.4000 ;
	    RECT 134.0000 105.6000 134.8000 106.4000 ;
	    RECT 130.8000 101.6000 131.6000 102.4000 ;
	    RECT 129.2000 97.6000 130.0000 98.4000 ;
	    RECT 124.4000 93.7000 126.7000 94.3000 ;
	    RECT 124.4000 93.6000 125.2000 93.7000 ;
	    RECT 129.3000 92.4000 129.9000 97.6000 ;
	    RECT 132.4000 95.6000 133.2000 96.4000 ;
	    RECT 132.4000 93.6000 133.2000 94.4000 ;
	    RECT 129.2000 91.6000 130.0000 92.4000 ;
	    RECT 126.0000 89.6000 126.8000 90.4000 ;
	    RECT 129.2000 89.6000 130.0000 90.4000 ;
	    RECT 129.3000 78.4000 129.9000 89.6000 ;
	    RECT 129.2000 77.6000 130.0000 78.4000 ;
	    RECT 130.8000 73.6000 131.6000 74.4000 ;
	    RECT 130.9000 70.4000 131.5000 73.6000 ;
	    RECT 132.5000 70.4000 133.1000 93.6000 ;
	    RECT 134.1000 92.4000 134.7000 105.6000 ;
	    RECT 135.7000 98.4000 136.3000 115.7000 ;
	    RECT 142.1000 114.4000 142.7000 133.6000 ;
	    RECT 143.6000 131.6000 144.4000 132.4000 ;
	    RECT 143.7000 128.4000 144.3000 131.6000 ;
	    RECT 143.6000 127.6000 144.4000 128.4000 ;
	    RECT 146.9000 126.3000 147.5000 169.7000 ;
	    RECT 148.5000 152.3000 149.1000 179.7000 ;
	    RECT 151.7000 174.4000 152.3000 181.7000 ;
	    RECT 154.9000 180.3000 155.5000 185.6000 ;
	    RECT 153.3000 179.7000 155.5000 180.3000 ;
	    RECT 153.3000 178.4000 153.9000 179.7000 ;
	    RECT 153.2000 177.6000 154.0000 178.4000 ;
	    RECT 151.6000 173.6000 152.4000 174.4000 ;
	    RECT 156.5000 172.4000 157.1000 193.6000 ;
	    RECT 158.1000 190.4000 158.7000 207.6000 ;
	    RECT 158.0000 189.6000 158.8000 190.4000 ;
	    RECT 159.7000 188.4000 160.3000 209.7000 ;
	    RECT 162.8000 209.6000 163.6000 210.4000 ;
	    RECT 167.6000 210.2000 168.4000 215.8000 ;
	    RECT 169.2000 213.6000 170.0000 214.4000 ;
	    RECT 162.9000 208.4000 163.5000 209.6000 ;
	    RECT 162.8000 207.6000 163.6000 208.4000 ;
	    RECT 170.8000 206.2000 171.6000 217.8000 ;
	    RECT 162.8000 201.6000 163.6000 202.4000 ;
	    RECT 161.2000 189.6000 162.0000 190.4000 ;
	    RECT 159.6000 187.6000 160.4000 188.4000 ;
	    RECT 158.0000 177.6000 158.8000 178.4000 ;
	    RECT 159.7000 172.4000 160.3000 187.6000 ;
	    RECT 162.9000 186.3000 163.5000 201.6000 ;
	    RECT 170.8000 195.6000 171.6000 196.4000 ;
	    RECT 170.9000 192.4000 171.5000 195.6000 ;
	    RECT 172.5000 192.4000 173.1000 225.7000 ;
	    RECT 174.0000 225.6000 174.8000 225.7000 ;
	    RECT 174.0000 213.6000 174.8000 214.4000 ;
	    RECT 174.1000 212.4000 174.7000 213.6000 ;
	    RECT 174.0000 211.6000 174.8000 212.4000 ;
	    RECT 175.7000 210.3000 176.3000 227.6000 ;
	    RECT 174.1000 209.7000 176.3000 210.3000 ;
	    RECT 164.4000 191.6000 165.2000 192.4000 ;
	    RECT 170.8000 191.6000 171.6000 192.4000 ;
	    RECT 172.4000 191.6000 173.2000 192.4000 ;
	    RECT 164.5000 186.4000 165.1000 191.6000 ;
	    RECT 174.1000 190.4000 174.7000 209.7000 ;
	    RECT 175.6000 203.6000 176.4000 204.4000 ;
	    RECT 169.2000 189.6000 170.0000 190.4000 ;
	    RECT 174.0000 189.6000 174.8000 190.4000 ;
	    RECT 161.3000 185.7000 163.5000 186.3000 ;
	    RECT 150.0000 171.6000 150.8000 172.4000 ;
	    RECT 156.4000 171.6000 157.2000 172.4000 ;
	    RECT 159.6000 171.6000 160.4000 172.4000 ;
	    RECT 159.6000 163.6000 160.4000 164.4000 ;
	    RECT 153.2000 159.6000 154.0000 160.4000 ;
	    RECT 153.3000 158.4000 153.9000 159.6000 ;
	    RECT 153.2000 157.6000 154.0000 158.4000 ;
	    RECT 156.4000 157.6000 157.2000 158.4000 ;
	    RECT 150.0000 152.3000 150.8000 152.4000 ;
	    RECT 148.5000 151.7000 150.8000 152.3000 ;
	    RECT 150.0000 151.6000 150.8000 151.7000 ;
	    RECT 150.1000 150.4000 150.7000 151.6000 ;
	    RECT 156.5000 150.4000 157.1000 157.6000 ;
	    RECT 150.0000 149.6000 150.8000 150.4000 ;
	    RECT 153.2000 150.3000 154.0000 150.4000 ;
	    RECT 153.2000 149.7000 155.5000 150.3000 ;
	    RECT 153.2000 149.6000 154.0000 149.7000 ;
	    RECT 154.9000 148.3000 155.5000 149.7000 ;
	    RECT 156.4000 149.6000 157.2000 150.4000 ;
	    RECT 158.0000 149.6000 158.8000 150.4000 ;
	    RECT 158.1000 148.4000 158.7000 149.6000 ;
	    RECT 154.9000 147.7000 157.1000 148.3000 ;
	    RECT 156.5000 146.3000 157.1000 147.7000 ;
	    RECT 158.0000 147.6000 158.8000 148.4000 ;
	    RECT 159.7000 146.4000 160.3000 163.6000 ;
	    RECT 161.3000 148.3000 161.9000 185.7000 ;
	    RECT 164.4000 185.6000 165.2000 186.4000 ;
	    RECT 166.0000 185.6000 166.8000 186.4000 ;
	    RECT 162.8000 183.6000 163.6000 184.4000 ;
	    RECT 164.5000 178.4000 165.1000 185.6000 ;
	    RECT 162.8000 166.2000 163.6000 177.8000 ;
	    RECT 164.4000 177.6000 165.2000 178.4000 ;
	    RECT 164.4000 173.6000 165.2000 174.4000 ;
	    RECT 164.5000 172.4000 165.1000 173.6000 ;
	    RECT 164.4000 171.6000 165.2000 172.4000 ;
	    RECT 164.4000 165.6000 165.2000 166.4000 ;
	    RECT 164.5000 164.3000 165.1000 165.6000 ;
	    RECT 166.1000 164.4000 166.7000 185.6000 ;
	    RECT 167.6000 183.6000 168.4000 184.4000 ;
	    RECT 167.7000 176.4000 168.3000 183.6000 ;
	    RECT 169.3000 176.4000 169.9000 189.6000 ;
	    RECT 170.8000 183.6000 171.6000 184.4000 ;
	    RECT 167.6000 175.6000 168.4000 176.4000 ;
	    RECT 169.2000 175.6000 170.0000 176.4000 ;
	    RECT 170.9000 172.6000 171.5000 183.6000 ;
	    RECT 174.1000 180.4000 174.7000 189.6000 ;
	    RECT 175.7000 188.4000 176.3000 203.6000 ;
	    RECT 177.3000 194.4000 177.9000 227.6000 ;
	    RECT 178.9000 226.4000 179.5000 229.6000 ;
	    RECT 186.9000 228.4000 187.5000 251.6000 ;
	    RECT 193.3000 250.4000 193.9000 257.6000 ;
	    RECT 190.0000 249.6000 190.8000 250.4000 ;
	    RECT 193.2000 249.6000 194.0000 250.4000 ;
	    RECT 188.4000 232.3000 189.2000 232.4000 ;
	    RECT 190.1000 232.3000 190.7000 249.6000 ;
	    RECT 194.9000 248.3000 195.5000 261.6000 ;
	    RECT 199.7000 258.4000 200.3000 265.6000 ;
	    RECT 199.6000 257.6000 200.4000 258.4000 ;
	    RECT 196.4000 255.6000 197.2000 256.4000 ;
	    RECT 198.0000 255.6000 198.8000 256.4000 ;
	    RECT 196.5000 252.4000 197.1000 255.6000 ;
	    RECT 198.1000 254.4000 198.7000 255.6000 ;
	    RECT 198.0000 253.6000 198.8000 254.4000 ;
	    RECT 198.1000 252.4000 198.7000 253.6000 ;
	    RECT 196.4000 251.6000 197.2000 252.4000 ;
	    RECT 198.0000 251.6000 198.8000 252.4000 ;
	    RECT 199.6000 251.6000 200.4000 252.4000 ;
	    RECT 196.4000 249.6000 197.2000 250.4000 ;
	    RECT 199.7000 250.3000 200.3000 251.6000 ;
	    RECT 198.1000 249.7000 200.3000 250.3000 ;
	    RECT 194.9000 247.7000 197.1000 248.3000 ;
	    RECT 196.5000 238.4000 197.1000 247.7000 ;
	    RECT 196.4000 237.6000 197.2000 238.4000 ;
	    RECT 193.2000 235.6000 194.0000 236.4000 ;
	    RECT 194.8000 235.6000 195.6000 236.4000 ;
	    RECT 194.9000 232.4000 195.5000 235.6000 ;
	    RECT 188.4000 231.7000 190.7000 232.3000 ;
	    RECT 188.4000 231.6000 189.2000 231.7000 ;
	    RECT 183.6000 227.6000 184.4000 228.4000 ;
	    RECT 186.8000 227.6000 187.6000 228.4000 ;
	    RECT 178.8000 225.6000 179.6000 226.4000 ;
	    RECT 178.8000 219.6000 179.6000 220.4000 ;
	    RECT 177.2000 193.6000 178.0000 194.4000 ;
	    RECT 177.2000 191.6000 178.0000 192.4000 ;
	    RECT 177.2000 189.6000 178.0000 190.4000 ;
	    RECT 175.6000 187.6000 176.4000 188.4000 ;
	    RECT 174.0000 179.6000 174.8000 180.4000 ;
	    RECT 177.3000 178.4000 177.9000 189.6000 ;
	    RECT 178.9000 182.3000 179.5000 219.6000 ;
	    RECT 180.4000 206.2000 181.2000 217.8000 ;
	    RECT 182.0000 209.6000 182.8000 210.4000 ;
	    RECT 180.4000 195.6000 181.2000 196.4000 ;
	    RECT 180.4000 189.6000 181.2000 190.4000 ;
	    RECT 180.5000 186.4000 181.1000 189.6000 ;
	    RECT 182.1000 188.4000 182.7000 209.6000 ;
	    RECT 183.7000 208.4000 184.3000 227.6000 ;
	    RECT 190.1000 226.4000 190.7000 231.7000 ;
	    RECT 194.8000 231.6000 195.6000 232.4000 ;
	    RECT 194.8000 230.3000 195.6000 230.4000 ;
	    RECT 194.8000 229.7000 197.1000 230.3000 ;
	    RECT 194.8000 229.6000 195.6000 229.7000 ;
	    RECT 194.8000 228.3000 195.6000 228.4000 ;
	    RECT 193.3000 227.7000 195.6000 228.3000 ;
	    RECT 190.0000 225.6000 190.8000 226.4000 ;
	    RECT 185.2000 219.6000 186.0000 220.4000 ;
	    RECT 186.8000 219.6000 187.6000 220.4000 ;
	    RECT 188.4000 219.6000 189.2000 220.4000 ;
	    RECT 185.3000 216.4000 185.9000 219.6000 ;
	    RECT 186.9000 218.4000 187.5000 219.6000 ;
	    RECT 186.8000 217.6000 187.6000 218.4000 ;
	    RECT 185.2000 215.6000 186.0000 216.4000 ;
	    RECT 183.6000 207.6000 184.4000 208.4000 ;
	    RECT 185.2000 203.6000 186.0000 204.4000 ;
	    RECT 185.3000 192.4000 185.9000 203.6000 ;
	    RECT 188.5000 202.4000 189.1000 219.6000 ;
	    RECT 190.0000 215.6000 190.8000 216.4000 ;
	    RECT 190.1000 212.4000 190.7000 215.6000 ;
	    RECT 190.0000 211.6000 190.8000 212.4000 ;
	    RECT 193.3000 204.4000 193.9000 227.7000 ;
	    RECT 194.8000 227.6000 195.6000 227.7000 ;
	    RECT 196.5000 226.4000 197.1000 229.7000 ;
	    RECT 198.1000 226.4000 198.7000 249.7000 ;
	    RECT 201.3000 244.4000 201.9000 269.7000 ;
	    RECT 202.8000 269.6000 203.6000 269.7000 ;
	    RECT 207.6000 269.6000 208.4000 270.4000 ;
	    RECT 210.9000 270.3000 211.5000 271.7000 ;
	    RECT 214.1000 270.4000 214.7000 271.7000 ;
	    RECT 215.7000 270.4000 216.3000 293.6000 ;
	    RECT 217.3000 290.4000 217.9000 297.6000 ;
	    RECT 217.2000 289.6000 218.0000 290.4000 ;
	    RECT 217.3000 286.4000 217.9000 289.6000 ;
	    RECT 217.2000 285.6000 218.0000 286.4000 ;
	    RECT 218.9000 284.3000 219.5000 323.6000 ;
	    RECT 226.9000 318.4000 227.5000 333.6000 ;
	    RECT 234.8000 331.6000 235.6000 332.4000 ;
	    RECT 241.2000 331.6000 242.0000 332.4000 ;
	    RECT 234.9000 330.4000 235.5000 331.6000 ;
	    RECT 234.8000 329.6000 235.6000 330.4000 ;
	    RECT 242.8000 329.6000 243.6000 330.4000 ;
	    RECT 233.2000 327.6000 234.0000 328.4000 ;
	    RECT 228.4000 323.6000 229.2000 324.4000 ;
	    RECT 220.4000 317.6000 221.2000 318.4000 ;
	    RECT 226.8000 317.6000 227.6000 318.4000 ;
	    RECT 223.6000 313.6000 224.4000 314.4000 ;
	    RECT 226.8000 312.3000 227.6000 312.4000 ;
	    RECT 228.5000 312.3000 229.1000 323.6000 ;
	    RECT 233.3000 314.4000 233.9000 327.6000 ;
	    RECT 233.2000 313.6000 234.0000 314.4000 ;
	    RECT 226.8000 311.7000 229.1000 312.3000 ;
	    RECT 226.8000 311.6000 227.6000 311.7000 ;
	    RECT 223.6000 309.6000 224.4000 310.4000 ;
	    RECT 222.0000 307.6000 222.8000 308.4000 ;
	    RECT 225.2000 307.6000 226.0000 308.4000 ;
	    RECT 222.1000 306.4000 222.7000 307.6000 ;
	    RECT 222.0000 305.6000 222.8000 306.4000 ;
	    RECT 225.3000 304.4000 225.9000 307.6000 ;
	    RECT 233.3000 306.4000 233.9000 313.6000 ;
	    RECT 234.9000 312.4000 235.5000 329.6000 ;
	    RECT 241.2000 321.6000 242.0000 322.4000 ;
	    RECT 236.4000 314.3000 237.2000 314.4000 ;
	    RECT 236.4000 313.7000 238.7000 314.3000 ;
	    RECT 236.4000 313.6000 237.2000 313.7000 ;
	    RECT 234.8000 311.6000 235.6000 312.4000 ;
	    RECT 236.4000 311.6000 237.2000 312.4000 ;
	    RECT 233.2000 305.6000 234.0000 306.4000 ;
	    RECT 225.2000 303.6000 226.0000 304.4000 ;
	    RECT 231.6000 303.6000 232.4000 304.4000 ;
	    RECT 225.2000 297.6000 226.0000 298.4000 ;
	    RECT 228.4000 297.6000 229.2000 298.4000 ;
	    RECT 223.6000 293.6000 224.4000 294.4000 ;
	    RECT 225.2000 293.6000 226.0000 294.4000 ;
	    RECT 220.4000 291.6000 221.2000 292.4000 ;
	    RECT 222.0000 291.6000 222.8000 292.4000 ;
	    RECT 220.5000 290.3000 221.1000 291.6000 ;
	    RECT 225.3000 290.3000 225.9000 293.6000 ;
	    RECT 220.5000 289.7000 225.9000 290.3000 ;
	    RECT 220.4000 285.6000 221.2000 286.4000 ;
	    RECT 217.3000 283.7000 219.5000 284.3000 ;
	    RECT 209.3000 269.7000 211.5000 270.3000 ;
	    RECT 204.4000 268.3000 205.2000 268.4000 ;
	    RECT 209.3000 268.3000 209.9000 269.7000 ;
	    RECT 212.4000 269.6000 213.2000 270.4000 ;
	    RECT 214.0000 269.6000 214.8000 270.4000 ;
	    RECT 215.6000 269.6000 216.4000 270.4000 ;
	    RECT 204.4000 267.7000 209.9000 268.3000 ;
	    RECT 204.4000 267.6000 205.2000 267.7000 ;
	    RECT 210.8000 267.6000 211.6000 268.4000 ;
	    RECT 214.0000 268.3000 214.8000 268.4000 ;
	    RECT 212.5000 267.7000 214.8000 268.3000 ;
	    RECT 210.9000 266.4000 211.5000 267.6000 ;
	    RECT 202.8000 265.6000 203.6000 266.4000 ;
	    RECT 204.4000 265.6000 205.2000 266.4000 ;
	    RECT 210.8000 265.6000 211.6000 266.4000 ;
	    RECT 202.9000 258.4000 203.5000 265.6000 ;
	    RECT 204.5000 264.4000 205.1000 265.6000 ;
	    RECT 204.4000 263.6000 205.2000 264.4000 ;
	    RECT 209.2000 261.6000 210.0000 262.4000 ;
	    RECT 204.4000 259.6000 205.2000 260.4000 ;
	    RECT 202.8000 257.6000 203.6000 258.4000 ;
	    RECT 201.2000 243.6000 202.0000 244.4000 ;
	    RECT 201.3000 230.4000 201.9000 243.6000 ;
	    RECT 199.6000 229.6000 200.4000 230.4000 ;
	    RECT 201.2000 229.6000 202.0000 230.4000 ;
	    RECT 202.8000 229.6000 203.6000 230.4000 ;
	    RECT 196.4000 225.6000 197.2000 226.4000 ;
	    RECT 198.0000 225.6000 198.8000 226.4000 ;
	    RECT 199.7000 216.3000 200.3000 229.6000 ;
	    RECT 201.2000 227.6000 202.0000 228.4000 ;
	    RECT 198.1000 215.7000 200.3000 216.3000 ;
	    RECT 196.4000 213.6000 197.2000 214.4000 ;
	    RECT 193.2000 203.6000 194.0000 204.4000 ;
	    RECT 194.8000 203.6000 195.6000 204.4000 ;
	    RECT 188.4000 201.6000 189.2000 202.4000 ;
	    RECT 194.9000 200.4000 195.5000 203.6000 ;
	    RECT 191.6000 199.6000 192.4000 200.4000 ;
	    RECT 194.8000 199.6000 195.6000 200.4000 ;
	    RECT 191.7000 198.4000 192.3000 199.6000 ;
	    RECT 191.6000 197.6000 192.4000 198.4000 ;
	    RECT 191.6000 195.6000 192.4000 196.4000 ;
	    RECT 183.6000 191.6000 184.4000 192.4000 ;
	    RECT 185.2000 191.6000 186.0000 192.4000 ;
	    RECT 188.4000 191.6000 189.2000 192.4000 ;
	    RECT 183.7000 188.4000 184.3000 191.6000 ;
	    RECT 188.5000 190.4000 189.1000 191.6000 ;
	    RECT 191.7000 190.4000 192.3000 195.6000 ;
	    RECT 196.5000 192.4000 197.1000 213.6000 ;
	    RECT 198.1000 198.3000 198.7000 215.7000 ;
	    RECT 199.6000 213.6000 200.4000 214.4000 ;
	    RECT 199.6000 209.6000 200.4000 210.4000 ;
	    RECT 199.7000 200.4000 200.3000 209.6000 ;
	    RECT 199.6000 199.6000 200.4000 200.4000 ;
	    RECT 198.1000 197.7000 200.3000 198.3000 ;
	    RECT 199.7000 196.4000 200.3000 197.7000 ;
	    RECT 198.0000 195.6000 198.8000 196.4000 ;
	    RECT 199.6000 195.6000 200.4000 196.4000 ;
	    RECT 201.3000 194.3000 201.9000 227.6000 ;
	    RECT 204.5000 226.4000 205.1000 259.6000 ;
	    RECT 207.6000 257.6000 208.4000 258.4000 ;
	    RECT 206.0000 251.6000 206.8000 252.4000 ;
	    RECT 206.1000 250.4000 206.7000 251.6000 ;
	    RECT 206.0000 249.6000 206.8000 250.4000 ;
	    RECT 207.7000 248.3000 208.3000 257.6000 ;
	    RECT 206.1000 247.7000 208.3000 248.3000 ;
	    RECT 206.1000 242.4000 206.7000 247.7000 ;
	    RECT 207.6000 243.6000 208.4000 244.4000 ;
	    RECT 206.0000 241.6000 206.8000 242.4000 ;
	    RECT 207.7000 230.4000 208.3000 243.6000 ;
	    RECT 207.6000 229.6000 208.4000 230.4000 ;
	    RECT 206.0000 227.6000 206.8000 228.4000 ;
	    RECT 202.8000 225.6000 203.6000 226.4000 ;
	    RECT 204.4000 225.6000 205.2000 226.4000 ;
	    RECT 202.9000 196.4000 203.5000 225.6000 ;
	    RECT 207.6000 223.6000 208.4000 224.4000 ;
	    RECT 207.7000 218.4000 208.3000 223.6000 ;
	    RECT 209.3000 222.3000 209.9000 261.6000 ;
	    RECT 210.8000 257.6000 211.6000 258.4000 ;
	    RECT 210.9000 252.4000 211.5000 257.6000 ;
	    RECT 212.5000 252.4000 213.1000 267.7000 ;
	    RECT 214.0000 267.6000 214.8000 267.7000 ;
	    RECT 215.6000 267.6000 216.4000 268.4000 ;
	    RECT 214.0000 266.3000 214.8000 266.4000 ;
	    RECT 215.7000 266.3000 216.3000 267.6000 ;
	    RECT 214.0000 265.7000 216.3000 266.3000 ;
	    RECT 214.0000 265.6000 214.8000 265.7000 ;
	    RECT 217.3000 258.4000 217.9000 283.7000 ;
	    RECT 220.5000 274.4000 221.1000 285.6000 ;
	    RECT 228.5000 284.3000 229.1000 297.6000 ;
	    RECT 230.0000 286.2000 230.8000 297.8000 ;
	    RECT 231.7000 292.4000 232.3000 303.6000 ;
	    RECT 234.9000 294.4000 235.5000 311.6000 ;
	    RECT 236.5000 310.4000 237.1000 311.6000 ;
	    RECT 238.1000 310.4000 238.7000 313.7000 ;
	    RECT 236.4000 309.6000 237.2000 310.4000 ;
	    RECT 238.0000 309.6000 238.8000 310.4000 ;
	    RECT 238.0000 307.6000 238.8000 308.4000 ;
	    RECT 238.1000 294.4000 238.7000 307.6000 ;
	    RECT 233.2000 293.6000 234.0000 294.4000 ;
	    RECT 234.8000 293.6000 235.6000 294.4000 ;
	    RECT 238.0000 293.6000 238.8000 294.4000 ;
	    RECT 233.3000 292.4000 233.9000 293.6000 ;
	    RECT 231.6000 291.6000 232.4000 292.4000 ;
	    RECT 233.2000 291.6000 234.0000 292.4000 ;
	    RECT 234.9000 290.4000 235.5000 293.6000 ;
	    RECT 234.8000 289.6000 235.6000 290.4000 ;
	    RECT 239.6000 286.2000 240.4000 297.8000 ;
	    RECT 241.3000 288.3000 241.9000 321.6000 ;
	    RECT 242.9000 310.4000 243.5000 329.6000 ;
	    RECT 247.6000 326.2000 248.4000 337.8000 ;
	    RECT 255.6000 333.6000 256.4000 334.4000 ;
	    RECT 255.7000 332.6000 256.3000 333.6000 ;
	    RECT 249.2000 331.6000 250.0000 332.4000 ;
	    RECT 255.6000 331.8000 256.4000 332.6000 ;
	    RECT 257.2000 326.2000 258.0000 337.8000 ;
	    RECT 263.6000 337.6000 264.4000 338.4000 ;
	    RECT 292.4000 337.6000 293.2000 338.4000 ;
	    RECT 260.4000 330.2000 261.2000 335.8000 ;
	    RECT 262.0000 335.6000 262.8000 336.4000 ;
	    RECT 262.1000 328.4000 262.7000 335.6000 ;
	    RECT 262.0000 327.6000 262.8000 328.4000 ;
	    RECT 244.4000 323.6000 245.2000 324.4000 ;
	    RECT 242.8000 309.6000 243.6000 310.4000 ;
	    RECT 244.5000 308.4000 245.1000 323.6000 ;
	    RECT 252.4000 319.6000 253.2000 320.4000 ;
	    RECT 247.6000 309.6000 248.4000 310.4000 ;
	    RECT 247.7000 308.4000 248.3000 309.6000 ;
	    RECT 252.5000 308.4000 253.1000 319.6000 ;
	    RECT 260.4000 311.6000 261.2000 312.4000 ;
	    RECT 260.5000 310.4000 261.1000 311.6000 ;
	    RECT 260.4000 310.3000 261.2000 310.4000 ;
	    RECT 260.4000 309.7000 262.7000 310.3000 ;
	    RECT 260.4000 309.6000 261.2000 309.7000 ;
	    RECT 244.4000 307.6000 245.2000 308.4000 ;
	    RECT 246.0000 307.6000 246.8000 308.4000 ;
	    RECT 247.6000 307.6000 248.4000 308.4000 ;
	    RECT 252.4000 307.6000 253.2000 308.4000 ;
	    RECT 242.8000 303.6000 243.6000 304.4000 ;
	    RECT 242.9000 302.4000 243.5000 303.6000 ;
	    RECT 242.8000 301.6000 243.6000 302.4000 ;
	    RECT 244.4000 301.6000 245.2000 302.4000 ;
	    RECT 242.8000 290.2000 243.6000 295.8000 ;
	    RECT 244.5000 294.4000 245.1000 301.6000 ;
	    RECT 246.1000 294.4000 246.7000 307.6000 ;
	    RECT 247.6000 303.6000 248.4000 304.4000 ;
	    RECT 249.2000 303.6000 250.0000 304.4000 ;
	    RECT 247.7000 300.4000 248.3000 303.6000 ;
	    RECT 247.6000 299.6000 248.4000 300.4000 ;
	    RECT 244.4000 293.6000 245.2000 294.4000 ;
	    RECT 246.0000 293.6000 246.8000 294.4000 ;
	    RECT 244.4000 291.6000 245.2000 292.4000 ;
	    RECT 246.0000 291.6000 246.8000 292.4000 ;
	    RECT 246.1000 290.3000 246.7000 291.6000 ;
	    RECT 244.5000 289.7000 246.7000 290.3000 ;
	    RECT 249.3000 290.3000 249.9000 303.6000 ;
	    RECT 252.4000 301.6000 253.2000 302.4000 ;
	    RECT 250.8000 297.6000 251.6000 298.4000 ;
	    RECT 250.9000 292.4000 251.5000 297.6000 ;
	    RECT 252.5000 294.4000 253.1000 301.6000 ;
	    RECT 252.4000 293.6000 253.2000 294.4000 ;
	    RECT 260.4000 293.6000 261.2000 294.4000 ;
	    RECT 250.8000 291.6000 251.6000 292.4000 ;
	    RECT 260.5000 290.4000 261.1000 293.6000 ;
	    RECT 249.3000 289.7000 251.5000 290.3000 ;
	    RECT 244.5000 288.3000 245.1000 289.7000 ;
	    RECT 241.3000 287.7000 245.1000 288.3000 ;
	    RECT 228.5000 283.7000 230.7000 284.3000 ;
	    RECT 225.2000 279.6000 226.0000 280.4000 ;
	    RECT 222.0000 275.6000 222.8000 276.4000 ;
	    RECT 225.3000 276.3000 225.9000 279.6000 ;
	    RECT 226.8000 277.6000 227.6000 278.4000 ;
	    RECT 225.3000 275.7000 227.5000 276.3000 ;
	    RECT 220.4000 273.6000 221.2000 274.4000 ;
	    RECT 220.4000 269.6000 221.2000 270.4000 ;
	    RECT 218.8000 267.6000 219.6000 268.4000 ;
	    RECT 218.9000 262.4000 219.5000 267.6000 ;
	    RECT 218.8000 261.6000 219.6000 262.4000 ;
	    RECT 220.5000 258.4000 221.1000 269.6000 ;
	    RECT 222.1000 268.4000 222.7000 275.6000 ;
	    RECT 223.6000 271.6000 224.4000 272.4000 ;
	    RECT 223.7000 270.4000 224.3000 271.6000 ;
	    RECT 223.6000 269.6000 224.4000 270.4000 ;
	    RECT 225.2000 269.6000 226.0000 270.4000 ;
	    RECT 222.0000 267.6000 222.8000 268.4000 ;
	    RECT 215.6000 257.6000 216.4000 258.4000 ;
	    RECT 217.2000 257.6000 218.0000 258.4000 ;
	    RECT 220.4000 257.6000 221.2000 258.4000 ;
	    RECT 215.7000 256.3000 216.3000 257.6000 ;
	    RECT 218.8000 256.3000 219.6000 256.4000 ;
	    RECT 215.7000 255.7000 219.6000 256.3000 ;
	    RECT 214.0000 253.6000 214.8000 254.4000 ;
	    RECT 214.1000 252.4000 214.7000 253.6000 ;
	    RECT 215.7000 252.4000 216.3000 255.7000 ;
	    RECT 218.8000 255.6000 219.6000 255.7000 ;
	    RECT 223.6000 253.6000 224.4000 254.4000 ;
	    RECT 210.8000 251.6000 211.6000 252.4000 ;
	    RECT 212.4000 251.6000 213.2000 252.4000 ;
	    RECT 214.0000 251.6000 214.8000 252.4000 ;
	    RECT 215.6000 251.6000 216.4000 252.4000 ;
	    RECT 220.4000 251.6000 221.2000 252.4000 ;
	    RECT 212.5000 250.3000 213.1000 251.6000 ;
	    RECT 220.5000 250.4000 221.1000 251.6000 ;
	    RECT 212.5000 249.7000 214.7000 250.3000 ;
	    RECT 214.1000 238.3000 214.7000 249.7000 ;
	    RECT 220.4000 249.6000 221.2000 250.4000 ;
	    RECT 223.7000 244.4000 224.3000 253.6000 ;
	    RECT 225.2000 251.6000 226.0000 252.4000 ;
	    RECT 226.9000 250.4000 227.5000 275.7000 ;
	    RECT 228.4000 273.6000 229.2000 274.4000 ;
	    RECT 228.5000 252.4000 229.1000 273.6000 ;
	    RECT 230.1000 270.4000 230.7000 283.7000 ;
	    RECT 247.6000 283.6000 248.4000 284.4000 ;
	    RECT 231.6000 279.6000 232.4000 280.4000 ;
	    RECT 246.0000 279.6000 246.8000 280.4000 ;
	    RECT 230.0000 269.6000 230.8000 270.4000 ;
	    RECT 231.7000 258.4000 232.3000 279.6000 ;
	    RECT 246.1000 278.4000 246.7000 279.6000 ;
	    RECT 239.6000 277.6000 240.4000 278.4000 ;
	    RECT 246.0000 277.6000 246.8000 278.4000 ;
	    RECT 233.2000 271.6000 234.0000 272.4000 ;
	    RECT 238.0000 271.6000 238.8000 272.4000 ;
	    RECT 233.3000 270.4000 233.9000 271.6000 ;
	    RECT 239.7000 270.4000 240.3000 277.6000 ;
	    RECT 242.8000 275.6000 243.6000 276.4000 ;
	    RECT 233.2000 269.6000 234.0000 270.4000 ;
	    RECT 234.8000 270.3000 235.6000 270.4000 ;
	    RECT 234.8000 269.7000 237.1000 270.3000 ;
	    RECT 234.8000 269.6000 235.6000 269.7000 ;
	    RECT 231.6000 257.6000 232.4000 258.4000 ;
	    RECT 233.3000 254.4000 233.9000 269.6000 ;
	    RECT 236.5000 266.4000 237.1000 269.7000 ;
	    RECT 239.6000 269.6000 240.4000 270.4000 ;
	    RECT 241.2000 269.6000 242.0000 270.4000 ;
	    RECT 241.3000 268.3000 241.9000 269.6000 ;
	    RECT 238.1000 267.7000 241.9000 268.3000 ;
	    RECT 236.4000 265.6000 237.2000 266.4000 ;
	    RECT 236.4000 263.6000 237.2000 264.4000 ;
	    RECT 233.2000 253.6000 234.0000 254.4000 ;
	    RECT 234.8000 253.6000 235.6000 254.4000 ;
	    RECT 228.4000 251.6000 229.2000 252.4000 ;
	    RECT 230.0000 251.6000 230.8000 252.4000 ;
	    RECT 226.8000 249.6000 227.6000 250.4000 ;
	    RECT 225.2000 247.6000 226.0000 248.4000 ;
	    RECT 226.8000 247.6000 227.6000 248.4000 ;
	    RECT 218.8000 243.6000 219.6000 244.4000 ;
	    RECT 222.0000 243.6000 222.8000 244.4000 ;
	    RECT 223.6000 243.6000 224.4000 244.4000 ;
	    RECT 214.1000 237.7000 216.3000 238.3000 ;
	    RECT 214.0000 231.6000 214.8000 232.4000 ;
	    RECT 210.8000 229.6000 211.6000 230.4000 ;
	    RECT 214.1000 228.4000 214.7000 231.6000 ;
	    RECT 215.7000 230.4000 216.3000 237.7000 ;
	    RECT 217.2000 235.6000 218.0000 236.4000 ;
	    RECT 217.3000 230.4000 217.9000 235.6000 ;
	    RECT 222.1000 230.4000 222.7000 243.6000 ;
	    RECT 223.7000 230.4000 224.3000 243.6000 ;
	    RECT 215.6000 229.6000 216.4000 230.4000 ;
	    RECT 217.2000 229.6000 218.0000 230.4000 ;
	    RECT 218.8000 229.6000 219.6000 230.4000 ;
	    RECT 220.4000 229.6000 221.2000 230.4000 ;
	    RECT 222.0000 229.6000 222.8000 230.4000 ;
	    RECT 223.6000 229.6000 224.4000 230.4000 ;
	    RECT 225.2000 229.6000 226.0000 230.4000 ;
	    RECT 214.0000 227.6000 214.8000 228.4000 ;
	    RECT 209.3000 221.7000 211.5000 222.3000 ;
	    RECT 209.2000 219.6000 210.0000 220.4000 ;
	    RECT 209.3000 218.4000 209.9000 219.6000 ;
	    RECT 207.6000 217.6000 208.4000 218.4000 ;
	    RECT 209.2000 217.6000 210.0000 218.4000 ;
	    RECT 207.6000 215.6000 208.4000 216.4000 ;
	    RECT 206.0000 213.6000 206.8000 214.4000 ;
	    RECT 210.9000 212.4000 211.5000 221.7000 ;
	    RECT 212.4000 219.6000 213.2000 220.4000 ;
	    RECT 212.5000 214.4000 213.1000 219.6000 ;
	    RECT 212.4000 213.6000 213.2000 214.4000 ;
	    RECT 204.4000 211.6000 205.2000 212.4000 ;
	    RECT 210.8000 211.6000 211.6000 212.4000 ;
	    RECT 204.5000 200.4000 205.1000 211.6000 ;
	    RECT 204.4000 199.6000 205.2000 200.4000 ;
	    RECT 214.1000 198.4000 214.7000 227.6000 ;
	    RECT 215.6000 221.6000 216.4000 222.4000 ;
	    RECT 215.7000 210.4000 216.3000 221.6000 ;
	    RECT 217.3000 220.4000 217.9000 229.6000 ;
	    RECT 220.5000 228.4000 221.1000 229.6000 ;
	    RECT 220.4000 228.3000 221.2000 228.4000 ;
	    RECT 218.9000 227.7000 221.2000 228.3000 ;
	    RECT 217.2000 219.6000 218.0000 220.4000 ;
	    RECT 218.9000 218.3000 219.5000 227.7000 ;
	    RECT 220.4000 227.6000 221.2000 227.7000 ;
	    RECT 222.0000 223.6000 222.8000 224.4000 ;
	    RECT 220.4000 221.6000 221.2000 222.4000 ;
	    RECT 217.3000 217.7000 219.5000 218.3000 ;
	    RECT 215.6000 209.6000 216.4000 210.4000 ;
	    RECT 217.3000 200.4000 217.9000 217.7000 ;
	    RECT 220.5000 212.4000 221.1000 221.6000 ;
	    RECT 222.1000 220.4000 222.7000 223.6000 ;
	    RECT 222.0000 219.6000 222.8000 220.4000 ;
	    RECT 222.0000 213.6000 222.8000 214.4000 ;
	    RECT 218.8000 211.6000 219.6000 212.4000 ;
	    RECT 220.4000 211.6000 221.2000 212.4000 ;
	    RECT 223.6000 210.2000 224.4000 215.8000 ;
	    RECT 225.3000 214.4000 225.9000 229.6000 ;
	    RECT 226.9000 228.4000 227.5000 247.6000 ;
	    RECT 228.4000 231.6000 229.2000 232.4000 ;
	    RECT 228.5000 230.4000 229.1000 231.6000 ;
	    RECT 228.4000 229.6000 229.2000 230.4000 ;
	    RECT 230.1000 228.4000 230.7000 251.6000 ;
	    RECT 231.6000 247.6000 232.4000 248.4000 ;
	    RECT 231.7000 244.4000 232.3000 247.6000 ;
	    RECT 231.6000 243.6000 232.4000 244.4000 ;
	    RECT 231.6000 241.6000 232.4000 242.4000 ;
	    RECT 226.8000 227.6000 227.6000 228.4000 ;
	    RECT 230.0000 227.6000 230.8000 228.4000 ;
	    RECT 230.0000 225.6000 230.8000 226.4000 ;
	    RECT 225.2000 213.6000 226.0000 214.4000 ;
	    RECT 220.4000 205.6000 221.2000 206.4000 ;
	    RECT 226.8000 206.2000 227.6000 217.8000 ;
	    RECT 228.4000 215.6000 229.2000 216.4000 ;
	    RECT 228.4000 211.6000 229.2000 212.6000 ;
	    RECT 230.1000 206.4000 230.7000 225.6000 ;
	    RECT 231.7000 224.4000 232.3000 241.6000 ;
	    RECT 233.3000 230.4000 233.9000 253.6000 ;
	    RECT 234.9000 252.4000 235.5000 253.6000 ;
	    RECT 234.8000 251.6000 235.6000 252.4000 ;
	    RECT 234.8000 235.6000 235.6000 236.4000 ;
	    RECT 233.2000 229.6000 234.0000 230.4000 ;
	    RECT 233.2000 228.3000 234.0000 228.4000 ;
	    RECT 234.9000 228.3000 235.5000 235.6000 ;
	    RECT 236.5000 230.4000 237.1000 263.6000 ;
	    RECT 238.1000 256.4000 238.7000 267.7000 ;
	    RECT 239.6000 259.6000 240.4000 260.4000 ;
	    RECT 238.0000 255.6000 238.8000 256.4000 ;
	    RECT 238.1000 254.4000 238.7000 255.6000 ;
	    RECT 238.0000 253.6000 238.8000 254.4000 ;
	    RECT 238.1000 248.4000 238.7000 253.6000 ;
	    RECT 239.7000 252.4000 240.3000 259.6000 ;
	    RECT 242.9000 254.3000 243.5000 275.6000 ;
	    RECT 244.4000 269.6000 245.2000 270.4000 ;
	    RECT 244.5000 266.4000 245.1000 269.6000 ;
	    RECT 244.4000 265.6000 245.2000 266.4000 ;
	    RECT 247.7000 256.3000 248.3000 283.6000 ;
	    RECT 249.2000 279.6000 250.0000 280.4000 ;
	    RECT 249.3000 278.4000 249.9000 279.6000 ;
	    RECT 249.2000 277.6000 250.0000 278.4000 ;
	    RECT 249.3000 270.4000 249.9000 277.6000 ;
	    RECT 250.9000 274.4000 251.5000 289.7000 ;
	    RECT 260.4000 289.6000 261.2000 290.4000 ;
	    RECT 257.2000 285.6000 258.0000 286.4000 ;
	    RECT 257.3000 278.4000 257.9000 285.6000 ;
	    RECT 257.2000 277.6000 258.0000 278.4000 ;
	    RECT 250.8000 273.6000 251.6000 274.4000 ;
	    RECT 250.8000 271.6000 251.6000 272.4000 ;
	    RECT 249.2000 269.6000 250.0000 270.4000 ;
	    RECT 250.9000 260.4000 251.5000 271.6000 ;
	    RECT 262.1000 264.4000 262.7000 309.7000 ;
	    RECT 263.7000 306.4000 264.3000 337.6000 ;
	    RECT 279.6000 335.6000 280.4000 336.4000 ;
	    RECT 284.4000 335.6000 285.2000 336.4000 ;
	    RECT 279.7000 334.4000 280.3000 335.6000 ;
	    RECT 274.8000 333.6000 275.6000 334.4000 ;
	    RECT 278.0000 333.6000 278.8000 334.4000 ;
	    RECT 279.6000 333.6000 280.4000 334.4000 ;
	    RECT 278.1000 332.4000 278.7000 333.6000 ;
	    RECT 284.5000 332.4000 285.1000 335.6000 ;
	    RECT 289.2000 333.6000 290.0000 334.4000 ;
	    RECT 289.3000 332.4000 289.9000 333.6000 ;
	    RECT 273.2000 331.6000 274.0000 332.4000 ;
	    RECT 278.0000 331.6000 278.8000 332.4000 ;
	    RECT 279.6000 331.6000 280.4000 332.4000 ;
	    RECT 284.4000 331.6000 285.2000 332.4000 ;
	    RECT 286.0000 331.6000 286.8000 332.4000 ;
	    RECT 289.2000 331.6000 290.0000 332.4000 ;
	    RECT 276.4000 329.6000 277.2000 330.4000 ;
	    RECT 274.8000 327.6000 275.6000 328.4000 ;
	    RECT 268.4000 319.6000 269.2000 320.4000 ;
	    RECT 268.5000 318.4000 269.1000 319.6000 ;
	    RECT 268.4000 317.6000 269.2000 318.4000 ;
	    RECT 266.8000 313.6000 267.6000 314.4000 ;
	    RECT 268.4000 313.6000 269.2000 314.4000 ;
	    RECT 265.2000 311.6000 266.0000 312.4000 ;
	    RECT 263.6000 305.6000 264.4000 306.4000 ;
	    RECT 263.6000 303.6000 264.4000 304.4000 ;
	    RECT 263.7000 296.4000 264.3000 303.6000 ;
	    RECT 263.6000 295.6000 264.4000 296.4000 ;
	    RECT 265.3000 294.4000 265.9000 311.6000 ;
	    RECT 266.9000 296.4000 267.5000 313.6000 ;
	    RECT 268.5000 310.4000 269.1000 313.6000 ;
	    RECT 268.4000 309.6000 269.2000 310.4000 ;
	    RECT 271.6000 309.6000 272.4000 310.4000 ;
	    RECT 268.5000 304.4000 269.1000 309.6000 ;
	    RECT 270.0000 307.6000 270.8000 308.4000 ;
	    RECT 268.4000 303.6000 269.2000 304.4000 ;
	    RECT 266.8000 295.6000 267.6000 296.4000 ;
	    RECT 265.2000 293.6000 266.0000 294.4000 ;
	    RECT 266.8000 293.6000 267.6000 294.4000 ;
	    RECT 263.6000 291.6000 264.4000 292.4000 ;
	    RECT 263.7000 286.4000 264.3000 291.6000 ;
	    RECT 266.9000 290.4000 267.5000 293.6000 ;
	    RECT 266.8000 290.3000 267.6000 290.4000 ;
	    RECT 265.3000 289.7000 267.6000 290.3000 ;
	    RECT 263.6000 285.6000 264.4000 286.4000 ;
	    RECT 263.6000 278.3000 264.4000 278.4000 ;
	    RECT 265.3000 278.3000 265.9000 289.7000 ;
	    RECT 266.8000 289.6000 267.6000 289.7000 ;
	    RECT 268.5000 286.4000 269.1000 303.6000 ;
	    RECT 270.1000 300.4000 270.7000 307.6000 ;
	    RECT 271.7000 302.4000 272.3000 309.6000 ;
	    RECT 273.2000 307.6000 274.0000 308.4000 ;
	    RECT 271.6000 301.6000 272.4000 302.4000 ;
	    RECT 270.0000 299.6000 270.8000 300.4000 ;
	    RECT 270.0000 295.6000 270.8000 296.4000 ;
	    RECT 271.6000 295.6000 272.4000 296.4000 ;
	    RECT 270.1000 292.4000 270.7000 295.6000 ;
	    RECT 271.7000 294.4000 272.3000 295.6000 ;
	    RECT 271.6000 293.6000 272.4000 294.4000 ;
	    RECT 270.0000 291.6000 270.8000 292.4000 ;
	    RECT 271.6000 291.6000 272.4000 292.4000 ;
	    RECT 271.7000 290.3000 272.3000 291.6000 ;
	    RECT 270.1000 289.7000 272.3000 290.3000 ;
	    RECT 270.1000 288.4000 270.7000 289.7000 ;
	    RECT 270.0000 287.6000 270.8000 288.4000 ;
	    RECT 268.4000 285.6000 269.2000 286.4000 ;
	    RECT 273.2000 283.6000 274.0000 284.4000 ;
	    RECT 263.6000 277.7000 265.9000 278.3000 ;
	    RECT 263.6000 277.6000 264.4000 277.7000 ;
	    RECT 265.2000 275.6000 266.0000 276.4000 ;
	    RECT 262.0000 263.6000 262.8000 264.4000 ;
	    RECT 250.8000 259.6000 251.6000 260.4000 ;
	    RECT 246.1000 255.7000 248.3000 256.3000 ;
	    RECT 244.4000 254.3000 245.2000 254.4000 ;
	    RECT 242.9000 253.7000 245.2000 254.3000 ;
	    RECT 244.4000 253.6000 245.2000 253.7000 ;
	    RECT 246.1000 252.4000 246.7000 255.7000 ;
	    RECT 258.8000 255.6000 259.6000 256.4000 ;
	    RECT 260.4000 255.6000 261.2000 256.4000 ;
	    RECT 250.8000 254.3000 251.6000 254.4000 ;
	    RECT 247.7000 253.7000 251.6000 254.3000 ;
	    RECT 239.6000 251.6000 240.4000 252.4000 ;
	    RECT 246.0000 251.6000 246.8000 252.4000 ;
	    RECT 247.7000 250.3000 248.3000 253.7000 ;
	    RECT 250.8000 253.6000 251.6000 253.7000 ;
	    RECT 250.8000 251.6000 251.6000 252.4000 ;
	    RECT 252.4000 252.3000 253.2000 252.4000 ;
	    RECT 252.4000 251.7000 254.7000 252.3000 ;
	    RECT 252.4000 251.6000 253.2000 251.7000 ;
	    RECT 242.9000 249.7000 248.3000 250.3000 ;
	    RECT 242.9000 248.4000 243.5000 249.7000 ;
	    RECT 249.2000 249.6000 250.0000 250.4000 ;
	    RECT 250.9000 250.3000 251.5000 251.6000 ;
	    RECT 250.9000 249.7000 253.1000 250.3000 ;
	    RECT 238.0000 247.6000 238.8000 248.4000 ;
	    RECT 239.6000 247.6000 240.4000 248.4000 ;
	    RECT 242.8000 247.6000 243.6000 248.4000 ;
	    RECT 244.4000 247.6000 245.2000 248.4000 ;
	    RECT 246.0000 247.6000 246.8000 248.4000 ;
	    RECT 244.5000 238.4000 245.1000 247.6000 ;
	    RECT 244.4000 237.6000 245.2000 238.4000 ;
	    RECT 238.0000 235.6000 238.8000 236.4000 ;
	    RECT 238.1000 230.4000 238.7000 235.6000 ;
	    RECT 236.4000 229.6000 237.2000 230.4000 ;
	    RECT 238.0000 229.6000 238.8000 230.4000 ;
	    RECT 242.8000 229.6000 243.6000 230.4000 ;
	    RECT 233.2000 227.7000 235.5000 228.3000 ;
	    RECT 233.2000 227.6000 234.0000 227.7000 ;
	    RECT 231.6000 223.6000 232.4000 224.4000 ;
	    RECT 233.3000 220.4000 233.9000 227.6000 ;
	    RECT 234.8000 225.6000 235.6000 226.4000 ;
	    RECT 238.0000 225.6000 238.8000 226.4000 ;
	    RECT 233.2000 219.6000 234.0000 220.4000 ;
	    RECT 233.2000 207.6000 234.0000 208.4000 ;
	    RECT 230.0000 205.6000 230.8000 206.4000 ;
	    RECT 231.6000 205.6000 232.4000 206.4000 ;
	    RECT 217.2000 199.6000 218.0000 200.4000 ;
	    RECT 214.0000 197.6000 214.8000 198.4000 ;
	    RECT 217.2000 197.6000 218.0000 198.4000 ;
	    RECT 202.8000 195.6000 203.6000 196.4000 ;
	    RECT 206.0000 195.6000 206.8000 196.4000 ;
	    RECT 210.8000 195.6000 211.6000 196.4000 ;
	    RECT 199.7000 193.7000 201.9000 194.3000 ;
	    RECT 196.4000 191.6000 197.2000 192.4000 ;
	    RECT 185.2000 189.6000 186.0000 190.4000 ;
	    RECT 188.4000 189.6000 189.2000 190.4000 ;
	    RECT 191.6000 189.6000 192.4000 190.4000 ;
	    RECT 194.8000 189.6000 195.6000 190.4000 ;
	    RECT 196.4000 189.6000 197.2000 190.4000 ;
	    RECT 198.0000 189.6000 198.8000 190.4000 ;
	    RECT 182.0000 187.6000 182.8000 188.4000 ;
	    RECT 183.6000 187.6000 184.4000 188.4000 ;
	    RECT 180.4000 185.6000 181.2000 186.4000 ;
	    RECT 182.0000 183.6000 182.8000 184.4000 ;
	    RECT 178.9000 181.7000 181.1000 182.3000 ;
	    RECT 170.8000 171.8000 171.6000 172.6000 ;
	    RECT 172.4000 166.2000 173.2000 177.8000 ;
	    RECT 177.2000 177.6000 178.0000 178.4000 ;
	    RECT 175.6000 170.2000 176.4000 175.8000 ;
	    RECT 180.5000 172.4000 181.1000 181.7000 ;
	    RECT 180.4000 171.6000 181.2000 172.4000 ;
	    RECT 180.5000 170.4000 181.1000 171.6000 ;
	    RECT 180.4000 169.6000 181.2000 170.4000 ;
	    RECT 162.9000 163.7000 165.1000 164.3000 ;
	    RECT 162.9000 158.4000 163.5000 163.7000 ;
	    RECT 166.0000 163.6000 166.8000 164.4000 ;
	    RECT 177.2000 163.6000 178.0000 164.4000 ;
	    RECT 167.6000 161.6000 168.4000 162.4000 ;
	    RECT 164.4000 159.6000 165.2000 160.4000 ;
	    RECT 162.8000 157.6000 163.6000 158.4000 ;
	    RECT 164.5000 152.3000 165.1000 159.6000 ;
	    RECT 162.9000 151.7000 165.1000 152.3000 ;
	    RECT 162.9000 150.4000 163.5000 151.7000 ;
	    RECT 162.8000 149.6000 163.6000 150.4000 ;
	    RECT 164.4000 149.6000 165.2000 150.4000 ;
	    RECT 167.7000 148.3000 168.3000 161.6000 ;
	    RECT 169.2000 155.6000 170.0000 156.4000 ;
	    RECT 170.8000 155.6000 171.6000 156.4000 ;
	    RECT 175.6000 155.6000 176.4000 156.4000 ;
	    RECT 169.3000 148.4000 169.9000 155.6000 ;
	    RECT 170.9000 152.4000 171.5000 155.6000 ;
	    RECT 170.8000 151.6000 171.6000 152.4000 ;
	    RECT 174.0000 151.6000 174.8000 152.4000 ;
	    RECT 175.7000 150.4000 176.3000 155.6000 ;
	    RECT 170.8000 149.6000 171.6000 150.4000 ;
	    RECT 172.4000 149.6000 173.2000 150.4000 ;
	    RECT 175.6000 149.6000 176.4000 150.4000 ;
	    RECT 161.3000 147.7000 165.1000 148.3000 ;
	    RECT 156.5000 145.7000 158.7000 146.3000 ;
	    RECT 158.1000 144.3000 158.7000 145.7000 ;
	    RECT 159.6000 145.6000 160.4000 146.4000 ;
	    RECT 162.8000 145.6000 163.6000 146.4000 ;
	    RECT 162.9000 144.3000 163.5000 145.6000 ;
	    RECT 158.1000 143.7000 163.5000 144.3000 ;
	    RECT 151.6000 137.6000 152.4000 138.4000 ;
	    RECT 150.0000 135.6000 150.8000 136.4000 ;
	    RECT 150.1000 134.4000 150.7000 135.6000 ;
	    RECT 148.4000 133.6000 149.2000 134.4000 ;
	    RECT 150.0000 133.6000 150.8000 134.4000 ;
	    RECT 148.5000 128.4000 149.1000 133.6000 ;
	    RECT 151.7000 132.4000 152.3000 137.6000 ;
	    RECT 161.2000 134.3000 162.0000 134.4000 ;
	    RECT 158.1000 133.7000 162.0000 134.3000 ;
	    RECT 150.0000 131.6000 150.8000 132.4000 ;
	    RECT 151.6000 131.6000 152.4000 132.4000 ;
	    RECT 158.1000 132.3000 158.7000 133.7000 ;
	    RECT 161.2000 133.6000 162.0000 133.7000 ;
	    RECT 153.3000 131.7000 158.7000 132.3000 ;
	    RECT 150.1000 130.3000 150.7000 131.6000 ;
	    RECT 153.3000 130.3000 153.9000 131.7000 ;
	    RECT 161.2000 131.6000 162.0000 132.4000 ;
	    RECT 150.1000 129.7000 153.9000 130.3000 ;
	    RECT 154.8000 129.6000 155.6000 130.4000 ;
	    RECT 148.4000 127.6000 149.2000 128.4000 ;
	    RECT 151.6000 127.6000 152.4000 128.4000 ;
	    RECT 146.9000 125.7000 149.1000 126.3000 ;
	    RECT 146.8000 121.6000 147.6000 122.4000 ;
	    RECT 137.2000 113.6000 138.0000 114.4000 ;
	    RECT 142.0000 113.6000 142.8000 114.4000 ;
	    RECT 137.3000 112.4000 137.9000 113.6000 ;
	    RECT 137.2000 111.6000 138.0000 112.4000 ;
	    RECT 137.2000 107.6000 138.0000 108.4000 ;
	    RECT 135.6000 97.6000 136.4000 98.4000 ;
	    RECT 137.3000 94.4000 137.9000 107.6000 ;
	    RECT 138.8000 103.6000 139.6000 104.4000 ;
	    RECT 142.0000 103.6000 142.8000 104.4000 ;
	    RECT 143.6000 104.2000 144.4000 115.8000 ;
	    RECT 145.2000 109.6000 146.0000 110.4000 ;
	    RECT 138.9000 98.4000 139.5000 103.6000 ;
	    RECT 138.8000 97.6000 139.6000 98.4000 ;
	    RECT 138.8000 95.6000 139.6000 96.4000 ;
	    RECT 138.9000 94.4000 139.5000 95.6000 ;
	    RECT 137.2000 93.6000 138.0000 94.4000 ;
	    RECT 138.8000 93.6000 139.6000 94.4000 ;
	    RECT 137.3000 92.4000 137.9000 93.6000 ;
	    RECT 142.1000 92.4000 142.7000 103.6000 ;
	    RECT 145.3000 102.3000 145.9000 109.6000 ;
	    RECT 143.7000 101.7000 145.9000 102.3000 ;
	    RECT 134.0000 91.6000 134.8000 92.4000 ;
	    RECT 135.6000 91.6000 136.4000 92.4000 ;
	    RECT 137.2000 91.6000 138.0000 92.4000 ;
	    RECT 138.8000 91.6000 139.6000 92.4000 ;
	    RECT 142.0000 91.6000 142.8000 92.4000 ;
	    RECT 134.0000 83.6000 134.8000 84.4000 ;
	    RECT 134.1000 72.4000 134.7000 83.6000 ;
	    RECT 135.7000 82.4000 136.3000 91.6000 ;
	    RECT 138.9000 90.4000 139.5000 91.6000 ;
	    RECT 138.8000 89.6000 139.6000 90.4000 ;
	    RECT 140.4000 89.6000 141.2000 90.4000 ;
	    RECT 140.5000 88.3000 141.1000 89.6000 ;
	    RECT 138.9000 87.7000 141.1000 88.3000 ;
	    RECT 135.6000 81.6000 136.4000 82.4000 ;
	    RECT 138.9000 78.4000 139.5000 87.7000 ;
	    RECT 138.8000 77.6000 139.6000 78.4000 ;
	    RECT 140.4000 73.6000 141.2000 74.4000 ;
	    RECT 134.0000 71.6000 134.8000 72.4000 ;
	    RECT 140.5000 70.4000 141.1000 73.6000 ;
	    RECT 124.4000 70.3000 125.2000 70.4000 ;
	    RECT 122.9000 69.7000 125.2000 70.3000 ;
	    RECT 124.4000 69.6000 125.2000 69.7000 ;
	    RECT 126.0000 69.6000 126.8000 70.4000 ;
	    RECT 127.6000 69.6000 128.4000 70.4000 ;
	    RECT 130.8000 69.6000 131.6000 70.4000 ;
	    RECT 132.4000 69.6000 133.2000 70.4000 ;
	    RECT 134.0000 69.6000 134.8000 70.4000 ;
	    RECT 135.6000 69.6000 136.4000 70.4000 ;
	    RECT 140.4000 69.6000 141.2000 70.4000 ;
	    RECT 126.1000 68.4000 126.7000 69.6000 ;
	    RECT 126.0000 67.6000 126.8000 68.4000 ;
	    RECT 122.8000 63.6000 123.6000 64.4000 ;
	    RECT 122.9000 58.4000 123.5000 63.6000 ;
	    RECT 127.7000 58.4000 128.3000 69.6000 ;
	    RECT 132.5000 66.4000 133.1000 69.6000 ;
	    RECT 135.7000 68.4000 136.3000 69.6000 ;
	    RECT 135.6000 67.6000 136.4000 68.4000 ;
	    RECT 142.0000 67.6000 142.8000 68.4000 ;
	    RECT 132.4000 65.6000 133.2000 66.4000 ;
	    RECT 134.0000 61.6000 134.8000 62.4000 ;
	    RECT 122.8000 57.6000 123.6000 58.4000 ;
	    RECT 127.6000 57.6000 128.4000 58.4000 ;
	    RECT 134.1000 54.4000 134.7000 61.6000 ;
	    RECT 135.7000 58.4000 136.3000 67.6000 ;
	    RECT 135.6000 57.6000 136.4000 58.4000 ;
	    RECT 134.0000 54.3000 134.8000 54.4000 ;
	    RECT 134.0000 53.7000 136.3000 54.3000 ;
	    RECT 134.0000 53.6000 134.8000 53.7000 ;
	    RECT 126.0000 51.6000 126.8000 52.4000 ;
	    RECT 134.0000 51.6000 134.8000 52.4000 ;
	    RECT 124.4000 39.6000 125.2000 40.4000 ;
	    RECT 124.5000 30.4000 125.1000 39.6000 ;
	    RECT 124.4000 29.6000 125.2000 30.4000 ;
	    RECT 126.1000 28.4000 126.7000 51.6000 ;
	    RECT 129.2000 49.6000 130.0000 50.4000 ;
	    RECT 129.3000 44.4000 129.9000 49.6000 ;
	    RECT 129.2000 43.6000 130.0000 44.4000 ;
	    RECT 132.4000 43.6000 133.2000 44.4000 ;
	    RECT 134.1000 40.3000 134.7000 51.6000 ;
	    RECT 132.5000 39.7000 134.7000 40.3000 ;
	    RECT 126.0000 27.6000 126.8000 28.4000 ;
	    RECT 124.4000 23.6000 125.2000 24.4000 ;
	    RECT 127.6000 24.2000 128.4000 35.8000 ;
	    RECT 132.5000 32.4000 133.1000 39.7000 ;
	    RECT 134.0000 37.6000 134.8000 38.4000 ;
	    RECT 130.8000 26.2000 131.6000 31.8000 ;
	    RECT 132.4000 31.6000 133.2000 32.4000 ;
	    RECT 134.0000 31.6000 134.8000 32.4000 ;
	    RECT 134.1000 30.4000 134.7000 31.6000 ;
	    RECT 135.7000 30.4000 136.3000 53.7000 ;
	    RECT 140.4000 46.2000 141.2000 57.8000 ;
	    RECT 143.7000 54.4000 144.3000 101.7000 ;
	    RECT 145.2000 91.6000 146.0000 92.4000 ;
	    RECT 145.3000 90.4000 145.9000 91.6000 ;
	    RECT 145.2000 89.6000 146.0000 90.4000 ;
	    RECT 146.9000 72.4000 147.5000 121.6000 ;
	    RECT 148.5000 118.4000 149.1000 125.7000 ;
	    RECT 148.4000 117.6000 149.2000 118.4000 ;
	    RECT 148.4000 115.6000 149.2000 116.4000 ;
	    RECT 148.5000 102.4000 149.1000 115.6000 ;
	    RECT 151.6000 109.4000 152.4000 110.4000 ;
	    RECT 151.6000 105.6000 152.4000 106.4000 ;
	    RECT 148.4000 101.6000 149.2000 102.4000 ;
	    RECT 151.7000 102.3000 152.3000 105.6000 ;
	    RECT 153.2000 104.2000 154.0000 115.8000 ;
	    RECT 154.9000 114.4000 155.5000 129.6000 ;
	    RECT 156.4000 123.6000 157.2000 124.4000 ;
	    RECT 156.5000 116.4000 157.1000 123.6000 ;
	    RECT 158.0000 119.6000 158.8000 120.4000 ;
	    RECT 158.1000 116.4000 158.7000 119.6000 ;
	    RECT 156.4000 115.6000 157.2000 116.4000 ;
	    RECT 158.0000 115.6000 158.8000 116.4000 ;
	    RECT 154.8000 113.6000 155.6000 114.4000 ;
	    RECT 159.6000 113.6000 160.4000 114.4000 ;
	    RECT 156.4000 106.2000 157.2000 111.8000 ;
	    RECT 158.0000 107.6000 158.8000 108.4000 ;
	    RECT 151.7000 101.7000 153.9000 102.3000 ;
	    RECT 148.5000 92.4000 149.1000 101.6000 ;
	    RECT 153.3000 98.4000 153.9000 101.7000 ;
	    RECT 158.1000 98.4000 158.7000 107.6000 ;
	    RECT 150.0000 97.6000 150.8000 98.4000 ;
	    RECT 153.2000 97.6000 154.0000 98.4000 ;
	    RECT 158.0000 97.6000 158.8000 98.4000 ;
	    RECT 150.1000 94.4000 150.7000 97.6000 ;
	    RECT 150.0000 93.6000 150.8000 94.4000 ;
	    RECT 151.6000 93.6000 152.4000 94.4000 ;
	    RECT 151.7000 92.4000 152.3000 93.6000 ;
	    RECT 159.7000 92.4000 160.3000 113.6000 ;
	    RECT 161.2000 111.6000 162.0000 112.4000 ;
	    RECT 161.2000 109.6000 162.0000 110.4000 ;
	    RECT 161.3000 108.4000 161.9000 109.6000 ;
	    RECT 161.2000 107.6000 162.0000 108.4000 ;
	    RECT 164.5000 100.3000 165.1000 147.7000 ;
	    RECT 166.1000 147.7000 168.3000 148.3000 ;
	    RECT 166.1000 136.4000 166.7000 147.7000 ;
	    RECT 169.2000 147.6000 170.0000 148.4000 ;
	    RECT 167.6000 145.6000 168.4000 146.4000 ;
	    RECT 167.7000 142.4000 168.3000 145.6000 ;
	    RECT 172.5000 142.4000 173.1000 149.6000 ;
	    RECT 167.6000 141.6000 168.4000 142.4000 ;
	    RECT 172.4000 141.6000 173.2000 142.4000 ;
	    RECT 172.4000 137.6000 173.2000 138.4000 ;
	    RECT 174.0000 137.6000 174.8000 138.4000 ;
	    RECT 174.1000 136.4000 174.7000 137.6000 ;
	    RECT 166.0000 135.6000 166.8000 136.4000 ;
	    RECT 174.0000 135.6000 174.8000 136.4000 ;
	    RECT 174.0000 133.6000 174.8000 134.4000 ;
	    RECT 177.3000 132.4000 177.9000 163.6000 ;
	    RECT 180.4000 159.6000 181.2000 160.4000 ;
	    RECT 180.5000 150.4000 181.1000 159.6000 ;
	    RECT 182.1000 152.4000 182.7000 183.6000 ;
	    RECT 185.3000 182.4000 185.9000 189.6000 ;
	    RECT 188.5000 184.4000 189.1000 189.6000 ;
	    RECT 194.9000 184.4000 195.5000 189.6000 ;
	    RECT 196.5000 188.4000 197.1000 189.6000 ;
	    RECT 196.4000 187.6000 197.2000 188.4000 ;
	    RECT 198.1000 186.3000 198.7000 189.6000 ;
	    RECT 196.5000 185.7000 198.7000 186.3000 ;
	    RECT 188.4000 183.6000 189.2000 184.4000 ;
	    RECT 194.8000 183.6000 195.6000 184.4000 ;
	    RECT 185.2000 181.6000 186.0000 182.4000 ;
	    RECT 194.8000 181.6000 195.6000 182.4000 ;
	    RECT 188.4000 177.6000 189.2000 178.4000 ;
	    RECT 183.6000 173.6000 184.4000 174.4000 ;
	    RECT 183.7000 172.4000 184.3000 173.6000 ;
	    RECT 188.5000 172.4000 189.1000 177.6000 ;
	    RECT 183.6000 171.6000 184.4000 172.4000 ;
	    RECT 188.4000 171.6000 189.2000 172.4000 ;
	    RECT 190.0000 171.6000 190.8000 172.4000 ;
	    RECT 193.2000 171.6000 194.0000 172.4000 ;
	    RECT 185.2000 163.6000 186.0000 164.4000 ;
	    RECT 185.3000 158.4000 185.9000 163.6000 ;
	    RECT 190.1000 160.4000 190.7000 171.6000 ;
	    RECT 191.6000 169.6000 192.4000 170.4000 ;
	    RECT 190.0000 159.6000 190.8000 160.4000 ;
	    RECT 185.2000 157.6000 186.0000 158.4000 ;
	    RECT 191.7000 156.4000 192.3000 169.6000 ;
	    RECT 194.9000 166.4000 195.5000 181.6000 ;
	    RECT 194.8000 165.6000 195.6000 166.4000 ;
	    RECT 194.8000 163.6000 195.6000 164.4000 ;
	    RECT 194.9000 158.4000 195.5000 163.6000 ;
	    RECT 194.8000 157.6000 195.6000 158.4000 ;
	    RECT 185.2000 155.6000 186.0000 156.4000 ;
	    RECT 191.6000 155.6000 192.4000 156.4000 ;
	    RECT 182.0000 151.6000 182.8000 152.4000 ;
	    RECT 183.6000 151.6000 184.4000 152.4000 ;
	    RECT 188.4000 151.6000 189.2000 152.4000 ;
	    RECT 194.8000 151.6000 195.6000 152.4000 ;
	    RECT 180.4000 149.6000 181.2000 150.4000 ;
	    RECT 182.1000 148.4000 182.7000 151.6000 ;
	    RECT 183.7000 150.4000 184.3000 151.6000 ;
	    RECT 194.9000 150.4000 195.5000 151.6000 ;
	    RECT 183.6000 149.6000 184.4000 150.4000 ;
	    RECT 188.4000 149.6000 189.2000 150.4000 ;
	    RECT 190.0000 149.6000 190.8000 150.4000 ;
	    RECT 191.6000 149.6000 192.4000 150.4000 ;
	    RECT 194.8000 149.6000 195.6000 150.4000 ;
	    RECT 182.0000 147.6000 182.8000 148.4000 ;
	    RECT 183.7000 146.4000 184.3000 149.6000 ;
	    RECT 183.6000 145.6000 184.4000 146.4000 ;
	    RECT 180.4000 143.6000 181.2000 144.4000 ;
	    RECT 180.5000 142.4000 181.1000 143.6000 ;
	    RECT 188.5000 142.4000 189.1000 149.6000 ;
	    RECT 191.7000 146.4000 192.3000 149.6000 ;
	    RECT 193.2000 147.6000 194.0000 148.4000 ;
	    RECT 191.6000 145.6000 192.4000 146.4000 ;
	    RECT 180.4000 141.6000 181.2000 142.4000 ;
	    RECT 188.4000 141.6000 189.2000 142.4000 ;
	    RECT 193.3000 138.4000 193.9000 147.6000 ;
	    RECT 194.8000 142.3000 195.6000 142.4000 ;
	    RECT 196.5000 142.3000 197.1000 185.7000 ;
	    RECT 199.7000 182.4000 200.3000 193.7000 ;
	    RECT 204.4000 191.6000 205.2000 192.4000 ;
	    RECT 204.5000 190.4000 205.1000 191.6000 ;
	    RECT 204.4000 189.6000 205.2000 190.4000 ;
	    RECT 202.8000 187.6000 203.6000 188.4000 ;
	    RECT 201.2000 185.6000 202.0000 186.4000 ;
	    RECT 199.6000 181.6000 200.4000 182.4000 ;
	    RECT 201.3000 180.4000 201.9000 185.6000 ;
	    RECT 201.2000 179.6000 202.0000 180.4000 ;
	    RECT 198.0000 177.6000 198.8000 178.4000 ;
	    RECT 198.1000 172.4000 198.7000 177.6000 ;
	    RECT 202.9000 172.4000 203.5000 187.6000 ;
	    RECT 206.1000 176.3000 206.7000 195.6000 ;
	    RECT 207.6000 191.6000 208.4000 192.4000 ;
	    RECT 210.9000 190.4000 211.5000 195.6000 ;
	    RECT 217.3000 192.4000 217.9000 197.6000 ;
	    RECT 218.8000 195.6000 219.6000 196.4000 ;
	    RECT 220.5000 192.4000 221.1000 205.6000 ;
	    RECT 230.0000 199.6000 230.8000 200.4000 ;
	    RECT 225.2000 195.6000 226.0000 196.4000 ;
	    RECT 217.2000 191.6000 218.0000 192.4000 ;
	    RECT 220.4000 191.6000 221.2000 192.4000 ;
	    RECT 228.4000 191.6000 229.2000 192.4000 ;
	    RECT 210.8000 189.6000 211.6000 190.4000 ;
	    RECT 214.0000 189.6000 214.8000 190.4000 ;
	    RECT 215.6000 189.6000 216.4000 190.4000 ;
	    RECT 214.1000 188.4000 214.7000 189.6000 ;
	    RECT 207.6000 187.6000 208.4000 188.4000 ;
	    RECT 212.4000 187.6000 213.2000 188.4000 ;
	    RECT 214.0000 187.6000 214.8000 188.4000 ;
	    RECT 207.7000 178.4000 208.3000 187.6000 ;
	    RECT 207.6000 177.6000 208.4000 178.4000 ;
	    RECT 212.5000 176.4000 213.1000 187.6000 ;
	    RECT 214.0000 177.6000 214.8000 178.4000 ;
	    RECT 204.5000 175.7000 206.7000 176.3000 ;
	    RECT 204.5000 172.4000 205.1000 175.7000 ;
	    RECT 212.4000 175.6000 213.2000 176.4000 ;
	    RECT 214.1000 174.4000 214.7000 177.6000 ;
	    RECT 206.0000 173.6000 206.8000 174.4000 ;
	    RECT 214.0000 173.6000 214.8000 174.4000 ;
	    RECT 198.0000 171.6000 198.8000 172.4000 ;
	    RECT 199.6000 171.6000 200.4000 172.4000 ;
	    RECT 202.8000 172.3000 203.6000 172.4000 ;
	    RECT 201.3000 171.7000 203.6000 172.3000 ;
	    RECT 199.7000 170.3000 200.3000 171.6000 ;
	    RECT 198.1000 169.7000 200.3000 170.3000 ;
	    RECT 198.1000 166.4000 198.7000 169.7000 ;
	    RECT 198.0000 165.6000 198.8000 166.4000 ;
	    RECT 201.3000 166.3000 201.9000 171.7000 ;
	    RECT 202.8000 171.6000 203.6000 171.7000 ;
	    RECT 204.4000 171.6000 205.2000 172.4000 ;
	    RECT 202.8000 169.6000 203.6000 170.4000 ;
	    RECT 199.7000 165.7000 201.9000 166.3000 ;
	    RECT 199.7000 160.4000 200.3000 165.7000 ;
	    RECT 201.2000 163.6000 202.0000 164.4000 ;
	    RECT 201.3000 160.4000 201.9000 163.6000 ;
	    RECT 199.6000 159.6000 200.4000 160.4000 ;
	    RECT 201.2000 159.6000 202.0000 160.4000 ;
	    RECT 198.0000 157.6000 198.8000 158.4000 ;
	    RECT 199.6000 153.6000 200.4000 154.4000 ;
	    RECT 201.2000 153.6000 202.0000 154.4000 ;
	    RECT 198.0000 149.6000 198.8000 150.4000 ;
	    RECT 199.7000 148.4000 200.3000 153.6000 ;
	    RECT 201.3000 152.4000 201.9000 153.6000 ;
	    RECT 201.2000 151.6000 202.0000 152.4000 ;
	    RECT 199.6000 147.6000 200.4000 148.4000 ;
	    RECT 201.2000 145.6000 202.0000 146.4000 ;
	    RECT 194.8000 141.7000 197.1000 142.3000 ;
	    RECT 194.8000 141.6000 195.6000 141.7000 ;
	    RECT 198.0000 141.6000 198.8000 142.4000 ;
	    RECT 194.9000 138.4000 195.5000 141.6000 ;
	    RECT 178.8000 137.6000 179.6000 138.4000 ;
	    RECT 193.2000 137.6000 194.0000 138.4000 ;
	    RECT 194.8000 137.6000 195.6000 138.4000 ;
	    RECT 178.9000 136.4000 179.5000 137.6000 ;
	    RECT 178.8000 135.6000 179.6000 136.4000 ;
	    RECT 180.4000 135.6000 181.2000 136.4000 ;
	    RECT 186.8000 135.6000 187.6000 136.4000 ;
	    RECT 169.2000 131.6000 170.0000 132.4000 ;
	    RECT 170.8000 131.6000 171.6000 132.4000 ;
	    RECT 174.0000 131.6000 174.8000 132.4000 ;
	    RECT 175.6000 131.6000 176.4000 132.4000 ;
	    RECT 177.2000 131.6000 178.0000 132.4000 ;
	    RECT 178.8000 131.6000 179.6000 132.4000 ;
	    RECT 167.6000 129.6000 168.4000 130.4000 ;
	    RECT 169.3000 112.4000 169.9000 131.6000 ;
	    RECT 166.0000 111.6000 166.8000 112.4000 ;
	    RECT 169.2000 111.6000 170.0000 112.4000 ;
	    RECT 166.1000 110.4000 166.7000 111.6000 ;
	    RECT 169.3000 110.4000 169.9000 111.6000 ;
	    RECT 174.1000 110.4000 174.7000 131.6000 ;
	    RECT 175.7000 112.4000 176.3000 131.6000 ;
	    RECT 178.9000 124.4000 179.5000 131.6000 ;
	    RECT 178.8000 123.6000 179.6000 124.4000 ;
	    RECT 180.4000 123.6000 181.2000 124.4000 ;
	    RECT 185.2000 123.6000 186.0000 124.4000 ;
	    RECT 177.2000 119.6000 178.0000 120.4000 ;
	    RECT 175.6000 111.6000 176.4000 112.4000 ;
	    RECT 166.0000 109.6000 166.8000 110.4000 ;
	    RECT 169.2000 109.6000 170.0000 110.4000 ;
	    RECT 174.0000 109.6000 174.8000 110.4000 ;
	    RECT 169.2000 107.6000 170.0000 108.4000 ;
	    RECT 166.0000 105.6000 166.8000 106.4000 ;
	    RECT 161.3000 99.7000 165.1000 100.3000 ;
	    RECT 148.4000 91.6000 149.2000 92.4000 ;
	    RECT 151.6000 91.6000 152.4000 92.4000 ;
	    RECT 153.2000 91.6000 154.0000 92.4000 ;
	    RECT 158.0000 91.6000 158.8000 92.4000 ;
	    RECT 159.6000 91.6000 160.4000 92.4000 ;
	    RECT 153.3000 90.4000 153.9000 91.6000 ;
	    RECT 153.2000 89.6000 154.0000 90.4000 ;
	    RECT 158.1000 88.3000 158.7000 91.6000 ;
	    RECT 159.7000 90.4000 160.3000 91.6000 ;
	    RECT 159.6000 89.6000 160.4000 90.4000 ;
	    RECT 161.3000 90.3000 161.9000 99.7000 ;
	    RECT 166.1000 98.4000 166.7000 105.6000 ;
	    RECT 162.8000 97.6000 163.6000 98.4000 ;
	    RECT 166.0000 97.6000 166.8000 98.4000 ;
	    RECT 162.9000 92.4000 163.5000 97.6000 ;
	    RECT 166.0000 95.6000 166.8000 96.4000 ;
	    RECT 167.6000 95.6000 168.4000 96.4000 ;
	    RECT 164.4000 93.6000 165.2000 94.4000 ;
	    RECT 162.8000 91.6000 163.6000 92.4000 ;
	    RECT 161.3000 89.7000 165.1000 90.3000 ;
	    RECT 162.8000 88.3000 163.6000 88.4000 ;
	    RECT 158.1000 87.7000 163.6000 88.3000 ;
	    RECT 162.8000 87.6000 163.6000 87.7000 ;
	    RECT 153.2000 85.6000 154.0000 86.4000 ;
	    RECT 146.8000 71.6000 147.6000 72.4000 ;
	    RECT 146.9000 70.4000 147.5000 71.6000 ;
	    RECT 146.8000 69.6000 147.6000 70.4000 ;
	    RECT 151.6000 69.6000 152.4000 70.4000 ;
	    RECT 153.3000 68.4000 153.9000 85.6000 ;
	    RECT 158.0000 73.6000 158.8000 74.4000 ;
	    RECT 158.1000 72.4000 158.7000 73.6000 ;
	    RECT 158.0000 71.6000 158.8000 72.4000 ;
	    RECT 159.6000 71.6000 160.4000 72.4000 ;
	    RECT 154.8000 69.6000 155.6000 70.4000 ;
	    RECT 153.2000 67.6000 154.0000 68.4000 ;
	    RECT 148.4000 63.6000 149.2000 64.4000 ;
	    RECT 143.6000 53.6000 144.4000 54.4000 ;
	    RECT 145.2000 53.6000 146.0000 54.4000 ;
	    RECT 142.0000 51.6000 142.8000 52.4000 ;
	    RECT 137.2000 31.6000 138.0000 32.4000 ;
	    RECT 134.0000 29.6000 134.8000 30.4000 ;
	    RECT 135.6000 29.6000 136.4000 30.4000 ;
	    RECT 135.7000 28.4000 136.3000 29.6000 ;
	    RECT 132.4000 27.6000 133.2000 28.4000 ;
	    RECT 135.6000 27.6000 136.4000 28.4000 ;
	    RECT 130.8000 23.6000 131.6000 24.4000 ;
	    RECT 124.5000 14.4000 125.1000 23.6000 ;
	    RECT 126.0000 17.6000 126.8000 18.4000 ;
	    RECT 129.2000 15.6000 130.0000 16.4000 ;
	    RECT 121.2000 13.6000 122.0000 14.4000 ;
	    RECT 124.4000 13.6000 125.2000 14.4000 ;
	    RECT 129.3000 12.4000 129.9000 15.6000 ;
	    RECT 130.9000 14.4000 131.5000 23.6000 ;
	    RECT 137.3000 18.4000 137.9000 31.6000 ;
	    RECT 140.4000 25.6000 141.2000 26.4000 ;
	    RECT 138.8000 24.3000 139.6000 24.4000 ;
	    RECT 140.5000 24.3000 141.1000 25.6000 ;
	    RECT 138.8000 23.7000 141.1000 24.3000 ;
	    RECT 143.6000 24.2000 144.4000 35.8000 ;
	    RECT 145.3000 30.4000 145.9000 53.6000 ;
	    RECT 148.5000 52.6000 149.1000 63.6000 ;
	    RECT 148.4000 51.8000 149.2000 52.6000 ;
	    RECT 150.0000 46.2000 150.8000 57.8000 ;
	    RECT 151.6000 51.6000 152.4000 52.4000 ;
	    RECT 145.2000 29.6000 146.0000 30.4000 ;
	    RECT 151.7000 30.2000 152.3000 51.6000 ;
	    RECT 153.2000 50.2000 154.0000 55.8000 ;
	    RECT 154.9000 54.4000 155.5000 69.6000 ;
	    RECT 158.1000 62.4000 158.7000 71.6000 ;
	    RECT 159.7000 70.4000 160.3000 71.6000 ;
	    RECT 159.6000 69.6000 160.4000 70.4000 ;
	    RECT 162.8000 69.6000 163.6000 70.4000 ;
	    RECT 164.5000 68.4000 165.1000 89.7000 ;
	    RECT 166.0000 88.3000 166.8000 88.4000 ;
	    RECT 167.7000 88.3000 168.3000 95.6000 ;
	    RECT 169.3000 88.4000 169.9000 107.6000 ;
	    RECT 177.3000 106.4000 177.9000 119.6000 ;
	    RECT 178.8000 109.6000 179.6000 110.4000 ;
	    RECT 172.4000 105.6000 173.2000 106.4000 ;
	    RECT 177.2000 105.6000 178.0000 106.4000 ;
	    RECT 178.8000 105.6000 179.6000 106.4000 ;
	    RECT 170.8000 103.6000 171.6000 104.4000 ;
	    RECT 172.4000 103.6000 173.2000 104.4000 ;
	    RECT 175.6000 103.6000 176.4000 104.4000 ;
	    RECT 172.5000 98.4000 173.1000 103.6000 ;
	    RECT 172.4000 97.6000 173.2000 98.4000 ;
	    RECT 174.0000 97.6000 174.8000 98.4000 ;
	    RECT 174.1000 92.4000 174.7000 97.6000 ;
	    RECT 175.7000 96.4000 176.3000 103.6000 ;
	    RECT 175.6000 95.6000 176.4000 96.4000 ;
	    RECT 175.6000 93.6000 176.4000 94.4000 ;
	    RECT 177.2000 93.6000 178.0000 94.4000 ;
	    RECT 177.3000 92.4000 177.9000 93.6000 ;
	    RECT 178.9000 92.4000 179.5000 105.6000 ;
	    RECT 170.8000 92.3000 171.6000 92.4000 ;
	    RECT 170.8000 91.7000 173.1000 92.3000 ;
	    RECT 170.8000 91.6000 171.6000 91.7000 ;
	    RECT 170.8000 89.6000 171.6000 90.4000 ;
	    RECT 172.5000 90.3000 173.1000 91.7000 ;
	    RECT 174.0000 91.6000 174.8000 92.4000 ;
	    RECT 177.2000 91.6000 178.0000 92.4000 ;
	    RECT 178.8000 91.6000 179.6000 92.4000 ;
	    RECT 178.8000 90.3000 179.6000 90.4000 ;
	    RECT 172.5000 89.7000 179.6000 90.3000 ;
	    RECT 178.8000 89.6000 179.6000 89.7000 ;
	    RECT 166.0000 87.7000 168.3000 88.3000 ;
	    RECT 166.0000 87.6000 166.8000 87.7000 ;
	    RECT 169.2000 87.6000 170.0000 88.4000 ;
	    RECT 167.6000 83.6000 168.4000 84.4000 ;
	    RECT 174.0000 83.6000 174.8000 84.4000 ;
	    RECT 167.7000 80.4000 168.3000 83.6000 ;
	    RECT 167.6000 79.6000 168.4000 80.4000 ;
	    RECT 169.2000 79.6000 170.0000 80.4000 ;
	    RECT 166.0000 71.6000 166.8000 72.4000 ;
	    RECT 169.3000 70.4000 169.9000 79.6000 ;
	    RECT 174.0000 75.6000 174.8000 76.4000 ;
	    RECT 175.6000 75.6000 176.4000 76.4000 ;
	    RECT 169.2000 69.6000 170.0000 70.4000 ;
	    RECT 174.0000 69.6000 174.8000 70.4000 ;
	    RECT 164.4000 67.6000 165.2000 68.4000 ;
	    RECT 166.0000 67.6000 166.8000 68.4000 ;
	    RECT 170.8000 67.6000 171.6000 68.4000 ;
	    RECT 172.4000 67.6000 173.2000 68.4000 ;
	    RECT 170.9000 66.4000 171.5000 67.6000 ;
	    RECT 170.8000 65.6000 171.6000 66.4000 ;
	    RECT 159.6000 63.6000 160.4000 64.4000 ;
	    RECT 166.0000 63.6000 166.8000 64.4000 ;
	    RECT 158.0000 61.6000 158.8000 62.4000 ;
	    RECT 159.6000 57.6000 160.4000 58.4000 ;
	    RECT 159.7000 54.4000 160.3000 57.6000 ;
	    RECT 166.1000 54.4000 166.7000 63.6000 ;
	    RECT 154.8000 53.6000 155.6000 54.4000 ;
	    RECT 159.6000 53.6000 160.4000 54.4000 ;
	    RECT 161.2000 53.6000 162.0000 54.4000 ;
	    RECT 162.8000 53.6000 163.6000 54.4000 ;
	    RECT 166.0000 53.6000 166.8000 54.4000 ;
	    RECT 170.9000 54.3000 171.5000 65.6000 ;
	    RECT 172.5000 58.4000 173.1000 67.6000 ;
	    RECT 174.1000 60.4000 174.7000 69.6000 ;
	    RECT 175.7000 68.4000 176.3000 75.6000 ;
	    RECT 177.2000 71.6000 178.0000 72.4000 ;
	    RECT 175.6000 67.6000 176.4000 68.4000 ;
	    RECT 177.3000 62.4000 177.9000 71.6000 ;
	    RECT 178.8000 69.6000 179.6000 70.4000 ;
	    RECT 180.5000 70.3000 181.1000 123.6000 ;
	    RECT 185.3000 114.4000 185.9000 123.6000 ;
	    RECT 182.0000 113.6000 182.8000 114.4000 ;
	    RECT 185.2000 113.6000 186.0000 114.4000 ;
	    RECT 182.1000 96.3000 182.7000 113.6000 ;
	    RECT 183.6000 111.6000 184.4000 112.4000 ;
	    RECT 183.7000 108.4000 184.3000 111.6000 ;
	    RECT 186.9000 110.4000 187.5000 135.6000 ;
	    RECT 196.4000 131.6000 197.2000 132.4000 ;
	    RECT 190.0000 123.6000 190.8000 124.4000 ;
	    RECT 194.8000 123.6000 195.6000 124.4000 ;
	    RECT 188.4000 113.6000 189.2000 114.4000 ;
	    RECT 188.5000 112.4000 189.1000 113.6000 ;
	    RECT 188.4000 111.6000 189.2000 112.4000 ;
	    RECT 186.8000 109.6000 187.6000 110.4000 ;
	    RECT 183.6000 107.6000 184.4000 108.4000 ;
	    RECT 186.8000 107.6000 187.6000 108.4000 ;
	    RECT 183.6000 105.6000 184.4000 106.4000 ;
	    RECT 185.2000 103.6000 186.0000 104.4000 ;
	    RECT 186.9000 96.3000 187.5000 107.6000 ;
	    RECT 188.5000 106.4000 189.1000 111.6000 ;
	    RECT 190.1000 108.4000 190.7000 123.6000 ;
	    RECT 193.2000 113.6000 194.0000 114.4000 ;
	    RECT 194.9000 110.4000 195.5000 123.6000 ;
	    RECT 196.5000 110.4000 197.1000 131.6000 ;
	    RECT 198.1000 126.4000 198.7000 141.6000 ;
	    RECT 199.6000 137.6000 200.4000 138.4000 ;
	    RECT 199.7000 134.4000 200.3000 137.6000 ;
	    RECT 199.6000 133.6000 200.4000 134.4000 ;
	    RECT 201.3000 132.4000 201.9000 145.6000 ;
	    RECT 199.6000 131.6000 200.4000 132.4000 ;
	    RECT 201.2000 131.6000 202.0000 132.4000 ;
	    RECT 199.7000 126.4000 200.3000 131.6000 ;
	    RECT 198.0000 125.6000 198.8000 126.4000 ;
	    RECT 199.6000 125.6000 200.4000 126.4000 ;
	    RECT 202.9000 124.4000 203.5000 169.6000 ;
	    RECT 206.1000 166.4000 206.7000 173.6000 ;
	    RECT 215.7000 172.4000 216.3000 189.6000 ;
	    RECT 217.3000 188.4000 217.9000 191.6000 ;
	    RECT 220.4000 189.6000 221.2000 190.4000 ;
	    RECT 217.2000 187.6000 218.0000 188.4000 ;
	    RECT 217.2000 185.6000 218.0000 186.4000 ;
	    RECT 217.3000 180.4000 217.9000 185.6000 ;
	    RECT 220.5000 182.4000 221.1000 189.6000 ;
	    RECT 223.6000 185.6000 224.4000 186.4000 ;
	    RECT 223.7000 182.4000 224.3000 185.6000 ;
	    RECT 228.5000 184.4000 229.1000 191.6000 ;
	    RECT 230.1000 190.4000 230.7000 199.6000 ;
	    RECT 231.7000 196.4000 232.3000 205.6000 ;
	    RECT 231.6000 195.6000 232.4000 196.4000 ;
	    RECT 231.7000 192.4000 232.3000 195.6000 ;
	    RECT 231.6000 191.6000 232.4000 192.4000 ;
	    RECT 230.0000 189.6000 230.8000 190.4000 ;
	    RECT 226.8000 183.6000 227.6000 184.4000 ;
	    RECT 228.4000 183.6000 229.2000 184.4000 ;
	    RECT 230.1000 182.4000 230.7000 189.6000 ;
	    RECT 231.7000 188.4000 232.3000 191.6000 ;
	    RECT 233.3000 190.4000 233.9000 207.6000 ;
	    RECT 236.4000 206.2000 237.2000 217.8000 ;
	    RECT 238.1000 216.4000 238.7000 225.6000 ;
	    RECT 239.6000 223.6000 240.4000 224.4000 ;
	    RECT 239.7000 222.4000 240.3000 223.6000 ;
	    RECT 242.9000 222.4000 243.5000 229.6000 ;
	    RECT 246.1000 224.4000 246.7000 247.6000 ;
	    RECT 249.3000 244.4000 249.9000 249.6000 ;
	    RECT 252.5000 248.4000 253.1000 249.7000 ;
	    RECT 252.4000 247.6000 253.2000 248.4000 ;
	    RECT 247.6000 243.6000 248.4000 244.4000 ;
	    RECT 249.2000 243.6000 250.0000 244.4000 ;
	    RECT 252.4000 243.6000 253.2000 244.4000 ;
	    RECT 247.7000 232.3000 248.3000 243.6000 ;
	    RECT 249.2000 235.6000 250.0000 236.4000 ;
	    RECT 247.7000 231.7000 249.9000 232.3000 ;
	    RECT 247.6000 229.6000 248.4000 230.4000 ;
	    RECT 247.7000 226.4000 248.3000 229.6000 ;
	    RECT 249.3000 228.4000 249.9000 231.7000 ;
	    RECT 250.8000 231.6000 251.6000 232.4000 ;
	    RECT 249.2000 227.6000 250.0000 228.4000 ;
	    RECT 247.6000 225.6000 248.4000 226.4000 ;
	    RECT 249.2000 225.6000 250.0000 226.4000 ;
	    RECT 246.0000 223.6000 246.8000 224.4000 ;
	    RECT 239.6000 221.6000 240.4000 222.4000 ;
	    RECT 242.8000 221.6000 243.6000 222.4000 ;
	    RECT 249.3000 220.4000 249.9000 225.6000 ;
	    RECT 241.2000 219.6000 242.0000 220.4000 ;
	    RECT 244.4000 219.6000 245.2000 220.4000 ;
	    RECT 247.6000 219.6000 248.4000 220.4000 ;
	    RECT 249.2000 219.6000 250.0000 220.4000 ;
	    RECT 241.3000 218.4000 241.9000 219.6000 ;
	    RECT 241.2000 217.6000 242.0000 218.4000 ;
	    RECT 238.0000 215.6000 238.8000 216.4000 ;
	    RECT 244.5000 212.4000 245.1000 219.6000 ;
	    RECT 244.4000 211.6000 245.2000 212.4000 ;
	    RECT 247.7000 210.3000 248.3000 219.6000 ;
	    RECT 249.2000 215.6000 250.0000 216.4000 ;
	    RECT 250.9000 216.3000 251.5000 231.6000 ;
	    RECT 252.5000 230.4000 253.1000 243.6000 ;
	    RECT 254.1000 234.4000 254.7000 251.7000 ;
	    RECT 255.6000 251.6000 256.4000 252.4000 ;
	    RECT 257.2000 251.6000 258.0000 252.4000 ;
	    RECT 257.3000 248.4000 257.9000 251.6000 ;
	    RECT 258.9000 248.4000 259.5000 255.6000 ;
	    RECT 260.5000 252.4000 261.1000 255.6000 ;
	    RECT 262.1000 252.4000 262.7000 263.6000 ;
	    RECT 263.6000 261.6000 264.4000 262.4000 ;
	    RECT 263.7000 256.4000 264.3000 261.6000 ;
	    RECT 265.3000 258.4000 265.9000 275.6000 ;
	    RECT 268.4000 264.2000 269.2000 275.8000 ;
	    RECT 270.0000 269.6000 270.8000 270.4000 ;
	    RECT 266.8000 261.6000 267.6000 262.4000 ;
	    RECT 265.2000 257.6000 266.0000 258.4000 ;
	    RECT 266.9000 256.4000 267.5000 261.6000 ;
	    RECT 268.5000 257.7000 272.3000 258.3000 ;
	    RECT 263.6000 255.6000 264.4000 256.4000 ;
	    RECT 266.8000 255.6000 267.6000 256.4000 ;
	    RECT 268.5000 254.3000 269.1000 257.7000 ;
	    RECT 271.7000 256.4000 272.3000 257.7000 ;
	    RECT 270.0000 255.6000 270.8000 256.4000 ;
	    RECT 271.6000 255.6000 272.4000 256.4000 ;
	    RECT 266.9000 253.7000 269.1000 254.3000 ;
	    RECT 266.9000 252.4000 267.5000 253.7000 ;
	    RECT 260.4000 251.6000 261.2000 252.4000 ;
	    RECT 262.0000 251.6000 262.8000 252.4000 ;
	    RECT 266.8000 251.6000 267.6000 252.4000 ;
	    RECT 270.1000 250.4000 270.7000 255.6000 ;
	    RECT 271.6000 251.6000 272.4000 252.4000 ;
	    RECT 273.2000 251.6000 274.0000 252.4000 ;
	    RECT 266.8000 249.6000 267.6000 250.4000 ;
	    RECT 270.0000 249.6000 270.8000 250.4000 ;
	    RECT 257.2000 247.6000 258.0000 248.4000 ;
	    RECT 258.8000 247.6000 259.6000 248.4000 ;
	    RECT 265.2000 247.6000 266.0000 248.4000 ;
	    RECT 265.3000 244.4000 265.9000 247.6000 ;
	    RECT 265.2000 243.6000 266.0000 244.4000 ;
	    RECT 254.0000 233.6000 254.8000 234.4000 ;
	    RECT 254.0000 231.6000 254.8000 232.4000 ;
	    RECT 252.4000 229.6000 253.2000 230.4000 ;
	    RECT 254.1000 226.4000 254.7000 231.6000 ;
	    RECT 262.0000 229.6000 262.8000 230.4000 ;
	    RECT 265.2000 229.6000 266.0000 230.4000 ;
	    RECT 260.4000 227.6000 261.2000 228.4000 ;
	    RECT 254.0000 225.6000 254.8000 226.4000 ;
	    RECT 262.1000 222.4000 262.7000 229.6000 ;
	    RECT 263.6000 227.6000 264.4000 228.4000 ;
	    RECT 252.4000 221.6000 253.2000 222.4000 ;
	    RECT 262.0000 221.6000 262.8000 222.4000 ;
	    RECT 252.5000 218.3000 253.1000 221.6000 ;
	    RECT 252.5000 217.7000 254.7000 218.3000 ;
	    RECT 250.9000 215.7000 253.1000 216.3000 ;
	    RECT 249.3000 212.4000 249.9000 215.6000 ;
	    RECT 252.5000 214.4000 253.1000 215.7000 ;
	    RECT 252.4000 213.6000 253.2000 214.4000 ;
	    RECT 249.2000 211.6000 250.0000 212.4000 ;
	    RECT 252.4000 210.3000 253.2000 210.4000 ;
	    RECT 247.7000 209.7000 253.2000 210.3000 ;
	    RECT 252.4000 209.6000 253.2000 209.7000 ;
	    RECT 242.8000 208.3000 243.6000 208.4000 ;
	    RECT 241.3000 207.7000 243.6000 208.3000 ;
	    RECT 241.3000 198.4000 241.9000 207.7000 ;
	    RECT 242.8000 207.6000 243.6000 207.7000 ;
	    RECT 247.6000 207.6000 248.4000 208.4000 ;
	    RECT 249.2000 207.6000 250.0000 208.4000 ;
	    RECT 246.0000 203.6000 246.8000 204.4000 ;
	    RECT 241.2000 197.6000 242.0000 198.4000 ;
	    RECT 242.8000 197.6000 243.6000 198.4000 ;
	    RECT 238.0000 195.6000 238.8000 196.4000 ;
	    RECT 233.2000 189.6000 234.0000 190.4000 ;
	    RECT 234.8000 189.6000 235.6000 190.4000 ;
	    RECT 236.4000 189.6000 237.2000 190.4000 ;
	    RECT 231.6000 187.6000 232.4000 188.4000 ;
	    RECT 234.9000 184.4000 235.5000 189.6000 ;
	    RECT 233.2000 183.6000 234.0000 184.4000 ;
	    RECT 234.8000 183.6000 235.6000 184.4000 ;
	    RECT 236.5000 182.4000 237.1000 189.6000 ;
	    RECT 238.1000 186.4000 238.7000 195.6000 ;
	    RECT 239.6000 191.6000 240.4000 192.4000 ;
	    RECT 242.9000 190.4000 243.5000 197.6000 ;
	    RECT 241.2000 189.6000 242.0000 190.4000 ;
	    RECT 242.8000 189.6000 243.6000 190.4000 ;
	    RECT 244.4000 189.6000 245.2000 190.4000 ;
	    RECT 241.3000 188.3000 241.9000 189.6000 ;
	    RECT 246.1000 188.4000 246.7000 203.6000 ;
	    RECT 247.7000 200.4000 248.3000 207.6000 ;
	    RECT 247.6000 199.6000 248.4000 200.4000 ;
	    RECT 249.3000 192.4000 249.9000 207.6000 ;
	    RECT 250.8000 197.6000 251.6000 198.4000 ;
	    RECT 249.2000 191.6000 250.0000 192.4000 ;
	    RECT 249.2000 189.6000 250.0000 190.4000 ;
	    RECT 250.9000 188.4000 251.5000 197.6000 ;
	    RECT 252.4000 195.6000 253.2000 196.4000 ;
	    RECT 254.1000 194.3000 254.7000 217.7000 ;
	    RECT 257.3000 213.7000 261.1000 214.3000 ;
	    RECT 257.3000 210.4000 257.9000 213.7000 ;
	    RECT 260.5000 212.4000 261.1000 213.7000 ;
	    RECT 263.7000 212.4000 264.3000 227.6000 ;
	    RECT 265.3000 226.4000 265.9000 229.6000 ;
	    RECT 265.2000 225.6000 266.0000 226.4000 ;
	    RECT 265.2000 215.6000 266.0000 216.4000 ;
	    RECT 265.3000 212.4000 265.9000 215.6000 ;
	    RECT 266.9000 214.4000 267.5000 249.6000 ;
	    RECT 271.7000 248.3000 272.3000 251.6000 ;
	    RECT 273.3000 248.4000 273.9000 251.6000 ;
	    RECT 270.1000 247.7000 272.3000 248.3000 ;
	    RECT 268.4000 231.6000 269.2000 232.4000 ;
	    RECT 270.1000 230.3000 270.7000 247.7000 ;
	    RECT 273.2000 247.6000 274.0000 248.4000 ;
	    RECT 271.6000 243.6000 272.4000 244.4000 ;
	    RECT 271.7000 232.3000 272.3000 243.6000 ;
	    RECT 274.9000 232.4000 275.5000 327.6000 ;
	    RECT 276.5000 320.4000 277.1000 329.6000 ;
	    RECT 276.4000 319.6000 277.2000 320.4000 ;
	    RECT 279.7000 314.4000 280.3000 331.6000 ;
	    RECT 290.8000 323.6000 291.6000 324.4000 ;
	    RECT 279.6000 313.6000 280.4000 314.4000 ;
	    RECT 282.8000 313.6000 283.6000 314.4000 ;
	    RECT 279.7000 310.4000 280.3000 313.6000 ;
	    RECT 282.9000 310.4000 283.5000 313.6000 ;
	    RECT 290.9000 310.4000 291.5000 323.6000 ;
	    RECT 292.5000 314.3000 293.1000 337.6000 ;
	    RECT 294.0000 335.6000 294.8000 336.4000 ;
	    RECT 294.1000 332.4000 294.7000 335.6000 ;
	    RECT 303.6000 333.6000 304.4000 334.4000 ;
	    RECT 313.2000 333.6000 314.0000 334.4000 ;
	    RECT 303.7000 332.4000 304.3000 333.6000 ;
	    RECT 313.3000 332.4000 313.9000 333.6000 ;
	    RECT 294.0000 331.6000 294.8000 332.4000 ;
	    RECT 295.6000 331.6000 296.4000 332.4000 ;
	    RECT 297.2000 331.6000 298.0000 332.4000 ;
	    RECT 298.8000 331.6000 299.6000 332.4000 ;
	    RECT 303.6000 331.6000 304.4000 332.4000 ;
	    RECT 305.2000 331.6000 306.0000 332.4000 ;
	    RECT 308.4000 331.6000 309.2000 332.4000 ;
	    RECT 313.2000 331.6000 314.0000 332.4000 ;
	    RECT 297.3000 330.4000 297.9000 331.6000 ;
	    RECT 297.2000 329.6000 298.0000 330.4000 ;
	    RECT 298.9000 328.4000 299.5000 331.6000 ;
	    RECT 298.8000 327.6000 299.6000 328.4000 ;
	    RECT 300.4000 323.6000 301.2000 324.4000 ;
	    RECT 302.0000 323.6000 302.8000 324.4000 ;
	    RECT 292.5000 313.7000 294.7000 314.3000 ;
	    RECT 292.4000 311.6000 293.2000 312.4000 ;
	    RECT 276.4000 309.6000 277.2000 310.4000 ;
	    RECT 278.0000 309.6000 278.8000 310.4000 ;
	    RECT 279.6000 309.6000 280.4000 310.4000 ;
	    RECT 281.2000 309.6000 282.0000 310.4000 ;
	    RECT 282.8000 309.6000 283.6000 310.4000 ;
	    RECT 289.2000 309.6000 290.0000 310.4000 ;
	    RECT 290.8000 309.6000 291.6000 310.4000 ;
	    RECT 292.4000 309.6000 293.2000 310.4000 ;
	    RECT 276.5000 292.4000 277.1000 309.6000 ;
	    RECT 278.1000 308.4000 278.7000 309.6000 ;
	    RECT 278.0000 307.6000 278.8000 308.4000 ;
	    RECT 281.3000 308.3000 281.9000 309.6000 ;
	    RECT 282.9000 308.4000 283.5000 309.6000 ;
	    RECT 279.7000 307.7000 281.9000 308.3000 ;
	    RECT 279.7000 294.4000 280.3000 307.7000 ;
	    RECT 282.8000 307.6000 283.6000 308.4000 ;
	    RECT 287.6000 307.6000 288.4000 308.4000 ;
	    RECT 282.8000 295.6000 283.6000 296.4000 ;
	    RECT 282.9000 294.4000 283.5000 295.6000 ;
	    RECT 278.0000 293.6000 278.8000 294.4000 ;
	    RECT 279.6000 293.6000 280.4000 294.4000 ;
	    RECT 282.8000 293.6000 283.6000 294.4000 ;
	    RECT 286.0000 293.6000 286.8000 294.4000 ;
	    RECT 276.4000 291.6000 277.2000 292.4000 ;
	    RECT 278.1000 286.4000 278.7000 293.6000 ;
	    RECT 279.7000 292.4000 280.3000 293.6000 ;
	    RECT 279.6000 291.6000 280.4000 292.4000 ;
	    RECT 281.2000 292.3000 282.0000 292.4000 ;
	    RECT 281.2000 291.7000 283.5000 292.3000 ;
	    RECT 281.2000 291.6000 282.0000 291.7000 ;
	    RECT 281.3000 290.4000 281.9000 291.6000 ;
	    RECT 281.2000 289.6000 282.0000 290.4000 ;
	    RECT 278.0000 285.6000 278.8000 286.4000 ;
	    RECT 276.4000 273.6000 277.2000 274.4000 ;
	    RECT 276.5000 270.2000 277.1000 273.6000 ;
	    RECT 276.4000 269.4000 277.2000 270.2000 ;
	    RECT 278.0000 264.2000 278.8000 275.8000 ;
	    RECT 281.2000 266.2000 282.0000 271.8000 ;
	    RECT 282.9000 268.4000 283.5000 291.7000 ;
	    RECT 284.4000 289.6000 285.2000 290.4000 ;
	    RECT 284.5000 286.4000 285.1000 289.6000 ;
	    RECT 286.1000 286.4000 286.7000 293.6000 ;
	    RECT 287.7000 292.4000 288.3000 307.6000 ;
	    RECT 289.3000 302.4000 289.9000 309.6000 ;
	    RECT 292.5000 308.4000 293.1000 309.6000 ;
	    RECT 290.8000 307.6000 291.6000 308.4000 ;
	    RECT 292.4000 307.6000 293.2000 308.4000 ;
	    RECT 289.2000 301.6000 290.0000 302.4000 ;
	    RECT 290.9000 296.4000 291.5000 307.6000 ;
	    RECT 294.1000 296.4000 294.7000 313.7000 ;
	    RECT 300.5000 312.4000 301.1000 323.6000 ;
	    RECT 295.6000 311.6000 296.4000 312.4000 ;
	    RECT 300.4000 311.6000 301.2000 312.4000 ;
	    RECT 295.7000 310.4000 296.3000 311.6000 ;
	    RECT 295.6000 309.6000 296.4000 310.4000 ;
	    RECT 298.8000 309.6000 299.6000 310.4000 ;
	    RECT 297.2000 307.6000 298.0000 308.4000 ;
	    RECT 298.8000 307.6000 299.6000 308.4000 ;
	    RECT 290.8000 295.6000 291.6000 296.4000 ;
	    RECT 294.0000 295.6000 294.8000 296.4000 ;
	    RECT 297.3000 294.4000 297.9000 307.6000 ;
	    RECT 302.1000 306.4000 302.7000 323.6000 ;
	    RECT 303.6000 313.6000 304.4000 314.4000 ;
	    RECT 302.0000 305.6000 302.8000 306.4000 ;
	    RECT 302.0000 299.6000 302.8000 300.4000 ;
	    RECT 294.0000 294.3000 294.8000 294.4000 ;
	    RECT 294.0000 293.7000 296.3000 294.3000 ;
	    RECT 294.0000 293.6000 294.8000 293.7000 ;
	    RECT 287.6000 291.6000 288.4000 292.4000 ;
	    RECT 287.6000 287.6000 288.4000 288.4000 ;
	    RECT 295.7000 288.3000 296.3000 293.7000 ;
	    RECT 297.2000 293.6000 298.0000 294.4000 ;
	    RECT 302.1000 292.4000 302.7000 299.6000 ;
	    RECT 303.6000 294.3000 304.4000 294.4000 ;
	    RECT 305.3000 294.3000 305.9000 331.6000 ;
	    RECT 308.5000 328.4000 309.1000 331.6000 ;
	    RECT 308.4000 327.6000 309.2000 328.4000 ;
	    RECT 310.0000 323.6000 310.8000 324.4000 ;
	    RECT 311.6000 323.6000 312.4000 324.4000 ;
	    RECT 306.8000 305.6000 307.6000 306.4000 ;
	    RECT 306.9000 298.4000 307.5000 305.6000 ;
	    RECT 308.4000 304.2000 309.2000 315.8000 ;
	    RECT 310.1000 302.3000 310.7000 323.6000 ;
	    RECT 308.5000 301.7000 310.7000 302.3000 ;
	    RECT 306.8000 297.6000 307.6000 298.4000 ;
	    RECT 308.5000 296.4000 309.1000 301.7000 ;
	    RECT 308.4000 295.6000 309.2000 296.4000 ;
	    RECT 308.4000 294.3000 309.2000 294.4000 ;
	    RECT 303.6000 293.7000 305.9000 294.3000 ;
	    RECT 306.9000 293.7000 309.2000 294.3000 ;
	    RECT 303.6000 293.6000 304.4000 293.7000 ;
	    RECT 303.7000 292.4000 304.3000 293.6000 ;
	    RECT 297.2000 291.6000 298.0000 292.4000 ;
	    RECT 300.4000 291.6000 301.2000 292.4000 ;
	    RECT 302.0000 291.6000 302.8000 292.4000 ;
	    RECT 303.6000 291.6000 304.4000 292.4000 ;
	    RECT 305.2000 291.6000 306.0000 292.4000 ;
	    RECT 297.3000 290.4000 297.9000 291.6000 ;
	    RECT 297.2000 289.6000 298.0000 290.4000 ;
	    RECT 298.8000 289.6000 299.6000 290.4000 ;
	    RECT 295.7000 287.7000 297.9000 288.3000 ;
	    RECT 284.4000 285.6000 285.2000 286.4000 ;
	    RECT 286.0000 285.6000 286.8000 286.4000 ;
	    RECT 294.0000 285.6000 294.8000 286.4000 ;
	    RECT 284.4000 275.6000 285.2000 276.4000 ;
	    RECT 284.5000 272.4000 285.1000 275.6000 ;
	    RECT 290.8000 273.6000 291.6000 274.4000 ;
	    RECT 284.4000 271.6000 285.2000 272.4000 ;
	    RECT 286.0000 271.6000 286.8000 272.4000 ;
	    RECT 290.8000 271.6000 291.6000 272.4000 ;
	    RECT 292.4000 271.6000 293.2000 272.4000 ;
	    RECT 290.9000 270.4000 291.5000 271.6000 ;
	    RECT 286.0000 269.6000 286.8000 270.4000 ;
	    RECT 290.8000 269.6000 291.6000 270.4000 ;
	    RECT 282.8000 267.6000 283.6000 268.4000 ;
	    RECT 278.0000 246.2000 278.8000 257.8000 ;
	    RECT 286.1000 256.4000 286.7000 269.6000 ;
	    RECT 290.9000 268.4000 291.5000 269.6000 ;
	    RECT 292.5000 268.4000 293.1000 271.6000 ;
	    RECT 294.1000 268.4000 294.7000 285.6000 ;
	    RECT 297.3000 284.4000 297.9000 287.7000 ;
	    RECT 298.9000 286.4000 299.5000 289.6000 ;
	    RECT 298.8000 285.6000 299.6000 286.4000 ;
	    RECT 300.5000 284.4000 301.1000 291.6000 ;
	    RECT 305.3000 290.4000 305.9000 291.6000 ;
	    RECT 306.9000 290.4000 307.5000 293.7000 ;
	    RECT 308.4000 293.6000 309.2000 293.7000 ;
	    RECT 311.7000 292.4000 312.3000 323.6000 ;
	    RECT 313.3000 312.4000 313.9000 331.6000 ;
	    RECT 316.4000 327.6000 317.2000 328.4000 ;
	    RECT 321.2000 326.2000 322.0000 337.8000 ;
	    RECT 329.2000 331.8000 330.0000 332.6000 ;
	    RECT 313.2000 311.6000 314.0000 312.4000 ;
	    RECT 316.4000 309.4000 317.2000 310.4000 ;
	    RECT 313.2000 307.6000 314.0000 308.4000 ;
	    RECT 313.3000 294.4000 313.9000 307.6000 ;
	    RECT 314.8000 305.6000 315.6000 306.4000 ;
	    RECT 316.4000 305.6000 317.2000 306.4000 ;
	    RECT 313.2000 293.6000 314.0000 294.4000 ;
	    RECT 314.9000 292.4000 315.5000 305.6000 ;
	    RECT 311.6000 291.6000 312.4000 292.4000 ;
	    RECT 314.8000 291.6000 315.6000 292.4000 ;
	    RECT 305.2000 289.6000 306.0000 290.4000 ;
	    RECT 306.8000 289.6000 307.6000 290.4000 ;
	    RECT 316.5000 290.3000 317.1000 305.6000 ;
	    RECT 318.0000 304.2000 318.8000 315.8000 ;
	    RECT 329.3000 314.4000 329.9000 331.8000 ;
	    RECT 330.8000 326.2000 331.6000 337.8000 ;
	    RECT 346.8000 337.6000 347.6000 338.4000 ;
	    RECT 346.9000 336.4000 347.5000 337.6000 ;
	    RECT 332.4000 333.6000 333.2000 334.4000 ;
	    RECT 334.0000 330.2000 334.8000 335.8000 ;
	    RECT 335.6000 335.6000 336.4000 336.4000 ;
	    RECT 346.8000 335.6000 347.6000 336.4000 ;
	    RECT 335.7000 334.4000 336.3000 335.6000 ;
	    RECT 335.6000 333.6000 336.4000 334.4000 ;
	    RECT 345.2000 333.6000 346.0000 334.4000 ;
	    RECT 345.3000 332.4000 345.9000 333.6000 ;
	    RECT 338.8000 331.6000 339.6000 332.4000 ;
	    RECT 343.6000 331.6000 344.4000 332.4000 ;
	    RECT 345.2000 331.6000 346.0000 332.4000 ;
	    RECT 338.9000 330.4000 339.5000 331.6000 ;
	    RECT 338.8000 329.6000 339.6000 330.4000 ;
	    RECT 334.0000 327.6000 334.8000 328.4000 ;
	    RECT 332.4000 317.6000 333.2000 318.4000 ;
	    RECT 322.8000 313.6000 323.6000 314.4000 ;
	    RECT 329.2000 313.6000 330.0000 314.4000 ;
	    RECT 321.2000 306.2000 322.0000 311.8000 ;
	    RECT 322.9000 308.4000 323.5000 313.6000 ;
	    RECT 326.0000 311.6000 326.8000 312.4000 ;
	    RECT 326.1000 310.4000 326.7000 311.6000 ;
	    RECT 326.0000 309.6000 326.8000 310.4000 ;
	    RECT 330.8000 309.6000 331.6000 310.4000 ;
	    RECT 322.8000 307.6000 323.6000 308.4000 ;
	    RECT 327.6000 307.6000 328.4000 308.4000 ;
	    RECT 327.6000 303.6000 328.4000 304.4000 ;
	    RECT 321.2000 295.6000 322.0000 296.4000 ;
	    RECT 321.3000 292.4000 321.9000 295.6000 ;
	    RECT 322.8000 293.6000 323.6000 294.4000 ;
	    RECT 324.4000 293.6000 325.2000 294.4000 ;
	    RECT 322.9000 292.4000 323.5000 293.6000 ;
	    RECT 321.2000 291.6000 322.0000 292.4000 ;
	    RECT 322.8000 291.6000 323.6000 292.4000 ;
	    RECT 324.5000 290.4000 325.1000 293.6000 ;
	    RECT 327.7000 292.4000 328.3000 303.6000 ;
	    RECT 329.2000 295.6000 330.0000 296.4000 ;
	    RECT 329.3000 294.4000 329.9000 295.6000 ;
	    RECT 329.2000 293.6000 330.0000 294.4000 ;
	    RECT 327.6000 291.6000 328.4000 292.4000 ;
	    RECT 329.2000 291.6000 330.0000 292.4000 ;
	    RECT 314.9000 289.7000 317.1000 290.3000 ;
	    RECT 295.6000 283.6000 296.4000 284.4000 ;
	    RECT 297.2000 283.6000 298.0000 284.4000 ;
	    RECT 300.4000 283.6000 301.2000 284.4000 ;
	    RECT 302.0000 283.6000 302.8000 284.4000 ;
	    RECT 295.7000 278.4000 296.3000 283.6000 ;
	    RECT 295.6000 277.6000 296.4000 278.4000 ;
	    RECT 302.1000 274.4000 302.7000 283.6000 ;
	    RECT 305.3000 274.4000 305.9000 289.6000 ;
	    RECT 306.9000 286.4000 307.5000 289.6000 ;
	    RECT 306.8000 285.6000 307.6000 286.4000 ;
	    RECT 298.8000 273.6000 299.6000 274.4000 ;
	    RECT 302.0000 273.6000 302.8000 274.4000 ;
	    RECT 305.2000 273.6000 306.0000 274.4000 ;
	    RECT 295.6000 271.6000 296.4000 272.4000 ;
	    RECT 295.7000 270.4000 296.3000 271.6000 ;
	    RECT 298.9000 270.4000 299.5000 273.6000 ;
	    RECT 306.9000 272.4000 307.5000 285.6000 ;
	    RECT 310.0000 283.6000 310.8000 284.4000 ;
	    RECT 313.2000 283.6000 314.0000 284.4000 ;
	    RECT 310.1000 278.4000 310.7000 283.6000 ;
	    RECT 308.4000 277.6000 309.2000 278.4000 ;
	    RECT 310.0000 277.6000 310.8000 278.4000 ;
	    RECT 311.6000 277.6000 312.4000 278.4000 ;
	    RECT 308.5000 276.3000 309.1000 277.6000 ;
	    RECT 308.5000 275.7000 310.7000 276.3000 ;
	    RECT 310.1000 274.4000 310.7000 275.7000 ;
	    RECT 308.4000 273.6000 309.2000 274.4000 ;
	    RECT 310.0000 273.6000 310.8000 274.4000 ;
	    RECT 303.6000 272.3000 304.4000 272.4000 ;
	    RECT 302.1000 271.7000 304.4000 272.3000 ;
	    RECT 302.1000 270.4000 302.7000 271.7000 ;
	    RECT 303.6000 271.6000 304.4000 271.7000 ;
	    RECT 306.8000 271.6000 307.6000 272.4000 ;
	    RECT 295.6000 269.6000 296.4000 270.4000 ;
	    RECT 298.8000 269.6000 299.6000 270.4000 ;
	    RECT 302.0000 269.6000 302.8000 270.4000 ;
	    RECT 303.6000 270.3000 304.4000 270.4000 ;
	    RECT 303.6000 269.7000 305.9000 270.3000 ;
	    RECT 303.6000 269.6000 304.4000 269.7000 ;
	    RECT 290.8000 267.6000 291.6000 268.4000 ;
	    RECT 292.4000 267.6000 293.2000 268.4000 ;
	    RECT 294.0000 267.6000 294.8000 268.4000 ;
	    RECT 300.4000 267.6000 301.2000 268.4000 ;
	    RECT 302.0000 267.6000 302.8000 268.4000 ;
	    RECT 297.2000 263.6000 298.0000 264.4000 ;
	    RECT 286.0000 255.6000 286.8000 256.4000 ;
	    RECT 279.6000 251.6000 280.4000 252.4000 ;
	    RECT 286.0000 251.8000 286.8000 252.6000 ;
	    RECT 271.7000 231.7000 273.9000 232.3000 ;
	    RECT 268.5000 229.7000 270.7000 230.3000 ;
	    RECT 266.8000 213.6000 267.6000 214.4000 ;
	    RECT 258.8000 211.6000 259.6000 212.4000 ;
	    RECT 260.4000 211.6000 261.2000 212.4000 ;
	    RECT 263.6000 211.6000 264.4000 212.4000 ;
	    RECT 265.2000 211.6000 266.0000 212.4000 ;
	    RECT 266.8000 211.6000 267.6000 212.4000 ;
	    RECT 257.2000 209.6000 258.0000 210.4000 ;
	    RECT 255.6000 199.6000 256.4000 200.4000 ;
	    RECT 252.5000 193.7000 254.7000 194.3000 ;
	    RECT 241.3000 187.7000 243.5000 188.3000 ;
	    RECT 238.0000 185.6000 238.8000 186.4000 ;
	    RECT 220.4000 181.6000 221.2000 182.4000 ;
	    RECT 223.6000 181.6000 224.4000 182.4000 ;
	    RECT 230.0000 181.6000 230.8000 182.4000 ;
	    RECT 234.8000 181.6000 235.6000 182.4000 ;
	    RECT 236.4000 181.6000 237.2000 182.4000 ;
	    RECT 242.9000 182.3000 243.5000 187.7000 ;
	    RECT 244.4000 187.6000 245.2000 188.4000 ;
	    RECT 246.0000 187.6000 246.8000 188.4000 ;
	    RECT 247.6000 187.6000 248.4000 188.4000 ;
	    RECT 249.2000 187.6000 250.0000 188.4000 ;
	    RECT 250.8000 187.6000 251.6000 188.4000 ;
	    RECT 244.5000 184.4000 245.1000 187.6000 ;
	    RECT 244.4000 183.6000 245.2000 184.4000 ;
	    RECT 242.9000 181.7000 245.1000 182.3000 ;
	    RECT 217.2000 179.6000 218.0000 180.4000 ;
	    RECT 225.2000 177.6000 226.0000 178.4000 ;
	    RECT 228.4000 177.6000 229.2000 178.4000 ;
	    RECT 223.6000 173.6000 224.4000 174.4000 ;
	    RECT 215.6000 171.6000 216.4000 172.4000 ;
	    RECT 217.2000 171.6000 218.0000 172.4000 ;
	    RECT 222.0000 171.6000 222.8000 172.4000 ;
	    RECT 217.3000 170.4000 217.9000 171.6000 ;
	    RECT 217.2000 169.6000 218.0000 170.4000 ;
	    RECT 206.0000 165.6000 206.8000 166.4000 ;
	    RECT 210.8000 163.6000 211.6000 164.4000 ;
	    RECT 204.4000 155.6000 205.2000 156.4000 ;
	    RECT 204.5000 134.4000 205.1000 155.6000 ;
	    RECT 206.0000 144.2000 206.8000 155.8000 ;
	    RECT 207.6000 145.6000 208.4000 146.4000 ;
	    RECT 206.0000 137.6000 206.8000 138.4000 ;
	    RECT 206.1000 134.4000 206.7000 137.6000 ;
	    RECT 204.4000 133.6000 205.2000 134.4000 ;
	    RECT 206.0000 133.6000 206.8000 134.4000 ;
	    RECT 207.7000 132.4000 208.3000 145.6000 ;
	    RECT 207.6000 131.6000 208.4000 132.4000 ;
	    RECT 210.9000 130.3000 211.5000 163.6000 ;
	    RECT 217.3000 160.4000 217.9000 169.6000 ;
	    RECT 222.0000 163.6000 222.8000 164.4000 ;
	    RECT 223.7000 162.3000 224.3000 173.6000 ;
	    RECT 225.2000 165.6000 226.0000 166.4000 ;
	    RECT 222.1000 161.7000 224.3000 162.3000 ;
	    RECT 217.2000 159.6000 218.0000 160.4000 ;
	    RECT 212.4000 157.6000 213.2000 158.4000 ;
	    RECT 217.2000 157.6000 218.0000 158.4000 ;
	    RECT 212.5000 150.4000 213.1000 157.6000 ;
	    RECT 212.4000 149.6000 213.2000 150.4000 ;
	    RECT 215.6000 144.2000 216.4000 155.8000 ;
	    RECT 217.3000 148.4000 217.9000 157.6000 ;
	    RECT 222.1000 154.4000 222.7000 161.7000 ;
	    RECT 223.6000 159.6000 224.4000 160.4000 ;
	    RECT 223.7000 158.4000 224.3000 159.6000 ;
	    RECT 223.6000 157.6000 224.4000 158.4000 ;
	    RECT 222.0000 153.6000 222.8000 154.4000 ;
	    RECT 223.7000 152.4000 224.3000 157.6000 ;
	    RECT 225.3000 152.4000 225.9000 165.6000 ;
	    RECT 217.2000 147.6000 218.0000 148.4000 ;
	    RECT 218.8000 146.2000 219.6000 151.8000 ;
	    RECT 223.6000 151.6000 224.4000 152.4000 ;
	    RECT 225.2000 151.6000 226.0000 152.4000 ;
	    RECT 228.5000 150.4000 229.1000 177.6000 ;
	    RECT 230.0000 166.2000 230.8000 177.8000 ;
	    RECT 234.9000 174.3000 235.5000 181.6000 ;
	    RECT 234.9000 173.7000 237.1000 174.3000 ;
	    RECT 234.8000 171.6000 235.6000 172.4000 ;
	    RECT 234.9000 164.4000 235.5000 171.6000 ;
	    RECT 234.8000 163.6000 235.6000 164.4000 ;
	    RECT 231.6000 157.6000 232.4000 158.4000 ;
	    RECT 228.4000 149.6000 229.2000 150.4000 ;
	    RECT 225.2000 145.6000 226.0000 146.4000 ;
	    RECT 228.4000 145.6000 229.2000 146.4000 ;
	    RECT 225.3000 138.3000 225.9000 145.6000 ;
	    RECT 226.8000 143.6000 227.6000 144.4000 ;
	    RECT 226.9000 140.4000 227.5000 143.6000 ;
	    RECT 226.8000 139.6000 227.6000 140.4000 ;
	    RECT 228.5000 138.4000 229.1000 145.6000 ;
	    RECT 218.8000 135.6000 219.6000 136.4000 ;
	    RECT 217.2000 134.3000 218.0000 134.4000 ;
	    RECT 209.3000 129.7000 211.5000 130.3000 ;
	    RECT 214.1000 133.7000 218.0000 134.3000 ;
	    RECT 204.4000 127.6000 205.2000 128.4000 ;
	    RECT 204.5000 126.3000 205.1000 127.6000 ;
	    RECT 209.3000 126.4000 209.9000 129.7000 ;
	    RECT 210.8000 127.6000 211.6000 128.4000 ;
	    RECT 204.5000 125.7000 206.7000 126.3000 ;
	    RECT 201.2000 123.6000 202.0000 124.4000 ;
	    RECT 202.8000 123.6000 203.6000 124.4000 ;
	    RECT 204.4000 123.6000 205.2000 124.4000 ;
	    RECT 191.6000 109.6000 192.4000 110.4000 ;
	    RECT 194.8000 109.6000 195.6000 110.4000 ;
	    RECT 196.4000 109.6000 197.2000 110.4000 ;
	    RECT 190.0000 107.6000 190.8000 108.4000 ;
	    RECT 188.4000 105.6000 189.2000 106.4000 ;
	    RECT 190.0000 103.6000 190.8000 104.4000 ;
	    RECT 198.0000 104.2000 198.8000 115.8000 ;
	    RECT 201.3000 112.4000 201.9000 123.6000 ;
	    RECT 201.2000 111.6000 202.0000 112.4000 ;
	    RECT 204.5000 110.4000 205.1000 123.6000 ;
	    RECT 206.1000 114.4000 206.7000 125.7000 ;
	    RECT 209.2000 125.6000 210.0000 126.4000 ;
	    RECT 206.0000 113.6000 206.8000 114.4000 ;
	    RECT 204.4000 109.6000 205.2000 110.4000 ;
	    RECT 202.8000 107.6000 203.6000 108.4000 ;
	    RECT 182.1000 95.7000 184.3000 96.3000 ;
	    RECT 183.7000 94.4000 184.3000 95.7000 ;
	    RECT 185.3000 95.7000 187.5000 96.3000 ;
	    RECT 185.3000 94.4000 185.9000 95.7000 ;
	    RECT 182.0000 93.6000 182.8000 94.4000 ;
	    RECT 183.6000 93.6000 184.4000 94.4000 ;
	    RECT 185.2000 93.6000 186.0000 94.4000 ;
	    RECT 186.8000 93.6000 187.6000 94.4000 ;
	    RECT 182.1000 92.4000 182.7000 93.6000 ;
	    RECT 185.3000 92.4000 185.9000 93.6000 ;
	    RECT 186.9000 92.4000 187.5000 93.6000 ;
	    RECT 190.1000 92.4000 190.7000 103.6000 ;
	    RECT 196.4000 101.6000 197.2000 102.4000 ;
	    RECT 202.9000 102.3000 203.5000 107.6000 ;
	    RECT 201.3000 101.7000 203.5000 102.3000 ;
	    RECT 194.8000 95.6000 195.6000 96.4000 ;
	    RECT 194.9000 92.4000 195.5000 95.6000 ;
	    RECT 196.5000 92.4000 197.1000 101.6000 ;
	    RECT 198.0000 95.6000 198.8000 96.4000 ;
	    RECT 198.1000 94.4000 198.7000 95.6000 ;
	    RECT 198.0000 93.6000 198.8000 94.4000 ;
	    RECT 182.0000 91.6000 182.8000 92.4000 ;
	    RECT 185.2000 91.6000 186.0000 92.4000 ;
	    RECT 186.8000 91.6000 187.6000 92.4000 ;
	    RECT 190.0000 91.6000 190.8000 92.4000 ;
	    RECT 193.2000 91.6000 194.0000 92.4000 ;
	    RECT 194.8000 91.6000 195.6000 92.4000 ;
	    RECT 196.4000 91.6000 197.2000 92.4000 ;
	    RECT 193.3000 90.4000 193.9000 91.6000 ;
	    RECT 186.8000 89.6000 187.6000 90.4000 ;
	    RECT 193.2000 89.6000 194.0000 90.4000 ;
	    RECT 199.6000 89.6000 200.4000 90.4000 ;
	    RECT 182.0000 70.3000 182.8000 70.4000 ;
	    RECT 180.5000 69.7000 182.8000 70.3000 ;
	    RECT 182.0000 69.6000 182.8000 69.7000 ;
	    RECT 183.6000 67.6000 184.4000 68.4000 ;
	    RECT 183.7000 66.4000 184.3000 67.6000 ;
	    RECT 183.6000 65.6000 184.4000 66.4000 ;
	    RECT 188.4000 65.6000 189.2000 66.4000 ;
	    RECT 178.8000 63.6000 179.6000 64.4000 ;
	    RECT 177.2000 61.6000 178.0000 62.4000 ;
	    RECT 174.0000 59.6000 174.8000 60.4000 ;
	    RECT 172.4000 57.6000 173.2000 58.4000 ;
	    RECT 178.9000 54.4000 179.5000 63.6000 ;
	    RECT 172.4000 54.3000 173.2000 54.4000 ;
	    RECT 170.9000 53.7000 173.2000 54.3000 ;
	    RECT 172.4000 53.6000 173.2000 53.7000 ;
	    RECT 178.8000 53.6000 179.6000 54.4000 ;
	    RECT 183.7000 54.3000 184.3000 65.6000 ;
	    RECT 185.2000 63.6000 186.0000 64.4000 ;
	    RECT 185.3000 56.4000 185.9000 63.6000 ;
	    RECT 185.2000 55.6000 186.0000 56.4000 ;
	    RECT 185.2000 54.3000 186.0000 54.4000 ;
	    RECT 183.7000 53.7000 186.0000 54.3000 ;
	    RECT 185.2000 53.6000 186.0000 53.7000 ;
	    RECT 186.8000 53.6000 187.6000 54.4000 ;
	    RECT 161.3000 52.4000 161.9000 53.6000 ;
	    RECT 159.6000 51.6000 160.4000 52.4000 ;
	    RECT 161.2000 51.6000 162.0000 52.4000 ;
	    RECT 154.8000 49.6000 155.6000 50.4000 ;
	    RECT 154.9000 46.4000 155.5000 49.6000 ;
	    RECT 158.0000 47.6000 158.8000 48.4000 ;
	    RECT 154.8000 45.6000 155.6000 46.4000 ;
	    RECT 151.6000 29.4000 152.4000 30.2000 ;
	    RECT 153.2000 24.2000 154.0000 35.8000 ;
	    RECT 154.8000 27.6000 155.6000 28.4000 ;
	    RECT 138.8000 23.6000 139.6000 23.7000 ;
	    RECT 135.6000 17.6000 136.4000 18.4000 ;
	    RECT 137.2000 17.6000 138.0000 18.4000 ;
	    RECT 130.8000 13.6000 131.6000 14.4000 ;
	    RECT 135.7000 12.4000 136.3000 17.6000 ;
	    RECT 140.5000 12.4000 141.1000 23.7000 ;
	    RECT 142.0000 17.6000 142.8000 18.4000 ;
	    RECT 124.4000 11.6000 125.2000 12.4000 ;
	    RECT 129.2000 11.6000 130.0000 12.4000 ;
	    RECT 135.6000 11.6000 136.4000 12.4000 ;
	    RECT 140.4000 11.6000 141.2000 12.4000 ;
	    RECT 113.2000 9.6000 114.0000 10.4000 ;
	    RECT 119.6000 9.6000 120.4000 10.4000 ;
	    RECT 100.4000 7.7000 102.7000 8.3000 ;
	    RECT 100.4000 7.6000 101.2000 7.7000 ;
	    RECT 124.5000 4.4000 125.1000 11.6000 ;
	    RECT 126.0000 9.6000 126.8000 10.4000 ;
	    RECT 146.8000 6.2000 147.6000 17.8000 ;
	    RECT 154.9000 16.4000 155.5000 27.6000 ;
	    RECT 156.4000 26.2000 157.2000 31.8000 ;
	    RECT 158.0000 31.6000 158.8000 32.4000 ;
	    RECT 158.1000 26.4000 158.7000 31.6000 ;
	    RECT 158.0000 25.6000 158.8000 26.4000 ;
	    RECT 159.7000 24.4000 160.3000 51.6000 ;
	    RECT 161.2000 49.6000 162.0000 50.4000 ;
	    RECT 161.3000 38.4000 161.9000 49.6000 ;
	    RECT 161.2000 37.6000 162.0000 38.4000 ;
	    RECT 161.2000 31.6000 162.0000 32.4000 ;
	    RECT 161.3000 30.4000 161.9000 31.6000 ;
	    RECT 162.9000 30.4000 163.5000 53.6000 ;
	    RECT 188.5000 52.4000 189.1000 65.6000 ;
	    RECT 190.0000 64.2000 190.8000 75.8000 ;
	    RECT 196.4000 71.6000 197.2000 72.4000 ;
	    RECT 196.5000 64.4000 197.1000 71.6000 ;
	    RECT 198.0000 69.4000 198.8000 70.4000 ;
	    RECT 196.4000 63.6000 197.2000 64.4000 ;
	    RECT 199.6000 64.2000 200.4000 75.8000 ;
	    RECT 201.3000 68.4000 201.9000 101.7000 ;
	    RECT 204.5000 94.4000 205.1000 109.6000 ;
	    RECT 206.0000 109.4000 206.8000 110.4000 ;
	    RECT 207.6000 104.2000 208.4000 115.8000 ;
	    RECT 209.3000 104.4000 209.9000 125.6000 ;
	    RECT 210.9000 120.4000 211.5000 127.6000 ;
	    RECT 210.8000 119.6000 211.6000 120.4000 ;
	    RECT 214.1000 114.4000 214.7000 133.7000 ;
	    RECT 217.2000 133.6000 218.0000 133.7000 ;
	    RECT 218.9000 132.4000 219.5000 135.6000 ;
	    RECT 215.6000 132.3000 216.4000 132.4000 ;
	    RECT 215.6000 131.7000 217.9000 132.3000 ;
	    RECT 215.6000 131.6000 216.4000 131.7000 ;
	    RECT 215.6000 125.6000 216.4000 126.4000 ;
	    RECT 214.0000 113.6000 214.8000 114.4000 ;
	    RECT 210.8000 106.2000 211.6000 111.8000 ;
	    RECT 212.4000 111.6000 213.2000 112.4000 ;
	    RECT 215.6000 111.6000 216.4000 112.4000 ;
	    RECT 212.4000 109.6000 213.2000 110.4000 ;
	    RECT 209.2000 103.6000 210.0000 104.4000 ;
	    RECT 214.0000 103.6000 214.8000 104.4000 ;
	    RECT 206.0000 101.6000 206.8000 102.4000 ;
	    RECT 204.4000 93.6000 205.2000 94.4000 ;
	    RECT 206.1000 92.4000 206.7000 101.6000 ;
	    RECT 210.8000 97.6000 211.6000 98.4000 ;
	    RECT 209.2000 95.6000 210.0000 96.4000 ;
	    RECT 209.3000 94.4000 209.9000 95.6000 ;
	    RECT 209.2000 93.6000 210.0000 94.4000 ;
	    RECT 202.8000 91.6000 203.6000 92.4000 ;
	    RECT 206.0000 91.6000 206.8000 92.4000 ;
	    RECT 207.6000 91.6000 208.4000 92.4000 ;
	    RECT 202.8000 83.6000 203.6000 84.4000 ;
	    RECT 202.9000 74.3000 203.5000 83.6000 ;
	    RECT 209.2000 79.6000 210.0000 80.4000 ;
	    RECT 202.9000 73.7000 205.1000 74.3000 ;
	    RECT 204.5000 72.4000 205.1000 73.7000 ;
	    RECT 201.2000 67.6000 202.0000 68.4000 ;
	    RECT 199.6000 61.6000 200.4000 62.4000 ;
	    RECT 190.0000 55.6000 190.8000 56.4000 ;
	    RECT 198.0000 55.6000 198.8000 56.4000 ;
	    RECT 170.8000 51.6000 171.6000 52.4000 ;
	    RECT 172.4000 51.6000 173.2000 52.4000 ;
	    RECT 185.2000 51.6000 186.0000 52.4000 ;
	    RECT 186.8000 51.6000 187.6000 52.4000 ;
	    RECT 188.4000 51.6000 189.2000 52.4000 ;
	    RECT 166.0000 49.6000 166.8000 50.4000 ;
	    RECT 167.6000 49.6000 168.4000 50.4000 ;
	    RECT 166.1000 38.4000 166.7000 49.6000 ;
	    RECT 167.7000 46.4000 168.3000 49.6000 ;
	    RECT 167.6000 45.6000 168.4000 46.4000 ;
	    RECT 172.5000 40.4000 173.1000 51.6000 ;
	    RECT 174.0000 49.6000 174.8000 50.4000 ;
	    RECT 180.4000 49.6000 181.2000 50.4000 ;
	    RECT 174.1000 44.4000 174.7000 49.6000 ;
	    RECT 180.5000 46.4000 181.1000 49.6000 ;
	    RECT 180.4000 45.6000 181.2000 46.4000 ;
	    RECT 174.0000 43.6000 174.8000 44.4000 ;
	    RECT 172.4000 39.6000 173.2000 40.4000 ;
	    RECT 177.2000 39.6000 178.0000 40.4000 ;
	    RECT 166.0000 37.6000 166.8000 38.4000 ;
	    RECT 169.2000 31.6000 170.0000 32.4000 ;
	    RECT 161.2000 29.6000 162.0000 30.4000 ;
	    RECT 162.8000 29.6000 163.6000 30.4000 ;
	    RECT 162.9000 28.4000 163.5000 29.6000 ;
	    RECT 162.8000 27.6000 163.6000 28.4000 ;
	    RECT 159.6000 23.6000 160.4000 24.4000 ;
	    RECT 169.3000 18.4000 169.9000 31.6000 ;
	    RECT 170.8000 26.2000 171.6000 31.8000 ;
	    RECT 172.4000 27.6000 173.2000 28.4000 ;
	    RECT 154.8000 15.6000 155.6000 16.4000 ;
	    RECT 154.8000 13.6000 155.6000 14.4000 ;
	    RECT 154.9000 12.6000 155.5000 13.6000 ;
	    RECT 154.8000 11.8000 155.6000 12.6000 ;
	    RECT 154.9000 11.7000 155.5000 11.8000 ;
	    RECT 156.4000 6.2000 157.2000 17.8000 ;
	    RECT 166.0000 17.6000 166.8000 18.4000 ;
	    RECT 169.2000 17.6000 170.0000 18.4000 ;
	    RECT 159.6000 10.2000 160.4000 15.8000 ;
	    RECT 170.8000 6.2000 171.6000 17.8000 ;
	    RECT 172.5000 12.4000 173.1000 27.6000 ;
	    RECT 174.0000 24.2000 174.8000 35.8000 ;
	    RECT 177.3000 30.4000 177.9000 39.6000 ;
	    RECT 177.2000 29.6000 178.0000 30.4000 ;
	    RECT 183.6000 24.2000 184.4000 35.8000 ;
	    RECT 185.3000 34.4000 185.9000 51.6000 ;
	    RECT 185.2000 33.6000 186.0000 34.4000 ;
	    RECT 186.9000 32.4000 187.5000 51.6000 ;
	    RECT 188.4000 37.6000 189.2000 38.4000 ;
	    RECT 186.8000 31.6000 187.6000 32.4000 ;
	    RECT 190.1000 32.3000 190.7000 55.6000 ;
	    RECT 198.1000 54.4000 198.7000 55.6000 ;
	    RECT 191.6000 53.6000 192.4000 54.4000 ;
	    RECT 196.4000 53.6000 197.2000 54.4000 ;
	    RECT 198.0000 53.6000 198.8000 54.4000 ;
	    RECT 191.7000 52.4000 192.3000 53.6000 ;
	    RECT 196.5000 52.4000 197.1000 53.6000 ;
	    RECT 191.6000 51.6000 192.4000 52.4000 ;
	    RECT 194.8000 51.6000 195.6000 52.4000 ;
	    RECT 196.4000 51.6000 197.2000 52.4000 ;
	    RECT 193.2000 49.6000 194.0000 50.4000 ;
	    RECT 191.6000 47.6000 192.4000 48.4000 ;
	    RECT 191.7000 38.4000 192.3000 47.6000 ;
	    RECT 191.6000 37.6000 192.4000 38.4000 ;
	    RECT 191.6000 32.3000 192.4000 32.4000 ;
	    RECT 190.1000 31.7000 192.4000 32.3000 ;
	    RECT 191.6000 31.6000 192.4000 31.7000 ;
	    RECT 191.7000 30.4000 192.3000 31.6000 ;
	    RECT 194.9000 30.4000 195.5000 51.6000 ;
	    RECT 199.7000 50.4000 200.3000 61.6000 ;
	    RECT 199.6000 49.6000 200.4000 50.4000 ;
	    RECT 201.3000 46.3000 201.9000 67.6000 ;
	    RECT 202.8000 66.2000 203.6000 71.8000 ;
	    RECT 204.4000 71.6000 205.2000 72.4000 ;
	    RECT 206.0000 69.6000 206.8000 70.4000 ;
	    RECT 207.6000 69.6000 208.4000 70.4000 ;
	    RECT 209.3000 68.4000 209.9000 79.6000 ;
	    RECT 210.9000 72.4000 211.5000 97.6000 ;
	    RECT 214.1000 96.4000 214.7000 103.6000 ;
	    RECT 215.7000 102.4000 216.3000 111.6000 ;
	    RECT 217.3000 110.4000 217.9000 131.7000 ;
	    RECT 218.8000 131.6000 219.6000 132.4000 ;
	    RECT 223.6000 126.2000 224.4000 137.8000 ;
	    RECT 225.3000 137.7000 227.5000 138.3000 ;
	    RECT 218.8000 123.6000 219.6000 124.4000 ;
	    RECT 218.9000 120.4000 219.5000 123.6000 ;
	    RECT 218.8000 119.6000 219.6000 120.4000 ;
	    RECT 217.2000 109.6000 218.0000 110.4000 ;
	    RECT 222.0000 109.6000 222.8000 110.4000 ;
	    RECT 217.2000 107.6000 218.0000 108.4000 ;
	    RECT 218.8000 107.6000 219.6000 108.4000 ;
	    RECT 215.6000 101.6000 216.4000 102.4000 ;
	    RECT 214.0000 95.6000 214.8000 96.4000 ;
	    RECT 215.6000 93.6000 216.4000 94.4000 ;
	    RECT 215.7000 92.4000 216.3000 93.6000 ;
	    RECT 215.6000 91.6000 216.4000 92.4000 ;
	    RECT 217.3000 80.4000 217.9000 107.6000 ;
	    RECT 218.9000 106.4000 219.5000 107.6000 ;
	    RECT 218.8000 105.6000 219.6000 106.4000 ;
	    RECT 220.4000 103.6000 221.2000 104.4000 ;
	    RECT 218.8000 89.6000 219.6000 90.4000 ;
	    RECT 220.5000 84.4000 221.1000 103.6000 ;
	    RECT 222.1000 96.4000 222.7000 109.6000 ;
	    RECT 223.6000 107.6000 224.4000 108.4000 ;
	    RECT 223.7000 106.4000 224.3000 107.6000 ;
	    RECT 226.9000 106.4000 227.5000 137.7000 ;
	    RECT 228.4000 137.6000 229.2000 138.4000 ;
	    RECT 231.7000 136.4000 232.3000 157.6000 ;
	    RECT 233.2000 153.6000 234.0000 154.4000 ;
	    RECT 233.3000 152.4000 233.9000 153.6000 ;
	    RECT 233.2000 151.6000 234.0000 152.4000 ;
	    RECT 234.8000 146.2000 235.6000 151.8000 ;
	    RECT 236.5000 138.3000 237.1000 173.7000 ;
	    RECT 239.6000 166.2000 240.4000 177.8000 ;
	    RECT 241.2000 173.6000 242.0000 174.4000 ;
	    RECT 239.6000 163.6000 240.4000 164.4000 ;
	    RECT 239.7000 160.4000 240.3000 163.6000 ;
	    RECT 239.6000 159.6000 240.4000 160.4000 ;
	    RECT 241.3000 158.4000 241.9000 173.6000 ;
	    RECT 242.8000 170.2000 243.6000 175.8000 ;
	    RECT 244.5000 174.4000 245.1000 181.7000 ;
	    RECT 247.7000 178.4000 248.3000 187.6000 ;
	    RECT 249.3000 180.4000 249.9000 187.6000 ;
	    RECT 249.2000 179.6000 250.0000 180.4000 ;
	    RECT 246.0000 177.6000 246.8000 178.4000 ;
	    RECT 247.6000 177.6000 248.4000 178.4000 ;
	    RECT 250.8000 177.6000 251.6000 178.4000 ;
	    RECT 252.5000 178.3000 253.1000 193.7000 ;
	    RECT 255.7000 190.4000 256.3000 199.6000 ;
	    RECT 255.6000 189.6000 256.4000 190.4000 ;
	    RECT 258.9000 184.4000 259.5000 211.6000 ;
	    RECT 266.9000 210.3000 267.5000 211.6000 ;
	    RECT 265.3000 209.7000 267.5000 210.3000 ;
	    RECT 263.6000 203.6000 264.4000 204.4000 ;
	    RECT 263.7000 200.4000 264.3000 203.6000 ;
	    RECT 263.6000 199.6000 264.4000 200.4000 ;
	    RECT 263.6000 192.3000 264.4000 192.4000 ;
	    RECT 262.1000 191.7000 264.4000 192.3000 ;
	    RECT 258.8000 183.6000 259.6000 184.4000 ;
	    RECT 252.5000 177.7000 254.7000 178.3000 ;
	    RECT 250.9000 174.4000 251.5000 177.6000 ;
	    RECT 254.1000 174.4000 254.7000 177.7000 ;
	    RECT 255.6000 177.6000 256.4000 178.4000 ;
	    RECT 255.7000 174.4000 256.3000 177.6000 ;
	    RECT 244.4000 173.6000 245.2000 174.4000 ;
	    RECT 249.2000 173.6000 250.0000 174.4000 ;
	    RECT 250.8000 173.6000 251.6000 174.4000 ;
	    RECT 252.4000 173.6000 253.2000 174.4000 ;
	    RECT 254.0000 173.6000 254.8000 174.4000 ;
	    RECT 255.6000 173.6000 256.4000 174.4000 ;
	    RECT 257.2000 173.6000 258.0000 174.4000 ;
	    RECT 258.8000 173.6000 259.6000 174.4000 ;
	    RECT 244.5000 168.3000 245.1000 173.6000 ;
	    RECT 249.3000 172.4000 249.9000 173.6000 ;
	    RECT 246.0000 171.6000 246.8000 172.4000 ;
	    RECT 249.2000 171.6000 250.0000 172.4000 ;
	    RECT 252.4000 172.3000 253.2000 172.4000 ;
	    RECT 252.4000 171.7000 254.7000 172.3000 ;
	    RECT 252.4000 171.6000 253.2000 171.7000 ;
	    RECT 242.9000 167.7000 246.7000 168.3000 ;
	    RECT 242.9000 164.4000 243.5000 167.7000 ;
	    RECT 242.8000 163.6000 243.6000 164.4000 ;
	    RECT 244.4000 163.6000 245.2000 164.4000 ;
	    RECT 242.8000 159.6000 243.6000 160.4000 ;
	    RECT 241.2000 157.6000 242.0000 158.4000 ;
	    RECT 238.0000 144.2000 238.8000 155.8000 ;
	    RECT 242.9000 150.4000 243.5000 159.6000 ;
	    RECT 242.8000 149.6000 243.6000 150.4000 ;
	    RECT 244.5000 146.3000 245.1000 163.6000 ;
	    RECT 246.1000 160.4000 246.7000 167.7000 ;
	    RECT 246.0000 159.6000 246.8000 160.4000 ;
	    RECT 249.2000 159.6000 250.0000 160.4000 ;
	    RECT 246.0000 157.6000 246.8000 158.4000 ;
	    RECT 246.1000 150.4000 246.7000 157.6000 ;
	    RECT 246.0000 149.6000 246.8000 150.4000 ;
	    RECT 244.5000 145.7000 246.7000 146.3000 ;
	    RECT 244.4000 143.6000 245.2000 144.4000 ;
	    RECT 241.2000 138.3000 242.0000 138.4000 ;
	    RECT 242.8000 138.3000 243.6000 138.4000 ;
	    RECT 231.6000 135.6000 232.4000 136.4000 ;
	    RECT 228.4000 131.6000 229.2000 132.4000 ;
	    RECT 228.5000 126.4000 229.1000 131.6000 ;
	    RECT 231.6000 127.6000 232.4000 128.4000 ;
	    RECT 228.4000 125.6000 229.2000 126.4000 ;
	    RECT 230.0000 125.6000 230.8000 126.4000 ;
	    RECT 228.4000 110.3000 229.2000 110.4000 ;
	    RECT 230.1000 110.3000 230.7000 125.6000 ;
	    RECT 231.7000 110.4000 232.3000 127.6000 ;
	    RECT 233.2000 126.2000 234.0000 137.8000 ;
	    RECT 236.5000 137.7000 238.7000 138.3000 ;
	    RECT 236.4000 130.2000 237.2000 135.8000 ;
	    RECT 238.1000 132.4000 238.7000 137.7000 ;
	    RECT 241.2000 137.7000 243.6000 138.3000 ;
	    RECT 241.2000 137.6000 242.0000 137.7000 ;
	    RECT 242.8000 137.6000 243.6000 137.7000 ;
	    RECT 238.0000 131.6000 238.8000 132.4000 ;
	    RECT 241.2000 123.6000 242.0000 124.4000 ;
	    RECT 242.8000 123.6000 243.6000 124.4000 ;
	    RECT 238.0000 121.6000 238.8000 122.4000 ;
	    RECT 233.2000 111.6000 234.0000 112.4000 ;
	    RECT 233.3000 110.4000 233.9000 111.6000 ;
	    RECT 228.4000 109.7000 230.7000 110.3000 ;
	    RECT 228.4000 109.6000 229.2000 109.7000 ;
	    RECT 231.6000 109.6000 232.4000 110.4000 ;
	    RECT 233.2000 109.6000 234.0000 110.4000 ;
	    RECT 236.4000 109.6000 237.2000 110.4000 ;
	    RECT 228.4000 107.6000 229.2000 108.4000 ;
	    RECT 228.5000 106.4000 229.1000 107.6000 ;
	    RECT 223.6000 105.6000 224.4000 106.4000 ;
	    RECT 226.8000 105.6000 227.6000 106.4000 ;
	    RECT 228.4000 105.6000 229.2000 106.4000 ;
	    RECT 231.6000 105.6000 232.4000 106.4000 ;
	    RECT 233.2000 105.6000 234.0000 106.4000 ;
	    RECT 236.4000 105.6000 237.2000 106.4000 ;
	    RECT 222.0000 95.6000 222.8000 96.4000 ;
	    RECT 223.7000 96.3000 224.3000 105.6000 ;
	    RECT 225.2000 103.6000 226.0000 104.4000 ;
	    RECT 225.3000 98.4000 225.9000 103.6000 ;
	    RECT 228.4000 101.6000 229.2000 102.4000 ;
	    RECT 225.2000 97.6000 226.0000 98.4000 ;
	    RECT 225.2000 96.3000 226.0000 96.4000 ;
	    RECT 223.7000 95.7000 226.0000 96.3000 ;
	    RECT 225.2000 95.6000 226.0000 95.7000 ;
	    RECT 228.5000 92.4000 229.1000 101.6000 ;
	    RECT 230.0000 95.6000 230.8000 96.4000 ;
	    RECT 230.1000 94.4000 230.7000 95.6000 ;
	    RECT 230.0000 93.6000 230.8000 94.4000 ;
	    RECT 230.1000 92.4000 230.7000 93.6000 ;
	    RECT 222.0000 91.6000 222.8000 92.4000 ;
	    RECT 223.6000 91.6000 224.4000 92.4000 ;
	    RECT 228.4000 91.6000 229.2000 92.4000 ;
	    RECT 230.0000 91.6000 230.8000 92.4000 ;
	    RECT 223.7000 84.4000 224.3000 91.6000 ;
	    RECT 226.8000 85.6000 227.6000 86.4000 ;
	    RECT 220.4000 83.6000 221.2000 84.4000 ;
	    RECT 223.6000 83.6000 224.4000 84.4000 ;
	    RECT 230.0000 83.6000 230.8000 84.4000 ;
	    RECT 217.2000 79.6000 218.0000 80.4000 ;
	    RECT 210.8000 71.6000 211.6000 72.4000 ;
	    RECT 215.6000 71.6000 216.4000 72.4000 ;
	    RECT 223.6000 71.6000 224.4000 72.4000 ;
	    RECT 225.3000 71.7000 229.1000 72.3000 ;
	    RECT 215.7000 70.4000 216.3000 71.6000 ;
	    RECT 215.6000 69.6000 216.4000 70.4000 ;
	    RECT 217.2000 69.6000 218.0000 70.4000 ;
	    RECT 223.6000 70.3000 224.4000 70.4000 ;
	    RECT 225.3000 70.3000 225.9000 71.7000 ;
	    RECT 228.5000 70.4000 229.1000 71.7000 ;
	    RECT 223.6000 69.7000 225.9000 70.3000 ;
	    RECT 223.6000 69.6000 224.4000 69.7000 ;
	    RECT 226.8000 69.6000 227.6000 70.4000 ;
	    RECT 228.4000 69.6000 229.2000 70.4000 ;
	    RECT 217.3000 68.4000 217.9000 69.6000 ;
	    RECT 226.9000 68.4000 227.5000 69.6000 ;
	    RECT 230.1000 68.4000 230.7000 83.6000 ;
	    RECT 231.7000 78.4000 232.3000 105.6000 ;
	    RECT 233.3000 94.3000 233.9000 105.6000 ;
	    RECT 233.3000 93.7000 235.5000 94.3000 ;
	    RECT 233.2000 91.6000 234.0000 92.4000 ;
	    RECT 233.3000 90.4000 233.9000 91.6000 ;
	    RECT 233.2000 89.6000 234.0000 90.4000 ;
	    RECT 234.9000 88.3000 235.5000 93.7000 ;
	    RECT 238.1000 92.4000 238.7000 121.6000 ;
	    RECT 244.5000 118.3000 245.1000 143.6000 ;
	    RECT 246.1000 132.4000 246.7000 145.7000 ;
	    RECT 247.6000 144.2000 248.4000 155.8000 ;
	    RECT 249.3000 150.4000 249.9000 159.6000 ;
	    RECT 254.1000 158.4000 254.7000 171.7000 ;
	    RECT 255.6000 171.6000 256.4000 172.4000 ;
	    RECT 254.0000 157.6000 254.8000 158.4000 ;
	    RECT 255.7000 152.4000 256.3000 171.6000 ;
	    RECT 257.3000 164.4000 257.9000 173.6000 ;
	    RECT 258.9000 166.4000 259.5000 173.6000 ;
	    RECT 262.1000 168.4000 262.7000 191.7000 ;
	    RECT 263.6000 191.6000 264.4000 191.7000 ;
	    RECT 265.3000 190.4000 265.9000 209.7000 ;
	    RECT 268.5000 208.3000 269.1000 229.7000 ;
	    RECT 271.6000 229.6000 272.4000 230.4000 ;
	    RECT 273.3000 228.4000 273.9000 231.7000 ;
	    RECT 274.8000 231.6000 275.6000 232.4000 ;
	    RECT 279.7000 230.4000 280.3000 251.6000 ;
	    RECT 286.1000 248.4000 286.7000 251.8000 ;
	    RECT 284.4000 247.6000 285.2000 248.4000 ;
	    RECT 286.0000 247.6000 286.8000 248.4000 ;
	    RECT 284.5000 242.4000 285.1000 247.6000 ;
	    RECT 287.6000 246.2000 288.4000 257.8000 ;
	    RECT 290.8000 250.2000 291.6000 255.8000 ;
	    RECT 292.4000 253.6000 293.2000 254.4000 ;
	    RECT 295.6000 254.3000 296.4000 254.4000 ;
	    RECT 294.1000 253.7000 296.4000 254.3000 ;
	    RECT 292.5000 252.4000 293.1000 253.6000 ;
	    RECT 292.4000 251.6000 293.2000 252.4000 ;
	    RECT 294.1000 248.4000 294.7000 253.7000 ;
	    RECT 295.6000 253.6000 296.4000 253.7000 ;
	    RECT 295.6000 251.6000 296.4000 252.4000 ;
	    RECT 295.7000 250.4000 296.3000 251.6000 ;
	    RECT 295.6000 249.6000 296.4000 250.4000 ;
	    RECT 294.0000 247.6000 294.8000 248.4000 ;
	    RECT 284.4000 241.6000 285.2000 242.4000 ;
	    RECT 282.8000 233.6000 283.6000 234.4000 ;
	    RECT 281.2000 231.6000 282.0000 232.4000 ;
	    RECT 281.3000 230.4000 281.9000 231.6000 ;
	    RECT 274.8000 229.6000 275.6000 230.4000 ;
	    RECT 279.6000 229.6000 280.4000 230.4000 ;
	    RECT 281.2000 229.6000 282.0000 230.4000 ;
	    RECT 274.9000 228.4000 275.5000 229.6000 ;
	    RECT 279.7000 228.4000 280.3000 229.6000 ;
	    RECT 273.2000 227.6000 274.0000 228.4000 ;
	    RECT 274.8000 227.6000 275.6000 228.4000 ;
	    RECT 279.6000 227.6000 280.4000 228.4000 ;
	    RECT 281.2000 227.6000 282.0000 228.4000 ;
	    RECT 274.8000 225.6000 275.6000 226.4000 ;
	    RECT 278.0000 225.6000 278.8000 226.4000 ;
	    RECT 270.0000 223.6000 270.8000 224.4000 ;
	    RECT 270.1000 208.4000 270.7000 223.6000 ;
	    RECT 278.0000 215.6000 278.8000 216.4000 ;
	    RECT 278.1000 214.4000 278.7000 215.6000 ;
	    RECT 281.3000 214.4000 281.9000 227.6000 ;
	    RECT 282.9000 222.4000 283.5000 233.6000 ;
	    RECT 284.4000 231.6000 285.2000 232.4000 ;
	    RECT 292.4000 231.6000 293.2000 232.4000 ;
	    RECT 284.5000 228.4000 285.1000 231.6000 ;
	    RECT 287.6000 229.6000 288.4000 230.4000 ;
	    RECT 284.4000 227.6000 285.2000 228.4000 ;
	    RECT 286.0000 227.6000 286.8000 228.4000 ;
	    RECT 286.1000 224.4000 286.7000 227.6000 ;
	    RECT 287.7000 224.4000 288.3000 229.6000 ;
	    RECT 292.5000 228.4000 293.1000 231.6000 ;
	    RECT 297.3000 230.4000 297.9000 263.6000 ;
	    RECT 300.5000 252.4000 301.1000 267.6000 ;
	    RECT 302.1000 260.4000 302.7000 267.6000 ;
	    RECT 305.3000 266.4000 305.9000 269.7000 ;
	    RECT 306.9000 268.3000 307.5000 271.6000 ;
	    RECT 308.5000 270.4000 309.1000 273.6000 ;
	    RECT 308.4000 270.3000 309.2000 270.4000 ;
	    RECT 308.4000 269.7000 310.7000 270.3000 ;
	    RECT 308.4000 269.6000 309.2000 269.7000 ;
	    RECT 306.9000 267.7000 309.1000 268.3000 ;
	    RECT 303.6000 265.6000 304.4000 266.4000 ;
	    RECT 305.2000 265.6000 306.0000 266.4000 ;
	    RECT 306.8000 265.6000 307.6000 266.4000 ;
	    RECT 303.7000 260.4000 304.3000 265.6000 ;
	    RECT 302.0000 259.6000 302.8000 260.4000 ;
	    RECT 303.6000 259.6000 304.4000 260.4000 ;
	    RECT 306.9000 258.4000 307.5000 265.6000 ;
	    RECT 308.5000 258.4000 309.1000 267.7000 ;
	    RECT 306.8000 257.6000 307.6000 258.4000 ;
	    RECT 308.4000 257.6000 309.2000 258.4000 ;
	    RECT 302.0000 253.6000 302.8000 254.4000 ;
	    RECT 300.4000 251.6000 301.2000 252.4000 ;
	    RECT 302.1000 250.3000 302.7000 253.6000 ;
	    RECT 302.1000 249.7000 304.3000 250.3000 ;
	    RECT 302.0000 241.6000 302.8000 242.4000 ;
	    RECT 298.8000 231.6000 299.6000 232.4000 ;
	    RECT 297.2000 229.6000 298.0000 230.4000 ;
	    RECT 289.2000 227.6000 290.0000 228.4000 ;
	    RECT 292.4000 227.6000 293.2000 228.4000 ;
	    RECT 286.0000 223.6000 286.8000 224.4000 ;
	    RECT 287.6000 223.6000 288.4000 224.4000 ;
	    RECT 282.8000 221.6000 283.6000 222.4000 ;
	    RECT 287.6000 221.6000 288.4000 222.4000 ;
	    RECT 287.7000 214.4000 288.3000 221.6000 ;
	    RECT 289.3000 220.4000 289.9000 227.6000 ;
	    RECT 294.0000 225.6000 294.8000 226.4000 ;
	    RECT 298.9000 226.3000 299.5000 231.6000 ;
	    RECT 302.1000 230.4000 302.7000 241.6000 ;
	    RECT 303.7000 238.4000 304.3000 249.7000 ;
	    RECT 305.2000 249.6000 306.0000 250.4000 ;
	    RECT 305.3000 242.4000 305.9000 249.6000 ;
	    RECT 310.1000 244.4000 310.7000 269.7000 ;
	    RECT 311.7000 266.4000 312.3000 277.6000 ;
	    RECT 313.3000 272.4000 313.9000 283.6000 ;
	    RECT 313.2000 271.6000 314.0000 272.4000 ;
	    RECT 314.9000 270.4000 315.5000 289.7000 ;
	    RECT 318.0000 289.6000 318.8000 290.4000 ;
	    RECT 322.8000 289.6000 323.6000 290.4000 ;
	    RECT 324.4000 289.6000 325.2000 290.4000 ;
	    RECT 316.4000 277.6000 317.2000 278.4000 ;
	    RECT 313.2000 269.6000 314.0000 270.4000 ;
	    RECT 314.8000 269.6000 315.6000 270.4000 ;
	    RECT 311.6000 265.6000 312.4000 266.4000 ;
	    RECT 313.3000 264.4000 313.9000 269.6000 ;
	    RECT 316.5000 266.4000 317.1000 277.6000 ;
	    RECT 319.6000 273.6000 320.4000 274.4000 ;
	    RECT 318.0000 271.6000 318.8000 272.4000 ;
	    RECT 318.1000 268.4000 318.7000 271.6000 ;
	    RECT 322.9000 270.4000 323.5000 289.6000 ;
	    RECT 319.6000 269.6000 320.4000 270.4000 ;
	    RECT 322.8000 269.6000 323.6000 270.4000 ;
	    RECT 318.0000 267.6000 318.8000 268.4000 ;
	    RECT 316.4000 265.6000 317.2000 266.4000 ;
	    RECT 313.2000 263.6000 314.0000 264.4000 ;
	    RECT 313.2000 257.6000 314.0000 258.4000 ;
	    RECT 313.3000 254.4000 313.9000 257.6000 ;
	    RECT 313.2000 253.6000 314.0000 254.4000 ;
	    RECT 318.0000 246.2000 318.8000 257.8000 ;
	    RECT 319.7000 252.4000 320.3000 269.6000 ;
	    RECT 324.5000 268.4000 325.1000 289.6000 ;
	    RECT 327.6000 285.6000 328.4000 286.4000 ;
	    RECT 326.0000 271.6000 326.8000 272.4000 ;
	    RECT 326.1000 268.4000 326.7000 271.6000 ;
	    RECT 329.3000 270.4000 329.9000 291.6000 ;
	    RECT 330.9000 274.4000 331.5000 309.6000 ;
	    RECT 332.5000 308.4000 333.1000 317.6000 ;
	    RECT 334.1000 308.4000 334.7000 327.6000 ;
	    RECT 338.9000 326.4000 339.5000 329.6000 ;
	    RECT 343.6000 327.6000 344.4000 328.4000 ;
	    RECT 338.8000 325.6000 339.6000 326.4000 ;
	    RECT 337.2000 311.6000 338.0000 312.4000 ;
	    RECT 337.3000 310.4000 337.9000 311.6000 ;
	    RECT 337.2000 309.6000 338.0000 310.4000 ;
	    RECT 332.4000 307.6000 333.2000 308.4000 ;
	    RECT 334.0000 307.6000 334.8000 308.4000 ;
	    RECT 332.4000 303.6000 333.2000 304.4000 ;
	    RECT 332.5000 292.4000 333.1000 303.6000 ;
	    RECT 334.0000 301.6000 334.8000 302.4000 ;
	    RECT 337.2000 301.6000 338.0000 302.4000 ;
	    RECT 332.4000 291.6000 333.2000 292.4000 ;
	    RECT 334.1000 284.4000 334.7000 301.6000 ;
	    RECT 337.3000 292.4000 337.9000 301.6000 ;
	    RECT 337.2000 291.6000 338.0000 292.4000 ;
	    RECT 335.6000 289.6000 336.4000 290.4000 ;
	    RECT 338.9000 286.4000 339.5000 325.6000 ;
	    RECT 340.4000 313.6000 341.2000 314.4000 ;
	    RECT 343.6000 313.6000 344.4000 314.4000 ;
	    RECT 340.5000 310.4000 341.1000 313.6000 ;
	    RECT 340.4000 309.6000 341.2000 310.4000 ;
	    RECT 342.0000 309.6000 342.8000 310.4000 ;
	    RECT 343.7000 308.4000 344.3000 313.6000 ;
	    RECT 345.3000 308.4000 345.9000 331.6000 ;
	    RECT 351.6000 326.2000 352.4000 337.8000 ;
	    RECT 353.2000 331.6000 354.0000 332.4000 ;
	    RECT 358.0000 331.6000 358.8000 332.4000 ;
	    RECT 343.6000 307.6000 344.4000 308.4000 ;
	    RECT 345.2000 307.6000 346.0000 308.4000 ;
	    RECT 342.0000 303.6000 342.8000 304.4000 ;
	    RECT 345.2000 303.6000 346.0000 304.4000 ;
	    RECT 350.0000 304.2000 350.8000 315.8000 ;
	    RECT 353.3000 310.4000 353.9000 331.6000 ;
	    RECT 358.1000 328.4000 358.7000 331.6000 ;
	    RECT 358.0000 327.6000 358.8000 328.4000 ;
	    RECT 361.2000 326.2000 362.0000 337.8000 ;
	    RECT 362.8000 333.6000 363.6000 334.4000 ;
	    RECT 364.4000 330.2000 365.2000 335.8000 ;
	    RECT 366.0000 331.6000 366.8000 332.4000 ;
	    RECT 353.2000 309.6000 354.0000 310.4000 ;
	    RECT 358.0000 309.4000 358.8000 310.2000 ;
	    RECT 358.1000 308.4000 358.7000 309.4000 ;
	    RECT 358.0000 307.6000 358.8000 308.4000 ;
	    RECT 359.6000 304.2000 360.4000 315.8000 ;
	    RECT 361.2000 307.6000 362.0000 308.4000 ;
	    RECT 342.1000 292.4000 342.7000 303.6000 ;
	    RECT 346.8000 301.6000 347.6000 302.4000 ;
	    RECT 346.9000 292.4000 347.5000 301.6000 ;
	    RECT 350.0000 299.6000 350.8000 300.4000 ;
	    RECT 350.1000 298.4000 350.7000 299.6000 ;
	    RECT 350.0000 297.6000 350.8000 298.4000 ;
	    RECT 340.4000 291.6000 341.2000 292.4000 ;
	    RECT 342.0000 291.6000 342.8000 292.4000 ;
	    RECT 346.8000 291.6000 347.6000 292.4000 ;
	    RECT 338.8000 285.6000 339.6000 286.4000 ;
	    RECT 342.0000 285.6000 342.8000 286.4000 ;
	    RECT 354.8000 286.2000 355.6000 297.8000 ;
	    RECT 361.3000 294.4000 361.9000 307.6000 ;
	    RECT 362.8000 306.2000 363.6000 311.8000 ;
	    RECT 364.4000 307.6000 365.2000 308.4000 ;
	    RECT 364.5000 304.4000 365.1000 307.6000 ;
	    RECT 364.4000 303.6000 365.2000 304.4000 ;
	    RECT 362.8000 295.6000 363.6000 296.4000 ;
	    RECT 361.2000 293.6000 362.0000 294.4000 ;
	    RECT 361.2000 291.6000 362.0000 292.4000 ;
	    RECT 334.0000 283.6000 334.8000 284.4000 ;
	    RECT 332.4000 278.3000 333.2000 278.4000 ;
	    RECT 334.1000 278.3000 334.7000 283.6000 ;
	    RECT 332.4000 277.7000 334.7000 278.3000 ;
	    RECT 332.4000 277.6000 333.2000 277.7000 ;
	    RECT 330.8000 273.6000 331.6000 274.4000 ;
	    RECT 329.2000 269.6000 330.0000 270.4000 ;
	    RECT 321.2000 267.6000 322.0000 268.4000 ;
	    RECT 324.4000 267.6000 325.2000 268.4000 ;
	    RECT 326.0000 267.6000 326.8000 268.4000 ;
	    RECT 330.8000 267.6000 331.6000 268.4000 ;
	    RECT 319.6000 251.6000 320.4000 252.4000 ;
	    RECT 310.0000 243.6000 310.8000 244.4000 ;
	    RECT 305.2000 241.6000 306.0000 242.4000 ;
	    RECT 321.3000 238.4000 321.9000 267.6000 ;
	    RECT 324.5000 266.4000 325.1000 267.6000 ;
	    RECT 324.4000 265.6000 325.2000 266.4000 ;
	    RECT 330.9000 264.4000 331.5000 267.6000 ;
	    RECT 330.8000 263.6000 331.6000 264.4000 ;
	    RECT 337.2000 264.2000 338.0000 275.8000 ;
	    RECT 340.4000 273.6000 341.2000 274.4000 ;
	    RECT 338.8000 269.6000 339.6000 270.4000 ;
	    RECT 326.0000 251.6000 326.8000 252.6000 ;
	    RECT 327.6000 246.2000 328.4000 257.8000 ;
	    RECT 330.8000 250.2000 331.6000 255.8000 ;
	    RECT 332.4000 253.6000 333.2000 254.4000 ;
	    RECT 337.2000 253.6000 338.0000 254.4000 ;
	    RECT 337.3000 252.4000 337.9000 253.6000 ;
	    RECT 337.2000 251.6000 338.0000 252.4000 ;
	    RECT 335.6000 249.6000 336.4000 250.4000 ;
	    RECT 303.6000 237.6000 304.4000 238.4000 ;
	    RECT 321.2000 237.6000 322.0000 238.4000 ;
	    RECT 305.2000 233.6000 306.0000 234.4000 ;
	    RECT 308.4000 233.6000 309.2000 234.4000 ;
	    RECT 318.0000 233.6000 318.8000 234.4000 ;
	    RECT 308.5000 230.4000 309.1000 233.6000 ;
	    RECT 318.1000 230.4000 318.7000 233.6000 ;
	    RECT 302.0000 229.6000 302.8000 230.4000 ;
	    RECT 303.6000 229.6000 304.4000 230.4000 ;
	    RECT 308.4000 229.6000 309.2000 230.4000 ;
	    RECT 311.6000 229.6000 312.4000 230.4000 ;
	    RECT 313.2000 229.6000 314.0000 230.4000 ;
	    RECT 318.0000 229.6000 318.8000 230.4000 ;
	    RECT 324.4000 229.6000 325.2000 230.4000 ;
	    RECT 303.7000 228.4000 304.3000 229.6000 ;
	    RECT 302.0000 227.6000 302.8000 228.4000 ;
	    RECT 303.6000 227.6000 304.4000 228.4000 ;
	    RECT 297.3000 225.7000 299.5000 226.3000 ;
	    RECT 290.8000 221.6000 291.6000 222.4000 ;
	    RECT 289.2000 219.6000 290.0000 220.4000 ;
	    RECT 289.2000 217.6000 290.0000 218.4000 ;
	    RECT 289.3000 216.4000 289.9000 217.6000 ;
	    RECT 289.2000 215.6000 290.0000 216.4000 ;
	    RECT 271.6000 213.6000 272.4000 214.4000 ;
	    RECT 278.0000 213.6000 278.8000 214.4000 ;
	    RECT 281.2000 213.6000 282.0000 214.4000 ;
	    RECT 282.8000 213.6000 283.6000 214.4000 ;
	    RECT 287.6000 213.6000 288.4000 214.4000 ;
	    RECT 271.7000 212.4000 272.3000 213.6000 ;
	    RECT 271.6000 211.6000 272.4000 212.4000 ;
	    RECT 281.2000 209.6000 282.0000 210.4000 ;
	    RECT 266.9000 207.7000 269.1000 208.3000 ;
	    RECT 266.9000 196.3000 267.5000 207.7000 ;
	    RECT 270.0000 207.6000 270.8000 208.4000 ;
	    RECT 268.4000 203.6000 269.2000 204.4000 ;
	    RECT 273.2000 203.6000 274.0000 204.4000 ;
	    RECT 268.5000 200.3000 269.1000 203.6000 ;
	    RECT 273.3000 200.4000 273.9000 203.6000 ;
	    RECT 274.8000 201.6000 275.6000 202.4000 ;
	    RECT 268.5000 199.7000 270.7000 200.3000 ;
	    RECT 268.4000 197.6000 269.2000 198.4000 ;
	    RECT 266.9000 195.7000 269.1000 196.3000 ;
	    RECT 266.8000 193.6000 267.6000 194.4000 ;
	    RECT 265.2000 189.6000 266.0000 190.4000 ;
	    RECT 263.6000 183.6000 264.4000 184.4000 ;
	    RECT 263.7000 182.4000 264.3000 183.6000 ;
	    RECT 263.6000 181.6000 264.4000 182.4000 ;
	    RECT 265.3000 180.4000 265.9000 189.6000 ;
	    RECT 266.9000 188.4000 267.5000 193.6000 ;
	    RECT 268.5000 190.3000 269.1000 195.7000 ;
	    RECT 270.1000 192.4000 270.7000 199.7000 ;
	    RECT 271.6000 199.6000 272.4000 200.4000 ;
	    RECT 273.2000 199.6000 274.0000 200.4000 ;
	    RECT 270.0000 191.6000 270.8000 192.4000 ;
	    RECT 268.5000 189.7000 270.7000 190.3000 ;
	    RECT 266.8000 187.6000 267.6000 188.4000 ;
	    RECT 265.2000 179.6000 266.0000 180.4000 ;
	    RECT 263.6000 177.6000 264.4000 178.4000 ;
	    RECT 263.7000 176.4000 264.3000 177.6000 ;
	    RECT 263.6000 175.6000 264.4000 176.4000 ;
	    RECT 265.3000 174.3000 265.9000 179.6000 ;
	    RECT 268.4000 177.6000 269.2000 178.4000 ;
	    RECT 270.1000 176.3000 270.7000 189.7000 ;
	    RECT 271.7000 176.4000 272.3000 199.6000 ;
	    RECT 273.2000 184.2000 274.0000 195.8000 ;
	    RECT 274.9000 192.4000 275.5000 201.6000 ;
	    RECT 281.3000 200.4000 281.9000 209.6000 ;
	    RECT 282.9000 202.4000 283.5000 213.6000 ;
	    RECT 287.6000 211.6000 288.4000 212.4000 ;
	    RECT 284.4000 209.6000 285.2000 210.4000 ;
	    RECT 286.0000 209.6000 286.8000 210.4000 ;
	    RECT 282.8000 201.6000 283.6000 202.4000 ;
	    RECT 278.0000 199.6000 278.8000 200.4000 ;
	    RECT 281.2000 199.6000 282.0000 200.4000 ;
	    RECT 274.8000 191.6000 275.6000 192.4000 ;
	    RECT 274.8000 189.6000 275.6000 190.4000 ;
	    RECT 274.9000 182.4000 275.5000 189.6000 ;
	    RECT 278.1000 184.4000 278.7000 199.6000 ;
	    RECT 284.5000 196.4000 285.1000 209.6000 ;
	    RECT 287.7000 202.4000 288.3000 211.6000 ;
	    RECT 287.6000 201.6000 288.4000 202.4000 ;
	    RECT 290.9000 200.3000 291.5000 221.6000 ;
	    RECT 294.0000 206.2000 294.8000 217.8000 ;
	    RECT 287.7000 199.7000 291.5000 200.3000 ;
	    RECT 287.7000 198.4000 288.3000 199.7000 ;
	    RECT 287.6000 197.6000 288.4000 198.4000 ;
	    RECT 289.2000 197.6000 290.0000 198.4000 ;
	    RECT 279.6000 189.6000 280.4000 190.4000 ;
	    RECT 278.0000 183.6000 278.8000 184.4000 ;
	    RECT 274.8000 181.6000 275.6000 182.4000 ;
	    RECT 263.7000 173.7000 265.9000 174.3000 ;
	    RECT 268.5000 175.7000 270.7000 176.3000 ;
	    RECT 263.7000 172.4000 264.3000 173.7000 ;
	    RECT 263.6000 171.6000 264.4000 172.4000 ;
	    RECT 266.8000 171.6000 267.6000 172.4000 ;
	    RECT 266.9000 168.4000 267.5000 171.6000 ;
	    RECT 262.0000 167.6000 262.8000 168.4000 ;
	    RECT 266.8000 167.6000 267.6000 168.4000 ;
	    RECT 258.8000 165.6000 259.6000 166.4000 ;
	    RECT 260.4000 165.6000 261.2000 166.4000 ;
	    RECT 268.5000 166.3000 269.1000 175.7000 ;
	    RECT 271.6000 175.6000 272.4000 176.4000 ;
	    RECT 266.9000 165.7000 269.1000 166.3000 ;
	    RECT 273.2000 166.2000 274.0000 177.8000 ;
	    RECT 274.8000 177.6000 275.6000 178.4000 ;
	    RECT 257.2000 163.6000 258.0000 164.4000 ;
	    RECT 258.8000 153.6000 259.6000 154.4000 ;
	    RECT 258.9000 152.4000 259.5000 153.6000 ;
	    RECT 255.6000 151.6000 256.4000 152.4000 ;
	    RECT 258.8000 151.6000 259.6000 152.4000 ;
	    RECT 249.2000 149.6000 250.0000 150.4000 ;
	    RECT 260.5000 146.4000 261.1000 165.6000 ;
	    RECT 265.2000 162.3000 266.0000 162.4000 ;
	    RECT 266.9000 162.3000 267.5000 165.7000 ;
	    RECT 268.4000 163.6000 269.2000 164.4000 ;
	    RECT 265.2000 161.7000 267.5000 162.3000 ;
	    RECT 265.2000 161.6000 266.0000 161.7000 ;
	    RECT 262.0000 157.6000 262.8000 158.4000 ;
	    RECT 260.4000 145.6000 261.2000 146.4000 ;
	    RECT 250.8000 143.6000 251.6000 144.4000 ;
	    RECT 252.4000 143.6000 253.2000 144.4000 ;
	    RECT 249.2000 141.6000 250.0000 142.4000 ;
	    RECT 249.3000 138.4000 249.9000 141.6000 ;
	    RECT 250.9000 140.4000 251.5000 143.6000 ;
	    RECT 250.8000 139.6000 251.6000 140.4000 ;
	    RECT 247.6000 137.6000 248.4000 138.4000 ;
	    RECT 249.2000 137.6000 250.0000 138.4000 ;
	    RECT 247.7000 134.4000 248.3000 137.6000 ;
	    RECT 247.6000 133.6000 248.4000 134.4000 ;
	    RECT 246.0000 131.6000 246.8000 132.4000 ;
	    RECT 249.2000 132.3000 250.0000 132.4000 ;
	    RECT 250.9000 132.3000 251.5000 139.6000 ;
	    RECT 249.2000 131.7000 251.5000 132.3000 ;
	    RECT 249.2000 131.6000 250.0000 131.7000 ;
	    RECT 252.5000 130.4000 253.1000 143.6000 ;
	    RECT 258.8000 133.6000 259.6000 134.4000 ;
	    RECT 260.4000 133.6000 261.2000 134.4000 ;
	    RECT 252.4000 129.6000 253.2000 130.4000 ;
	    RECT 252.5000 126.4000 253.1000 129.6000 ;
	    RECT 258.9000 128.4000 259.5000 133.6000 ;
	    RECT 260.5000 128.4000 261.1000 133.6000 ;
	    RECT 258.8000 127.6000 259.6000 128.4000 ;
	    RECT 260.4000 127.6000 261.2000 128.4000 ;
	    RECT 252.4000 125.6000 253.2000 126.4000 ;
	    RECT 247.6000 119.6000 248.4000 120.4000 ;
	    RECT 242.9000 117.7000 245.1000 118.3000 ;
	    RECT 239.6000 111.6000 240.4000 112.4000 ;
	    RECT 239.7000 98.4000 240.3000 111.6000 ;
	    RECT 242.9000 110.4000 243.5000 117.7000 ;
	    RECT 246.0000 117.6000 246.8000 118.4000 ;
	    RECT 246.1000 116.3000 246.7000 117.6000 ;
	    RECT 244.5000 115.7000 246.7000 116.3000 ;
	    RECT 241.2000 109.6000 242.0000 110.4000 ;
	    RECT 242.8000 109.6000 243.6000 110.4000 ;
	    RECT 241.3000 108.4000 241.9000 109.6000 ;
	    RECT 241.2000 107.6000 242.0000 108.4000 ;
	    RECT 242.8000 108.3000 243.6000 108.4000 ;
	    RECT 244.5000 108.3000 245.1000 115.7000 ;
	    RECT 247.7000 114.3000 248.3000 119.6000 ;
	    RECT 246.1000 113.7000 248.3000 114.3000 ;
	    RECT 246.1000 112.4000 246.7000 113.7000 ;
	    RECT 246.0000 111.6000 246.8000 112.4000 ;
	    RECT 247.6000 111.6000 248.4000 112.4000 ;
	    RECT 246.0000 109.6000 246.8000 110.4000 ;
	    RECT 242.8000 107.7000 245.1000 108.3000 ;
	    RECT 242.8000 107.6000 243.6000 107.7000 ;
	    RECT 239.6000 97.6000 240.4000 98.4000 ;
	    RECT 241.2000 97.6000 242.0000 98.4000 ;
	    RECT 241.3000 96.4000 241.9000 97.6000 ;
	    RECT 241.2000 95.6000 242.0000 96.4000 ;
	    RECT 239.6000 93.6000 240.4000 94.4000 ;
	    RECT 238.0000 91.6000 238.8000 92.4000 ;
	    RECT 238.0000 89.6000 238.8000 90.4000 ;
	    RECT 233.3000 87.7000 235.5000 88.3000 ;
	    RECT 233.3000 78.4000 233.9000 87.7000 ;
	    RECT 234.8000 85.6000 235.6000 86.4000 ;
	    RECT 231.6000 77.6000 232.4000 78.4000 ;
	    RECT 233.2000 77.6000 234.0000 78.4000 ;
	    RECT 234.9000 72.4000 235.5000 85.6000 ;
	    RECT 239.7000 80.4000 240.3000 93.6000 ;
	    RECT 239.6000 79.6000 240.4000 80.4000 ;
	    RECT 238.0000 77.6000 238.8000 78.4000 ;
	    RECT 236.4000 75.6000 237.2000 76.4000 ;
	    RECT 234.8000 71.6000 235.6000 72.4000 ;
	    RECT 231.6000 69.6000 232.4000 70.4000 ;
	    RECT 233.2000 69.6000 234.0000 70.4000 ;
	    RECT 209.2000 67.6000 210.0000 68.4000 ;
	    RECT 217.2000 67.6000 218.0000 68.4000 ;
	    RECT 226.8000 67.6000 227.6000 68.4000 ;
	    RECT 230.0000 67.6000 230.8000 68.4000 ;
	    RECT 202.8000 63.6000 203.6000 64.4000 ;
	    RECT 202.9000 52.4000 203.5000 63.6000 ;
	    RECT 209.3000 62.4000 209.9000 67.6000 ;
	    RECT 217.2000 65.6000 218.0000 66.4000 ;
	    RECT 230.0000 65.6000 230.8000 66.4000 ;
	    RECT 207.6000 61.6000 208.4000 62.4000 ;
	    RECT 209.2000 61.6000 210.0000 62.4000 ;
	    RECT 210.8000 61.6000 211.6000 62.4000 ;
	    RECT 204.4000 57.6000 205.2000 58.4000 ;
	    RECT 204.5000 54.4000 205.1000 57.6000 ;
	    RECT 204.4000 53.6000 205.2000 54.4000 ;
	    RECT 202.8000 51.6000 203.6000 52.4000 ;
	    RECT 204.4000 51.6000 205.2000 52.4000 ;
	    RECT 206.0000 51.6000 206.8000 52.4000 ;
	    RECT 202.8000 47.6000 203.6000 48.4000 ;
	    RECT 201.3000 45.7000 203.5000 46.3000 ;
	    RECT 201.2000 31.6000 202.0000 32.4000 ;
	    RECT 201.3000 30.4000 201.9000 31.6000 ;
	    RECT 191.6000 29.6000 192.4000 30.4000 ;
	    RECT 194.8000 29.6000 195.6000 30.4000 ;
	    RECT 196.4000 29.6000 197.2000 30.4000 ;
	    RECT 198.0000 29.6000 198.8000 30.4000 ;
	    RECT 201.2000 29.6000 202.0000 30.4000 ;
	    RECT 194.8000 27.6000 195.6000 28.4000 ;
	    RECT 194.9000 26.4000 195.5000 27.6000 ;
	    RECT 196.5000 26.4000 197.1000 29.6000 ;
	    RECT 201.2000 27.6000 202.0000 28.4000 ;
	    RECT 185.2000 25.6000 186.0000 26.4000 ;
	    RECT 190.0000 25.6000 190.8000 26.4000 ;
	    RECT 194.8000 25.6000 195.6000 26.4000 ;
	    RECT 196.4000 25.6000 197.2000 26.4000 ;
	    RECT 172.4000 11.6000 173.2000 12.4000 ;
	    RECT 178.8000 11.6000 179.6000 12.6000 ;
	    RECT 180.4000 6.2000 181.2000 17.8000 ;
	    RECT 182.0000 13.6000 182.8000 14.4000 ;
	    RECT 182.1000 12.4000 182.7000 13.6000 ;
	    RECT 182.0000 11.6000 182.8000 12.4000 ;
	    RECT 183.6000 10.2000 184.4000 15.8000 ;
	    RECT 185.3000 12.4000 185.9000 25.6000 ;
	    RECT 190.1000 18.4000 190.7000 25.6000 ;
	    RECT 190.0000 17.6000 190.8000 18.4000 ;
	    RECT 185.2000 11.6000 186.0000 12.4000 ;
	    RECT 194.8000 6.2000 195.6000 17.8000 ;
	    RECT 196.4000 11.6000 197.2000 12.4000 ;
	    RECT 196.5000 8.4000 197.1000 11.6000 ;
	    RECT 201.3000 10.4000 201.9000 27.6000 ;
	    RECT 202.9000 16.4000 203.5000 45.7000 ;
	    RECT 204.5000 40.4000 205.1000 51.6000 ;
	    RECT 206.1000 50.4000 206.7000 51.6000 ;
	    RECT 207.7000 50.4000 208.3000 61.6000 ;
	    RECT 210.9000 54.4000 211.5000 61.6000 ;
	    RECT 220.4000 59.6000 221.2000 60.4000 ;
	    RECT 217.2000 57.6000 218.0000 58.4000 ;
	    RECT 212.4000 55.6000 213.2000 56.4000 ;
	    RECT 217.3000 54.4000 217.9000 57.6000 ;
	    RECT 210.8000 53.6000 211.6000 54.4000 ;
	    RECT 217.2000 53.6000 218.0000 54.4000 ;
	    RECT 218.8000 53.6000 219.6000 54.4000 ;
	    RECT 218.9000 52.4000 219.5000 53.6000 ;
	    RECT 210.8000 51.6000 211.6000 52.4000 ;
	    RECT 215.6000 51.6000 216.4000 52.4000 ;
	    RECT 218.8000 51.6000 219.6000 52.4000 ;
	    RECT 206.0000 49.6000 206.8000 50.4000 ;
	    RECT 207.6000 49.6000 208.4000 50.4000 ;
	    RECT 212.4000 49.6000 213.2000 50.4000 ;
	    RECT 215.7000 40.4000 216.3000 51.6000 ;
	    RECT 220.5000 50.4000 221.1000 59.6000 ;
	    RECT 230.1000 58.4000 230.7000 65.6000 ;
	    RECT 223.6000 57.6000 224.4000 58.4000 ;
	    RECT 230.0000 57.6000 230.8000 58.4000 ;
	    RECT 222.0000 55.6000 222.8000 56.4000 ;
	    RECT 222.1000 52.4000 222.7000 55.6000 ;
	    RECT 223.7000 54.4000 224.3000 57.6000 ;
	    RECT 231.7000 56.4000 232.3000 69.6000 ;
	    RECT 234.9000 68.4000 235.5000 71.6000 ;
	    RECT 236.4000 70.3000 237.2000 70.4000 ;
	    RECT 238.1000 70.3000 238.7000 77.6000 ;
	    RECT 239.6000 71.6000 240.4000 72.4000 ;
	    RECT 239.7000 70.4000 240.3000 71.6000 ;
	    RECT 236.4000 69.7000 238.7000 70.3000 ;
	    RECT 236.4000 69.6000 237.2000 69.7000 ;
	    RECT 239.6000 69.6000 240.4000 70.4000 ;
	    RECT 242.9000 68.4000 243.5000 107.6000 ;
	    RECT 247.6000 105.6000 248.4000 106.4000 ;
	    RECT 255.6000 106.2000 256.4000 111.8000 ;
	    RECT 244.4000 99.6000 245.2000 100.4000 ;
	    RECT 244.5000 94.4000 245.1000 99.6000 ;
	    RECT 244.4000 93.6000 245.2000 94.4000 ;
	    RECT 246.0000 86.2000 246.8000 97.8000 ;
	    RECT 246.0000 82.3000 246.8000 82.4000 ;
	    RECT 247.7000 82.3000 248.3000 105.6000 ;
	    RECT 258.8000 104.2000 259.6000 115.8000 ;
	    RECT 260.4000 109.4000 261.2000 110.4000 ;
	    RECT 262.1000 108.4000 262.7000 157.6000 ;
	    RECT 265.3000 150.4000 265.9000 161.6000 ;
	    RECT 268.5000 160.3000 269.1000 163.6000 ;
	    RECT 268.5000 159.7000 270.7000 160.3000 ;
	    RECT 270.1000 154.4000 270.7000 159.7000 ;
	    RECT 270.0000 153.6000 270.8000 154.4000 ;
	    RECT 274.9000 150.4000 275.5000 177.6000 ;
	    RECT 276.4000 151.6000 277.2000 152.4000 ;
	    RECT 276.5000 150.4000 277.1000 151.6000 ;
	    RECT 265.2000 149.6000 266.0000 150.4000 ;
	    RECT 266.8000 149.6000 267.6000 150.4000 ;
	    RECT 270.0000 149.6000 270.8000 150.4000 ;
	    RECT 274.8000 149.6000 275.6000 150.4000 ;
	    RECT 276.4000 149.6000 277.2000 150.4000 ;
	    RECT 265.2000 147.6000 266.0000 148.4000 ;
	    RECT 263.6000 145.6000 264.4000 146.4000 ;
	    RECT 263.7000 132.4000 264.3000 145.6000 ;
	    RECT 265.3000 136.4000 265.9000 147.6000 ;
	    RECT 266.9000 144.4000 267.5000 149.6000 ;
	    RECT 271.6000 147.6000 272.4000 148.4000 ;
	    RECT 266.8000 143.6000 267.6000 144.4000 ;
	    RECT 266.8000 139.6000 267.6000 140.4000 ;
	    RECT 265.2000 135.6000 266.0000 136.4000 ;
	    RECT 265.2000 134.3000 266.0000 134.4000 ;
	    RECT 266.9000 134.3000 267.5000 139.6000 ;
	    RECT 278.1000 138.4000 278.7000 183.6000 ;
	    RECT 279.7000 182.4000 280.3000 189.6000 ;
	    RECT 281.2000 185.6000 282.0000 186.4000 ;
	    RECT 279.6000 181.6000 280.4000 182.4000 ;
	    RECT 281.3000 174.4000 281.9000 185.6000 ;
	    RECT 282.8000 184.2000 283.6000 195.8000 ;
	    RECT 284.4000 195.6000 285.2000 196.4000 ;
	    RECT 284.4000 187.6000 285.2000 188.4000 ;
	    RECT 284.5000 184.4000 285.1000 187.6000 ;
	    RECT 286.0000 186.2000 286.8000 191.8000 ;
	    RECT 284.4000 183.6000 285.2000 184.4000 ;
	    RECT 287.6000 183.6000 288.4000 184.4000 ;
	    RECT 284.4000 179.6000 285.2000 180.4000 ;
	    RECT 281.2000 173.6000 282.0000 174.4000 ;
	    RECT 279.6000 171.6000 280.4000 172.4000 ;
	    RECT 279.7000 158.4000 280.3000 171.6000 ;
	    RECT 281.3000 158.4000 281.9000 173.6000 ;
	    RECT 282.8000 166.2000 283.6000 177.8000 ;
	    RECT 284.5000 170.4000 285.1000 179.6000 ;
	    RECT 284.4000 169.6000 285.2000 170.4000 ;
	    RECT 286.0000 170.2000 286.8000 175.8000 ;
	    RECT 287.7000 174.4000 288.3000 183.6000 ;
	    RECT 287.6000 173.6000 288.4000 174.4000 ;
	    RECT 289.3000 172.4000 289.9000 197.6000 ;
	    RECT 292.4000 191.6000 293.2000 192.4000 ;
	    RECT 292.5000 190.4000 293.1000 191.6000 ;
	    RECT 297.3000 190.4000 297.9000 225.7000 ;
	    RECT 298.8000 223.6000 299.6000 224.4000 ;
	    RECT 298.9000 204.4000 299.5000 223.6000 ;
	    RECT 300.4000 211.6000 301.2000 212.4000 ;
	    RECT 300.5000 210.4000 301.1000 211.6000 ;
	    RECT 302.1000 210.4000 302.7000 227.6000 ;
	    RECT 300.4000 209.6000 301.2000 210.4000 ;
	    RECT 302.0000 209.6000 302.8000 210.4000 ;
	    RECT 303.6000 206.2000 304.4000 217.8000 ;
	    RECT 305.2000 213.6000 306.0000 214.4000 ;
	    RECT 306.8000 210.2000 307.6000 215.8000 ;
	    RECT 308.4000 215.6000 309.2000 216.4000 ;
	    RECT 310.0000 215.6000 310.8000 216.4000 ;
	    RECT 308.5000 212.4000 309.1000 215.6000 ;
	    RECT 310.1000 212.4000 310.7000 215.6000 ;
	    RECT 308.4000 211.6000 309.2000 212.4000 ;
	    RECT 310.0000 211.6000 310.8000 212.4000 ;
	    RECT 311.7000 210.4000 312.3000 229.6000 ;
	    RECT 313.3000 228.4000 313.9000 229.6000 ;
	    RECT 313.2000 227.6000 314.0000 228.4000 ;
	    RECT 314.8000 223.6000 315.6000 224.4000 ;
	    RECT 316.4000 223.6000 317.2000 224.4000 ;
	    RECT 322.8000 223.6000 323.6000 224.4000 ;
	    RECT 316.5000 212.4000 317.1000 223.6000 ;
	    RECT 319.6000 215.6000 320.4000 216.4000 ;
	    RECT 319.7000 212.4000 320.3000 215.6000 ;
	    RECT 316.4000 211.6000 317.2000 212.4000 ;
	    RECT 318.0000 211.6000 318.8000 212.4000 ;
	    RECT 319.6000 211.6000 320.4000 212.4000 ;
	    RECT 322.9000 212.3000 323.5000 223.6000 ;
	    RECT 324.5000 214.3000 325.1000 229.6000 ;
	    RECT 326.0000 225.6000 326.8000 226.4000 ;
	    RECT 326.1000 224.4000 326.7000 225.6000 ;
	    RECT 326.0000 223.6000 326.8000 224.4000 ;
	    RECT 330.8000 224.2000 331.6000 235.8000 ;
	    RECT 337.2000 229.6000 338.0000 230.4000 ;
	    RECT 338.9000 228.4000 339.5000 269.6000 ;
	    RECT 340.5000 252.4000 341.1000 273.6000 ;
	    RECT 342.1000 254.4000 342.7000 285.6000 ;
	    RECT 343.6000 283.6000 344.4000 284.4000 ;
	    RECT 351.6000 283.6000 352.4000 284.4000 ;
	    RECT 361.2000 283.6000 362.0000 284.4000 ;
	    RECT 343.7000 272.4000 344.3000 283.6000 ;
	    RECT 343.6000 271.6000 344.4000 272.4000 ;
	    RECT 345.2000 271.6000 346.0000 272.4000 ;
	    RECT 345.3000 270.2000 345.9000 271.6000 ;
	    RECT 345.2000 269.4000 346.0000 270.2000 ;
	    RECT 346.8000 264.2000 347.6000 275.8000 ;
	    RECT 351.7000 272.4000 352.3000 283.6000 ;
	    RECT 356.4000 281.6000 357.2000 282.4000 ;
	    RECT 358.0000 281.6000 358.8000 282.4000 ;
	    RECT 350.0000 266.2000 350.8000 271.8000 ;
	    RECT 351.6000 271.6000 352.4000 272.4000 ;
	    RECT 356.5000 270.4000 357.1000 281.6000 ;
	    RECT 358.1000 278.4000 358.7000 281.6000 ;
	    RECT 358.0000 277.6000 358.8000 278.4000 ;
	    RECT 358.0000 271.6000 358.8000 272.4000 ;
	    RECT 359.6000 271.6000 360.4000 272.4000 ;
	    RECT 353.2000 269.6000 354.0000 270.4000 ;
	    RECT 354.8000 269.6000 355.6000 270.4000 ;
	    RECT 356.4000 269.6000 357.2000 270.4000 ;
	    RECT 351.6000 265.6000 352.4000 266.4000 ;
	    RECT 350.0000 261.6000 350.8000 262.4000 ;
	    RECT 342.0000 253.6000 342.8000 254.4000 ;
	    RECT 348.4000 253.6000 349.2000 254.4000 ;
	    RECT 340.4000 251.6000 341.2000 252.4000 ;
	    RECT 340.5000 250.4000 341.1000 251.6000 ;
	    RECT 340.4000 249.6000 341.2000 250.4000 ;
	    RECT 342.1000 240.4000 342.7000 253.6000 ;
	    RECT 350.1000 252.4000 350.7000 261.6000 ;
	    RECT 351.7000 254.4000 352.3000 265.6000 ;
	    RECT 354.9000 264.4000 355.5000 269.6000 ;
	    RECT 356.4000 267.6000 357.2000 268.4000 ;
	    RECT 356.5000 266.4000 357.1000 267.6000 ;
	    RECT 356.4000 265.6000 357.2000 266.4000 ;
	    RECT 354.8000 263.6000 355.6000 264.4000 ;
	    RECT 353.2000 261.6000 354.0000 262.4000 ;
	    RECT 353.3000 256.4000 353.9000 261.6000 ;
	    RECT 354.9000 258.4000 355.5000 263.6000 ;
	    RECT 354.8000 257.6000 355.6000 258.4000 ;
	    RECT 353.2000 255.6000 354.0000 256.4000 ;
	    RECT 351.6000 253.6000 352.4000 254.4000 ;
	    RECT 343.6000 251.6000 344.4000 252.4000 ;
	    RECT 350.0000 251.6000 350.8000 252.4000 ;
	    RECT 353.3000 250.4000 353.9000 255.6000 ;
	    RECT 356.5000 250.4000 357.1000 265.6000 ;
	    RECT 358.1000 264.4000 358.7000 271.6000 ;
	    RECT 359.7000 270.4000 360.3000 271.6000 ;
	    RECT 361.3000 270.4000 361.9000 283.6000 ;
	    RECT 359.6000 269.6000 360.4000 270.4000 ;
	    RECT 361.2000 269.6000 362.0000 270.4000 ;
	    RECT 358.0000 263.6000 358.8000 264.4000 ;
	    RECT 346.8000 249.6000 347.6000 250.4000 ;
	    RECT 353.2000 250.3000 354.0000 250.4000 ;
	    RECT 353.2000 249.7000 355.5000 250.3000 ;
	    RECT 353.2000 249.6000 354.0000 249.7000 ;
	    RECT 346.9000 248.4000 347.5000 249.6000 ;
	    RECT 346.8000 247.6000 347.6000 248.4000 ;
	    RECT 346.8000 243.6000 347.6000 244.4000 ;
	    RECT 342.0000 239.6000 342.8000 240.4000 ;
	    RECT 345.2000 237.6000 346.0000 238.4000 ;
	    RECT 338.8000 227.6000 339.6000 228.4000 ;
	    RECT 324.5000 213.7000 326.7000 214.3000 ;
	    RECT 324.4000 212.3000 325.2000 212.4000 ;
	    RECT 322.9000 211.7000 325.2000 212.3000 ;
	    RECT 324.4000 211.6000 325.2000 211.7000 ;
	    RECT 318.1000 210.4000 318.7000 211.6000 ;
	    RECT 310.0000 209.6000 310.8000 210.4000 ;
	    RECT 311.6000 209.6000 312.4000 210.4000 ;
	    RECT 318.0000 209.6000 318.8000 210.4000 ;
	    RECT 298.8000 203.6000 299.6000 204.4000 ;
	    RECT 302.0000 203.6000 302.8000 204.4000 ;
	    RECT 298.8000 199.6000 299.6000 200.4000 ;
	    RECT 298.9000 198.4000 299.5000 199.6000 ;
	    RECT 298.8000 197.6000 299.6000 198.4000 ;
	    RECT 302.1000 190.4000 302.7000 203.6000 ;
	    RECT 303.6000 197.6000 304.4000 198.4000 ;
	    RECT 308.4000 197.6000 309.2000 198.4000 ;
	    RECT 306.8000 193.6000 307.6000 194.4000 ;
	    RECT 306.9000 190.4000 307.5000 193.6000 ;
	    RECT 290.8000 189.6000 291.6000 190.4000 ;
	    RECT 292.4000 189.6000 293.2000 190.4000 ;
	    RECT 295.6000 189.6000 296.4000 190.4000 ;
	    RECT 297.2000 189.6000 298.0000 190.4000 ;
	    RECT 302.0000 189.6000 302.8000 190.4000 ;
	    RECT 306.8000 189.6000 307.6000 190.4000 ;
	    RECT 290.9000 178.4000 291.5000 189.6000 ;
	    RECT 292.4000 183.6000 293.2000 184.4000 ;
	    RECT 292.5000 182.4000 293.1000 183.6000 ;
	    RECT 292.4000 181.6000 293.2000 182.4000 ;
	    RECT 292.4000 179.6000 293.2000 180.4000 ;
	    RECT 294.0000 179.6000 294.8000 180.4000 ;
	    RECT 290.8000 177.6000 291.6000 178.4000 ;
	    RECT 292.5000 174.3000 293.1000 179.6000 ;
	    RECT 294.1000 178.4000 294.7000 179.6000 ;
	    RECT 295.7000 178.4000 296.3000 189.6000 ;
	    RECT 297.3000 188.4000 297.9000 189.6000 ;
	    RECT 308.5000 188.4000 309.1000 197.6000 ;
	    RECT 297.2000 187.6000 298.0000 188.4000 ;
	    RECT 308.4000 187.6000 309.2000 188.4000 ;
	    RECT 297.2000 185.6000 298.0000 186.4000 ;
	    RECT 294.0000 177.6000 294.8000 178.4000 ;
	    RECT 295.6000 177.6000 296.4000 178.4000 ;
	    RECT 290.9000 173.7000 293.1000 174.3000 ;
	    RECT 289.2000 171.6000 290.0000 172.4000 ;
	    RECT 289.3000 168.4000 289.9000 171.6000 ;
	    RECT 284.4000 167.6000 285.2000 168.4000 ;
	    RECT 286.0000 167.6000 286.8000 168.4000 ;
	    RECT 289.2000 167.6000 290.0000 168.4000 ;
	    RECT 279.6000 157.6000 280.4000 158.4000 ;
	    RECT 281.2000 157.6000 282.0000 158.4000 ;
	    RECT 284.5000 150.4000 285.1000 167.6000 ;
	    RECT 279.6000 149.6000 280.4000 150.4000 ;
	    RECT 284.4000 149.6000 285.2000 150.4000 ;
	    RECT 281.2000 147.6000 282.0000 148.4000 ;
	    RECT 281.3000 140.4000 281.9000 147.6000 ;
	    RECT 281.2000 139.6000 282.0000 140.4000 ;
	    RECT 268.4000 137.6000 269.2000 138.4000 ;
	    RECT 271.6000 137.6000 272.4000 138.4000 ;
	    RECT 278.0000 137.6000 278.8000 138.4000 ;
	    RECT 265.2000 133.7000 267.5000 134.3000 ;
	    RECT 265.2000 133.6000 266.0000 133.7000 ;
	    RECT 268.5000 132.4000 269.1000 137.6000 ;
	    RECT 270.0000 135.6000 270.8000 136.4000 ;
	    RECT 271.7000 134.4000 272.3000 137.6000 ;
	    RECT 270.0000 133.6000 270.8000 134.4000 ;
	    RECT 271.6000 133.6000 272.4000 134.4000 ;
	    RECT 263.6000 131.6000 264.4000 132.4000 ;
	    RECT 265.2000 131.6000 266.0000 132.4000 ;
	    RECT 266.8000 131.6000 267.6000 132.4000 ;
	    RECT 268.4000 131.6000 269.2000 132.4000 ;
	    RECT 265.3000 112.4000 265.9000 131.6000 ;
	    RECT 263.6000 111.6000 264.4000 112.4000 ;
	    RECT 265.2000 111.6000 266.0000 112.4000 ;
	    RECT 262.0000 107.6000 262.8000 108.4000 ;
	    RECT 262.0000 99.6000 262.8000 100.4000 ;
	    RECT 254.0000 93.6000 254.8000 94.4000 ;
	    RECT 252.4000 91.6000 253.2000 92.4000 ;
	    RECT 252.5000 90.4000 253.1000 91.6000 ;
	    RECT 252.4000 89.6000 253.2000 90.4000 ;
	    RECT 249.2000 85.6000 250.0000 86.4000 ;
	    RECT 246.0000 81.7000 248.3000 82.3000 ;
	    RECT 246.0000 81.6000 246.8000 81.7000 ;
	    RECT 249.3000 72.4000 249.9000 85.6000 ;
	    RECT 247.6000 71.6000 248.4000 72.4000 ;
	    RECT 249.2000 71.6000 250.0000 72.4000 ;
	    RECT 254.1000 72.3000 254.7000 93.6000 ;
	    RECT 255.6000 86.2000 256.4000 97.8000 ;
	    RECT 258.8000 90.2000 259.6000 95.8000 ;
	    RECT 262.1000 94.4000 262.7000 99.6000 ;
	    RECT 263.7000 98.4000 264.3000 111.6000 ;
	    RECT 265.2000 107.6000 266.0000 108.4000 ;
	    RECT 265.3000 104.4000 265.9000 107.6000 ;
	    RECT 265.2000 103.6000 266.0000 104.4000 ;
	    RECT 263.6000 97.6000 264.4000 98.4000 ;
	    RECT 266.9000 94.4000 267.5000 131.6000 ;
	    RECT 268.4000 104.2000 269.2000 115.8000 ;
	    RECT 270.1000 112.4000 270.7000 133.6000 ;
	    RECT 273.2000 128.3000 274.0000 128.4000 ;
	    RECT 273.2000 127.7000 275.5000 128.3000 ;
	    RECT 273.2000 127.6000 274.0000 127.7000 ;
	    RECT 270.0000 111.6000 270.8000 112.4000 ;
	    RECT 271.6000 111.6000 272.4000 112.4000 ;
	    RECT 270.0000 105.6000 270.8000 106.4000 ;
	    RECT 270.1000 94.4000 270.7000 105.6000 ;
	    RECT 271.7000 98.4000 272.3000 111.6000 ;
	    RECT 274.9000 110.4000 275.5000 127.7000 ;
	    RECT 278.0000 127.6000 278.8000 128.4000 ;
	    RECT 281.3000 128.3000 281.9000 139.6000 ;
	    RECT 282.8000 137.6000 283.6000 138.4000 ;
	    RECT 282.9000 134.4000 283.5000 137.6000 ;
	    RECT 282.8000 133.6000 283.6000 134.4000 ;
	    RECT 282.9000 130.4000 283.5000 133.6000 ;
	    RECT 284.5000 132.4000 285.1000 149.6000 ;
	    RECT 286.1000 144.4000 286.7000 167.6000 ;
	    RECT 290.9000 152.4000 291.5000 173.7000 ;
	    RECT 297.3000 172.4000 297.9000 185.6000 ;
	    RECT 305.2000 179.6000 306.0000 180.4000 ;
	    RECT 298.8000 173.6000 299.6000 174.4000 ;
	    RECT 297.2000 171.6000 298.0000 172.4000 ;
	    RECT 300.4000 170.2000 301.2000 175.8000 ;
	    RECT 292.4000 167.6000 293.2000 168.4000 ;
	    RECT 292.5000 164.4000 293.1000 167.6000 ;
	    RECT 303.6000 166.2000 304.4000 177.8000 ;
	    RECT 305.3000 172.6000 305.9000 179.6000 ;
	    RECT 305.2000 171.8000 306.0000 172.6000 ;
	    RECT 292.4000 163.6000 293.2000 164.4000 ;
	    RECT 302.0000 163.6000 302.8000 164.4000 ;
	    RECT 290.8000 151.6000 291.6000 152.4000 ;
	    RECT 287.6000 149.6000 288.4000 150.4000 ;
	    RECT 289.2000 149.6000 290.0000 150.4000 ;
	    RECT 292.5000 150.3000 293.1000 163.6000 ;
	    RECT 302.1000 156.4000 302.7000 163.6000 ;
	    RECT 294.0000 155.6000 294.8000 156.4000 ;
	    RECT 295.6000 155.6000 296.4000 156.4000 ;
	    RECT 302.0000 155.6000 302.8000 156.4000 ;
	    RECT 303.6000 155.6000 304.4000 156.4000 ;
	    RECT 295.7000 154.3000 296.3000 155.6000 ;
	    RECT 294.1000 153.7000 296.3000 154.3000 ;
	    RECT 294.1000 150.4000 294.7000 153.7000 ;
	    RECT 295.6000 151.6000 296.4000 152.4000 ;
	    RECT 300.4000 151.6000 301.2000 152.4000 ;
	    RECT 290.9000 149.7000 293.1000 150.3000 ;
	    RECT 287.6000 147.6000 288.4000 148.4000 ;
	    RECT 286.0000 143.6000 286.8000 144.4000 ;
	    RECT 287.6000 143.6000 288.4000 144.4000 ;
	    RECT 287.7000 140.4000 288.3000 143.6000 ;
	    RECT 289.3000 142.4000 289.9000 149.6000 ;
	    RECT 290.9000 146.4000 291.5000 149.7000 ;
	    RECT 294.0000 149.6000 294.8000 150.4000 ;
	    RECT 292.4000 147.6000 293.2000 148.4000 ;
	    RECT 294.0000 147.6000 294.8000 148.4000 ;
	    RECT 290.8000 145.6000 291.6000 146.4000 ;
	    RECT 292.5000 142.4000 293.1000 147.6000 ;
	    RECT 289.2000 141.6000 290.0000 142.4000 ;
	    RECT 292.4000 141.6000 293.2000 142.4000 ;
	    RECT 287.6000 139.6000 288.4000 140.4000 ;
	    RECT 287.7000 136.4000 288.3000 139.6000 ;
	    RECT 287.6000 135.6000 288.4000 136.4000 ;
	    RECT 289.3000 132.4000 289.9000 141.6000 ;
	    RECT 292.4000 139.6000 293.2000 140.4000 ;
	    RECT 292.5000 136.4000 293.1000 139.6000 ;
	    RECT 292.4000 135.6000 293.2000 136.4000 ;
	    RECT 294.1000 134.4000 294.7000 147.6000 ;
	    RECT 295.7000 142.4000 296.3000 151.6000 ;
	    RECT 297.2000 149.6000 298.0000 150.4000 ;
	    RECT 300.5000 148.4000 301.1000 151.6000 ;
	    RECT 298.8000 147.6000 299.6000 148.4000 ;
	    RECT 300.4000 147.6000 301.2000 148.4000 ;
	    RECT 295.6000 141.6000 296.4000 142.4000 ;
	    RECT 297.2000 141.6000 298.0000 142.4000 ;
	    RECT 295.6000 139.6000 296.4000 140.4000 ;
	    RECT 294.0000 133.6000 294.8000 134.4000 ;
	    RECT 295.7000 132.4000 296.3000 139.6000 ;
	    RECT 297.3000 134.4000 297.9000 141.6000 ;
	    RECT 297.2000 133.6000 298.0000 134.4000 ;
	    RECT 298.9000 132.4000 299.5000 147.6000 ;
	    RECT 300.4000 133.6000 301.2000 134.4000 ;
	    RECT 302.1000 132.4000 302.7000 155.6000 ;
	    RECT 303.7000 136.4000 304.3000 155.6000 ;
	    RECT 306.8000 151.6000 307.6000 152.4000 ;
	    RECT 308.5000 152.3000 309.1000 187.6000 ;
	    RECT 310.1000 170.4000 310.7000 209.6000 ;
	    RECT 321.2000 207.6000 322.0000 208.4000 ;
	    RECT 311.6000 205.6000 312.4000 206.4000 ;
	    RECT 326.1000 198.4000 326.7000 213.7000 ;
	    RECT 327.6000 205.6000 328.4000 206.4000 ;
	    RECT 332.4000 206.2000 333.2000 217.8000 ;
	    RECT 338.9000 214.4000 339.5000 227.6000 ;
	    RECT 340.4000 224.2000 341.2000 235.8000 ;
	    RECT 343.6000 226.2000 344.4000 231.8000 ;
	    RECT 345.3000 228.4000 345.9000 237.6000 ;
	    RECT 346.9000 230.4000 347.5000 243.6000 ;
	    RECT 351.6000 231.6000 352.4000 232.4000 ;
	    RECT 346.8000 229.6000 347.6000 230.4000 ;
	    RECT 348.4000 229.6000 349.2000 230.4000 ;
	    RECT 345.2000 227.6000 346.0000 228.4000 ;
	    RECT 338.8000 213.6000 339.6000 214.4000 ;
	    RECT 340.4000 211.8000 341.2000 212.6000 ;
	    RECT 340.5000 210.4000 341.1000 211.8000 ;
	    RECT 340.4000 209.6000 341.2000 210.4000 ;
	    RECT 338.8000 207.6000 339.6000 208.4000 ;
	    RECT 319.6000 197.6000 320.4000 198.4000 ;
	    RECT 326.0000 197.6000 326.8000 198.4000 ;
	    RECT 311.6000 191.6000 312.4000 192.4000 ;
	    RECT 316.4000 192.3000 317.2000 192.4000 ;
	    RECT 316.4000 191.7000 318.7000 192.3000 ;
	    RECT 316.4000 191.6000 317.2000 191.7000 ;
	    RECT 311.7000 190.4000 312.3000 191.6000 ;
	    RECT 318.1000 190.4000 318.7000 191.7000 ;
	    RECT 311.6000 189.6000 312.4000 190.4000 ;
	    RECT 316.4000 189.6000 317.2000 190.4000 ;
	    RECT 318.0000 189.6000 318.8000 190.4000 ;
	    RECT 314.8000 187.6000 315.6000 188.4000 ;
	    RECT 311.6000 171.6000 312.4000 172.4000 ;
	    RECT 311.7000 170.4000 312.3000 171.6000 ;
	    RECT 310.0000 169.6000 310.8000 170.4000 ;
	    RECT 311.6000 169.6000 312.4000 170.4000 ;
	    RECT 311.7000 158.4000 312.3000 169.6000 ;
	    RECT 313.2000 166.2000 314.0000 177.8000 ;
	    RECT 314.9000 160.3000 315.5000 187.6000 ;
	    RECT 316.5000 178.4000 317.1000 189.6000 ;
	    RECT 318.0000 187.6000 318.8000 188.4000 ;
	    RECT 324.4000 184.2000 325.2000 195.8000 ;
	    RECT 327.7000 184.4000 328.3000 205.6000 ;
	    RECT 338.9000 198.4000 339.5000 207.6000 ;
	    RECT 342.0000 206.2000 342.8000 217.8000 ;
	    RECT 346.9000 216.3000 347.5000 229.6000 ;
	    RECT 351.7000 226.4000 352.3000 231.6000 ;
	    RECT 354.9000 230.4000 355.5000 249.7000 ;
	    RECT 356.4000 249.6000 357.2000 250.4000 ;
	    RECT 359.6000 246.2000 360.4000 257.8000 ;
	    RECT 361.3000 254.4000 361.9000 269.6000 ;
	    RECT 362.9000 268.4000 363.5000 295.6000 ;
	    RECT 364.4000 286.2000 365.2000 297.8000 ;
	    RECT 366.1000 296.4000 366.7000 331.6000 ;
	    RECT 369.2000 327.6000 370.0000 328.4000 ;
	    RECT 374.0000 326.2000 374.8000 337.8000 ;
	    RECT 378.8000 333.6000 379.6000 334.4000 ;
	    RECT 378.9000 314.4000 379.5000 333.6000 ;
	    RECT 382.0000 331.8000 382.8000 332.6000 ;
	    RECT 382.1000 330.4000 382.7000 331.8000 ;
	    RECT 382.0000 329.6000 382.8000 330.4000 ;
	    RECT 383.6000 326.2000 384.4000 337.8000 ;
	    RECT 430.0000 337.6000 430.8000 338.4000 ;
	    RECT 439.6000 337.6000 440.4000 338.4000 ;
	    RECT 430.1000 336.4000 430.7000 337.6000 ;
	    RECT 386.8000 330.2000 387.6000 335.8000 ;
	    RECT 388.4000 335.6000 389.2000 336.4000 ;
	    RECT 430.0000 335.6000 430.8000 336.4000 ;
	    RECT 388.5000 328.4000 389.1000 335.6000 ;
	    RECT 438.0000 333.6000 438.8000 334.4000 ;
	    RECT 393.2000 331.6000 394.0000 332.4000 ;
	    RECT 399.6000 331.6000 400.4000 332.4000 ;
	    RECT 412.4000 331.6000 413.2000 332.4000 ;
	    RECT 418.8000 331.6000 419.6000 332.4000 ;
	    RECT 425.2000 331.6000 426.0000 332.4000 ;
	    RECT 434.8000 331.6000 435.6000 332.4000 ;
	    RECT 393.2000 329.6000 394.0000 330.4000 ;
	    RECT 396.4000 329.6000 397.2000 330.4000 ;
	    RECT 388.4000 327.6000 389.2000 328.4000 ;
	    RECT 398.0000 327.6000 398.8000 328.4000 ;
	    RECT 396.4000 325.6000 397.2000 326.4000 ;
	    RECT 374.0000 313.6000 374.8000 314.4000 ;
	    RECT 378.8000 313.6000 379.6000 314.4000 ;
	    RECT 367.6000 311.6000 368.4000 312.4000 ;
	    RECT 367.7000 310.4000 368.3000 311.6000 ;
	    RECT 367.6000 309.6000 368.4000 310.4000 ;
	    RECT 372.4000 309.6000 373.2000 310.4000 ;
	    RECT 367.6000 307.6000 368.4000 308.4000 ;
	    RECT 372.5000 306.3000 373.1000 309.6000 ;
	    RECT 374.1000 308.4000 374.7000 313.6000 ;
	    RECT 374.0000 307.6000 374.8000 308.4000 ;
	    RECT 372.5000 305.7000 374.7000 306.3000 ;
	    RECT 369.2000 299.6000 370.0000 300.4000 ;
	    RECT 366.0000 295.6000 366.8000 296.4000 ;
	    RECT 366.0000 293.6000 366.8000 294.4000 ;
	    RECT 364.4000 269.6000 365.2000 270.4000 ;
	    RECT 364.5000 268.4000 365.1000 269.6000 ;
	    RECT 362.8000 267.6000 363.6000 268.4000 ;
	    RECT 364.4000 267.6000 365.2000 268.4000 ;
	    RECT 366.1000 254.4000 366.7000 293.6000 ;
	    RECT 367.6000 290.2000 368.4000 295.8000 ;
	    RECT 369.3000 294.4000 369.9000 299.6000 ;
	    RECT 369.2000 293.6000 370.0000 294.4000 ;
	    RECT 372.4000 289.6000 373.2000 290.4000 ;
	    RECT 374.1000 272.4000 374.7000 305.7000 ;
	    RECT 375.6000 303.6000 376.4000 304.4000 ;
	    RECT 380.4000 304.2000 381.2000 315.8000 ;
	    RECT 388.4000 309.4000 389.2000 310.4000 ;
	    RECT 390.0000 304.2000 390.8000 315.8000 ;
	    RECT 391.6000 307.6000 392.4000 308.4000 ;
	    RECT 375.7000 298.4000 376.3000 303.6000 ;
	    RECT 375.6000 297.6000 376.4000 298.4000 ;
	    RECT 378.8000 295.6000 379.6000 296.4000 ;
	    RECT 378.9000 294.4000 379.5000 295.6000 ;
	    RECT 378.8000 293.6000 379.6000 294.4000 ;
	    RECT 375.6000 291.6000 376.4000 292.4000 ;
	    RECT 378.8000 291.6000 379.6000 292.4000 ;
	    RECT 378.9000 290.4000 379.5000 291.6000 ;
	    RECT 378.8000 289.6000 379.6000 290.4000 ;
	    RECT 378.9000 276.4000 379.5000 289.6000 ;
	    RECT 380.4000 285.6000 381.2000 286.4000 ;
	    RECT 388.4000 286.2000 389.2000 297.8000 ;
	    RECT 391.7000 294.4000 392.3000 307.6000 ;
	    RECT 393.2000 306.2000 394.0000 311.8000 ;
	    RECT 396.5000 310.4000 397.1000 325.6000 ;
	    RECT 398.1000 314.4000 398.7000 327.6000 ;
	    RECT 399.7000 326.4000 400.3000 331.6000 ;
	    RECT 401.2000 327.6000 402.0000 328.4000 ;
	    RECT 412.5000 326.4000 413.1000 331.6000 ;
	    RECT 415.6000 329.6000 416.4000 330.4000 ;
	    RECT 430.0000 329.6000 430.8000 330.4000 ;
	    RECT 414.0000 327.6000 414.8000 328.4000 ;
	    RECT 417.2000 327.6000 418.0000 328.4000 ;
	    RECT 425.2000 327.6000 426.0000 328.4000 ;
	    RECT 426.8000 327.6000 427.6000 328.4000 ;
	    RECT 399.6000 325.6000 400.4000 326.4000 ;
	    RECT 412.4000 325.6000 413.2000 326.4000 ;
	    RECT 399.6000 323.6000 400.4000 324.4000 ;
	    RECT 399.7000 322.4000 400.3000 323.6000 ;
	    RECT 399.6000 321.6000 400.4000 322.4000 ;
	    RECT 399.6000 319.6000 400.4000 320.4000 ;
	    RECT 399.7000 318.4000 400.3000 319.6000 ;
	    RECT 399.6000 317.6000 400.4000 318.4000 ;
	    RECT 398.0000 313.6000 398.8000 314.4000 ;
	    RECT 399.6000 313.6000 400.4000 314.4000 ;
	    RECT 407.6000 313.6000 408.4000 314.4000 ;
	    RECT 396.4000 309.6000 397.2000 310.4000 ;
	    RECT 391.6000 293.6000 392.4000 294.4000 ;
	    RECT 394.8000 293.6000 395.6000 294.4000 ;
	    RECT 394.9000 286.4000 395.5000 293.6000 ;
	    RECT 396.4000 291.8000 397.2000 292.6000 ;
	    RECT 394.8000 285.6000 395.6000 286.4000 ;
	    RECT 383.6000 283.6000 384.4000 284.4000 ;
	    RECT 383.7000 282.4000 384.3000 283.6000 ;
	    RECT 383.6000 281.6000 384.4000 282.4000 ;
	    RECT 391.6000 281.6000 392.4000 282.4000 ;
	    RECT 378.8000 275.6000 379.6000 276.4000 ;
	    RECT 390.0000 275.6000 390.8000 276.4000 ;
	    RECT 375.6000 273.6000 376.4000 274.4000 ;
	    RECT 367.6000 271.6000 368.4000 272.4000 ;
	    RECT 374.0000 271.6000 374.8000 272.4000 ;
	    RECT 367.7000 268.4000 368.3000 271.6000 ;
	    RECT 372.4000 269.6000 373.2000 270.4000 ;
	    RECT 374.0000 269.6000 374.8000 270.4000 ;
	    RECT 378.8000 269.6000 379.6000 270.4000 ;
	    RECT 380.4000 269.6000 381.2000 270.4000 ;
	    RECT 388.4000 269.6000 389.2000 270.4000 ;
	    RECT 372.5000 268.4000 373.1000 269.6000 ;
	    RECT 374.1000 268.4000 374.7000 269.6000 ;
	    RECT 367.6000 267.6000 368.4000 268.4000 ;
	    RECT 372.4000 267.6000 373.2000 268.4000 ;
	    RECT 374.0000 267.6000 374.8000 268.4000 ;
	    RECT 374.0000 265.6000 374.8000 266.4000 ;
	    RECT 369.2000 263.6000 370.0000 264.4000 ;
	    RECT 369.3000 260.3000 369.9000 263.6000 ;
	    RECT 374.1000 260.4000 374.7000 265.6000 ;
	    RECT 378.9000 260.4000 379.5000 269.6000 ;
	    RECT 367.7000 259.7000 369.9000 260.3000 ;
	    RECT 361.2000 253.6000 362.0000 254.4000 ;
	    RECT 366.0000 253.6000 366.8000 254.4000 ;
	    RECT 367.7000 252.6000 368.3000 259.7000 ;
	    RECT 374.0000 259.6000 374.8000 260.4000 ;
	    RECT 378.8000 259.6000 379.6000 260.4000 ;
	    RECT 374.1000 258.4000 374.7000 259.6000 ;
	    RECT 367.6000 251.8000 368.4000 252.6000 ;
	    RECT 361.2000 249.6000 362.0000 250.4000 ;
	    RECT 356.4000 239.6000 357.2000 240.4000 ;
	    RECT 354.8000 229.6000 355.6000 230.4000 ;
	    RECT 356.5000 228.4000 357.1000 239.6000 ;
	    RECT 361.3000 238.4000 361.9000 249.6000 ;
	    RECT 369.2000 246.2000 370.0000 257.8000 ;
	    RECT 374.0000 257.6000 374.8000 258.4000 ;
	    RECT 370.8000 253.6000 371.6000 254.4000 ;
	    RECT 370.9000 250.4000 371.5000 253.6000 ;
	    RECT 370.8000 249.6000 371.6000 250.4000 ;
	    RECT 372.4000 250.2000 373.2000 255.8000 ;
	    RECT 361.2000 237.6000 362.0000 238.4000 ;
	    RECT 366.0000 231.6000 366.8000 232.4000 ;
	    RECT 358.0000 229.6000 358.8000 230.4000 ;
	    RECT 356.4000 227.6000 357.2000 228.4000 ;
	    RECT 351.6000 225.6000 352.4000 226.4000 ;
	    RECT 350.0000 221.6000 350.8000 222.4000 ;
	    RECT 345.2000 210.2000 346.0000 215.8000 ;
	    RECT 346.9000 215.7000 349.1000 216.3000 ;
	    RECT 346.8000 213.6000 347.6000 214.4000 ;
	    RECT 348.5000 212.4000 349.1000 215.7000 ;
	    RECT 350.1000 214.4000 350.7000 221.6000 ;
	    RECT 350.0000 213.6000 350.8000 214.4000 ;
	    RECT 356.5000 214.3000 357.1000 227.6000 ;
	    RECT 358.1000 216.3000 358.7000 229.6000 ;
	    RECT 362.8000 223.6000 363.6000 224.4000 ;
	    RECT 361.2000 221.6000 362.0000 222.4000 ;
	    RECT 359.6000 219.6000 360.4000 220.4000 ;
	    RECT 359.7000 218.4000 360.3000 219.6000 ;
	    RECT 359.6000 217.6000 360.4000 218.4000 ;
	    RECT 358.1000 215.7000 360.3000 216.3000 ;
	    RECT 358.0000 214.3000 358.8000 214.4000 ;
	    RECT 356.5000 213.7000 358.8000 214.3000 ;
	    RECT 358.0000 213.6000 358.8000 213.7000 ;
	    RECT 348.4000 212.3000 349.2000 212.4000 ;
	    RECT 348.4000 211.7000 350.7000 212.3000 ;
	    RECT 348.4000 211.6000 349.2000 211.7000 ;
	    RECT 348.4000 209.6000 349.2000 210.4000 ;
	    RECT 343.6000 203.6000 344.4000 204.4000 ;
	    RECT 338.8000 197.6000 339.6000 198.4000 ;
	    RECT 330.8000 189.6000 331.6000 190.4000 ;
	    RECT 329.2000 187.6000 330.0000 188.4000 ;
	    RECT 329.3000 184.4000 329.9000 187.6000 ;
	    RECT 332.4000 185.6000 333.2000 186.4000 ;
	    RECT 327.6000 183.6000 328.4000 184.4000 ;
	    RECT 329.2000 183.6000 330.0000 184.4000 ;
	    RECT 319.6000 179.6000 320.4000 180.4000 ;
	    RECT 316.4000 177.6000 317.2000 178.4000 ;
	    RECT 318.0000 164.3000 318.8000 164.4000 ;
	    RECT 316.5000 163.7000 318.8000 164.3000 ;
	    RECT 316.5000 162.4000 317.1000 163.7000 ;
	    RECT 318.0000 163.6000 318.8000 163.7000 ;
	    RECT 316.4000 161.6000 317.2000 162.4000 ;
	    RECT 314.9000 159.7000 317.1000 160.3000 ;
	    RECT 311.6000 157.6000 312.4000 158.4000 ;
	    RECT 314.8000 157.6000 315.6000 158.4000 ;
	    RECT 310.0000 154.3000 310.8000 154.4000 ;
	    RECT 310.0000 153.7000 313.9000 154.3000 ;
	    RECT 310.0000 153.6000 310.8000 153.7000 ;
	    RECT 308.5000 151.7000 312.3000 152.3000 ;
	    RECT 305.2000 149.6000 306.0000 150.4000 ;
	    RECT 306.9000 148.4000 307.5000 151.6000 ;
	    RECT 308.5000 150.4000 309.1000 151.7000 ;
	    RECT 308.4000 149.6000 309.2000 150.4000 ;
	    RECT 310.0000 149.6000 310.8000 150.4000 ;
	    RECT 305.2000 147.6000 306.0000 148.4000 ;
	    RECT 306.8000 147.6000 307.6000 148.4000 ;
	    RECT 305.3000 138.4000 305.9000 147.6000 ;
	    RECT 305.2000 137.6000 306.0000 138.4000 ;
	    RECT 303.6000 135.6000 304.4000 136.4000 ;
	    RECT 305.2000 135.6000 306.0000 136.4000 ;
	    RECT 305.2000 133.6000 306.0000 134.4000 ;
	    RECT 284.4000 131.6000 285.2000 132.4000 ;
	    RECT 289.2000 131.6000 290.0000 132.4000 ;
	    RECT 295.6000 131.6000 296.4000 132.4000 ;
	    RECT 297.2000 131.6000 298.0000 132.4000 ;
	    RECT 298.8000 131.6000 299.6000 132.4000 ;
	    RECT 300.4000 131.6000 301.2000 132.4000 ;
	    RECT 302.0000 131.6000 302.8000 132.4000 ;
	    RECT 282.8000 129.6000 283.6000 130.4000 ;
	    RECT 284.5000 128.4000 285.1000 131.6000 ;
	    RECT 287.6000 129.6000 288.4000 130.4000 ;
	    RECT 290.8000 129.6000 291.6000 130.4000 ;
	    RECT 298.8000 129.6000 299.6000 130.4000 ;
	    RECT 300.5000 130.3000 301.1000 131.6000 ;
	    RECT 306.9000 130.4000 307.5000 147.6000 ;
	    RECT 310.1000 132.4000 310.7000 149.6000 ;
	    RECT 311.7000 148.4000 312.3000 151.7000 ;
	    RECT 313.3000 148.4000 313.9000 153.7000 ;
	    RECT 314.9000 150.4000 315.5000 157.6000 ;
	    RECT 314.8000 149.6000 315.6000 150.4000 ;
	    RECT 311.6000 147.6000 312.4000 148.4000 ;
	    RECT 313.2000 147.6000 314.0000 148.4000 ;
	    RECT 311.6000 139.6000 312.4000 140.4000 ;
	    RECT 313.2000 139.6000 314.0000 140.4000 ;
	    RECT 311.7000 134.4000 312.3000 139.6000 ;
	    RECT 313.3000 136.4000 313.9000 139.6000 ;
	    RECT 316.5000 138.3000 317.1000 159.7000 ;
	    RECT 318.0000 150.3000 318.8000 150.4000 ;
	    RECT 319.7000 150.3000 320.3000 179.6000 ;
	    RECT 329.3000 174.4000 329.9000 183.6000 ;
	    RECT 329.2000 173.6000 330.0000 174.4000 ;
	    RECT 322.8000 171.6000 323.6000 172.4000 ;
	    RECT 322.9000 164.4000 323.5000 171.6000 ;
	    RECT 332.5000 170.4000 333.1000 185.6000 ;
	    RECT 334.0000 184.2000 334.8000 195.8000 ;
	    RECT 337.2000 186.2000 338.0000 191.8000 ;
	    RECT 338.9000 190.4000 339.5000 197.6000 ;
	    RECT 343.7000 190.4000 344.3000 203.6000 ;
	    RECT 345.2000 199.6000 346.0000 200.4000 ;
	    RECT 338.8000 189.6000 339.6000 190.4000 ;
	    RECT 343.6000 189.6000 344.4000 190.4000 ;
	    RECT 342.0000 183.6000 342.8000 184.4000 ;
	    RECT 335.6000 181.6000 336.4000 182.4000 ;
	    RECT 338.8000 181.6000 339.6000 182.4000 ;
	    RECT 335.7000 178.4000 336.3000 181.6000 ;
	    RECT 335.6000 177.6000 336.4000 178.4000 ;
	    RECT 334.0000 173.6000 334.8000 174.4000 ;
	    RECT 334.1000 172.4000 334.7000 173.6000 ;
	    RECT 338.9000 172.4000 339.5000 181.6000 ;
	    RECT 342.1000 178.4000 342.7000 183.6000 ;
	    RECT 342.0000 177.6000 342.8000 178.4000 ;
	    RECT 343.6000 173.6000 344.4000 174.4000 ;
	    RECT 343.7000 172.4000 344.3000 173.6000 ;
	    RECT 334.0000 171.6000 334.8000 172.4000 ;
	    RECT 338.8000 171.6000 339.6000 172.4000 ;
	    RECT 340.4000 171.6000 341.2000 172.4000 ;
	    RECT 343.6000 172.3000 344.4000 172.4000 ;
	    RECT 345.3000 172.3000 345.9000 199.6000 ;
	    RECT 346.8000 193.6000 347.6000 194.4000 ;
	    RECT 348.4000 189.6000 349.2000 190.4000 ;
	    RECT 346.8000 179.6000 347.6000 180.4000 ;
	    RECT 346.9000 178.4000 347.5000 179.6000 ;
	    RECT 346.8000 177.6000 347.6000 178.4000 ;
	    RECT 348.5000 176.4000 349.1000 189.6000 ;
	    RECT 350.1000 186.4000 350.7000 211.7000 ;
	    RECT 356.4000 211.6000 357.2000 212.4000 ;
	    RECT 353.2000 207.6000 354.0000 208.4000 ;
	    RECT 353.3000 206.4000 353.9000 207.6000 ;
	    RECT 356.5000 206.4000 357.1000 211.6000 ;
	    RECT 353.2000 205.6000 354.0000 206.4000 ;
	    RECT 356.4000 205.6000 357.2000 206.4000 ;
	    RECT 356.4000 201.6000 357.2000 202.4000 ;
	    RECT 351.6000 197.6000 352.4000 198.4000 ;
	    RECT 356.5000 194.4000 357.1000 201.6000 ;
	    RECT 358.1000 198.4000 358.7000 213.6000 ;
	    RECT 358.0000 197.6000 358.8000 198.4000 ;
	    RECT 359.7000 196.4000 360.3000 215.7000 ;
	    RECT 359.6000 195.6000 360.4000 196.4000 ;
	    RECT 356.4000 193.6000 357.2000 194.4000 ;
	    RECT 356.5000 192.4000 357.1000 193.6000 ;
	    RECT 356.4000 191.6000 357.2000 192.4000 ;
	    RECT 353.2000 189.6000 354.0000 190.4000 ;
	    RECT 353.3000 188.4000 353.9000 189.6000 ;
	    RECT 353.2000 187.6000 354.0000 188.4000 ;
	    RECT 359.6000 187.6000 360.4000 188.4000 ;
	    RECT 350.0000 185.6000 350.8000 186.4000 ;
	    RECT 353.3000 182.4000 353.9000 187.6000 ;
	    RECT 350.0000 181.6000 350.8000 182.4000 ;
	    RECT 353.2000 181.6000 354.0000 182.4000 ;
	    RECT 348.4000 175.6000 349.2000 176.4000 ;
	    RECT 343.6000 171.7000 345.9000 172.3000 ;
	    RECT 348.4000 172.3000 349.2000 172.4000 ;
	    RECT 350.1000 172.3000 350.7000 181.6000 ;
	    RECT 361.3000 180.4000 361.9000 221.6000 ;
	    RECT 364.4000 219.6000 365.2000 220.4000 ;
	    RECT 364.5000 218.4000 365.1000 219.6000 ;
	    RECT 364.4000 217.6000 365.2000 218.4000 ;
	    RECT 364.5000 216.4000 365.1000 217.6000 ;
	    RECT 366.1000 216.4000 366.7000 231.6000 ;
	    RECT 367.6000 224.2000 368.4000 235.8000 ;
	    RECT 370.9000 230.4000 371.5000 249.6000 ;
	    RECT 378.8000 246.2000 379.6000 257.8000 ;
	    RECT 380.5000 244.4000 381.1000 269.6000 ;
	    RECT 383.6000 268.3000 384.4000 268.4000 ;
	    RECT 382.1000 267.7000 384.4000 268.3000 ;
	    RECT 380.4000 243.6000 381.2000 244.4000 ;
	    RECT 382.1000 240.4000 382.7000 267.7000 ;
	    RECT 383.6000 267.6000 384.4000 267.7000 ;
	    RECT 385.2000 265.6000 386.0000 266.4000 ;
	    RECT 385.3000 262.4000 385.9000 265.6000 ;
	    RECT 388.5000 262.4000 389.1000 269.6000 ;
	    RECT 385.2000 261.6000 386.0000 262.4000 ;
	    RECT 388.4000 261.6000 389.2000 262.4000 ;
	    RECT 386.8000 255.6000 387.6000 256.4000 ;
	    RECT 383.6000 253.6000 384.4000 254.4000 ;
	    RECT 383.7000 250.4000 384.3000 253.6000 ;
	    RECT 386.9000 252.6000 387.5000 255.6000 ;
	    RECT 386.8000 251.8000 387.6000 252.6000 ;
	    RECT 383.6000 249.6000 384.4000 250.4000 ;
	    RECT 388.4000 246.2000 389.2000 257.8000 ;
	    RECT 390.1000 248.3000 390.7000 275.6000 ;
	    RECT 391.7000 274.4000 392.3000 281.6000 ;
	    RECT 396.5000 278.4000 397.1000 291.8000 ;
	    RECT 398.0000 286.2000 398.8000 297.8000 ;
	    RECT 396.4000 277.6000 397.2000 278.4000 ;
	    RECT 391.6000 273.6000 392.4000 274.4000 ;
	    RECT 393.2000 273.6000 394.0000 274.4000 ;
	    RECT 393.3000 258.4000 393.9000 273.6000 ;
	    RECT 399.7000 270.4000 400.3000 313.6000 ;
	    RECT 407.7000 312.4000 408.3000 313.6000 ;
	    RECT 407.6000 311.6000 408.4000 312.4000 ;
	    RECT 402.8000 309.6000 403.6000 310.4000 ;
	    RECT 402.9000 298.4000 403.5000 309.6000 ;
	    RECT 412.4000 304.2000 413.2000 315.8000 ;
	    RECT 415.6000 313.6000 416.4000 314.4000 ;
	    RECT 402.8000 297.6000 403.6000 298.4000 ;
	    RECT 401.2000 290.2000 402.0000 295.8000 ;
	    RECT 415.7000 294.4000 416.3000 313.6000 ;
	    RECT 417.3000 300.4000 417.9000 327.6000 ;
	    RECT 420.5000 310.2000 421.1000 310.3000 ;
	    RECT 420.4000 309.4000 421.2000 310.2000 ;
	    RECT 418.8000 307.6000 419.6000 308.4000 ;
	    RECT 417.2000 299.6000 418.0000 300.4000 ;
	    RECT 407.6000 293.6000 408.4000 294.4000 ;
	    RECT 415.6000 293.6000 416.4000 294.4000 ;
	    RECT 406.0000 291.6000 406.8000 292.4000 ;
	    RECT 402.8000 289.6000 403.6000 290.4000 ;
	    RECT 402.9000 278.3000 403.5000 289.6000 ;
	    RECT 406.1000 284.4000 406.7000 291.6000 ;
	    RECT 407.7000 288.4000 408.3000 293.6000 ;
	    RECT 407.6000 287.6000 408.4000 288.4000 ;
	    RECT 407.7000 284.4000 408.3000 287.6000 ;
	    RECT 418.9000 286.4000 419.5000 307.6000 ;
	    RECT 420.5000 298.4000 421.1000 309.4000 ;
	    RECT 422.0000 304.2000 422.8000 315.8000 ;
	    RECT 425.3000 314.3000 425.9000 327.6000 ;
	    RECT 434.9000 322.4000 435.5000 331.6000 ;
	    RECT 438.0000 329.6000 438.8000 330.4000 ;
	    RECT 444.4000 326.2000 445.2000 337.8000 ;
	    RECT 450.8000 333.6000 451.6000 334.4000 ;
	    RECT 452.4000 333.6000 453.2000 334.4000 ;
	    RECT 450.9000 332.4000 451.5000 333.6000 ;
	    RECT 450.8000 331.6000 451.6000 332.4000 ;
	    RECT 431.6000 321.6000 432.4000 322.4000 ;
	    RECT 434.8000 321.6000 435.6000 322.4000 ;
	    RECT 425.3000 313.7000 427.5000 314.3000 ;
	    RECT 426.9000 312.4000 427.5000 313.7000 ;
	    RECT 425.2000 306.2000 426.0000 311.8000 ;
	    RECT 426.8000 311.6000 427.6000 312.4000 ;
	    RECT 428.4000 311.6000 429.2000 312.4000 ;
	    RECT 430.0000 311.6000 430.8000 312.4000 ;
	    RECT 420.4000 297.6000 421.2000 298.4000 ;
	    RECT 425.2000 293.6000 426.0000 294.4000 ;
	    RECT 426.8000 291.6000 427.6000 292.4000 ;
	    RECT 426.9000 290.4000 427.5000 291.6000 ;
	    RECT 420.4000 289.6000 421.2000 290.4000 ;
	    RECT 426.8000 289.6000 427.6000 290.4000 ;
	    RECT 420.5000 288.4000 421.1000 289.6000 ;
	    RECT 420.4000 287.6000 421.2000 288.4000 ;
	    RECT 418.8000 285.6000 419.6000 286.4000 ;
	    RECT 406.0000 283.6000 406.8000 284.4000 ;
	    RECT 407.6000 283.6000 408.4000 284.4000 ;
	    RECT 415.6000 283.6000 416.4000 284.4000 ;
	    RECT 422.0000 284.3000 422.8000 284.4000 ;
	    RECT 422.0000 283.7000 424.3000 284.3000 ;
	    RECT 422.0000 283.6000 422.8000 283.7000 ;
	    RECT 402.9000 277.7000 405.1000 278.3000 ;
	    RECT 402.8000 271.6000 403.6000 272.4000 ;
	    RECT 396.4000 269.6000 397.2000 270.4000 ;
	    RECT 399.6000 269.6000 400.4000 270.4000 ;
	    RECT 399.6000 267.6000 400.4000 268.4000 ;
	    RECT 399.7000 266.4000 400.3000 267.6000 ;
	    RECT 399.6000 265.6000 400.4000 266.4000 ;
	    RECT 393.2000 257.6000 394.0000 258.4000 ;
	    RECT 391.6000 250.2000 392.4000 255.8000 ;
	    RECT 390.1000 247.7000 392.3000 248.3000 ;
	    RECT 390.0000 243.6000 390.8000 244.4000 ;
	    RECT 382.0000 239.6000 382.8000 240.4000 ;
	    RECT 375.6000 231.6000 376.4000 232.4000 ;
	    RECT 370.8000 229.6000 371.6000 230.4000 ;
	    RECT 375.7000 230.2000 376.3000 231.6000 ;
	    RECT 364.4000 215.6000 365.2000 216.4000 ;
	    RECT 366.0000 215.6000 366.8000 216.4000 ;
	    RECT 362.8000 211.6000 363.6000 212.4000 ;
	    RECT 362.9000 204.4000 363.5000 211.6000 ;
	    RECT 369.2000 206.2000 370.0000 217.8000 ;
	    RECT 370.9000 212.4000 371.5000 229.6000 ;
	    RECT 375.6000 229.4000 376.4000 230.2000 ;
	    RECT 377.2000 224.2000 378.0000 235.8000 ;
	    RECT 390.1000 232.4000 390.7000 243.6000 ;
	    RECT 391.7000 238.4000 392.3000 247.7000 ;
	    RECT 398.0000 246.2000 398.8000 257.8000 ;
	    RECT 391.6000 237.6000 392.4000 238.4000 ;
	    RECT 402.9000 232.4000 403.5000 271.6000 ;
	    RECT 404.5000 270.4000 405.1000 277.7000 ;
	    RECT 414.0000 271.6000 414.8000 272.4000 ;
	    RECT 414.1000 270.4000 414.7000 271.6000 ;
	    RECT 404.4000 269.6000 405.2000 270.4000 ;
	    RECT 414.0000 269.6000 414.8000 270.4000 ;
	    RECT 415.7000 268.4000 416.3000 283.6000 ;
	    RECT 420.4000 275.6000 421.2000 276.4000 ;
	    RECT 417.2000 273.6000 418.0000 274.4000 ;
	    RECT 417.3000 268.4000 417.9000 273.6000 ;
	    RECT 420.5000 272.4000 421.1000 275.6000 ;
	    RECT 420.4000 271.6000 421.2000 272.4000 ;
	    RECT 422.0000 271.6000 422.8000 272.4000 ;
	    RECT 415.6000 267.6000 416.4000 268.4000 ;
	    RECT 417.2000 267.6000 418.0000 268.4000 ;
	    RECT 404.4000 263.6000 405.2000 264.4000 ;
	    RECT 418.8000 263.6000 419.6000 264.4000 ;
	    RECT 404.5000 256.4000 405.1000 263.6000 ;
	    RECT 404.4000 255.6000 405.2000 256.4000 ;
	    RECT 406.0000 251.8000 406.8000 252.6000 ;
	    RECT 406.1000 250.4000 406.7000 251.8000 ;
	    RECT 406.0000 249.6000 406.8000 250.4000 ;
	    RECT 407.6000 246.2000 408.4000 257.8000 ;
	    RECT 409.2000 255.6000 410.0000 256.4000 ;
	    RECT 418.9000 256.3000 419.5000 263.6000 ;
	    RECT 409.3000 254.4000 409.9000 255.6000 ;
	    RECT 409.2000 253.6000 410.0000 254.4000 ;
	    RECT 410.8000 250.2000 411.6000 255.8000 ;
	    RECT 417.3000 255.7000 419.5000 256.3000 ;
	    RECT 417.3000 250.4000 417.9000 255.7000 ;
	    RECT 418.8000 253.6000 419.6000 254.4000 ;
	    RECT 418.9000 250.4000 419.5000 253.6000 ;
	    RECT 420.5000 252.3000 421.1000 271.6000 ;
	    RECT 422.0000 269.6000 422.8000 270.4000 ;
	    RECT 423.7000 254.4000 424.3000 283.7000 ;
	    RECT 426.9000 276.4000 427.5000 289.6000 ;
	    RECT 426.8000 275.6000 427.6000 276.4000 ;
	    RECT 428.5000 272.4000 429.1000 311.6000 ;
	    RECT 430.1000 310.4000 430.7000 311.6000 ;
	    RECT 431.7000 310.4000 432.3000 321.6000 ;
	    RECT 434.8000 315.6000 435.6000 316.4000 ;
	    RECT 434.9000 314.4000 435.5000 315.6000 ;
	    RECT 434.8000 313.6000 435.6000 314.4000 ;
	    RECT 430.0000 309.6000 430.8000 310.4000 ;
	    RECT 431.6000 309.6000 432.4000 310.4000 ;
	    RECT 434.9000 306.4000 435.5000 313.6000 ;
	    RECT 434.8000 305.6000 435.6000 306.4000 ;
	    RECT 441.2000 304.2000 442.0000 315.8000 ;
	    RECT 446.0000 309.6000 446.8000 310.4000 ;
	    RECT 450.8000 304.2000 451.6000 315.8000 ;
	    RECT 452.5000 308.4000 453.1000 333.6000 ;
	    RECT 454.0000 326.2000 454.8000 337.8000 ;
	    RECT 457.2000 330.2000 458.0000 335.8000 ;
	    RECT 479.6000 335.6000 480.4000 336.4000 ;
	    RECT 462.0000 333.6000 462.8000 334.4000 ;
	    RECT 462.1000 332.4000 462.7000 333.6000 ;
	    RECT 462.0000 331.6000 462.8000 332.4000 ;
	    RECT 466.8000 331.6000 467.6000 332.4000 ;
	    RECT 473.2000 331.6000 474.0000 332.4000 ;
	    RECT 474.8000 331.6000 475.6000 332.4000 ;
	    RECT 458.8000 329.6000 459.6000 330.4000 ;
	    RECT 452.4000 307.6000 453.2000 308.4000 ;
	    RECT 436.4000 297.6000 437.2000 298.4000 ;
	    RECT 434.8000 296.3000 435.6000 296.4000 ;
	    RECT 436.5000 296.3000 437.1000 297.6000 ;
	    RECT 434.8000 295.7000 437.1000 296.3000 ;
	    RECT 434.8000 295.6000 435.6000 295.7000 ;
	    RECT 434.9000 294.4000 435.5000 295.6000 ;
	    RECT 431.6000 294.3000 432.4000 294.4000 ;
	    RECT 431.6000 293.7000 433.9000 294.3000 ;
	    RECT 431.6000 293.6000 432.4000 293.7000 ;
	    RECT 433.3000 292.3000 433.9000 293.7000 ;
	    RECT 434.8000 293.6000 435.6000 294.4000 ;
	    RECT 434.8000 292.3000 435.6000 292.4000 ;
	    RECT 433.3000 291.7000 435.6000 292.3000 ;
	    RECT 434.8000 291.6000 435.6000 291.7000 ;
	    RECT 431.6000 289.6000 432.4000 290.4000 ;
	    RECT 430.0000 287.6000 430.8000 288.4000 ;
	    RECT 428.4000 271.6000 429.2000 272.4000 ;
	    RECT 430.1000 270.4000 430.7000 287.6000 ;
	    RECT 434.8000 285.6000 435.6000 286.4000 ;
	    RECT 441.2000 286.2000 442.0000 297.8000 ;
	    RECT 444.4000 291.6000 445.2000 292.4000 ;
	    RECT 450.8000 286.2000 451.6000 297.8000 ;
	    RECT 452.5000 294.4000 453.1000 307.6000 ;
	    RECT 454.0000 306.2000 454.8000 311.8000 ;
	    RECT 462.1000 306.4000 462.7000 331.6000 ;
	    RECT 466.9000 326.4000 467.5000 331.6000 ;
	    RECT 471.6000 329.6000 472.4000 330.4000 ;
	    RECT 468.4000 327.6000 469.2000 328.4000 ;
	    RECT 466.8000 325.6000 467.6000 326.4000 ;
	    RECT 466.8000 321.6000 467.6000 322.4000 ;
	    RECT 457.2000 305.6000 458.0000 306.4000 ;
	    RECT 462.0000 305.6000 462.8000 306.4000 ;
	    RECT 455.6000 303.6000 456.4000 304.4000 ;
	    RECT 452.4000 293.6000 453.2000 294.4000 ;
	    RECT 454.0000 290.2000 454.8000 295.8000 ;
	    RECT 455.7000 294.4000 456.3000 303.6000 ;
	    RECT 455.6000 293.6000 456.4000 294.4000 ;
	    RECT 457.3000 292.4000 457.9000 305.6000 ;
	    RECT 458.8000 303.6000 459.6000 304.4000 ;
	    RECT 463.6000 304.2000 464.4000 315.8000 ;
	    RECT 465.2000 307.6000 466.0000 308.4000 ;
	    RECT 458.8000 299.6000 459.6000 300.4000 ;
	    RECT 457.2000 291.6000 458.0000 292.4000 ;
	    RECT 458.9000 288.4000 459.5000 299.6000 ;
	    RECT 462.0000 297.6000 462.8000 298.4000 ;
	    RECT 462.1000 296.4000 462.7000 297.6000 ;
	    RECT 462.0000 295.6000 462.8000 296.4000 ;
	    RECT 466.9000 292.4000 467.5000 321.6000 ;
	    RECT 466.8000 291.6000 467.6000 292.4000 ;
	    RECT 458.8000 287.6000 459.6000 288.4000 ;
	    RECT 462.0000 287.6000 462.8000 288.4000 ;
	    RECT 425.2000 269.6000 426.0000 270.4000 ;
	    RECT 430.0000 269.6000 430.8000 270.4000 ;
	    RECT 431.6000 269.6000 432.4000 270.4000 ;
	    RECT 425.3000 262.4000 425.9000 269.6000 ;
	    RECT 426.8000 267.6000 427.6000 268.4000 ;
	    RECT 426.9000 264.4000 427.5000 267.6000 ;
	    RECT 426.8000 263.6000 427.6000 264.4000 ;
	    RECT 431.7000 262.4000 432.3000 269.6000 ;
	    RECT 434.9000 268.4000 435.5000 285.6000 ;
	    RECT 457.2000 275.6000 458.0000 276.4000 ;
	    RECT 457.3000 274.4000 457.9000 275.6000 ;
	    RECT 458.9000 274.4000 459.5000 287.6000 ;
	    RECT 454.0000 273.6000 454.8000 274.4000 ;
	    RECT 457.2000 273.6000 458.0000 274.4000 ;
	    RECT 458.8000 273.6000 459.6000 274.4000 ;
	    RECT 462.0000 273.6000 462.8000 274.4000 ;
	    RECT 454.1000 272.4000 454.7000 273.6000 ;
	    RECT 454.0000 271.6000 454.8000 272.4000 ;
	    RECT 457.2000 271.6000 458.0000 272.4000 ;
	    RECT 457.3000 270.4000 457.9000 271.6000 ;
	    RECT 450.8000 269.6000 451.6000 270.4000 ;
	    RECT 457.2000 269.6000 458.0000 270.4000 ;
	    RECT 465.2000 269.6000 466.0000 270.4000 ;
	    RECT 433.2000 267.6000 434.0000 268.4000 ;
	    RECT 434.8000 267.6000 435.6000 268.4000 ;
	    RECT 449.2000 267.6000 450.0000 268.4000 ;
	    RECT 433.3000 264.4000 433.9000 267.6000 ;
	    RECT 433.2000 263.6000 434.0000 264.4000 ;
	    RECT 425.2000 261.6000 426.0000 262.4000 ;
	    RECT 431.6000 261.6000 432.4000 262.4000 ;
	    RECT 428.4000 257.6000 429.2000 258.4000 ;
	    RECT 428.5000 256.4000 429.1000 257.6000 ;
	    RECT 428.4000 255.6000 429.2000 256.4000 ;
	    RECT 423.6000 253.6000 424.4000 254.4000 ;
	    RECT 422.0000 252.3000 422.8000 252.4000 ;
	    RECT 420.5000 251.7000 422.8000 252.3000 ;
	    RECT 422.0000 251.6000 422.8000 251.7000 ;
	    RECT 417.2000 249.6000 418.0000 250.4000 ;
	    RECT 418.8000 249.6000 419.6000 250.4000 ;
	    RECT 428.5000 246.4000 429.1000 255.6000 ;
	    RECT 430.0000 249.6000 430.8000 250.4000 ;
	    RECT 428.4000 245.6000 429.2000 246.4000 ;
	    RECT 425.2000 243.6000 426.0000 244.4000 ;
	    RECT 425.3000 242.4000 425.9000 243.6000 ;
	    RECT 412.4000 241.6000 413.2000 242.4000 ;
	    RECT 425.2000 241.6000 426.0000 242.4000 ;
	    RECT 412.5000 238.4000 413.1000 241.6000 ;
	    RECT 412.4000 237.6000 413.2000 238.4000 ;
	    RECT 380.4000 226.2000 381.2000 231.8000 ;
	    RECT 386.8000 231.6000 387.6000 232.4000 ;
	    RECT 390.0000 231.6000 390.8000 232.4000 ;
	    RECT 399.6000 232.3000 400.4000 232.4000 ;
	    RECT 398.1000 231.7000 400.4000 232.3000 ;
	    RECT 386.8000 229.6000 387.6000 230.4000 ;
	    RECT 394.8000 229.6000 395.6000 230.4000 ;
	    RECT 382.0000 225.6000 382.8000 226.4000 ;
	    RECT 382.1000 224.4000 382.7000 225.6000 ;
	    RECT 382.0000 223.6000 382.8000 224.4000 ;
	    RECT 383.6000 219.6000 384.4000 220.4000 ;
	    RECT 370.8000 211.6000 371.6000 212.4000 ;
	    RECT 377.2000 211.8000 378.0000 212.6000 ;
	    RECT 377.3000 210.4000 377.9000 211.8000 ;
	    RECT 377.2000 209.6000 378.0000 210.4000 ;
	    RECT 378.8000 206.2000 379.6000 217.8000 ;
	    RECT 382.0000 210.2000 382.8000 215.8000 ;
	    RECT 383.7000 214.4000 384.3000 219.6000 ;
	    RECT 383.6000 213.6000 384.4000 214.4000 ;
	    RECT 386.9000 212.4000 387.5000 229.6000 ;
	    RECT 394.9000 222.3000 395.5000 229.6000 ;
	    RECT 396.4000 227.6000 397.2000 228.4000 ;
	    RECT 396.5000 226.4000 397.1000 227.6000 ;
	    RECT 396.4000 225.6000 397.2000 226.4000 ;
	    RECT 396.4000 223.6000 397.2000 224.4000 ;
	    RECT 396.5000 222.3000 397.1000 223.6000 ;
	    RECT 394.9000 221.7000 397.1000 222.3000 ;
	    RECT 393.2000 215.6000 394.0000 216.4000 ;
	    RECT 393.3000 214.4000 393.9000 215.6000 ;
	    RECT 388.4000 213.6000 389.2000 214.4000 ;
	    RECT 393.2000 213.6000 394.0000 214.4000 ;
	    RECT 386.8000 211.6000 387.6000 212.4000 ;
	    RECT 388.5000 210.4000 389.1000 213.6000 ;
	    RECT 391.6000 211.6000 392.4000 212.4000 ;
	    RECT 394.8000 211.6000 395.6000 212.4000 ;
	    RECT 386.8000 209.6000 387.6000 210.4000 ;
	    RECT 388.4000 209.6000 389.2000 210.4000 ;
	    RECT 362.8000 203.6000 363.6000 204.4000 ;
	    RECT 386.9000 202.4000 387.5000 209.6000 ;
	    RECT 391.7000 202.4000 392.3000 211.6000 ;
	    RECT 394.9000 204.4000 395.5000 211.6000 ;
	    RECT 396.5000 210.4000 397.1000 221.7000 ;
	    RECT 398.1000 218.4000 398.7000 231.7000 ;
	    RECT 399.6000 231.6000 400.4000 231.7000 ;
	    RECT 402.8000 231.6000 403.6000 232.4000 ;
	    RECT 404.4000 231.6000 405.2000 232.4000 ;
	    RECT 404.5000 230.4000 405.1000 231.6000 ;
	    RECT 402.8000 229.6000 403.6000 230.4000 ;
	    RECT 404.4000 229.6000 405.2000 230.4000 ;
	    RECT 412.5000 228.4000 413.1000 237.6000 ;
	    RECT 412.4000 227.6000 413.2000 228.4000 ;
	    RECT 414.0000 225.6000 414.8000 226.4000 ;
	    RECT 414.1000 224.4000 414.7000 225.6000 ;
	    RECT 414.0000 223.6000 414.8000 224.4000 ;
	    RECT 418.8000 224.2000 419.6000 235.8000 ;
	    RECT 425.2000 229.6000 426.0000 230.4000 ;
	    RECT 428.4000 224.2000 429.2000 235.8000 ;
	    RECT 430.1000 228.4000 430.7000 249.6000 ;
	    RECT 433.2000 246.2000 434.0000 257.8000 ;
	    RECT 433.2000 243.6000 434.0000 244.4000 ;
	    RECT 433.3000 238.4000 433.9000 243.6000 ;
	    RECT 433.2000 237.6000 434.0000 238.4000 ;
	    RECT 430.0000 227.6000 430.8000 228.4000 ;
	    RECT 431.6000 226.2000 432.4000 231.8000 ;
	    RECT 398.0000 217.6000 398.8000 218.4000 ;
	    RECT 399.6000 217.6000 400.4000 218.4000 ;
	    RECT 417.2000 217.6000 418.0000 218.4000 ;
	    RECT 434.9000 218.3000 435.5000 267.6000 ;
	    RECT 439.6000 263.6000 440.4000 264.4000 ;
	    RECT 439.7000 252.4000 440.3000 263.6000 ;
	    RECT 449.3000 258.4000 449.9000 267.6000 ;
	    RECT 454.0000 263.6000 454.8000 264.4000 ;
	    RECT 465.3000 260.4000 465.9000 269.6000 ;
	    RECT 452.4000 259.6000 453.2000 260.4000 ;
	    RECT 465.2000 259.6000 466.0000 260.4000 ;
	    RECT 441.2000 253.6000 442.0000 254.4000 ;
	    RECT 439.6000 251.6000 440.4000 252.4000 ;
	    RECT 441.3000 250.4000 441.9000 253.6000 ;
	    RECT 441.2000 249.6000 442.0000 250.4000 ;
	    RECT 442.8000 246.2000 443.6000 257.8000 ;
	    RECT 449.2000 257.6000 450.0000 258.4000 ;
	    RECT 450.8000 257.6000 451.6000 258.4000 ;
	    RECT 446.0000 250.2000 446.8000 255.8000 ;
	    RECT 447.6000 255.6000 448.4000 256.4000 ;
	    RECT 450.9000 252.4000 451.5000 257.6000 ;
	    RECT 450.8000 251.6000 451.6000 252.4000 ;
	    RECT 442.8000 243.6000 443.6000 244.4000 ;
	    RECT 436.4000 233.6000 437.2000 234.4000 ;
	    RECT 441.2000 233.6000 442.0000 234.4000 ;
	    RECT 442.9000 230.4000 443.5000 243.6000 ;
	    RECT 452.5000 232.4000 453.1000 259.6000 ;
	    RECT 454.0000 251.6000 454.8000 252.4000 ;
	    RECT 449.2000 231.6000 450.0000 232.4000 ;
	    RECT 450.8000 231.6000 451.6000 232.4000 ;
	    RECT 452.4000 231.6000 453.2000 232.4000 ;
	    RECT 449.3000 230.4000 449.9000 231.6000 ;
	    RECT 450.9000 230.4000 451.5000 231.6000 ;
	    RECT 436.4000 229.6000 437.2000 230.4000 ;
	    RECT 441.2000 229.6000 442.0000 230.4000 ;
	    RECT 442.8000 229.6000 443.6000 230.4000 ;
	    RECT 449.2000 229.6000 450.0000 230.4000 ;
	    RECT 450.8000 229.6000 451.6000 230.4000 ;
	    RECT 436.5000 228.4000 437.1000 229.6000 ;
	    RECT 441.3000 228.4000 441.9000 229.6000 ;
	    RECT 436.4000 227.6000 437.2000 228.4000 ;
	    RECT 441.2000 227.6000 442.0000 228.4000 ;
	    RECT 439.6000 223.6000 440.4000 224.4000 ;
	    RECT 439.7000 218.4000 440.3000 223.6000 ;
	    RECT 399.7000 214.4000 400.3000 217.6000 ;
	    RECT 399.6000 213.6000 400.4000 214.4000 ;
	    RECT 412.4000 213.6000 413.2000 214.4000 ;
	    RECT 415.6000 213.6000 416.4000 214.4000 ;
	    RECT 396.4000 209.6000 397.2000 210.4000 ;
	    RECT 394.8000 203.6000 395.6000 204.4000 ;
	    RECT 362.8000 201.6000 363.6000 202.4000 ;
	    RECT 386.8000 201.6000 387.6000 202.4000 ;
	    RECT 391.6000 201.6000 392.4000 202.4000 ;
	    RECT 362.9000 190.4000 363.5000 201.6000 ;
	    RECT 367.6000 197.6000 368.4000 198.4000 ;
	    RECT 364.4000 193.6000 365.2000 194.4000 ;
	    RECT 364.5000 190.4000 365.1000 193.6000 ;
	    RECT 362.8000 189.6000 363.6000 190.4000 ;
	    RECT 364.4000 189.6000 365.2000 190.4000 ;
	    RECT 362.8000 187.6000 363.6000 188.4000 ;
	    RECT 362.9000 184.4000 363.5000 187.6000 ;
	    RECT 362.8000 183.6000 363.6000 184.4000 ;
	    RECT 353.2000 179.6000 354.0000 180.4000 ;
	    RECT 361.2000 179.6000 362.0000 180.4000 ;
	    RECT 353.3000 172.4000 353.9000 179.6000 ;
	    RECT 358.0000 173.6000 358.8000 174.4000 ;
	    RECT 358.1000 172.4000 358.7000 173.6000 ;
	    RECT 361.3000 172.4000 361.9000 179.6000 ;
	    RECT 367.7000 174.4000 368.3000 197.6000 ;
	    RECT 394.9000 196.4000 395.5000 203.6000 ;
	    RECT 399.7000 198.4000 400.3000 213.6000 ;
	    RECT 402.8000 209.6000 403.6000 210.4000 ;
	    RECT 402.9000 206.4000 403.5000 209.6000 ;
	    RECT 402.8000 205.6000 403.6000 206.4000 ;
	    RECT 402.9000 202.4000 403.5000 205.6000 ;
	    RECT 412.5000 204.3000 413.1000 213.6000 ;
	    RECT 415.6000 211.6000 416.4000 212.4000 ;
	    RECT 414.0000 209.6000 414.8000 210.4000 ;
	    RECT 415.7000 206.4000 416.3000 211.6000 ;
	    RECT 418.8000 207.6000 419.6000 208.4000 ;
	    RECT 415.6000 205.6000 416.4000 206.4000 ;
	    RECT 412.5000 203.7000 414.7000 204.3000 ;
	    RECT 402.8000 201.6000 403.6000 202.4000 ;
	    RECT 414.1000 198.4000 414.7000 203.7000 ;
	    RECT 417.2000 201.6000 418.0000 202.4000 ;
	    RECT 399.6000 197.6000 400.4000 198.4000 ;
	    RECT 414.0000 197.6000 414.8000 198.4000 ;
	    RECT 369.2000 184.2000 370.0000 195.8000 ;
	    RECT 375.6000 189.6000 376.4000 190.4000 ;
	    RECT 375.7000 188.4000 376.3000 189.6000 ;
	    RECT 375.6000 187.6000 376.4000 188.4000 ;
	    RECT 377.2000 185.6000 378.0000 186.4000 ;
	    RECT 377.3000 178.4000 377.9000 185.6000 ;
	    RECT 378.8000 184.2000 379.6000 195.8000 ;
	    RECT 382.0000 186.2000 382.8000 191.8000 ;
	    RECT 385.2000 189.6000 386.0000 190.4000 ;
	    RECT 383.6000 187.6000 384.4000 188.4000 ;
	    RECT 386.8000 187.6000 387.6000 188.4000 ;
	    RECT 383.7000 186.4000 384.3000 187.6000 ;
	    RECT 383.6000 185.6000 384.4000 186.4000 ;
	    RECT 380.4000 183.6000 381.2000 184.4000 ;
	    RECT 375.6000 177.6000 376.4000 178.4000 ;
	    RECT 377.2000 177.6000 378.0000 178.4000 ;
	    RECT 370.8000 175.6000 371.6000 176.4000 ;
	    RECT 367.6000 173.6000 368.4000 174.4000 ;
	    RECT 367.7000 172.4000 368.3000 173.6000 ;
	    RECT 370.9000 172.4000 371.5000 175.6000 ;
	    RECT 348.4000 171.7000 350.7000 172.3000 ;
	    RECT 343.6000 171.6000 344.4000 171.7000 ;
	    RECT 348.4000 171.6000 349.2000 171.7000 ;
	    RECT 351.6000 171.6000 352.4000 172.4000 ;
	    RECT 353.2000 171.6000 354.0000 172.4000 ;
	    RECT 358.0000 171.6000 358.8000 172.4000 ;
	    RECT 359.6000 171.6000 360.4000 172.4000 ;
	    RECT 361.2000 171.6000 362.0000 172.4000 ;
	    RECT 367.6000 171.6000 368.4000 172.4000 ;
	    RECT 369.2000 171.6000 370.0000 172.4000 ;
	    RECT 370.8000 171.6000 371.6000 172.4000 ;
	    RECT 372.4000 171.6000 373.2000 172.4000 ;
	    RECT 332.4000 169.6000 333.2000 170.4000 ;
	    RECT 321.2000 163.6000 322.0000 164.4000 ;
	    RECT 322.8000 163.6000 323.6000 164.4000 ;
	    RECT 324.4000 163.6000 325.2000 164.4000 ;
	    RECT 329.2000 163.6000 330.0000 164.4000 ;
	    RECT 321.3000 158.4000 321.9000 163.6000 ;
	    RECT 321.2000 157.6000 322.0000 158.4000 ;
	    RECT 324.5000 150.4000 325.1000 163.6000 ;
	    RECT 326.0000 157.6000 326.8000 158.4000 ;
	    RECT 318.0000 149.7000 320.3000 150.3000 ;
	    RECT 318.0000 149.6000 318.8000 149.7000 ;
	    RECT 321.2000 149.6000 322.0000 150.4000 ;
	    RECT 324.4000 149.6000 325.2000 150.4000 ;
	    RECT 319.6000 147.6000 320.4000 148.4000 ;
	    RECT 318.0000 143.6000 318.8000 144.4000 ;
	    RECT 318.1000 142.4000 318.7000 143.6000 ;
	    RECT 318.0000 141.6000 318.8000 142.4000 ;
	    RECT 314.9000 137.7000 317.1000 138.3000 ;
	    RECT 313.2000 135.6000 314.0000 136.4000 ;
	    RECT 311.6000 133.6000 312.4000 134.4000 ;
	    RECT 310.0000 131.6000 310.8000 132.4000 ;
	    RECT 300.5000 129.7000 302.7000 130.3000 ;
	    RECT 281.3000 127.7000 283.5000 128.3000 ;
	    RECT 278.1000 118.4000 278.7000 127.6000 ;
	    RECT 281.2000 125.6000 282.0000 126.4000 ;
	    RECT 278.0000 117.6000 278.8000 118.4000 ;
	    RECT 281.3000 110.4000 281.9000 125.6000 ;
	    RECT 282.9000 118.4000 283.5000 127.7000 ;
	    RECT 284.4000 127.6000 285.2000 128.4000 ;
	    RECT 286.0000 125.6000 286.8000 126.4000 ;
	    RECT 284.4000 123.6000 285.2000 124.4000 ;
	    RECT 282.8000 117.6000 283.6000 118.4000 ;
	    RECT 274.8000 109.6000 275.6000 110.4000 ;
	    RECT 281.2000 109.6000 282.0000 110.4000 ;
	    RECT 273.2000 105.6000 274.0000 106.4000 ;
	    RECT 273.3000 104.4000 273.9000 105.6000 ;
	    RECT 273.2000 103.6000 274.0000 104.4000 ;
	    RECT 271.6000 97.6000 272.4000 98.4000 ;
	    RECT 260.4000 93.6000 261.2000 94.4000 ;
	    RECT 262.0000 93.6000 262.8000 94.4000 ;
	    RECT 266.8000 93.6000 267.6000 94.4000 ;
	    RECT 270.0000 93.6000 270.8000 94.4000 ;
	    RECT 255.6000 83.6000 256.4000 84.4000 ;
	    RECT 252.5000 71.7000 254.7000 72.3000 ;
	    RECT 247.7000 70.4000 248.3000 71.6000 ;
	    RECT 244.4000 69.6000 245.2000 70.4000 ;
	    RECT 247.6000 69.6000 248.4000 70.4000 ;
	    RECT 250.8000 69.6000 251.6000 70.4000 ;
	    RECT 234.8000 67.6000 235.6000 68.4000 ;
	    RECT 238.0000 67.6000 238.8000 68.4000 ;
	    RECT 241.2000 67.6000 242.0000 68.4000 ;
	    RECT 242.8000 67.6000 243.6000 68.4000 ;
	    RECT 249.2000 67.6000 250.0000 68.4000 ;
	    RECT 236.4000 63.6000 237.2000 64.4000 ;
	    RECT 226.8000 55.6000 227.6000 56.4000 ;
	    RECT 231.6000 55.6000 232.4000 56.4000 ;
	    RECT 223.6000 53.6000 224.4000 54.4000 ;
	    RECT 225.2000 53.6000 226.0000 54.4000 ;
	    RECT 222.0000 51.6000 222.8000 52.4000 ;
	    RECT 218.8000 49.6000 219.6000 50.4000 ;
	    RECT 220.4000 49.6000 221.2000 50.4000 ;
	    RECT 225.3000 46.4000 225.9000 53.6000 ;
	    RECT 236.5000 52.4000 237.1000 63.6000 ;
	    RECT 238.1000 54.4000 238.7000 67.6000 ;
	    RECT 247.6000 64.3000 248.4000 64.4000 ;
	    RECT 247.6000 63.7000 249.9000 64.3000 ;
	    RECT 247.6000 63.6000 248.4000 63.7000 ;
	    RECT 239.6000 57.6000 240.4000 58.4000 ;
	    RECT 247.6000 57.6000 248.4000 58.4000 ;
	    RECT 239.7000 56.4000 240.3000 57.6000 ;
	    RECT 239.6000 55.6000 240.4000 56.4000 ;
	    RECT 249.3000 56.3000 249.9000 63.7000 ;
	    RECT 250.9000 58.4000 251.5000 69.6000 ;
	    RECT 250.8000 57.6000 251.6000 58.4000 ;
	    RECT 247.7000 55.7000 249.9000 56.3000 ;
	    RECT 238.0000 53.6000 238.8000 54.4000 ;
	    RECT 226.8000 51.6000 227.6000 52.4000 ;
	    RECT 231.6000 51.6000 232.4000 52.4000 ;
	    RECT 233.2000 51.6000 234.0000 52.4000 ;
	    RECT 236.4000 51.6000 237.2000 52.4000 ;
	    RECT 222.0000 45.6000 222.8000 46.4000 ;
	    RECT 225.2000 45.6000 226.0000 46.4000 ;
	    RECT 217.2000 43.6000 218.0000 44.4000 ;
	    RECT 204.4000 39.6000 205.2000 40.4000 ;
	    RECT 215.6000 39.6000 216.4000 40.4000 ;
	    RECT 214.0000 31.6000 214.8000 32.4000 ;
	    RECT 214.1000 30.4000 214.7000 31.6000 ;
	    RECT 206.0000 29.6000 206.8000 30.4000 ;
	    RECT 207.6000 29.6000 208.4000 30.4000 ;
	    RECT 214.0000 29.6000 214.8000 30.4000 ;
	    RECT 215.6000 29.6000 216.4000 30.4000 ;
	    RECT 206.1000 26.4000 206.7000 29.6000 ;
	    RECT 206.0000 25.6000 206.8000 26.4000 ;
	    RECT 207.7000 18.4000 208.3000 29.6000 ;
	    RECT 215.7000 28.4000 216.3000 29.6000 ;
	    RECT 215.6000 27.6000 216.4000 28.4000 ;
	    RECT 209.2000 25.6000 210.0000 26.4000 ;
	    RECT 202.8000 15.6000 203.6000 16.4000 ;
	    RECT 202.8000 13.6000 203.6000 14.4000 ;
	    RECT 202.9000 12.6000 203.5000 13.6000 ;
	    RECT 202.8000 11.8000 203.6000 12.6000 ;
	    RECT 202.9000 11.7000 203.5000 11.8000 ;
	    RECT 201.2000 9.6000 202.0000 10.4000 ;
	    RECT 196.4000 7.6000 197.2000 8.4000 ;
	    RECT 204.4000 6.2000 205.2000 17.8000 ;
	    RECT 207.6000 17.6000 208.4000 18.4000 ;
	    RECT 207.6000 10.2000 208.4000 15.8000 ;
	    RECT 209.3000 14.4000 209.9000 25.6000 ;
	    RECT 215.6000 23.6000 216.4000 24.4000 ;
	    RECT 209.2000 13.6000 210.0000 14.4000 ;
	    RECT 214.0000 13.6000 214.8000 14.4000 ;
	    RECT 217.3000 12.4000 217.9000 43.6000 ;
	    RECT 222.1000 32.4000 222.7000 45.6000 ;
	    RECT 231.7000 38.4000 232.3000 51.6000 ;
	    RECT 233.2000 49.6000 234.0000 50.4000 ;
	    RECT 233.3000 46.4000 233.9000 49.6000 ;
	    RECT 233.2000 45.6000 234.0000 46.4000 ;
	    RECT 231.6000 37.6000 232.4000 38.4000 ;
	    RECT 233.3000 34.4000 233.9000 45.6000 ;
	    RECT 233.2000 33.6000 234.0000 34.4000 ;
	    RECT 222.0000 31.6000 222.8000 32.4000 ;
	    RECT 236.5000 30.4000 237.1000 51.6000 ;
	    RECT 238.1000 38.4000 238.7000 53.6000 ;
	    RECT 239.6000 51.6000 240.4000 52.4000 ;
	    RECT 242.8000 51.6000 243.6000 52.4000 ;
	    RECT 238.0000 37.6000 238.8000 38.4000 ;
	    RECT 242.9000 30.4000 243.5000 51.6000 ;
	    RECT 246.0000 47.6000 246.8000 48.4000 ;
	    RECT 246.1000 38.4000 246.7000 47.6000 ;
	    RECT 246.0000 37.6000 246.8000 38.4000 ;
	    RECT 218.8000 29.6000 219.6000 30.4000 ;
	    RECT 225.2000 29.6000 226.0000 30.4000 ;
	    RECT 230.0000 29.6000 230.8000 30.4000 ;
	    RECT 234.8000 29.6000 235.6000 30.4000 ;
	    RECT 236.4000 29.6000 237.2000 30.4000 ;
	    RECT 242.8000 29.6000 243.6000 30.4000 ;
	    RECT 244.4000 29.6000 245.2000 30.4000 ;
	    RECT 218.9000 24.4000 219.5000 29.6000 ;
	    RECT 230.1000 28.4000 230.7000 29.6000 ;
	    RECT 226.8000 27.6000 227.6000 28.4000 ;
	    RECT 230.0000 27.6000 230.8000 28.4000 ;
	    RECT 220.4000 25.6000 221.2000 26.4000 ;
	    RECT 218.8000 23.6000 219.6000 24.4000 ;
	    RECT 218.8000 19.6000 219.6000 20.4000 ;
	    RECT 218.9000 14.4000 219.5000 19.6000 ;
	    RECT 220.5000 14.4000 221.1000 25.6000 ;
	    RECT 222.0000 15.6000 222.8000 16.4000 ;
	    RECT 218.8000 13.6000 219.6000 14.4000 ;
	    RECT 220.4000 13.6000 221.2000 14.4000 ;
	    RECT 226.9000 12.4000 227.5000 27.6000 ;
	    RECT 228.4000 25.6000 229.2000 26.4000 ;
	    RECT 212.4000 11.6000 213.2000 12.4000 ;
	    RECT 217.2000 11.6000 218.0000 12.4000 ;
	    RECT 222.0000 11.6000 222.8000 12.4000 ;
	    RECT 225.2000 11.6000 226.0000 12.4000 ;
	    RECT 226.8000 11.6000 227.6000 12.4000 ;
	    RECT 212.5000 10.4000 213.1000 11.6000 ;
	    RECT 222.1000 10.4000 222.7000 11.6000 ;
	    RECT 225.3000 10.4000 225.9000 11.6000 ;
	    RECT 228.5000 10.4000 229.1000 25.6000 ;
	    RECT 234.9000 16.4000 235.5000 29.6000 ;
	    RECT 238.0000 25.6000 238.8000 26.4000 ;
	    RECT 242.9000 26.3000 243.5000 29.6000 ;
	    RECT 244.5000 28.4000 245.1000 29.6000 ;
	    RECT 244.4000 27.6000 245.2000 28.4000 ;
	    RECT 242.9000 25.7000 245.1000 26.3000 ;
	    RECT 236.4000 19.6000 237.2000 20.4000 ;
	    RECT 236.5000 18.4000 237.1000 19.6000 ;
	    RECT 238.1000 18.4000 238.7000 25.6000 ;
	    RECT 239.6000 23.6000 240.4000 24.4000 ;
	    RECT 236.4000 17.6000 237.2000 18.4000 ;
	    RECT 238.0000 17.6000 238.8000 18.4000 ;
	    RECT 234.8000 15.6000 235.6000 16.4000 ;
	    RECT 233.2000 13.6000 234.0000 14.4000 ;
	    RECT 234.8000 14.3000 235.6000 14.4000 ;
	    RECT 236.5000 14.3000 237.1000 17.6000 ;
	    RECT 238.1000 16.4000 238.7000 17.6000 ;
	    RECT 238.0000 15.6000 238.8000 16.4000 ;
	    RECT 234.8000 13.7000 237.1000 14.3000 ;
	    RECT 234.8000 13.6000 235.6000 13.7000 ;
	    RECT 233.3000 12.4000 233.9000 13.6000 ;
	    RECT 231.6000 11.6000 232.4000 12.4000 ;
	    RECT 233.2000 11.6000 234.0000 12.4000 ;
	    RECT 212.4000 9.6000 213.2000 10.4000 ;
	    RECT 222.0000 9.6000 222.8000 10.4000 ;
	    RECT 225.2000 9.6000 226.0000 10.4000 ;
	    RECT 228.4000 9.6000 229.2000 10.4000 ;
	    RECT 234.8000 9.6000 235.6000 10.4000 ;
	    RECT 239.6000 10.2000 240.4000 15.8000 ;
	    RECT 241.2000 13.6000 242.0000 14.4000 ;
	    RECT 234.9000 8.4000 235.5000 9.6000 ;
	    RECT 241.3000 8.4000 241.9000 13.6000 ;
	    RECT 234.8000 7.6000 235.6000 8.4000 ;
	    RECT 241.2000 7.6000 242.0000 8.4000 ;
	    RECT 242.8000 6.2000 243.6000 17.8000 ;
	    RECT 244.5000 10.4000 245.1000 25.7000 ;
	    RECT 247.7000 12.4000 248.3000 55.7000 ;
	    RECT 252.5000 54.4000 253.1000 71.7000 ;
	    RECT 255.7000 68.4000 256.3000 83.6000 ;
	    RECT 257.2000 71.6000 258.0000 72.4000 ;
	    RECT 257.3000 70.4000 257.9000 71.6000 ;
	    RECT 257.2000 69.6000 258.0000 70.4000 ;
	    RECT 258.8000 69.6000 259.6000 70.4000 ;
	    RECT 258.9000 68.4000 259.5000 69.6000 ;
	    RECT 255.6000 67.6000 256.4000 68.4000 ;
	    RECT 258.8000 67.6000 259.6000 68.4000 ;
	    RECT 260.5000 68.3000 261.1000 93.6000 ;
	    RECT 274.9000 92.4000 275.5000 109.6000 ;
	    RECT 281.3000 108.4000 281.9000 109.6000 ;
	    RECT 281.2000 107.6000 282.0000 108.4000 ;
	    RECT 282.8000 103.6000 283.6000 104.4000 ;
	    RECT 281.2000 93.6000 282.0000 94.4000 ;
	    RECT 274.8000 91.6000 275.6000 92.4000 ;
	    RECT 278.0000 91.6000 278.8000 92.4000 ;
	    RECT 266.8000 89.6000 267.6000 90.4000 ;
	    RECT 266.9000 80.4000 267.5000 89.6000 ;
	    RECT 271.6000 83.6000 272.4000 84.4000 ;
	    RECT 276.4000 83.6000 277.2000 84.4000 ;
	    RECT 266.8000 79.6000 267.6000 80.4000 ;
	    RECT 268.4000 79.6000 269.2000 80.4000 ;
	    RECT 263.6000 78.3000 264.4000 78.4000 ;
	    RECT 268.5000 78.3000 269.1000 79.6000 ;
	    RECT 263.6000 77.7000 269.1000 78.3000 ;
	    RECT 263.6000 77.6000 264.4000 77.7000 ;
	    RECT 262.0000 75.6000 262.8000 76.4000 ;
	    RECT 262.1000 70.4000 262.7000 75.6000 ;
	    RECT 266.8000 71.6000 267.6000 72.4000 ;
	    RECT 268.4000 71.6000 269.2000 72.4000 ;
	    RECT 262.0000 69.6000 262.8000 70.4000 ;
	    RECT 266.9000 68.4000 267.5000 71.6000 ;
	    RECT 260.5000 67.7000 262.7000 68.3000 ;
	    RECT 262.1000 58.4000 262.7000 67.7000 ;
	    RECT 263.6000 67.6000 264.4000 68.4000 ;
	    RECT 266.8000 67.6000 267.6000 68.4000 ;
	    RECT 263.7000 58.4000 264.3000 67.6000 ;
	    RECT 268.5000 66.4000 269.1000 71.6000 ;
	    RECT 271.7000 70.4000 272.3000 83.6000 ;
	    RECT 273.2000 81.6000 274.0000 82.4000 ;
	    RECT 270.0000 69.6000 270.8000 70.4000 ;
	    RECT 271.6000 69.6000 272.4000 70.4000 ;
	    RECT 270.1000 68.4000 270.7000 69.6000 ;
	    RECT 273.3000 68.4000 273.9000 81.6000 ;
	    RECT 276.5000 80.4000 277.1000 83.6000 ;
	    RECT 278.1000 80.4000 278.7000 91.6000 ;
	    RECT 281.3000 90.4000 281.9000 93.6000 ;
	    RECT 282.9000 92.4000 283.5000 103.6000 ;
	    RECT 284.5000 96.3000 285.1000 123.6000 ;
	    RECT 286.1000 112.4000 286.7000 125.6000 ;
	    RECT 286.0000 111.6000 286.8000 112.4000 ;
	    RECT 287.7000 110.4000 288.3000 129.6000 ;
	    RECT 298.9000 120.4000 299.5000 129.6000 ;
	    RECT 302.1000 128.4000 302.7000 129.7000 ;
	    RECT 306.8000 129.6000 307.6000 130.4000 ;
	    RECT 302.0000 127.6000 302.8000 128.4000 ;
	    RECT 313.2000 127.6000 314.0000 128.4000 ;
	    RECT 313.3000 120.4000 313.9000 127.6000 ;
	    RECT 298.8000 119.6000 299.6000 120.4000 ;
	    RECT 303.6000 119.6000 304.4000 120.4000 ;
	    RECT 313.2000 119.6000 314.0000 120.4000 ;
	    RECT 300.4000 115.6000 301.2000 116.4000 ;
	    RECT 294.0000 113.6000 294.8000 114.4000 ;
	    RECT 300.4000 113.6000 301.2000 114.4000 ;
	    RECT 289.2000 111.6000 290.0000 112.4000 ;
	    RECT 289.3000 110.4000 289.9000 111.6000 ;
	    RECT 300.5000 110.4000 301.1000 113.6000 ;
	    RECT 303.7000 110.4000 304.3000 119.6000 ;
	    RECT 306.8000 111.6000 307.6000 112.4000 ;
	    RECT 311.6000 111.6000 312.4000 112.4000 ;
	    RECT 306.9000 110.4000 307.5000 111.6000 ;
	    RECT 311.7000 110.4000 312.3000 111.6000 ;
	    RECT 313.3000 110.4000 313.9000 119.6000 ;
	    RECT 314.9000 118.4000 315.5000 137.7000 ;
	    RECT 318.0000 137.6000 318.8000 138.4000 ;
	    RECT 316.4000 135.6000 317.2000 136.4000 ;
	    RECT 316.5000 132.4000 317.1000 135.6000 ;
	    RECT 318.1000 134.4000 318.7000 137.6000 ;
	    RECT 321.3000 136.4000 321.9000 149.6000 ;
	    RECT 326.1000 148.4000 326.7000 157.6000 ;
	    RECT 327.6000 155.6000 328.4000 156.4000 ;
	    RECT 329.3000 154.4000 329.9000 163.6000 ;
	    RECT 332.5000 158.4000 333.1000 169.6000 ;
	    RECT 332.4000 157.6000 333.2000 158.4000 ;
	    RECT 334.0000 155.6000 334.8000 156.4000 ;
	    RECT 329.2000 153.6000 330.0000 154.4000 ;
	    RECT 330.8000 153.6000 331.6000 154.4000 ;
	    RECT 329.2000 152.3000 330.0000 152.4000 ;
	    RECT 330.9000 152.3000 331.5000 153.6000 ;
	    RECT 329.2000 151.7000 331.5000 152.3000 ;
	    RECT 329.2000 151.6000 330.0000 151.7000 ;
	    RECT 326.0000 147.6000 326.8000 148.4000 ;
	    RECT 324.4000 145.6000 325.2000 146.4000 ;
	    RECT 324.5000 144.4000 325.1000 145.6000 ;
	    RECT 324.4000 143.6000 325.2000 144.4000 ;
	    RECT 326.0000 137.6000 326.8000 138.4000 ;
	    RECT 327.6000 137.6000 328.4000 138.4000 ;
	    RECT 321.2000 135.6000 322.0000 136.4000 ;
	    RECT 318.0000 133.6000 318.8000 134.4000 ;
	    RECT 324.4000 133.6000 325.2000 134.4000 ;
	    RECT 324.5000 132.4000 325.1000 133.6000 ;
	    RECT 316.4000 132.3000 317.2000 132.4000 ;
	    RECT 316.4000 131.7000 318.7000 132.3000 ;
	    RECT 316.4000 131.6000 317.2000 131.7000 ;
	    RECT 316.4000 127.6000 317.2000 128.4000 ;
	    RECT 318.1000 120.4000 318.7000 131.7000 ;
	    RECT 319.6000 131.6000 320.4000 132.4000 ;
	    RECT 322.8000 131.6000 323.6000 132.4000 ;
	    RECT 324.4000 131.6000 325.2000 132.4000 ;
	    RECT 319.7000 128.4000 320.3000 131.6000 ;
	    RECT 319.6000 127.6000 320.4000 128.4000 ;
	    RECT 322.9000 126.4000 323.5000 131.6000 ;
	    RECT 324.5000 130.3000 325.1000 131.6000 ;
	    RECT 326.0000 130.3000 326.8000 130.4000 ;
	    RECT 324.5000 129.7000 326.8000 130.3000 ;
	    RECT 326.0000 129.6000 326.8000 129.7000 ;
	    RECT 327.7000 128.4000 328.3000 137.6000 ;
	    RECT 329.3000 132.4000 329.9000 151.6000 ;
	    RECT 330.8000 149.6000 331.6000 150.4000 ;
	    RECT 330.9000 142.4000 331.5000 149.6000 ;
	    RECT 334.1000 148.4000 334.7000 155.6000 ;
	    RECT 337.2000 151.6000 338.0000 152.4000 ;
	    RECT 337.3000 150.4000 337.9000 151.6000 ;
	    RECT 337.2000 149.6000 338.0000 150.4000 ;
	    RECT 332.4000 147.6000 333.2000 148.4000 ;
	    RECT 334.0000 147.6000 334.8000 148.4000 ;
	    RECT 337.2000 147.6000 338.0000 148.4000 ;
	    RECT 338.8000 148.3000 339.6000 148.4000 ;
	    RECT 340.5000 148.3000 341.1000 171.6000 ;
	    RECT 351.7000 170.4000 352.3000 171.6000 ;
	    RECT 369.3000 170.4000 369.9000 171.6000 ;
	    RECT 351.6000 169.6000 352.4000 170.4000 ;
	    RECT 354.8000 170.3000 355.6000 170.4000 ;
	    RECT 353.3000 169.7000 355.6000 170.3000 ;
	    RECT 348.4000 165.6000 349.2000 166.4000 ;
	    RECT 342.0000 163.6000 342.8000 164.4000 ;
	    RECT 342.1000 150.3000 342.7000 163.6000 ;
	    RECT 343.6000 153.6000 344.4000 154.4000 ;
	    RECT 343.7000 152.3000 344.3000 153.6000 ;
	    RECT 343.7000 151.7000 345.9000 152.3000 ;
	    RECT 345.3000 150.4000 345.9000 151.7000 ;
	    RECT 346.8000 151.6000 347.6000 152.4000 ;
	    RECT 343.6000 150.3000 344.4000 150.4000 ;
	    RECT 342.1000 149.7000 344.4000 150.3000 ;
	    RECT 343.6000 149.6000 344.4000 149.7000 ;
	    RECT 345.2000 149.6000 346.0000 150.4000 ;
	    RECT 338.8000 147.7000 341.1000 148.3000 ;
	    RECT 338.8000 147.6000 339.6000 147.7000 ;
	    RECT 332.5000 146.3000 333.1000 147.6000 ;
	    RECT 332.5000 145.7000 334.7000 146.3000 ;
	    RECT 330.8000 141.6000 331.6000 142.4000 ;
	    RECT 330.8000 133.6000 331.6000 134.4000 ;
	    RECT 329.2000 131.6000 330.0000 132.4000 ;
	    RECT 332.4000 131.6000 333.2000 132.4000 ;
	    RECT 332.4000 130.3000 333.2000 130.4000 ;
	    RECT 334.1000 130.3000 334.7000 145.7000 ;
	    RECT 337.3000 134.4000 337.9000 147.6000 ;
	    RECT 338.9000 134.4000 339.5000 147.6000 ;
	    RECT 340.4000 145.6000 341.2000 146.4000 ;
	    RECT 340.5000 144.4000 341.1000 145.6000 ;
	    RECT 340.4000 143.6000 341.2000 144.4000 ;
	    RECT 335.6000 133.6000 336.4000 134.4000 ;
	    RECT 337.2000 133.6000 338.0000 134.4000 ;
	    RECT 338.8000 133.6000 339.6000 134.4000 ;
	    RECT 335.7000 132.4000 336.3000 133.6000 ;
	    RECT 335.6000 131.6000 336.4000 132.4000 ;
	    RECT 338.8000 131.6000 339.6000 132.4000 ;
	    RECT 332.4000 129.7000 334.7000 130.3000 ;
	    RECT 332.4000 129.6000 333.2000 129.7000 ;
	    RECT 327.6000 127.6000 328.4000 128.4000 ;
	    RECT 322.8000 125.6000 323.6000 126.4000 ;
	    RECT 319.6000 123.6000 320.4000 124.4000 ;
	    RECT 318.0000 119.6000 318.8000 120.4000 ;
	    RECT 332.5000 118.4000 333.1000 129.6000 ;
	    RECT 334.0000 127.6000 334.8000 128.4000 ;
	    RECT 334.1000 118.4000 334.7000 127.6000 ;
	    RECT 338.9000 120.3000 339.5000 131.6000 ;
	    RECT 340.5000 128.4000 341.1000 143.6000 ;
	    RECT 343.7000 138.3000 344.3000 149.6000 ;
	    RECT 345.2000 147.6000 346.0000 148.4000 ;
	    RECT 345.3000 144.4000 345.9000 147.6000 ;
	    RECT 345.2000 143.6000 346.0000 144.4000 ;
	    RECT 343.7000 137.7000 345.9000 138.3000 ;
	    RECT 343.6000 135.6000 344.4000 136.4000 ;
	    RECT 343.7000 134.4000 344.3000 135.6000 ;
	    RECT 343.6000 133.6000 344.4000 134.4000 ;
	    RECT 345.3000 132.4000 345.9000 137.7000 ;
	    RECT 343.6000 131.6000 344.4000 132.4000 ;
	    RECT 345.2000 131.6000 346.0000 132.4000 ;
	    RECT 343.7000 130.3000 344.3000 131.6000 ;
	    RECT 343.7000 129.7000 345.9000 130.3000 ;
	    RECT 345.3000 128.4000 345.9000 129.7000 ;
	    RECT 340.4000 127.6000 341.2000 128.4000 ;
	    RECT 345.2000 127.6000 346.0000 128.4000 ;
	    RECT 340.4000 123.6000 341.2000 124.4000 ;
	    RECT 337.3000 119.7000 339.5000 120.3000 ;
	    RECT 314.8000 117.6000 315.6000 118.4000 ;
	    RECT 316.4000 117.6000 317.2000 118.4000 ;
	    RECT 332.4000 117.6000 333.2000 118.4000 ;
	    RECT 334.0000 117.6000 334.8000 118.4000 ;
	    RECT 286.0000 109.6000 286.8000 110.4000 ;
	    RECT 287.6000 109.6000 288.4000 110.4000 ;
	    RECT 289.2000 109.6000 290.0000 110.4000 ;
	    RECT 290.8000 109.6000 291.6000 110.4000 ;
	    RECT 295.6000 109.6000 296.4000 110.4000 ;
	    RECT 297.2000 109.6000 298.0000 110.4000 ;
	    RECT 300.4000 109.6000 301.2000 110.4000 ;
	    RECT 303.6000 109.6000 304.4000 110.4000 ;
	    RECT 306.8000 109.6000 307.6000 110.4000 ;
	    RECT 311.6000 109.6000 312.4000 110.4000 ;
	    RECT 313.2000 109.6000 314.0000 110.4000 ;
	    RECT 286.1000 106.4000 286.7000 109.6000 ;
	    RECT 295.7000 108.4000 296.3000 109.6000 ;
	    RECT 297.3000 108.4000 297.9000 109.6000 ;
	    RECT 295.6000 107.6000 296.4000 108.4000 ;
	    RECT 297.2000 107.6000 298.0000 108.4000 ;
	    RECT 305.2000 107.6000 306.0000 108.4000 ;
	    RECT 306.8000 107.6000 307.6000 108.4000 ;
	    RECT 310.0000 107.6000 310.8000 108.4000 ;
	    RECT 286.0000 105.6000 286.8000 106.4000 ;
	    RECT 295.6000 105.6000 296.4000 106.4000 ;
	    RECT 295.7000 100.4000 296.3000 105.6000 ;
	    RECT 295.6000 99.6000 296.4000 100.4000 ;
	    RECT 284.5000 95.7000 286.7000 96.3000 ;
	    RECT 284.4000 93.6000 285.2000 94.4000 ;
	    RECT 286.1000 92.4000 286.7000 95.7000 ;
	    RECT 287.6000 93.6000 288.4000 94.4000 ;
	    RECT 290.8000 94.3000 291.6000 94.4000 ;
	    RECT 290.8000 93.7000 294.7000 94.3000 ;
	    RECT 290.8000 93.6000 291.6000 93.7000 ;
	    RECT 282.8000 91.6000 283.6000 92.4000 ;
	    RECT 286.0000 91.6000 286.8000 92.4000 ;
	    RECT 289.2000 91.6000 290.0000 92.4000 ;
	    RECT 279.6000 89.6000 280.4000 90.4000 ;
	    RECT 281.2000 89.6000 282.0000 90.4000 ;
	    RECT 279.7000 84.3000 280.3000 89.6000 ;
	    RECT 281.3000 86.4000 281.9000 89.6000 ;
	    RECT 289.3000 86.4000 289.9000 91.6000 ;
	    RECT 294.1000 90.3000 294.7000 93.7000 ;
	    RECT 295.7000 92.4000 296.3000 99.6000 ;
	    RECT 295.6000 91.6000 296.4000 92.4000 ;
	    RECT 295.6000 90.3000 296.4000 90.4000 ;
	    RECT 294.1000 89.7000 296.4000 90.3000 ;
	    RECT 295.6000 89.6000 296.4000 89.7000 ;
	    RECT 290.9000 87.7000 294.7000 88.3000 ;
	    RECT 281.2000 85.6000 282.0000 86.4000 ;
	    RECT 289.2000 85.6000 290.0000 86.4000 ;
	    RECT 290.9000 84.3000 291.5000 87.7000 ;
	    RECT 292.4000 85.6000 293.2000 86.4000 ;
	    RECT 294.1000 84.4000 294.7000 87.7000 ;
	    RECT 279.7000 83.7000 291.5000 84.3000 ;
	    RECT 294.0000 83.6000 294.8000 84.4000 ;
	    RECT 297.3000 82.4000 297.9000 107.6000 ;
	    RECT 305.3000 104.4000 305.9000 107.6000 ;
	    RECT 306.9000 106.4000 307.5000 107.6000 ;
	    RECT 306.8000 105.6000 307.6000 106.4000 ;
	    RECT 308.4000 105.6000 309.2000 106.4000 ;
	    RECT 305.2000 103.6000 306.0000 104.4000 ;
	    RECT 302.0000 99.6000 302.8000 100.4000 ;
	    RECT 300.4000 93.6000 301.2000 94.4000 ;
	    RECT 298.8000 90.3000 299.6000 90.4000 ;
	    RECT 300.5000 90.3000 301.1000 93.6000 ;
	    RECT 302.1000 92.4000 302.7000 99.6000 ;
	    RECT 308.5000 92.4000 309.1000 105.6000 ;
	    RECT 310.1000 104.4000 310.7000 107.6000 ;
	    RECT 316.5000 106.4000 317.1000 117.6000 ;
	    RECT 324.4000 113.6000 325.2000 114.4000 ;
	    RECT 324.5000 112.4000 325.1000 113.6000 ;
	    RECT 319.6000 111.6000 320.4000 112.4000 ;
	    RECT 322.8000 111.6000 323.6000 112.4000 ;
	    RECT 324.4000 111.6000 325.2000 112.4000 ;
	    RECT 319.7000 110.4000 320.3000 111.6000 ;
	    RECT 322.9000 110.4000 323.5000 111.6000 ;
	    RECT 319.6000 109.6000 320.4000 110.4000 ;
	    RECT 322.8000 109.6000 323.6000 110.4000 ;
	    RECT 326.0000 109.6000 326.8000 110.4000 ;
	    RECT 318.0000 107.6000 318.8000 108.4000 ;
	    RECT 321.2000 107.6000 322.0000 108.4000 ;
	    RECT 313.2000 105.6000 314.0000 106.4000 ;
	    RECT 316.4000 105.6000 317.2000 106.4000 ;
	    RECT 310.0000 103.6000 310.8000 104.4000 ;
	    RECT 311.6000 103.6000 312.4000 104.4000 ;
	    RECT 310.0000 95.6000 310.8000 96.4000 ;
	    RECT 302.0000 91.6000 302.8000 92.4000 ;
	    RECT 308.4000 91.6000 309.2000 92.4000 ;
	    RECT 310.1000 90.4000 310.7000 95.6000 ;
	    RECT 311.7000 92.4000 312.3000 103.6000 ;
	    RECT 316.5000 96.3000 317.1000 105.6000 ;
	    RECT 318.1000 104.4000 318.7000 107.6000 ;
	    RECT 318.0000 103.6000 318.8000 104.4000 ;
	    RECT 318.0000 96.3000 318.8000 96.4000 ;
	    RECT 316.5000 95.7000 318.8000 96.3000 ;
	    RECT 318.0000 95.6000 318.8000 95.7000 ;
	    RECT 313.2000 93.6000 314.0000 94.4000 ;
	    RECT 314.8000 93.6000 315.6000 94.4000 ;
	    RECT 319.6000 94.3000 320.4000 94.4000 ;
	    RECT 321.3000 94.3000 321.9000 107.6000 ;
	    RECT 326.1000 94.4000 326.7000 109.6000 ;
	    RECT 337.3000 106.4000 337.9000 119.7000 ;
	    RECT 337.2000 105.6000 338.0000 106.4000 ;
	    RECT 338.8000 104.2000 339.6000 115.8000 ;
	    RECT 340.5000 108.4000 341.1000 123.6000 ;
	    RECT 346.9000 122.4000 347.5000 151.6000 ;
	    RECT 348.5000 142.4000 349.1000 165.6000 ;
	    RECT 350.0000 155.6000 350.8000 156.4000 ;
	    RECT 350.1000 150.4000 350.7000 155.6000 ;
	    RECT 351.7000 150.4000 352.3000 169.6000 ;
	    RECT 353.3000 166.4000 353.9000 169.7000 ;
	    RECT 354.8000 169.6000 355.6000 169.7000 ;
	    RECT 369.2000 169.6000 370.0000 170.4000 ;
	    RECT 354.8000 167.6000 355.6000 168.4000 ;
	    RECT 361.2000 167.6000 362.0000 168.4000 ;
	    RECT 362.8000 167.6000 363.6000 168.4000 ;
	    RECT 353.2000 165.6000 354.0000 166.4000 ;
	    RECT 350.0000 149.6000 350.8000 150.4000 ;
	    RECT 351.6000 149.6000 352.4000 150.4000 ;
	    RECT 351.6000 147.6000 352.4000 148.4000 ;
	    RECT 348.4000 141.6000 349.2000 142.4000 ;
	    RECT 348.4000 135.6000 349.2000 136.4000 ;
	    RECT 350.0000 135.6000 350.8000 136.4000 ;
	    RECT 348.5000 124.4000 349.1000 135.6000 ;
	    RECT 350.0000 130.3000 350.8000 130.4000 ;
	    RECT 351.7000 130.3000 352.3000 147.6000 ;
	    RECT 353.2000 143.6000 354.0000 144.4000 ;
	    RECT 354.9000 136.4000 355.5000 167.6000 ;
	    RECT 359.6000 165.6000 360.4000 166.4000 ;
	    RECT 356.4000 149.6000 357.2000 150.4000 ;
	    RECT 358.0000 149.6000 358.8000 150.4000 ;
	    RECT 356.5000 142.4000 357.1000 149.6000 ;
	    RECT 358.1000 148.4000 358.7000 149.6000 ;
	    RECT 359.7000 148.4000 360.3000 165.6000 ;
	    RECT 361.3000 150.4000 361.9000 167.6000 ;
	    RECT 362.9000 150.4000 363.5000 167.6000 ;
	    RECT 364.4000 163.6000 365.2000 164.4000 ;
	    RECT 364.5000 156.4000 365.1000 163.6000 ;
	    RECT 364.4000 155.6000 365.2000 156.4000 ;
	    RECT 366.0000 155.6000 366.8000 156.4000 ;
	    RECT 366.1000 154.4000 366.7000 155.6000 ;
	    RECT 366.0000 153.6000 366.8000 154.4000 ;
	    RECT 364.4000 151.6000 365.2000 152.4000 ;
	    RECT 369.2000 151.6000 370.0000 152.4000 ;
	    RECT 361.2000 149.6000 362.0000 150.4000 ;
	    RECT 362.8000 149.6000 363.6000 150.4000 ;
	    RECT 358.0000 147.6000 358.8000 148.4000 ;
	    RECT 359.6000 147.6000 360.4000 148.4000 ;
	    RECT 356.4000 141.6000 357.2000 142.4000 ;
	    RECT 354.8000 135.6000 355.6000 136.4000 ;
	    RECT 354.8000 133.6000 355.6000 134.4000 ;
	    RECT 350.0000 129.7000 352.3000 130.3000 ;
	    RECT 350.0000 129.6000 350.8000 129.7000 ;
	    RECT 354.9000 126.4000 355.5000 133.6000 ;
	    RECT 356.5000 132.4000 357.1000 141.6000 ;
	    RECT 359.7000 138.3000 360.3000 147.6000 ;
	    RECT 364.5000 140.4000 365.1000 151.6000 ;
	    RECT 372.5000 150.4000 373.1000 171.6000 ;
	    RECT 375.7000 170.4000 376.3000 177.6000 ;
	    RECT 375.6000 169.6000 376.4000 170.4000 ;
	    RECT 374.0000 165.6000 374.8000 166.4000 ;
	    RECT 375.7000 152.4000 376.3000 169.6000 ;
	    RECT 380.5000 166.4000 381.1000 183.6000 ;
	    RECT 380.4000 165.6000 381.2000 166.4000 ;
	    RECT 377.2000 163.6000 378.0000 164.4000 ;
	    RECT 377.3000 158.4000 377.9000 163.6000 ;
	    RECT 377.2000 157.6000 378.0000 158.4000 ;
	    RECT 377.2000 153.6000 378.0000 154.4000 ;
	    RECT 375.6000 151.6000 376.4000 152.4000 ;
	    RECT 375.7000 150.4000 376.3000 151.6000 ;
	    RECT 377.3000 150.4000 377.9000 153.6000 ;
	    RECT 366.0000 149.6000 366.8000 150.4000 ;
	    RECT 372.4000 149.6000 373.2000 150.4000 ;
	    RECT 375.6000 149.6000 376.4000 150.4000 ;
	    RECT 377.2000 149.6000 378.0000 150.4000 ;
	    RECT 366.1000 148.4000 366.7000 149.6000 ;
	    RECT 366.0000 147.6000 366.8000 148.4000 ;
	    RECT 375.6000 147.6000 376.4000 148.4000 ;
	    RECT 374.0000 145.6000 374.8000 146.4000 ;
	    RECT 369.2000 141.6000 370.0000 142.4000 ;
	    RECT 372.4000 141.6000 373.2000 142.4000 ;
	    RECT 364.4000 139.6000 365.2000 140.4000 ;
	    RECT 359.7000 137.7000 361.9000 138.3000 ;
	    RECT 361.3000 136.4000 361.9000 137.7000 ;
	    RECT 359.6000 135.6000 360.4000 136.4000 ;
	    RECT 361.2000 135.6000 362.0000 136.4000 ;
	    RECT 359.7000 132.4000 360.3000 135.6000 ;
	    RECT 361.3000 134.4000 361.9000 135.6000 ;
	    RECT 361.2000 133.6000 362.0000 134.4000 ;
	    RECT 362.8000 133.6000 363.6000 134.4000 ;
	    RECT 362.9000 132.4000 363.5000 133.6000 ;
	    RECT 356.4000 131.6000 357.2000 132.4000 ;
	    RECT 358.0000 131.6000 358.8000 132.4000 ;
	    RECT 359.6000 131.6000 360.4000 132.4000 ;
	    RECT 362.8000 131.6000 363.6000 132.4000 ;
	    RECT 364.4000 131.6000 365.2000 132.4000 ;
	    RECT 356.4000 127.6000 357.2000 128.4000 ;
	    RECT 354.8000 125.6000 355.6000 126.4000 ;
	    RECT 348.4000 123.6000 349.2000 124.4000 ;
	    RECT 356.4000 123.6000 357.2000 124.4000 ;
	    RECT 346.8000 121.6000 347.6000 122.4000 ;
	    RECT 346.8000 111.6000 347.6000 112.4000 ;
	    RECT 346.9000 110.2000 347.5000 111.6000 ;
	    RECT 346.8000 109.4000 347.6000 110.2000 ;
	    RECT 340.4000 107.6000 341.2000 108.4000 ;
	    RECT 346.8000 107.6000 347.6000 108.4000 ;
	    RECT 348.4000 104.2000 349.2000 115.8000 ;
	    RECT 351.6000 106.2000 352.4000 111.8000 ;
	    RECT 354.8000 111.6000 355.6000 112.4000 ;
	    RECT 354.8000 109.6000 355.6000 110.4000 ;
	    RECT 353.2000 107.6000 354.0000 108.4000 ;
	    RECT 353.3000 100.4000 353.9000 107.6000 ;
	    RECT 345.2000 99.6000 346.0000 100.4000 ;
	    RECT 353.2000 99.6000 354.0000 100.4000 ;
	    RECT 345.3000 98.4000 345.9000 99.6000 ;
	    RECT 345.2000 97.6000 346.0000 98.4000 ;
	    RECT 335.6000 95.6000 336.4000 96.4000 ;
	    RECT 351.6000 95.6000 352.4000 96.4000 ;
	    RECT 354.8000 96.3000 355.6000 96.4000 ;
	    RECT 356.5000 96.3000 357.1000 123.6000 ;
	    RECT 358.1000 112.4000 358.7000 131.6000 ;
	    RECT 361.2000 115.6000 362.0000 116.4000 ;
	    RECT 358.0000 111.6000 358.8000 112.4000 ;
	    RECT 359.6000 111.6000 360.4000 112.4000 ;
	    RECT 359.7000 110.4000 360.3000 111.6000 ;
	    RECT 361.3000 110.4000 361.9000 115.6000 ;
	    RECT 362.9000 112.4000 363.5000 131.6000 ;
	    RECT 367.6000 125.6000 368.4000 126.4000 ;
	    RECT 366.0000 123.6000 366.8000 124.4000 ;
	    RECT 366.1000 122.4000 366.7000 123.6000 ;
	    RECT 366.0000 121.6000 366.8000 122.4000 ;
	    RECT 366.0000 113.6000 366.8000 114.4000 ;
	    RECT 362.8000 111.6000 363.6000 112.4000 ;
	    RECT 366.1000 110.4000 366.7000 113.6000 ;
	    RECT 359.6000 109.6000 360.4000 110.4000 ;
	    RECT 361.2000 109.6000 362.0000 110.4000 ;
	    RECT 366.0000 109.6000 366.8000 110.4000 ;
	    RECT 362.8000 103.6000 363.6000 104.4000 ;
	    RECT 362.9000 96.3000 363.5000 103.6000 ;
	    RECT 354.8000 95.7000 357.1000 96.3000 ;
	    RECT 361.3000 95.7000 363.5000 96.3000 ;
	    RECT 354.8000 95.6000 355.6000 95.7000 ;
	    RECT 335.7000 94.4000 336.3000 95.6000 ;
	    RECT 319.6000 93.7000 321.9000 94.3000 ;
	    RECT 319.6000 93.6000 320.4000 93.7000 ;
	    RECT 324.4000 93.6000 325.2000 94.4000 ;
	    RECT 326.0000 93.6000 326.8000 94.4000 ;
	    RECT 330.8000 93.6000 331.6000 94.4000 ;
	    RECT 335.6000 93.6000 336.4000 94.4000 ;
	    RECT 343.6000 93.6000 344.4000 94.4000 ;
	    RECT 311.6000 91.6000 312.4000 92.4000 ;
	    RECT 298.8000 89.7000 301.1000 90.3000 ;
	    RECT 298.8000 89.6000 299.6000 89.7000 ;
	    RECT 308.4000 89.6000 309.2000 90.4000 ;
	    RECT 310.0000 89.6000 310.8000 90.4000 ;
	    RECT 313.3000 86.4000 313.9000 93.6000 ;
	    RECT 314.9000 92.4000 315.5000 93.6000 ;
	    RECT 324.5000 92.4000 325.1000 93.6000 ;
	    RECT 314.8000 91.6000 315.6000 92.4000 ;
	    RECT 322.8000 91.6000 323.6000 92.4000 ;
	    RECT 324.4000 91.6000 325.2000 92.4000 ;
	    RECT 326.0000 91.6000 326.8000 92.4000 ;
	    RECT 330.9000 92.3000 331.5000 93.6000 ;
	    RECT 343.7000 92.4000 344.3000 93.6000 ;
	    RECT 351.7000 92.4000 352.3000 95.6000 ;
	    RECT 356.4000 93.6000 357.2000 94.4000 ;
	    RECT 356.5000 92.4000 357.1000 93.6000 ;
	    RECT 361.3000 92.4000 361.9000 95.7000 ;
	    RECT 362.8000 93.6000 363.6000 94.4000 ;
	    RECT 364.4000 93.6000 365.2000 94.4000 ;
	    RECT 364.5000 92.4000 365.1000 93.6000 ;
	    RECT 367.7000 92.4000 368.3000 125.6000 ;
	    RECT 369.3000 110.4000 369.9000 141.6000 ;
	    RECT 370.8000 137.6000 371.6000 138.4000 ;
	    RECT 370.9000 132.4000 371.5000 137.6000 ;
	    RECT 372.5000 132.4000 373.1000 141.6000 ;
	    RECT 374.1000 132.4000 374.7000 145.6000 ;
	    RECT 375.7000 142.4000 376.3000 147.6000 ;
	    RECT 375.6000 141.6000 376.4000 142.4000 ;
	    RECT 370.8000 131.6000 371.6000 132.4000 ;
	    RECT 372.4000 131.6000 373.2000 132.4000 ;
	    RECT 374.0000 131.6000 374.8000 132.4000 ;
	    RECT 375.7000 130.3000 376.3000 141.6000 ;
	    RECT 377.2000 139.6000 378.0000 140.4000 ;
	    RECT 377.3000 138.4000 377.9000 139.6000 ;
	    RECT 377.2000 137.6000 378.0000 138.4000 ;
	    RECT 378.8000 137.6000 379.6000 138.4000 ;
	    RECT 378.9000 132.4000 379.5000 137.6000 ;
	    RECT 378.8000 131.6000 379.6000 132.4000 ;
	    RECT 374.1000 129.7000 376.3000 130.3000 ;
	    RECT 370.8000 115.6000 371.6000 116.4000 ;
	    RECT 370.9000 110.4000 371.5000 115.6000 ;
	    RECT 369.2000 109.6000 370.0000 110.4000 ;
	    RECT 370.8000 109.6000 371.6000 110.4000 ;
	    RECT 372.4000 105.6000 373.2000 106.4000 ;
	    RECT 374.1000 100.4000 374.7000 129.7000 ;
	    RECT 377.2000 129.6000 378.0000 130.4000 ;
	    RECT 375.6000 113.6000 376.4000 114.4000 ;
	    RECT 375.7000 110.4000 376.3000 113.6000 ;
	    RECT 375.6000 109.6000 376.4000 110.4000 ;
	    RECT 375.6000 107.6000 376.4000 108.4000 ;
	    RECT 374.0000 99.6000 374.8000 100.4000 ;
	    RECT 375.7000 94.4000 376.3000 107.6000 ;
	    RECT 369.2000 93.6000 370.0000 94.4000 ;
	    RECT 375.6000 93.6000 376.4000 94.4000 ;
	    RECT 332.4000 92.3000 333.2000 92.4000 ;
	    RECT 330.9000 91.7000 333.2000 92.3000 ;
	    RECT 332.4000 91.6000 333.2000 91.7000 ;
	    RECT 334.0000 91.6000 334.8000 92.4000 ;
	    RECT 338.8000 91.6000 339.6000 92.4000 ;
	    RECT 343.6000 91.6000 344.4000 92.4000 ;
	    RECT 348.4000 91.6000 349.2000 92.4000 ;
	    RECT 350.0000 91.6000 350.8000 92.4000 ;
	    RECT 351.6000 91.6000 352.4000 92.4000 ;
	    RECT 356.4000 91.6000 357.2000 92.4000 ;
	    RECT 361.2000 91.6000 362.0000 92.4000 ;
	    RECT 364.4000 91.6000 365.2000 92.4000 ;
	    RECT 367.6000 91.6000 368.4000 92.4000 ;
	    RECT 313.2000 85.6000 314.0000 86.4000 ;
	    RECT 302.0000 83.6000 302.8000 84.4000 ;
	    RECT 303.6000 83.6000 304.4000 84.4000 ;
	    RECT 297.2000 81.6000 298.0000 82.4000 ;
	    RECT 274.8000 79.6000 275.6000 80.4000 ;
	    RECT 276.4000 79.6000 277.2000 80.4000 ;
	    RECT 278.0000 79.6000 278.8000 80.4000 ;
	    RECT 274.9000 78.3000 275.5000 79.6000 ;
	    RECT 274.9000 77.7000 280.3000 78.3000 ;
	    RECT 279.7000 76.4000 280.3000 77.7000 ;
	    RECT 278.0000 75.6000 278.8000 76.4000 ;
	    RECT 279.6000 75.6000 280.4000 76.4000 ;
	    RECT 290.8000 76.3000 291.6000 76.4000 ;
	    RECT 274.8000 71.6000 275.6000 72.4000 ;
	    RECT 276.4000 71.6000 277.2000 72.4000 ;
	    RECT 274.8000 70.3000 275.6000 70.4000 ;
	    RECT 276.5000 70.3000 277.1000 71.6000 ;
	    RECT 274.8000 69.7000 277.1000 70.3000 ;
	    RECT 274.8000 69.6000 275.6000 69.7000 ;
	    RECT 278.1000 68.4000 278.7000 75.6000 ;
	    RECT 284.4000 69.6000 285.2000 70.4000 ;
	    RECT 270.0000 67.6000 270.8000 68.4000 ;
	    RECT 271.6000 67.6000 272.4000 68.4000 ;
	    RECT 273.2000 67.6000 274.0000 68.4000 ;
	    RECT 278.0000 67.6000 278.8000 68.4000 ;
	    RECT 279.6000 67.6000 280.4000 68.4000 ;
	    RECT 265.2000 65.6000 266.0000 66.4000 ;
	    RECT 268.4000 65.6000 269.2000 66.4000 ;
	    RECT 274.8000 65.6000 275.6000 66.4000 ;
	    RECT 278.0000 65.6000 278.8000 66.4000 ;
	    RECT 265.3000 60.4000 265.9000 65.6000 ;
	    RECT 266.8000 63.6000 267.6000 64.4000 ;
	    RECT 265.2000 59.6000 266.0000 60.4000 ;
	    RECT 262.0000 57.6000 262.8000 58.4000 ;
	    RECT 263.6000 57.6000 264.4000 58.4000 ;
	    RECT 266.9000 56.4000 267.5000 63.6000 ;
	    RECT 260.4000 55.6000 261.2000 56.4000 ;
	    RECT 266.8000 55.6000 267.6000 56.4000 ;
	    RECT 260.5000 54.4000 261.1000 55.6000 ;
	    RECT 252.4000 53.6000 253.2000 54.4000 ;
	    RECT 254.0000 53.6000 254.8000 54.4000 ;
	    RECT 260.4000 53.6000 261.2000 54.4000 ;
	    RECT 265.2000 53.6000 266.0000 54.4000 ;
	    RECT 250.8000 51.6000 251.6000 52.4000 ;
	    RECT 249.2000 49.6000 250.0000 50.4000 ;
	    RECT 249.3000 46.4000 249.9000 49.6000 ;
	    RECT 249.2000 45.6000 250.0000 46.4000 ;
	    RECT 250.9000 30.4000 251.5000 51.6000 ;
	    RECT 254.1000 42.4000 254.7000 53.6000 ;
	    RECT 263.6000 49.6000 264.4000 50.4000 ;
	    RECT 257.2000 47.6000 258.0000 48.4000 ;
	    RECT 254.0000 41.6000 254.8000 42.4000 ;
	    RECT 257.3000 34.4000 257.9000 47.6000 ;
	    RECT 263.7000 46.4000 264.3000 49.6000 ;
	    RECT 265.3000 48.4000 265.9000 53.6000 ;
	    RECT 266.8000 51.6000 267.6000 52.4000 ;
	    RECT 270.0000 51.6000 270.8000 52.4000 ;
	    RECT 265.2000 47.6000 266.0000 48.4000 ;
	    RECT 263.6000 45.6000 264.4000 46.4000 ;
	    RECT 262.0000 41.6000 262.8000 42.4000 ;
	    RECT 263.6000 41.6000 264.4000 42.4000 ;
	    RECT 260.4000 35.6000 261.2000 36.4000 ;
	    RECT 257.2000 33.6000 258.0000 34.4000 ;
	    RECT 260.4000 33.6000 261.2000 34.4000 ;
	    RECT 249.2000 29.6000 250.0000 30.4000 ;
	    RECT 250.8000 29.6000 251.6000 30.4000 ;
	    RECT 249.3000 16.4000 249.9000 29.6000 ;
	    RECT 250.9000 20.4000 251.5000 29.6000 ;
	    RECT 257.3000 28.4000 257.9000 33.6000 ;
	    RECT 260.5000 30.4000 261.1000 33.6000 ;
	    RECT 260.4000 29.6000 261.2000 30.4000 ;
	    RECT 257.2000 27.6000 258.0000 28.4000 ;
	    RECT 262.1000 22.4000 262.7000 41.6000 ;
	    RECT 263.7000 34.4000 264.3000 41.6000 ;
	    RECT 266.9000 36.4000 267.5000 51.6000 ;
	    RECT 270.1000 50.4000 270.7000 51.6000 ;
	    RECT 268.4000 49.6000 269.2000 50.4000 ;
	    RECT 270.0000 49.6000 270.8000 50.4000 ;
	    RECT 273.2000 49.6000 274.0000 50.4000 ;
	    RECT 273.3000 48.4000 273.9000 49.6000 ;
	    RECT 271.6000 47.6000 272.4000 48.4000 ;
	    RECT 273.2000 47.6000 274.0000 48.4000 ;
	    RECT 266.8000 35.6000 267.6000 36.4000 ;
	    RECT 263.6000 33.6000 264.4000 34.4000 ;
	    RECT 265.2000 33.6000 266.0000 34.4000 ;
	    RECT 270.0000 33.6000 270.8000 34.4000 ;
	    RECT 263.6000 29.6000 264.4000 30.4000 ;
	    RECT 265.3000 28.4000 265.9000 33.6000 ;
	    RECT 270.1000 30.4000 270.7000 33.6000 ;
	    RECT 271.7000 32.4000 272.3000 47.6000 ;
	    RECT 274.9000 44.3000 275.5000 65.6000 ;
	    RECT 276.4000 61.6000 277.2000 62.4000 ;
	    RECT 276.5000 52.4000 277.1000 61.6000 ;
	    RECT 278.1000 54.4000 278.7000 65.6000 ;
	    RECT 279.7000 58.4000 280.3000 67.6000 ;
	    RECT 284.5000 66.4000 285.1000 69.6000 ;
	    RECT 281.2000 65.6000 282.0000 66.4000 ;
	    RECT 284.4000 65.6000 285.2000 66.4000 ;
	    RECT 286.0000 66.2000 286.8000 71.8000 ;
	    RECT 287.6000 67.6000 288.4000 68.4000 ;
	    RECT 281.3000 64.4000 281.9000 65.6000 ;
	    RECT 281.2000 63.6000 282.0000 64.4000 ;
	    RECT 281.3000 60.4000 281.9000 63.6000 ;
	    RECT 281.2000 59.6000 282.0000 60.4000 ;
	    RECT 279.6000 57.6000 280.4000 58.4000 ;
	    RECT 282.8000 57.6000 283.6000 58.4000 ;
	    RECT 278.0000 53.6000 278.8000 54.4000 ;
	    RECT 282.9000 52.4000 283.5000 57.6000 ;
	    RECT 276.4000 51.6000 277.2000 52.4000 ;
	    RECT 278.1000 51.7000 281.9000 52.3000 ;
	    RECT 278.1000 50.4000 278.7000 51.7000 ;
	    RECT 278.0000 49.6000 278.8000 50.4000 ;
	    RECT 279.6000 49.6000 280.4000 50.4000 ;
	    RECT 281.3000 50.3000 281.9000 51.7000 ;
	    RECT 282.8000 51.6000 283.6000 52.4000 ;
	    RECT 284.5000 52.3000 285.1000 65.6000 ;
	    RECT 287.7000 64.3000 288.3000 67.6000 ;
	    RECT 286.1000 63.7000 288.3000 64.3000 ;
	    RECT 289.2000 64.2000 290.0000 75.8000 ;
	    RECT 290.8000 75.7000 294.7000 76.3000 ;
	    RECT 290.8000 75.6000 291.6000 75.7000 ;
	    RECT 294.1000 72.4000 294.7000 75.7000 ;
	    RECT 294.0000 71.6000 294.8000 72.4000 ;
	    RECT 290.9000 70.2000 291.5000 70.3000 ;
	    RECT 290.8000 69.4000 291.6000 70.2000 ;
	    RECT 286.1000 54.4000 286.7000 63.7000 ;
	    RECT 290.9000 56.4000 291.5000 69.4000 ;
	    RECT 294.0000 67.6000 294.8000 68.4000 ;
	    RECT 289.2000 55.6000 290.0000 56.4000 ;
	    RECT 290.8000 55.6000 291.6000 56.4000 ;
	    RECT 286.0000 53.6000 286.8000 54.4000 ;
	    RECT 286.0000 52.3000 286.8000 52.4000 ;
	    RECT 284.5000 51.7000 286.8000 52.3000 ;
	    RECT 286.0000 51.6000 286.8000 51.7000 ;
	    RECT 286.1000 50.3000 286.7000 51.6000 ;
	    RECT 281.3000 49.7000 285.1000 50.3000 ;
	    RECT 286.1000 49.7000 288.3000 50.3000 ;
	    RECT 284.5000 48.3000 285.1000 49.7000 ;
	    RECT 286.0000 48.3000 286.8000 48.4000 ;
	    RECT 284.5000 47.7000 286.8000 48.3000 ;
	    RECT 286.0000 47.6000 286.8000 47.7000 ;
	    RECT 281.2000 45.6000 282.0000 46.4000 ;
	    RECT 274.9000 43.7000 277.1000 44.3000 ;
	    RECT 271.6000 31.6000 272.4000 32.4000 ;
	    RECT 276.5000 30.4000 277.1000 43.7000 ;
	    RECT 279.6000 33.6000 280.4000 34.4000 ;
	    RECT 266.8000 29.6000 267.6000 30.4000 ;
	    RECT 268.4000 29.6000 269.2000 30.4000 ;
	    RECT 270.0000 29.6000 270.8000 30.4000 ;
	    RECT 274.8000 29.6000 275.6000 30.4000 ;
	    RECT 276.4000 29.6000 277.2000 30.4000 ;
	    RECT 265.2000 27.6000 266.0000 28.4000 ;
	    RECT 263.6000 25.6000 264.4000 26.4000 ;
	    RECT 262.0000 21.6000 262.8000 22.4000 ;
	    RECT 250.8000 19.6000 251.6000 20.4000 ;
	    RECT 262.1000 18.4000 262.7000 21.6000 ;
	    RECT 263.7000 18.4000 264.3000 25.6000 ;
	    RECT 249.2000 15.6000 250.0000 16.4000 ;
	    RECT 247.6000 11.6000 248.4000 12.4000 ;
	    RECT 244.4000 9.6000 245.2000 10.4000 ;
	    RECT 252.4000 6.2000 253.2000 17.8000 ;
	    RECT 262.0000 17.6000 262.8000 18.4000 ;
	    RECT 263.6000 17.6000 264.4000 18.4000 ;
	    RECT 266.9000 10.4000 267.5000 29.6000 ;
	    RECT 276.4000 27.6000 277.2000 28.4000 ;
	    RECT 278.0000 27.6000 278.8000 28.4000 ;
	    RECT 270.0000 25.6000 270.8000 26.4000 ;
	    RECT 270.1000 20.4000 270.7000 25.6000 ;
	    RECT 270.0000 19.6000 270.8000 20.4000 ;
	    RECT 270.0000 17.6000 270.8000 18.4000 ;
	    RECT 270.1000 16.4000 270.7000 17.6000 ;
	    RECT 270.0000 15.6000 270.8000 16.4000 ;
	    RECT 266.8000 9.6000 267.6000 10.4000 ;
	    RECT 274.8000 6.2000 275.6000 17.8000 ;
	    RECT 124.4000 3.6000 125.2000 4.4000 ;
	    RECT 276.5000 2.4000 277.1000 27.6000 ;
	    RECT 278.1000 24.4000 278.7000 27.6000 ;
	    RECT 278.0000 23.6000 278.8000 24.4000 ;
	    RECT 278.0000 15.6000 278.8000 16.4000 ;
	    RECT 278.1000 12.4000 278.7000 15.6000 ;
	    RECT 278.0000 11.6000 278.8000 12.4000 ;
	    RECT 278.1000 8.4000 278.7000 11.6000 ;
	    RECT 279.7000 10.4000 280.3000 33.6000 ;
	    RECT 281.3000 32.4000 281.9000 45.6000 ;
	    RECT 281.2000 31.6000 282.0000 32.4000 ;
	    RECT 282.8000 24.2000 283.6000 35.8000 ;
	    RECT 287.7000 34.4000 288.3000 49.7000 ;
	    RECT 289.3000 34.4000 289.9000 55.6000 ;
	    RECT 294.1000 54.4000 294.7000 67.6000 ;
	    RECT 295.6000 59.6000 296.4000 60.4000 ;
	    RECT 290.8000 53.6000 291.6000 54.4000 ;
	    RECT 294.0000 53.6000 294.8000 54.4000 ;
	    RECT 290.9000 50.4000 291.5000 53.6000 ;
	    RECT 295.7000 52.4000 296.3000 59.6000 ;
	    RECT 292.4000 52.3000 293.2000 52.4000 ;
	    RECT 292.4000 51.7000 294.7000 52.3000 ;
	    RECT 292.4000 51.6000 293.2000 51.7000 ;
	    RECT 290.8000 49.6000 291.6000 50.4000 ;
	    RECT 290.8000 45.6000 291.6000 46.4000 ;
	    RECT 287.6000 33.6000 288.4000 34.4000 ;
	    RECT 289.2000 33.6000 290.0000 34.4000 ;
	    RECT 286.0000 29.6000 286.8000 30.4000 ;
	    RECT 289.2000 29.6000 290.0000 30.4000 ;
	    RECT 282.8000 11.8000 283.6000 12.6000 ;
	    RECT 279.6000 9.6000 280.4000 10.4000 ;
	    RECT 282.9000 8.4000 283.5000 11.8000 ;
	    RECT 278.0000 7.6000 278.8000 8.4000 ;
	    RECT 282.8000 7.6000 283.6000 8.4000 ;
	    RECT 284.4000 6.2000 285.2000 17.8000 ;
	    RECT 286.1000 16.4000 286.7000 29.6000 ;
	    RECT 290.9000 28.4000 291.5000 45.6000 ;
	    RECT 292.4000 43.6000 293.2000 44.4000 ;
	    RECT 292.5000 40.4000 293.1000 43.6000 ;
	    RECT 294.1000 40.4000 294.7000 51.7000 ;
	    RECT 295.6000 51.6000 296.4000 52.4000 ;
	    RECT 297.3000 50.4000 297.9000 81.6000 ;
	    RECT 303.7000 80.4000 304.3000 83.6000 ;
	    RECT 303.6000 79.6000 304.4000 80.4000 ;
	    RECT 298.8000 64.2000 299.6000 75.8000 ;
	    RECT 305.2000 71.6000 306.0000 72.4000 ;
	    RECT 306.8000 71.6000 307.6000 72.4000 ;
	    RECT 305.3000 68.4000 305.9000 71.6000 ;
	    RECT 306.9000 70.4000 307.5000 71.6000 ;
	    RECT 313.3000 70.4000 313.9000 85.6000 ;
	    RECT 314.8000 79.6000 315.6000 80.4000 ;
	    RECT 314.9000 72.4000 315.5000 79.6000 ;
	    RECT 318.0000 75.6000 318.8000 76.4000 ;
	    RECT 314.8000 71.6000 315.6000 72.4000 ;
	    RECT 316.4000 71.6000 317.2000 72.4000 ;
	    RECT 321.2000 71.6000 322.0000 72.4000 ;
	    RECT 314.9000 70.4000 315.5000 71.6000 ;
	    RECT 306.8000 69.6000 307.6000 70.4000 ;
	    RECT 311.6000 69.6000 312.4000 70.4000 ;
	    RECT 313.2000 69.6000 314.0000 70.4000 ;
	    RECT 314.8000 69.6000 315.6000 70.4000 ;
	    RECT 311.7000 68.4000 312.3000 69.6000 ;
	    RECT 316.5000 68.4000 317.1000 71.6000 ;
	    RECT 321.3000 70.4000 321.9000 71.6000 ;
	    RECT 326.1000 70.4000 326.7000 91.6000 ;
	    RECT 327.6000 77.6000 328.4000 78.4000 ;
	    RECT 321.2000 69.6000 322.0000 70.4000 ;
	    RECT 322.8000 69.6000 323.6000 70.4000 ;
	    RECT 326.0000 69.6000 326.8000 70.4000 ;
	    RECT 326.1000 68.4000 326.7000 69.6000 ;
	    RECT 303.6000 67.6000 304.4000 68.4000 ;
	    RECT 305.2000 67.6000 306.0000 68.4000 ;
	    RECT 311.6000 67.6000 312.4000 68.4000 ;
	    RECT 316.4000 67.6000 317.2000 68.4000 ;
	    RECT 324.4000 67.6000 325.2000 68.4000 ;
	    RECT 326.0000 67.6000 326.8000 68.4000 ;
	    RECT 303.7000 64.4000 304.3000 67.6000 ;
	    RECT 311.6000 65.6000 312.4000 66.4000 ;
	    RECT 303.6000 63.6000 304.4000 64.4000 ;
	    RECT 300.4000 61.6000 301.2000 62.4000 ;
	    RECT 297.2000 50.3000 298.0000 50.4000 ;
	    RECT 298.8000 50.3000 299.6000 50.4000 ;
	    RECT 297.2000 49.7000 299.6000 50.3000 ;
	    RECT 297.2000 49.6000 298.0000 49.7000 ;
	    RECT 298.8000 49.6000 299.6000 49.7000 ;
	    RECT 292.4000 39.6000 293.2000 40.4000 ;
	    RECT 294.0000 39.6000 294.8000 40.4000 ;
	    RECT 300.5000 36.4000 301.1000 61.6000 ;
	    RECT 306.8000 59.6000 307.6000 60.4000 ;
	    RECT 308.4000 59.6000 309.2000 60.4000 ;
	    RECT 306.9000 58.4000 307.5000 59.6000 ;
	    RECT 302.0000 57.6000 302.8000 58.4000 ;
	    RECT 306.8000 57.6000 307.6000 58.4000 ;
	    RECT 302.1000 54.4000 302.7000 57.6000 ;
	    RECT 308.5000 56.4000 309.1000 59.6000 ;
	    RECT 303.6000 55.6000 304.4000 56.4000 ;
	    RECT 305.2000 55.6000 306.0000 56.4000 ;
	    RECT 308.4000 55.6000 309.2000 56.4000 ;
	    RECT 302.0000 53.6000 302.8000 54.4000 ;
	    RECT 302.1000 52.4000 302.7000 53.6000 ;
	    RECT 303.7000 52.4000 304.3000 55.6000 ;
	    RECT 305.3000 54.4000 305.9000 55.6000 ;
	    RECT 305.2000 53.6000 306.0000 54.4000 ;
	    RECT 310.0000 53.6000 310.8000 54.4000 ;
	    RECT 310.1000 52.4000 310.7000 53.6000 ;
	    RECT 311.7000 52.4000 312.3000 65.6000 ;
	    RECT 321.2000 57.6000 322.0000 58.4000 ;
	    RECT 327.7000 58.3000 328.3000 77.6000 ;
	    RECT 330.8000 71.6000 331.6000 72.4000 ;
	    RECT 330.9000 68.4000 331.5000 71.6000 ;
	    RECT 332.5000 70.4000 333.1000 91.6000 ;
	    RECT 334.1000 74.4000 334.7000 91.6000 ;
	    RECT 334.0000 73.6000 334.8000 74.4000 ;
	    RECT 335.6000 73.6000 336.4000 74.4000 ;
	    RECT 335.7000 72.4000 336.3000 73.6000 ;
	    RECT 335.6000 71.6000 336.4000 72.4000 ;
	    RECT 332.4000 70.3000 333.2000 70.4000 ;
	    RECT 332.4000 69.7000 334.7000 70.3000 ;
	    RECT 332.4000 69.6000 333.2000 69.7000 ;
	    RECT 330.8000 67.6000 331.6000 68.4000 ;
	    RECT 332.4000 67.6000 333.2000 68.4000 ;
	    RECT 329.2000 66.3000 330.0000 66.4000 ;
	    RECT 332.5000 66.3000 333.1000 67.6000 ;
	    RECT 329.2000 65.7000 333.1000 66.3000 ;
	    RECT 329.2000 65.6000 330.0000 65.7000 ;
	    RECT 332.4000 59.6000 333.2000 60.4000 ;
	    RECT 327.7000 57.7000 329.9000 58.3000 ;
	    RECT 318.0000 55.6000 318.8000 56.4000 ;
	    RECT 318.1000 52.4000 318.7000 55.6000 ;
	    RECT 321.3000 52.4000 321.9000 57.6000 ;
	    RECT 324.4000 56.3000 325.2000 56.4000 ;
	    RECT 322.9000 55.7000 325.2000 56.3000 ;
	    RECT 302.0000 51.6000 302.8000 52.4000 ;
	    RECT 303.6000 51.6000 304.4000 52.4000 ;
	    RECT 310.0000 51.6000 310.8000 52.4000 ;
	    RECT 311.6000 51.6000 312.4000 52.4000 ;
	    RECT 318.0000 51.6000 318.8000 52.4000 ;
	    RECT 321.2000 51.6000 322.0000 52.4000 ;
	    RECT 311.7000 48.4000 312.3000 51.6000 ;
	    RECT 314.8000 49.6000 315.6000 50.4000 ;
	    RECT 318.0000 49.6000 318.8000 50.4000 ;
	    RECT 302.0000 47.6000 302.8000 48.4000 ;
	    RECT 311.6000 47.6000 312.4000 48.4000 ;
	    RECT 290.8000 27.6000 291.6000 28.4000 ;
	    RECT 292.4000 24.2000 293.2000 35.8000 ;
	    RECT 300.4000 35.6000 301.2000 36.4000 ;
	    RECT 295.6000 26.2000 296.4000 31.8000 ;
	    RECT 300.4000 31.6000 301.2000 32.4000 ;
	    RECT 300.5000 30.4000 301.1000 31.6000 ;
	    RECT 298.8000 29.6000 299.6000 30.4000 ;
	    RECT 300.4000 29.6000 301.2000 30.4000 ;
	    RECT 297.2000 27.6000 298.0000 28.4000 ;
	    RECT 286.0000 15.6000 286.8000 16.4000 ;
	    RECT 286.0000 11.6000 286.8000 12.4000 ;
	    RECT 286.1000 8.4000 286.7000 11.6000 ;
	    RECT 287.6000 10.2000 288.4000 15.8000 ;
	    RECT 289.2000 13.6000 290.0000 14.4000 ;
	    RECT 294.0000 13.6000 294.8000 14.4000 ;
	    RECT 297.3000 14.3000 297.9000 27.6000 ;
	    RECT 302.1000 16.4000 302.7000 47.6000 ;
	    RECT 313.2000 45.6000 314.0000 46.4000 ;
	    RECT 308.4000 39.6000 309.2000 40.4000 ;
	    RECT 303.6000 31.6000 304.4000 32.4000 ;
	    RECT 306.8000 31.6000 307.6000 32.4000 ;
	    RECT 303.7000 28.4000 304.3000 31.6000 ;
	    RECT 306.9000 30.4000 307.5000 31.6000 ;
	    RECT 306.8000 29.6000 307.6000 30.4000 ;
	    RECT 308.5000 30.3000 309.1000 39.6000 ;
	    RECT 311.6000 35.6000 312.4000 36.4000 ;
	    RECT 311.7000 30.4000 312.3000 35.6000 ;
	    RECT 308.5000 29.7000 310.7000 30.3000 ;
	    RECT 310.1000 28.4000 310.7000 29.7000 ;
	    RECT 311.6000 29.6000 312.4000 30.4000 ;
	    RECT 303.6000 27.6000 304.4000 28.4000 ;
	    RECT 308.4000 27.6000 309.2000 28.4000 ;
	    RECT 310.0000 27.6000 310.8000 28.4000 ;
	    RECT 308.5000 24.4000 309.1000 27.6000 ;
	    RECT 308.4000 23.6000 309.2000 24.4000 ;
	    RECT 302.0000 15.6000 302.8000 16.4000 ;
	    RECT 298.8000 14.3000 299.6000 14.4000 ;
	    RECT 297.3000 13.7000 299.6000 14.3000 ;
	    RECT 298.8000 13.6000 299.6000 13.7000 ;
	    RECT 292.4000 11.6000 293.2000 12.4000 ;
	    RECT 297.2000 11.6000 298.0000 12.4000 ;
	    RECT 300.4000 11.6000 301.2000 12.4000 ;
	    RECT 292.5000 10.4000 293.1000 11.6000 ;
	    RECT 292.4000 9.6000 293.2000 10.4000 ;
	    RECT 300.5000 8.4000 301.1000 11.6000 ;
	    RECT 286.0000 7.6000 286.8000 8.4000 ;
	    RECT 300.4000 7.6000 301.2000 8.4000 ;
	    RECT 305.2000 6.2000 306.0000 17.8000 ;
	    RECT 313.3000 16.4000 313.9000 45.6000 ;
	    RECT 314.9000 26.4000 315.5000 49.6000 ;
	    RECT 322.9000 34.4000 323.5000 55.7000 ;
	    RECT 324.4000 55.6000 325.2000 55.7000 ;
	    RECT 326.0000 55.6000 326.8000 56.4000 ;
	    RECT 327.6000 55.6000 328.4000 56.4000 ;
	    RECT 324.4000 53.6000 325.2000 54.4000 ;
	    RECT 316.5000 33.7000 321.9000 34.3000 ;
	    RECT 316.5000 32.4000 317.1000 33.7000 ;
	    RECT 316.4000 31.6000 317.2000 32.4000 ;
	    RECT 318.0000 31.6000 318.8000 32.4000 ;
	    RECT 321.3000 32.3000 321.9000 33.7000 ;
	    RECT 322.8000 33.6000 323.6000 34.4000 ;
	    RECT 324.5000 32.4000 325.1000 53.6000 ;
	    RECT 327.7000 52.4000 328.3000 55.6000 ;
	    RECT 327.6000 51.6000 328.4000 52.4000 ;
	    RECT 329.3000 50.4000 329.9000 57.7000 ;
	    RECT 332.5000 56.4000 333.1000 59.6000 ;
	    RECT 332.4000 55.6000 333.2000 56.4000 ;
	    RECT 334.1000 54.4000 334.7000 69.7000 ;
	    RECT 338.9000 62.4000 339.5000 91.6000 ;
	    RECT 340.4000 64.2000 341.2000 75.8000 ;
	    RECT 348.5000 74.4000 349.1000 91.6000 ;
	    RECT 350.1000 86.4000 350.7000 91.6000 ;
	    RECT 350.0000 85.6000 350.8000 86.4000 ;
	    RECT 348.4000 73.6000 349.2000 74.4000 ;
	    RECT 343.6000 69.6000 344.4000 70.4000 ;
	    RECT 343.7000 68.4000 344.3000 69.6000 ;
	    RECT 343.6000 67.6000 344.4000 68.4000 ;
	    RECT 346.8000 67.6000 347.6000 68.4000 ;
	    RECT 337.2000 61.6000 338.0000 62.4000 ;
	    RECT 338.8000 61.6000 339.6000 62.4000 ;
	    RECT 337.3000 58.4000 337.9000 61.6000 ;
	    RECT 335.6000 57.6000 336.4000 58.4000 ;
	    RECT 337.2000 57.6000 338.0000 58.4000 ;
	    RECT 334.0000 53.6000 334.8000 54.4000 ;
	    RECT 334.1000 52.4000 334.7000 53.6000 ;
	    RECT 335.7000 52.4000 336.3000 57.6000 ;
	    RECT 334.0000 51.6000 334.8000 52.4000 ;
	    RECT 335.6000 51.6000 336.4000 52.4000 ;
	    RECT 329.2000 49.6000 330.0000 50.4000 ;
	    RECT 329.2000 43.6000 330.0000 44.4000 ;
	    RECT 329.3000 34.3000 329.9000 43.6000 ;
	    RECT 326.1000 33.7000 329.9000 34.3000 ;
	    RECT 321.3000 31.7000 323.5000 32.3000 ;
	    RECT 318.1000 30.4000 318.7000 31.6000 ;
	    RECT 316.4000 29.6000 317.2000 30.4000 ;
	    RECT 318.0000 29.6000 318.8000 30.4000 ;
	    RECT 321.2000 29.6000 322.0000 30.4000 ;
	    RECT 314.8000 25.6000 315.6000 26.4000 ;
	    RECT 313.2000 15.6000 314.0000 16.4000 ;
	    RECT 313.2000 11.8000 314.0000 12.6000 ;
	    RECT 313.3000 8.4000 313.9000 11.8000 ;
	    RECT 313.2000 7.6000 314.0000 8.4000 ;
	    RECT 314.8000 6.2000 315.6000 17.8000 ;
	    RECT 316.5000 8.4000 317.1000 29.6000 ;
	    RECT 319.6000 27.6000 320.4000 28.4000 ;
	    RECT 321.3000 22.4000 321.9000 29.6000 ;
	    RECT 322.9000 22.4000 323.5000 31.7000 ;
	    RECT 324.4000 31.6000 325.2000 32.4000 ;
	    RECT 324.5000 26.4000 325.1000 31.6000 ;
	    RECT 326.1000 30.4000 326.7000 33.7000 ;
	    RECT 334.1000 32.4000 334.7000 51.6000 ;
	    RECT 338.9000 44.4000 339.5000 61.6000 ;
	    RECT 342.0000 53.6000 342.8000 54.4000 ;
	    RECT 345.2000 51.6000 346.0000 52.4000 ;
	    RECT 345.3000 50.4000 345.9000 51.6000 ;
	    RECT 345.2000 49.6000 346.0000 50.4000 ;
	    RECT 346.9000 46.4000 347.5000 67.6000 ;
	    RECT 350.0000 64.2000 350.8000 75.8000 ;
	    RECT 350.0000 57.6000 350.8000 58.4000 ;
	    RECT 350.1000 52.4000 350.7000 57.6000 ;
	    RECT 351.7000 56.4000 352.3000 91.6000 ;
	    RECT 369.3000 86.4000 369.9000 93.6000 ;
	    RECT 374.0000 91.6000 374.8000 92.4000 ;
	    RECT 369.2000 85.6000 370.0000 86.4000 ;
	    RECT 358.0000 83.6000 358.8000 84.4000 ;
	    RECT 370.8000 83.6000 371.6000 84.4000 ;
	    RECT 361.2000 81.6000 362.0000 82.4000 ;
	    RECT 359.6000 73.6000 360.4000 74.4000 ;
	    RECT 359.7000 72.4000 360.3000 73.6000 ;
	    RECT 353.2000 66.2000 354.0000 71.8000 ;
	    RECT 359.6000 71.6000 360.4000 72.4000 ;
	    RECT 354.8000 69.6000 355.6000 70.4000 ;
	    RECT 359.6000 67.6000 360.4000 68.4000 ;
	    RECT 359.7000 66.4000 360.3000 67.6000 ;
	    RECT 359.6000 65.6000 360.4000 66.4000 ;
	    RECT 358.0000 63.6000 358.8000 64.4000 ;
	    RECT 351.6000 55.6000 352.4000 56.4000 ;
	    RECT 350.0000 51.6000 350.8000 52.4000 ;
	    RECT 351.6000 51.6000 352.4000 52.4000 ;
	    RECT 353.2000 49.6000 354.0000 50.4000 ;
	    RECT 346.8000 45.6000 347.6000 46.4000 ;
	    RECT 338.8000 43.6000 339.6000 44.4000 ;
	    RECT 337.2000 41.6000 338.0000 42.4000 ;
	    RECT 337.3000 38.4000 337.9000 41.6000 ;
	    RECT 337.2000 37.6000 338.0000 38.4000 ;
	    RECT 343.6000 35.6000 344.4000 36.4000 ;
	    RECT 346.9000 34.4000 347.5000 45.6000 ;
	    RECT 353.3000 36.4000 353.9000 49.6000 ;
	    RECT 358.1000 48.4000 358.7000 63.6000 ;
	    RECT 359.6000 53.6000 360.4000 54.4000 ;
	    RECT 361.3000 52.4000 361.9000 81.6000 ;
	    RECT 362.8000 71.6000 363.6000 72.4000 ;
	    RECT 362.8000 67.6000 363.6000 68.4000 ;
	    RECT 364.4000 65.6000 365.2000 66.4000 ;
	    RECT 364.5000 64.4000 365.1000 65.6000 ;
	    RECT 364.4000 63.6000 365.2000 64.4000 ;
	    RECT 369.2000 64.2000 370.0000 75.8000 ;
	    RECT 370.9000 62.4000 371.5000 83.6000 ;
	    RECT 370.8000 61.6000 371.6000 62.4000 ;
	    RECT 361.2000 51.6000 362.0000 52.4000 ;
	    RECT 369.2000 51.6000 370.0000 52.4000 ;
	    RECT 364.4000 49.6000 365.2000 50.4000 ;
	    RECT 358.0000 47.6000 358.8000 48.4000 ;
	    RECT 361.2000 47.6000 362.0000 48.4000 ;
	    RECT 356.4000 43.6000 357.2000 44.4000 ;
	    RECT 356.5000 36.4000 357.1000 43.6000 ;
	    RECT 346.8000 33.6000 347.6000 34.4000 ;
	    RECT 327.6000 31.6000 328.4000 32.4000 ;
	    RECT 334.0000 31.6000 334.8000 32.4000 ;
	    RECT 326.0000 29.6000 326.8000 30.4000 ;
	    RECT 324.4000 25.6000 325.2000 26.4000 ;
	    RECT 327.7000 22.4000 328.3000 31.6000 ;
	    RECT 334.1000 30.4000 334.7000 31.6000 ;
	    RECT 330.8000 30.3000 331.6000 30.4000 ;
	    RECT 329.3000 29.7000 331.6000 30.3000 ;
	    RECT 329.3000 22.4000 329.9000 29.7000 ;
	    RECT 330.8000 29.6000 331.6000 29.7000 ;
	    RECT 334.0000 29.6000 334.8000 30.4000 ;
	    RECT 335.6000 29.6000 336.4000 30.4000 ;
	    RECT 342.0000 29.6000 342.8000 30.4000 ;
	    RECT 330.8000 27.6000 331.6000 28.4000 ;
	    RECT 332.4000 27.6000 333.2000 28.4000 ;
	    RECT 321.2000 21.6000 322.0000 22.4000 ;
	    RECT 322.8000 21.6000 323.6000 22.4000 ;
	    RECT 327.6000 21.6000 328.4000 22.4000 ;
	    RECT 329.2000 21.6000 330.0000 22.4000 ;
	    RECT 318.0000 10.2000 318.8000 15.8000 ;
	    RECT 330.9000 14.4000 331.5000 27.6000 ;
	    RECT 332.5000 26.4000 333.1000 27.6000 ;
	    RECT 335.7000 26.4000 336.3000 29.6000 ;
	    RECT 332.4000 25.6000 333.2000 26.4000 ;
	    RECT 335.6000 25.6000 336.4000 26.4000 ;
	    RECT 332.5000 14.4000 333.1000 25.6000 ;
	    RECT 342.1000 24.4000 342.7000 29.6000 ;
	    RECT 342.0000 23.6000 342.8000 24.4000 ;
	    RECT 348.4000 24.2000 349.2000 35.8000 ;
	    RECT 353.2000 35.6000 354.0000 36.4000 ;
	    RECT 356.4000 35.6000 357.2000 36.4000 ;
	    RECT 356.4000 31.6000 357.2000 32.4000 ;
	    RECT 356.5000 30.2000 357.1000 31.6000 ;
	    RECT 356.4000 29.4000 357.2000 30.2000 ;
	    RECT 350.0000 25.6000 350.8000 26.4000 ;
	    RECT 353.2000 25.6000 354.0000 26.4000 ;
	    RECT 335.6000 21.6000 336.4000 22.4000 ;
	    RECT 346.8000 21.6000 347.6000 22.4000 ;
	    RECT 348.4000 21.6000 349.2000 22.4000 ;
	    RECT 335.7000 18.4000 336.3000 21.6000 ;
	    RECT 335.6000 17.6000 336.4000 18.4000 ;
	    RECT 345.2000 16.3000 346.0000 16.4000 ;
	    RECT 342.1000 15.7000 346.0000 16.3000 ;
	    RECT 319.6000 13.6000 320.4000 14.4000 ;
	    RECT 324.4000 13.6000 325.2000 14.4000 ;
	    RECT 329.2000 13.6000 330.0000 14.4000 ;
	    RECT 330.8000 13.6000 331.6000 14.4000 ;
	    RECT 332.4000 13.6000 333.2000 14.4000 ;
	    RECT 337.2000 13.6000 338.0000 14.4000 ;
	    RECT 319.7000 12.4000 320.3000 13.6000 ;
	    RECT 330.9000 12.4000 331.5000 13.6000 ;
	    RECT 342.1000 12.4000 342.7000 15.7000 ;
	    RECT 345.2000 15.6000 346.0000 15.7000 ;
	    RECT 343.6000 13.6000 344.4000 14.4000 ;
	    RECT 345.2000 14.3000 346.0000 14.4000 ;
	    RECT 346.9000 14.3000 347.5000 21.6000 ;
	    RECT 348.5000 20.4000 349.1000 21.6000 ;
	    RECT 348.4000 19.6000 349.2000 20.4000 ;
	    RECT 348.5000 16.4000 349.1000 19.6000 ;
	    RECT 348.4000 15.6000 349.2000 16.4000 ;
	    RECT 345.2000 13.7000 347.5000 14.3000 ;
	    RECT 345.2000 13.6000 346.0000 13.7000 ;
	    RECT 343.7000 12.4000 344.3000 13.6000 ;
	    RECT 350.1000 12.4000 350.7000 25.6000 ;
	    RECT 353.3000 18.4000 353.9000 25.6000 ;
	    RECT 358.0000 24.2000 358.8000 35.8000 ;
	    RECT 362.8000 35.6000 363.6000 36.4000 ;
	    RECT 362.9000 32.4000 363.5000 35.6000 ;
	    RECT 359.6000 27.6000 360.4000 28.4000 ;
	    RECT 359.7000 20.4000 360.3000 27.6000 ;
	    RECT 361.2000 26.2000 362.0000 31.8000 ;
	    RECT 362.8000 31.6000 363.6000 32.4000 ;
	    RECT 364.4000 31.6000 365.2000 32.4000 ;
	    RECT 364.5000 30.4000 365.1000 31.6000 ;
	    RECT 369.3000 30.4000 369.9000 51.6000 ;
	    RECT 370.8000 46.2000 371.6000 57.8000 ;
	    RECT 375.7000 54.4000 376.3000 93.6000 ;
	    RECT 377.3000 92.4000 377.9000 129.6000 ;
	    RECT 380.5000 120.4000 381.1000 165.6000 ;
	    RECT 383.7000 162.4000 384.3000 185.6000 ;
	    RECT 386.9000 184.4000 387.5000 187.6000 ;
	    RECT 386.8000 183.6000 387.6000 184.4000 ;
	    RECT 391.6000 184.2000 392.4000 195.8000 ;
	    RECT 394.8000 195.6000 395.6000 196.4000 ;
	    RECT 399.6000 189.4000 400.4000 190.2000 ;
	    RECT 399.7000 182.4000 400.3000 189.4000 ;
	    RECT 401.2000 184.2000 402.0000 195.8000 ;
	    RECT 417.3000 192.4000 417.9000 201.6000 ;
	    RECT 402.8000 187.6000 403.6000 188.4000 ;
	    RECT 399.6000 181.6000 400.4000 182.4000 ;
	    RECT 393.2000 173.6000 394.0000 174.4000 ;
	    RECT 388.4000 171.6000 389.2000 172.4000 ;
	    RECT 383.6000 161.6000 384.4000 162.4000 ;
	    RECT 383.6000 157.6000 384.4000 158.4000 ;
	    RECT 382.0000 144.2000 382.8000 155.8000 ;
	    RECT 383.7000 150.4000 384.3000 157.6000 ;
	    RECT 388.5000 150.4000 389.1000 171.6000 ;
	    RECT 390.0000 169.6000 390.8000 170.4000 ;
	    RECT 391.6000 169.6000 392.4000 170.4000 ;
	    RECT 393.3000 168.4000 393.9000 173.6000 ;
	    RECT 393.2000 167.6000 394.0000 168.4000 ;
	    RECT 396.4000 167.6000 397.2000 168.4000 ;
	    RECT 383.6000 149.6000 384.4000 150.4000 ;
	    RECT 388.4000 149.6000 389.2000 150.4000 ;
	    RECT 383.6000 147.6000 384.4000 148.4000 ;
	    RECT 382.0000 123.6000 382.8000 124.4000 ;
	    RECT 380.4000 119.6000 381.2000 120.4000 ;
	    RECT 378.8000 117.6000 379.6000 118.4000 ;
	    RECT 380.5000 106.4000 381.1000 119.6000 ;
	    RECT 382.1000 108.4000 382.7000 123.6000 ;
	    RECT 383.7000 118.3000 384.3000 147.6000 ;
	    RECT 390.0000 145.6000 390.8000 146.4000 ;
	    RECT 385.2000 143.6000 386.0000 144.4000 ;
	    RECT 385.3000 132.4000 385.9000 143.6000 ;
	    RECT 385.2000 131.6000 386.0000 132.4000 ;
	    RECT 386.8000 127.6000 387.6000 128.4000 ;
	    RECT 386.9000 118.4000 387.5000 127.6000 ;
	    RECT 390.1000 126.3000 390.7000 145.6000 ;
	    RECT 391.6000 144.2000 392.4000 155.8000 ;
	    RECT 393.3000 154.4000 393.9000 167.6000 ;
	    RECT 393.2000 153.6000 394.0000 154.4000 ;
	    RECT 396.5000 152.4000 397.1000 167.6000 ;
	    RECT 399.6000 166.2000 400.4000 177.8000 ;
	    RECT 402.9000 174.4000 403.5000 187.6000 ;
	    RECT 404.4000 186.2000 405.2000 191.8000 ;
	    RECT 417.2000 191.6000 418.0000 192.4000 ;
	    RECT 418.9000 190.4000 419.5000 207.6000 ;
	    RECT 422.0000 206.2000 422.8000 217.8000 ;
	    RECT 428.4000 211.6000 429.2000 212.4000 ;
	    RECT 428.5000 210.4000 429.1000 211.6000 ;
	    RECT 428.4000 209.6000 429.2000 210.4000 ;
	    RECT 430.0000 207.6000 430.8000 208.4000 ;
	    RECT 430.1000 198.4000 430.7000 207.6000 ;
	    RECT 431.6000 206.2000 432.4000 217.8000 ;
	    RECT 433.3000 217.7000 435.5000 218.3000 ;
	    RECT 433.3000 214.4000 433.9000 217.7000 ;
	    RECT 439.6000 217.6000 440.4000 218.4000 ;
	    RECT 433.2000 213.6000 434.0000 214.4000 ;
	    RECT 434.8000 210.2000 435.6000 215.8000 ;
	    RECT 436.4000 215.6000 437.2000 216.4000 ;
	    RECT 441.2000 215.6000 442.0000 216.4000 ;
	    RECT 439.6000 209.6000 440.4000 210.4000 ;
	    RECT 439.7000 198.4000 440.3000 209.6000 ;
	    RECT 430.0000 197.6000 430.8000 198.4000 ;
	    RECT 431.6000 197.6000 432.4000 198.4000 ;
	    RECT 439.6000 197.6000 440.4000 198.4000 ;
	    RECT 423.6000 195.6000 424.4000 196.4000 ;
	    RECT 423.7000 190.4000 424.3000 195.6000 ;
	    RECT 431.7000 194.4000 432.3000 197.6000 ;
	    RECT 438.0000 195.6000 438.8000 196.4000 ;
	    RECT 426.8000 193.6000 427.6000 194.4000 ;
	    RECT 430.0000 193.6000 430.8000 194.4000 ;
	    RECT 431.6000 193.6000 432.4000 194.4000 ;
	    RECT 410.8000 189.6000 411.6000 190.4000 ;
	    RECT 414.0000 189.6000 414.8000 190.4000 ;
	    RECT 418.8000 189.6000 419.6000 190.4000 ;
	    RECT 423.6000 189.6000 424.4000 190.4000 ;
	    RECT 410.9000 188.4000 411.5000 189.6000 ;
	    RECT 410.8000 187.6000 411.6000 188.4000 ;
	    RECT 417.2000 183.6000 418.0000 184.4000 ;
	    RECT 422.0000 183.6000 422.8000 184.4000 ;
	    RECT 417.3000 182.4000 417.9000 183.6000 ;
	    RECT 417.2000 181.6000 418.0000 182.4000 ;
	    RECT 402.8000 173.6000 403.6000 174.4000 ;
	    RECT 407.6000 171.6000 408.4000 172.6000 ;
	    RECT 401.2000 167.6000 402.0000 168.4000 ;
	    RECT 394.8000 146.2000 395.6000 151.8000 ;
	    RECT 396.4000 151.6000 397.2000 152.4000 ;
	    RECT 398.0000 149.6000 398.8000 150.4000 ;
	    RECT 401.3000 148.4000 401.9000 167.6000 ;
	    RECT 409.2000 166.2000 410.0000 177.8000 ;
	    RECT 410.8000 173.6000 411.6000 174.4000 ;
	    RECT 410.9000 166.3000 411.5000 173.6000 ;
	    RECT 412.4000 170.2000 413.2000 175.8000 ;
	    RECT 414.0000 173.6000 414.8000 174.4000 ;
	    RECT 414.1000 172.4000 414.7000 173.6000 ;
	    RECT 414.0000 171.6000 414.8000 172.4000 ;
	    RECT 422.1000 172.3000 422.7000 183.6000 ;
	    RECT 426.9000 178.4000 427.5000 193.6000 ;
	    RECT 430.1000 192.3000 430.7000 193.6000 ;
	    RECT 430.1000 191.7000 432.3000 192.3000 ;
	    RECT 426.8000 177.6000 427.6000 178.4000 ;
	    RECT 425.2000 173.6000 426.0000 174.4000 ;
	    RECT 430.0000 173.6000 430.8000 174.4000 ;
	    RECT 423.6000 172.3000 424.4000 172.4000 ;
	    RECT 422.1000 171.7000 424.4000 172.3000 ;
	    RECT 420.4000 169.6000 421.2000 170.4000 ;
	    RECT 410.9000 165.7000 413.1000 166.3000 ;
	    RECT 409.2000 155.6000 410.0000 156.4000 ;
	    RECT 412.5000 154.4000 413.1000 165.7000 ;
	    RECT 412.4000 153.6000 413.2000 154.4000 ;
	    RECT 402.8000 149.6000 403.6000 150.4000 ;
	    RECT 401.2000 147.6000 402.0000 148.4000 ;
	    RECT 391.6000 135.6000 392.4000 136.4000 ;
	    RECT 391.7000 134.4000 392.3000 135.6000 ;
	    RECT 401.3000 134.4000 401.9000 147.6000 ;
	    RECT 391.6000 133.6000 392.4000 134.4000 ;
	    RECT 401.2000 133.6000 402.0000 134.4000 ;
	    RECT 402.9000 132.4000 403.5000 149.6000 ;
	    RECT 414.0000 144.2000 414.8000 155.8000 ;
	    RECT 420.4000 149.6000 421.2000 150.4000 ;
	    RECT 422.1000 140.4000 422.7000 171.7000 ;
	    RECT 423.6000 171.6000 424.4000 171.7000 ;
	    RECT 425.3000 168.4000 425.9000 173.6000 ;
	    RECT 426.8000 169.6000 427.6000 170.4000 ;
	    RECT 430.0000 169.6000 430.8000 170.4000 ;
	    RECT 425.2000 167.6000 426.0000 168.4000 ;
	    RECT 423.6000 144.2000 424.4000 155.8000 ;
	    RECT 431.7000 152.4000 432.3000 191.7000 ;
	    RECT 438.1000 190.4000 438.7000 195.6000 ;
	    RECT 439.7000 194.4000 440.3000 197.6000 ;
	    RECT 439.6000 193.6000 440.4000 194.4000 ;
	    RECT 438.0000 189.6000 438.8000 190.4000 ;
	    RECT 434.8000 183.6000 435.6000 184.4000 ;
	    RECT 436.4000 183.6000 437.2000 184.4000 ;
	    RECT 434.9000 176.4000 435.5000 183.6000 ;
	    RECT 436.5000 178.4000 437.1000 183.6000 ;
	    RECT 436.4000 177.6000 437.2000 178.4000 ;
	    RECT 439.7000 176.4000 440.3000 193.6000 ;
	    RECT 441.3000 192.4000 441.9000 215.6000 ;
	    RECT 442.9000 214.4000 443.5000 229.6000 ;
	    RECT 450.8000 225.6000 451.6000 226.4000 ;
	    RECT 446.0000 223.6000 446.8000 224.4000 ;
	    RECT 442.8000 213.6000 443.6000 214.4000 ;
	    RECT 446.1000 208.4000 446.7000 223.6000 ;
	    RECT 452.5000 218.4000 453.1000 231.6000 ;
	    RECT 454.1000 230.4000 454.7000 251.6000 ;
	    RECT 455.6000 246.2000 456.4000 257.8000 ;
	    RECT 463.6000 255.6000 464.4000 256.4000 ;
	    RECT 457.2000 251.6000 458.0000 252.4000 ;
	    RECT 463.6000 251.8000 464.4000 252.6000 ;
	    RECT 457.3000 250.4000 457.9000 251.6000 ;
	    RECT 463.7000 250.4000 464.3000 251.8000 ;
	    RECT 457.2000 249.6000 458.0000 250.4000 ;
	    RECT 463.6000 249.6000 464.4000 250.4000 ;
	    RECT 465.2000 246.2000 466.0000 257.8000 ;
	    RECT 466.9000 252.4000 467.5000 291.6000 ;
	    RECT 468.5000 286.3000 469.1000 327.6000 ;
	    RECT 470.0000 323.6000 470.8000 324.4000 ;
	    RECT 470.1000 312.4000 470.7000 323.6000 ;
	    RECT 474.9000 322.4000 475.5000 331.6000 ;
	    RECT 479.7000 328.4000 480.3000 335.6000 ;
	    RECT 479.6000 327.6000 480.4000 328.4000 ;
	    RECT 479.7000 324.4000 480.3000 327.6000 ;
	    RECT 486.0000 326.2000 486.8000 337.8000 ;
	    RECT 492.4000 333.6000 493.2000 334.4000 ;
	    RECT 490.8000 331.6000 491.6000 332.4000 ;
	    RECT 479.6000 323.6000 480.4000 324.4000 ;
	    RECT 474.8000 321.6000 475.6000 322.4000 ;
	    RECT 492.5000 318.4000 493.1000 333.6000 ;
	    RECT 495.6000 326.2000 496.4000 337.8000 ;
	    RECT 498.8000 330.2000 499.6000 335.8000 ;
	    RECT 500.4000 335.6000 501.2000 336.4000 ;
	    RECT 498.8000 325.6000 499.6000 326.4000 ;
	    RECT 492.4000 317.6000 493.2000 318.4000 ;
	    RECT 470.0000 311.6000 470.8000 312.4000 ;
	    RECT 471.6000 309.4000 472.4000 310.4000 ;
	    RECT 473.2000 304.2000 474.0000 315.8000 ;
	    RECT 474.8000 307.6000 475.6000 308.4000 ;
	    RECT 471.6000 297.6000 472.4000 298.4000 ;
	    RECT 470.0000 293.6000 470.8000 294.4000 ;
	    RECT 470.0000 289.6000 470.8000 290.4000 ;
	    RECT 470.1000 288.4000 470.7000 289.6000 ;
	    RECT 474.9000 288.4000 475.5000 307.6000 ;
	    RECT 476.4000 306.2000 477.2000 311.8000 ;
	    RECT 478.0000 311.6000 478.8000 312.4000 ;
	    RECT 478.0000 309.6000 478.8000 310.4000 ;
	    RECT 482.8000 309.6000 483.6000 310.4000 ;
	    RECT 495.6000 309.6000 496.4000 310.4000 ;
	    RECT 486.0000 305.6000 486.8000 306.4000 ;
	    RECT 487.6000 305.6000 488.4000 306.4000 ;
	    RECT 486.1000 304.4000 486.7000 305.6000 ;
	    RECT 486.0000 303.6000 486.8000 304.4000 ;
	    RECT 470.0000 287.6000 470.8000 288.4000 ;
	    RECT 474.8000 287.6000 475.6000 288.4000 ;
	    RECT 470.0000 286.3000 470.8000 286.4000 ;
	    RECT 468.5000 285.7000 470.8000 286.3000 ;
	    RECT 476.4000 286.2000 477.2000 297.8000 ;
	    RECT 484.4000 297.6000 485.2000 298.4000 ;
	    RECT 482.8000 293.6000 483.6000 294.4000 ;
	    RECT 482.9000 292.4000 483.5000 293.6000 ;
	    RECT 479.6000 291.6000 480.4000 292.4000 ;
	    RECT 482.8000 291.6000 483.6000 292.4000 ;
	    RECT 470.0000 285.6000 470.8000 285.7000 ;
	    RECT 470.1000 278.4000 470.7000 285.6000 ;
	    RECT 470.0000 277.6000 470.8000 278.4000 ;
	    RECT 471.6000 277.6000 472.4000 278.4000 ;
	    RECT 478.0000 277.6000 478.8000 278.4000 ;
	    RECT 471.7000 274.4000 472.3000 277.6000 ;
	    RECT 471.6000 273.6000 472.4000 274.4000 ;
	    RECT 476.4000 264.2000 477.2000 275.8000 ;
	    RECT 476.4000 259.6000 477.2000 260.4000 ;
	    RECT 470.0000 257.6000 470.8000 258.4000 ;
	    RECT 470.1000 256.4000 470.7000 257.6000 ;
	    RECT 476.5000 256.4000 477.1000 259.6000 ;
	    RECT 466.8000 251.6000 467.6000 252.4000 ;
	    RECT 468.4000 250.2000 469.2000 255.8000 ;
	    RECT 470.0000 255.6000 470.8000 256.4000 ;
	    RECT 476.4000 255.6000 477.2000 256.4000 ;
	    RECT 474.8000 251.6000 475.6000 252.4000 ;
	    RECT 474.8000 249.6000 475.6000 250.4000 ;
	    RECT 458.8000 235.6000 459.6000 236.4000 ;
	    RECT 458.9000 234.4000 459.5000 235.6000 ;
	    RECT 458.8000 233.6000 459.6000 234.4000 ;
	    RECT 454.0000 229.6000 454.8000 230.4000 ;
	    RECT 452.4000 217.6000 453.2000 218.4000 ;
	    RECT 447.6000 213.6000 448.4000 214.4000 ;
	    RECT 450.8000 213.6000 451.6000 214.4000 ;
	    RECT 447.7000 212.4000 448.3000 213.6000 ;
	    RECT 447.6000 211.6000 448.4000 212.4000 ;
	    RECT 446.0000 207.6000 446.8000 208.4000 ;
	    RECT 446.1000 206.4000 446.7000 207.6000 ;
	    RECT 446.0000 205.6000 446.8000 206.4000 ;
	    RECT 446.0000 203.6000 446.8000 204.4000 ;
	    RECT 446.1000 202.4000 446.7000 203.6000 ;
	    RECT 446.0000 201.6000 446.8000 202.4000 ;
	    RECT 450.8000 193.6000 451.6000 194.4000 ;
	    RECT 450.9000 192.4000 451.5000 193.6000 ;
	    RECT 441.2000 191.6000 442.0000 192.4000 ;
	    RECT 442.8000 191.6000 443.6000 192.4000 ;
	    RECT 450.8000 191.6000 451.6000 192.4000 ;
	    RECT 442.9000 188.4000 443.5000 191.6000 ;
	    RECT 454.1000 190.4000 454.7000 229.6000 ;
	    RECT 458.9000 226.4000 459.5000 233.6000 ;
	    RECT 458.8000 225.6000 459.6000 226.4000 ;
	    RECT 465.2000 224.2000 466.0000 235.8000 ;
	    RECT 471.6000 229.6000 472.4000 230.4000 ;
	    RECT 471.7000 226.4000 472.3000 229.6000 ;
	    RECT 471.6000 225.6000 472.4000 226.4000 ;
	    RECT 474.8000 224.2000 475.6000 235.8000 ;
	    RECT 476.5000 228.4000 477.1000 255.6000 ;
	    RECT 478.1000 250.4000 478.7000 277.6000 ;
	    RECT 479.7000 270.4000 480.3000 291.6000 ;
	    RECT 484.5000 276.4000 485.1000 297.6000 ;
	    RECT 486.0000 286.2000 486.8000 297.8000 ;
	    RECT 487.7000 296.4000 488.3000 305.6000 ;
	    RECT 489.2000 303.6000 490.0000 304.4000 ;
	    RECT 492.4000 303.6000 493.2000 304.4000 ;
	    RECT 489.3000 298.4000 489.9000 303.6000 ;
	    RECT 489.2000 297.6000 490.0000 298.4000 ;
	    RECT 487.6000 295.6000 488.4000 296.4000 ;
	    RECT 487.6000 293.6000 488.4000 294.4000 ;
	    RECT 489.2000 290.2000 490.0000 295.8000 ;
	    RECT 490.8000 295.6000 491.6000 296.4000 ;
	    RECT 484.4000 275.6000 485.2000 276.4000 ;
	    RECT 479.6000 269.6000 480.4000 270.4000 ;
	    RECT 479.7000 260.4000 480.3000 269.6000 ;
	    RECT 484.4000 269.4000 485.2000 270.2000 ;
	    RECT 484.5000 266.4000 485.1000 269.4000 ;
	    RECT 484.4000 265.6000 485.2000 266.4000 ;
	    RECT 486.0000 264.2000 486.8000 275.8000 ;
	    RECT 487.6000 275.6000 488.4000 276.4000 ;
	    RECT 490.9000 276.3000 491.5000 295.6000 ;
	    RECT 492.5000 294.4000 493.1000 303.6000 ;
	    RECT 492.4000 293.6000 493.2000 294.4000 ;
	    RECT 492.4000 291.6000 493.2000 292.4000 ;
	    RECT 494.0000 287.6000 494.8000 288.4000 ;
	    RECT 494.1000 286.4000 494.7000 287.6000 ;
	    RECT 494.0000 285.6000 494.8000 286.4000 ;
	    RECT 492.4000 283.6000 493.2000 284.4000 ;
	    RECT 492.5000 278.4000 493.1000 283.6000 ;
	    RECT 492.4000 277.6000 493.2000 278.4000 ;
	    RECT 490.9000 275.7000 493.1000 276.3000 ;
	    RECT 479.6000 259.6000 480.4000 260.4000 ;
	    RECT 486.0000 259.6000 486.8000 260.4000 ;
	    RECT 479.6000 257.6000 480.4000 258.4000 ;
	    RECT 479.7000 256.4000 480.3000 257.6000 ;
	    RECT 479.6000 255.6000 480.4000 256.4000 ;
	    RECT 478.0000 249.6000 478.8000 250.4000 ;
	    RECT 484.4000 246.2000 485.2000 257.8000 ;
	    RECT 486.1000 252.4000 486.7000 259.6000 ;
	    RECT 486.0000 251.6000 486.8000 252.4000 ;
	    RECT 482.8000 235.6000 483.6000 236.4000 ;
	    RECT 481.2000 233.6000 482.0000 234.4000 ;
	    RECT 482.9000 232.4000 483.5000 235.6000 ;
	    RECT 476.4000 227.6000 477.2000 228.4000 ;
	    RECT 478.0000 226.2000 478.8000 231.8000 ;
	    RECT 482.8000 231.6000 483.6000 232.4000 ;
	    RECT 486.0000 231.6000 486.8000 232.4000 ;
	    RECT 482.8000 229.6000 483.6000 230.4000 ;
	    RECT 486.0000 229.6000 486.8000 230.4000 ;
	    RECT 458.8000 217.6000 459.6000 218.4000 ;
	    RECT 458.9000 216.4000 459.5000 217.6000 ;
	    RECT 458.8000 215.6000 459.6000 216.4000 ;
	    RECT 457.2000 205.6000 458.0000 206.4000 ;
	    RECT 463.6000 206.2000 464.4000 217.8000 ;
	    RECT 471.6000 211.8000 472.4000 212.6000 ;
	    RECT 471.7000 210.4000 472.3000 211.8000 ;
	    RECT 471.6000 209.6000 472.4000 210.4000 ;
	    RECT 465.2000 207.6000 466.0000 208.4000 ;
	    RECT 455.6000 203.6000 456.4000 204.4000 ;
	    RECT 447.6000 189.6000 448.4000 190.4000 ;
	    RECT 454.0000 189.6000 454.8000 190.4000 ;
	    RECT 442.8000 187.6000 443.6000 188.4000 ;
	    RECT 444.4000 183.6000 445.2000 184.4000 ;
	    RECT 444.5000 180.4000 445.1000 183.6000 ;
	    RECT 444.4000 179.6000 445.2000 180.4000 ;
	    RECT 434.8000 175.6000 435.6000 176.4000 ;
	    RECT 436.4000 175.6000 437.2000 176.4000 ;
	    RECT 439.6000 175.6000 440.4000 176.4000 ;
	    RECT 436.5000 168.4000 437.1000 175.6000 ;
	    RECT 447.7000 174.4000 448.3000 189.6000 ;
	    RECT 452.4000 183.6000 453.2000 184.4000 ;
	    RECT 450.8000 175.6000 451.6000 176.4000 ;
	    RECT 439.6000 173.6000 440.4000 174.4000 ;
	    RECT 447.6000 173.6000 448.4000 174.4000 ;
	    RECT 455.7000 174.3000 456.3000 203.6000 ;
	    RECT 457.3000 194.4000 457.9000 205.6000 ;
	    RECT 465.3000 198.4000 465.9000 207.6000 ;
	    RECT 471.6000 205.6000 472.4000 206.4000 ;
	    RECT 473.2000 206.2000 474.0000 217.8000 ;
	    RECT 474.8000 213.6000 475.6000 214.4000 ;
	    RECT 476.4000 210.2000 477.2000 215.8000 ;
	    RECT 484.4000 215.6000 485.2000 216.4000 ;
	    RECT 487.7000 214.4000 488.3000 275.6000 ;
	    RECT 490.8000 273.6000 491.6000 274.4000 ;
	    RECT 489.2000 266.2000 490.0000 271.8000 ;
	    RECT 490.9000 266.4000 491.5000 273.6000 ;
	    RECT 490.8000 265.6000 491.6000 266.4000 ;
	    RECT 490.8000 257.6000 491.6000 258.4000 ;
	    RECT 490.9000 252.4000 491.5000 257.6000 ;
	    RECT 490.8000 251.6000 491.6000 252.4000 ;
	    RECT 490.8000 243.6000 491.6000 244.4000 ;
	    RECT 489.2000 235.6000 490.0000 236.4000 ;
	    RECT 489.3000 230.4000 489.9000 235.6000 ;
	    RECT 489.2000 229.6000 490.0000 230.4000 ;
	    RECT 487.6000 213.6000 488.4000 214.4000 ;
	    RECT 489.3000 212.4000 489.9000 229.6000 ;
	    RECT 490.9000 224.4000 491.5000 243.6000 ;
	    RECT 490.8000 223.6000 491.6000 224.4000 ;
	    RECT 492.5000 220.4000 493.1000 275.7000 ;
	    RECT 495.7000 270.4000 496.3000 309.6000 ;
	    RECT 498.9000 292.4000 499.5000 325.6000 ;
	    RECT 500.5000 296.4000 501.1000 335.6000 ;
	    RECT 503.6000 333.6000 504.4000 334.4000 ;
	    RECT 508.4000 333.6000 509.2000 334.4000 ;
	    RECT 506.8000 331.6000 507.6000 332.4000 ;
	    RECT 502.0000 323.6000 502.8000 324.4000 ;
	    RECT 500.4000 295.6000 501.2000 296.4000 ;
	    RECT 498.8000 291.6000 499.6000 292.4000 ;
	    RECT 497.2000 287.6000 498.0000 288.4000 ;
	    RECT 498.9000 288.3000 499.5000 291.6000 ;
	    RECT 498.9000 287.7000 501.1000 288.3000 ;
	    RECT 497.3000 286.4000 497.9000 287.6000 ;
	    RECT 497.2000 285.6000 498.0000 286.4000 ;
	    RECT 497.3000 270.4000 497.9000 285.6000 ;
	    RECT 498.8000 283.6000 499.6000 284.4000 ;
	    RECT 498.9000 272.4000 499.5000 283.6000 ;
	    RECT 500.5000 278.4000 501.1000 287.7000 ;
	    RECT 500.4000 277.6000 501.2000 278.4000 ;
	    RECT 498.8000 271.6000 499.6000 272.4000 ;
	    RECT 495.6000 269.6000 496.4000 270.4000 ;
	    RECT 497.2000 269.6000 498.0000 270.4000 ;
	    RECT 500.4000 269.6000 501.2000 270.4000 ;
	    RECT 494.0000 246.2000 494.8000 257.8000 ;
	    RECT 494.0000 237.6000 494.8000 238.4000 ;
	    RECT 494.1000 234.4000 494.7000 237.6000 ;
	    RECT 495.7000 236.4000 496.3000 269.6000 ;
	    RECT 497.2000 267.6000 498.0000 268.4000 ;
	    RECT 497.3000 266.4000 497.9000 267.6000 ;
	    RECT 497.2000 265.6000 498.0000 266.4000 ;
	    RECT 497.2000 250.2000 498.0000 255.8000 ;
	    RECT 500.5000 248.4000 501.1000 269.6000 ;
	    RECT 502.1000 260.4000 502.7000 323.6000 ;
	    RECT 505.2000 309.6000 506.0000 310.4000 ;
	    RECT 505.3000 308.4000 505.9000 309.6000 ;
	    RECT 506.9000 308.4000 507.5000 331.6000 ;
	    RECT 508.5000 328.4000 509.1000 333.6000 ;
	    RECT 510.0000 331.6000 510.8000 332.4000 ;
	    RECT 508.4000 327.6000 509.2000 328.4000 ;
	    RECT 505.2000 307.6000 506.0000 308.4000 ;
	    RECT 506.8000 307.6000 507.6000 308.4000 ;
	    RECT 508.4000 303.6000 509.2000 304.4000 ;
	    RECT 505.2000 291.6000 506.0000 292.4000 ;
	    RECT 505.3000 290.4000 505.9000 291.6000 ;
	    RECT 505.2000 289.6000 506.0000 290.4000 ;
	    RECT 506.8000 287.6000 507.6000 288.4000 ;
	    RECT 503.6000 269.6000 504.4000 270.4000 ;
	    RECT 503.7000 268.4000 504.3000 269.6000 ;
	    RECT 503.6000 267.6000 504.4000 268.4000 ;
	    RECT 502.0000 259.6000 502.8000 260.4000 ;
	    RECT 505.2000 257.6000 506.0000 258.4000 ;
	    RECT 502.0000 253.6000 502.8000 254.4000 ;
	    RECT 502.1000 252.4000 502.7000 253.6000 ;
	    RECT 502.0000 251.6000 502.8000 252.4000 ;
	    RECT 506.9000 250.4000 507.5000 287.6000 ;
	    RECT 508.5000 286.4000 509.1000 303.6000 ;
	    RECT 508.4000 285.6000 509.2000 286.4000 ;
	    RECT 508.4000 283.6000 509.2000 284.4000 ;
	    RECT 505.2000 249.6000 506.0000 250.4000 ;
	    RECT 506.8000 249.6000 507.6000 250.4000 ;
	    RECT 500.4000 247.6000 501.2000 248.4000 ;
	    RECT 505.3000 246.4000 505.9000 249.6000 ;
	    RECT 502.0000 245.6000 502.8000 246.4000 ;
	    RECT 505.2000 245.6000 506.0000 246.4000 ;
	    RECT 508.5000 238.4000 509.1000 283.6000 ;
	    RECT 510.1000 278.4000 510.7000 331.6000 ;
	    RECT 513.2000 323.6000 514.0000 324.4000 ;
	    RECT 513.3000 310.4000 513.9000 323.6000 ;
	    RECT 513.2000 309.6000 514.0000 310.4000 ;
	    RECT 511.6000 307.6000 512.4000 308.4000 ;
	    RECT 510.0000 277.6000 510.8000 278.4000 ;
	    RECT 510.1000 272.4000 510.7000 277.6000 ;
	    RECT 510.0000 271.6000 510.8000 272.4000 ;
	    RECT 510.0000 251.6000 510.8000 252.4000 ;
	    RECT 503.6000 237.6000 504.4000 238.4000 ;
	    RECT 508.4000 237.6000 509.2000 238.4000 ;
	    RECT 495.6000 235.6000 496.4000 236.4000 ;
	    RECT 494.0000 233.6000 494.8000 234.4000 ;
	    RECT 494.1000 226.4000 494.7000 233.6000 ;
	    RECT 494.0000 225.6000 494.8000 226.4000 ;
	    RECT 495.6000 226.2000 496.4000 231.8000 ;
	    RECT 497.2000 227.6000 498.0000 228.4000 ;
	    RECT 494.0000 223.6000 494.8000 224.4000 ;
	    RECT 498.8000 224.2000 499.6000 235.8000 ;
	    RECT 500.4000 229.4000 501.2000 230.4000 ;
	    RECT 492.4000 219.6000 493.2000 220.4000 ;
	    RECT 492.5000 214.3000 493.1000 219.6000 ;
	    RECT 494.1000 218.4000 494.7000 223.6000 ;
	    RECT 494.0000 217.6000 494.8000 218.4000 ;
	    RECT 492.5000 213.7000 494.7000 214.3000 ;
	    RECT 479.6000 211.6000 480.4000 212.4000 ;
	    RECT 481.2000 211.6000 482.0000 212.4000 ;
	    RECT 489.2000 211.6000 490.0000 212.4000 ;
	    RECT 492.4000 211.6000 493.2000 212.4000 ;
	    RECT 479.7000 210.4000 480.3000 211.6000 ;
	    RECT 478.0000 209.6000 478.8000 210.4000 ;
	    RECT 479.6000 209.6000 480.4000 210.4000 ;
	    RECT 478.1000 208.4000 478.7000 209.6000 ;
	    RECT 478.0000 207.6000 478.8000 208.4000 ;
	    RECT 471.7000 198.4000 472.3000 205.6000 ;
	    RECT 474.8000 199.6000 475.6000 200.4000 ;
	    RECT 465.2000 197.6000 466.0000 198.4000 ;
	    RECT 471.6000 197.6000 472.4000 198.4000 ;
	    RECT 458.8000 195.6000 459.6000 196.4000 ;
	    RECT 474.9000 194.4000 475.5000 199.6000 ;
	    RECT 457.2000 193.6000 458.0000 194.4000 ;
	    RECT 463.6000 193.6000 464.4000 194.4000 ;
	    RECT 470.0000 193.6000 470.8000 194.4000 ;
	    RECT 474.8000 193.6000 475.6000 194.4000 ;
	    RECT 458.8000 191.6000 459.6000 192.4000 ;
	    RECT 465.2000 191.6000 466.0000 192.4000 ;
	    RECT 471.6000 191.6000 472.4000 192.4000 ;
	    RECT 458.9000 190.4000 459.5000 191.6000 ;
	    RECT 465.3000 190.4000 465.9000 191.6000 ;
	    RECT 471.7000 190.4000 472.3000 191.6000 ;
	    RECT 458.8000 189.6000 459.6000 190.4000 ;
	    RECT 465.2000 189.6000 466.0000 190.4000 ;
	    RECT 471.6000 189.6000 472.4000 190.4000 ;
	    RECT 474.9000 186.4000 475.5000 193.6000 ;
	    RECT 479.6000 190.3000 480.4000 190.4000 ;
	    RECT 481.3000 190.3000 481.9000 211.6000 ;
	    RECT 492.4000 209.6000 493.2000 210.4000 ;
	    RECT 492.5000 206.4000 493.1000 209.6000 ;
	    RECT 492.4000 205.6000 493.2000 206.4000 ;
	    RECT 482.8000 195.6000 483.6000 196.4000 ;
	    RECT 482.9000 192.4000 483.5000 195.6000 ;
	    RECT 484.4000 193.6000 485.2000 194.4000 ;
	    RECT 487.6000 193.6000 488.4000 194.4000 ;
	    RECT 482.8000 191.6000 483.6000 192.4000 ;
	    RECT 479.6000 189.7000 481.9000 190.3000 ;
	    RECT 479.6000 189.6000 480.4000 189.7000 ;
	    RECT 474.8000 185.6000 475.6000 186.4000 ;
	    RECT 481.3000 184.4000 481.9000 189.7000 ;
	    RECT 482.8000 189.6000 483.6000 190.4000 ;
	    RECT 481.2000 183.6000 482.0000 184.4000 ;
	    RECT 465.2000 175.6000 466.0000 176.4000 ;
	    RECT 454.1000 173.7000 456.3000 174.3000 ;
	    RECT 439.7000 172.4000 440.3000 173.6000 ;
	    RECT 454.1000 172.4000 454.7000 173.7000 ;
	    RECT 455.7000 172.4000 456.3000 173.7000 ;
	    RECT 465.3000 172.4000 465.9000 175.6000 ;
	    RECT 481.2000 173.6000 482.0000 174.4000 ;
	    RECT 481.3000 172.4000 481.9000 173.6000 ;
	    RECT 438.0000 171.6000 438.8000 172.4000 ;
	    RECT 439.6000 171.6000 440.4000 172.4000 ;
	    RECT 447.6000 171.6000 448.4000 172.4000 ;
	    RECT 454.0000 171.6000 454.8000 172.4000 ;
	    RECT 455.6000 171.6000 456.4000 172.4000 ;
	    RECT 460.4000 171.6000 461.2000 172.4000 ;
	    RECT 465.2000 171.6000 466.0000 172.4000 ;
	    RECT 470.0000 171.6000 470.8000 172.4000 ;
	    RECT 478.0000 171.6000 478.8000 172.4000 ;
	    RECT 481.2000 171.6000 482.0000 172.4000 ;
	    RECT 486.0000 171.6000 486.8000 172.4000 ;
	    RECT 438.1000 170.4000 438.7000 171.6000 ;
	    RECT 447.7000 170.4000 448.3000 171.6000 ;
	    RECT 460.5000 170.4000 461.1000 171.6000 ;
	    RECT 478.1000 170.4000 478.7000 171.6000 ;
	    RECT 438.0000 169.6000 438.8000 170.4000 ;
	    RECT 447.6000 169.6000 448.4000 170.4000 ;
	    RECT 460.4000 169.6000 461.2000 170.4000 ;
	    RECT 468.4000 169.6000 469.2000 170.4000 ;
	    RECT 478.0000 169.6000 478.8000 170.4000 ;
	    RECT 468.5000 168.4000 469.1000 169.6000 ;
	    RECT 486.1000 168.4000 486.7000 171.6000 ;
	    RECT 487.7000 168.4000 488.3000 193.6000 ;
	    RECT 489.2000 184.2000 490.0000 195.8000 ;
	    RECT 492.4000 189.6000 493.2000 190.4000 ;
	    RECT 489.2000 169.6000 490.0000 170.4000 ;
	    RECT 436.4000 167.6000 437.2000 168.4000 ;
	    RECT 457.2000 167.6000 458.0000 168.4000 ;
	    RECT 462.0000 167.6000 462.8000 168.4000 ;
	    RECT 468.4000 167.6000 469.2000 168.4000 ;
	    RECT 473.2000 167.6000 474.0000 168.4000 ;
	    RECT 476.4000 167.6000 477.2000 168.4000 ;
	    RECT 486.0000 167.6000 486.8000 168.4000 ;
	    RECT 487.6000 167.6000 488.4000 168.4000 ;
	    RECT 425.2000 147.6000 426.0000 148.4000 ;
	    RECT 422.0000 139.6000 422.8000 140.4000 ;
	    RECT 412.4000 137.6000 413.2000 138.4000 ;
	    RECT 412.5000 136.4000 413.1000 137.6000 ;
	    RECT 412.4000 135.6000 413.2000 136.4000 ;
	    RECT 404.4000 133.6000 405.2000 134.4000 ;
	    RECT 391.6000 131.6000 392.4000 132.4000 ;
	    RECT 401.2000 131.6000 402.0000 132.4000 ;
	    RECT 402.8000 131.6000 403.6000 132.4000 ;
	    RECT 391.7000 130.4000 392.3000 131.6000 ;
	    RECT 391.6000 129.6000 392.4000 130.4000 ;
	    RECT 398.0000 127.6000 398.8000 128.4000 ;
	    RECT 390.1000 125.7000 392.3000 126.3000 ;
	    RECT 390.0000 123.6000 390.8000 124.4000 ;
	    RECT 383.7000 117.7000 385.9000 118.3000 ;
	    RECT 382.0000 107.6000 382.8000 108.4000 ;
	    RECT 380.4000 105.6000 381.2000 106.4000 ;
	    RECT 383.6000 104.2000 384.4000 115.8000 ;
	    RECT 385.3000 92.4000 385.9000 117.7000 ;
	    RECT 386.8000 117.6000 387.6000 118.4000 ;
	    RECT 390.1000 112.4000 390.7000 123.6000 ;
	    RECT 390.0000 111.6000 390.8000 112.4000 ;
	    RECT 390.0000 109.6000 390.8000 110.4000 ;
	    RECT 390.1000 108.4000 390.7000 109.6000 ;
	    RECT 391.7000 108.4000 392.3000 125.7000 ;
	    RECT 398.1000 124.4000 398.7000 127.6000 ;
	    RECT 398.0000 123.6000 398.8000 124.4000 ;
	    RECT 398.1000 118.4000 398.7000 123.6000 ;
	    RECT 398.0000 117.6000 398.8000 118.4000 ;
	    RECT 390.0000 107.6000 390.8000 108.4000 ;
	    RECT 391.6000 107.6000 392.4000 108.4000 ;
	    RECT 386.8000 105.6000 387.6000 106.4000 ;
	    RECT 386.9000 94.4000 387.5000 105.6000 ;
	    RECT 393.2000 104.2000 394.0000 115.8000 ;
	    RECT 401.3000 112.4000 401.9000 131.6000 ;
	    RECT 396.4000 106.2000 397.2000 111.8000 ;
	    RECT 398.0000 111.6000 398.8000 112.4000 ;
	    RECT 401.2000 111.6000 402.0000 112.4000 ;
	    RECT 401.2000 110.3000 402.0000 110.4000 ;
	    RECT 402.9000 110.3000 403.5000 131.6000 ;
	    RECT 417.2000 126.2000 418.0000 137.8000 ;
	    RECT 425.3000 136.4000 425.9000 147.6000 ;
	    RECT 426.8000 146.2000 427.6000 151.8000 ;
	    RECT 431.6000 151.6000 432.4000 152.4000 ;
	    RECT 428.4000 143.6000 429.2000 144.4000 ;
	    RECT 425.2000 135.6000 426.0000 136.4000 ;
	    RECT 425.2000 131.6000 426.0000 132.6000 ;
	    RECT 426.8000 126.2000 427.6000 137.8000 ;
	    RECT 430.0000 130.2000 430.8000 135.8000 ;
	    RECT 431.7000 130.4000 432.3000 151.6000 ;
	    RECT 433.2000 144.2000 434.0000 155.8000 ;
	    RECT 441.2000 149.4000 442.0000 150.4000 ;
	    RECT 442.8000 144.2000 443.6000 155.8000 ;
	    RECT 444.4000 147.6000 445.2000 148.4000 ;
	    RECT 446.0000 146.2000 446.8000 151.8000 ;
	    RECT 450.8000 151.6000 451.6000 152.4000 ;
	    RECT 455.6000 151.6000 456.4000 152.4000 ;
	    RECT 455.7000 150.4000 456.3000 151.6000 ;
	    RECT 450.8000 149.6000 451.6000 150.4000 ;
	    RECT 455.6000 149.6000 456.4000 150.4000 ;
	    RECT 450.9000 148.4000 451.5000 149.6000 ;
	    RECT 457.3000 148.4000 457.9000 167.6000 ;
	    RECT 460.4000 163.6000 461.2000 164.4000 ;
	    RECT 447.6000 147.6000 448.4000 148.4000 ;
	    RECT 450.8000 147.6000 451.6000 148.4000 ;
	    RECT 457.2000 147.6000 458.0000 148.4000 ;
	    RECT 447.7000 144.4000 448.3000 147.6000 ;
	    RECT 447.6000 143.6000 448.4000 144.4000 ;
	    RECT 450.8000 143.6000 451.6000 144.4000 ;
	    RECT 458.8000 143.6000 459.6000 144.4000 ;
	    RECT 433.2000 139.6000 434.0000 140.4000 ;
	    RECT 444.4000 139.6000 445.2000 140.4000 ;
	    RECT 431.6000 129.6000 432.4000 130.4000 ;
	    RECT 412.4000 123.6000 413.2000 124.4000 ;
	    RECT 404.4000 117.6000 405.2000 118.4000 ;
	    RECT 412.5000 116.4000 413.1000 123.6000 ;
	    RECT 412.4000 115.6000 413.2000 116.4000 ;
	    RECT 401.2000 109.7000 403.5000 110.3000 ;
	    RECT 401.2000 109.6000 402.0000 109.7000 ;
	    RECT 398.0000 107.6000 398.8000 108.4000 ;
	    RECT 407.6000 107.6000 408.4000 108.4000 ;
	    RECT 394.8000 99.6000 395.6000 100.4000 ;
	    RECT 386.8000 93.6000 387.6000 94.4000 ;
	    RECT 377.2000 91.6000 378.0000 92.4000 ;
	    RECT 383.6000 91.6000 384.4000 92.4000 ;
	    RECT 385.2000 91.6000 386.0000 92.4000 ;
	    RECT 377.3000 82.4000 377.9000 91.6000 ;
	    RECT 380.4000 89.6000 381.2000 90.4000 ;
	    RECT 377.2000 81.6000 378.0000 82.4000 ;
	    RECT 380.5000 80.4000 381.1000 89.6000 ;
	    RECT 385.3000 86.4000 385.9000 91.6000 ;
	    RECT 385.2000 85.6000 386.0000 86.4000 ;
	    RECT 393.2000 86.2000 394.0000 97.8000 ;
	    RECT 394.9000 90.3000 395.5000 99.6000 ;
	    RECT 396.4000 91.6000 397.2000 92.4000 ;
	    RECT 394.9000 89.7000 397.1000 90.3000 ;
	    RECT 388.4000 83.6000 389.2000 84.4000 ;
	    RECT 388.5000 80.4000 389.1000 83.6000 ;
	    RECT 380.4000 79.6000 381.2000 80.4000 ;
	    RECT 388.4000 79.6000 389.2000 80.4000 ;
	    RECT 377.2000 71.6000 378.0000 72.4000 ;
	    RECT 377.3000 70.2000 377.9000 71.6000 ;
	    RECT 377.2000 69.4000 378.0000 70.2000 ;
	    RECT 377.2000 65.6000 378.0000 66.4000 ;
	    RECT 377.3000 54.4000 377.9000 65.6000 ;
	    RECT 378.8000 64.2000 379.6000 75.8000 ;
	    RECT 394.8000 73.6000 395.6000 74.4000 ;
	    RECT 382.0000 66.2000 382.8000 71.8000 ;
	    RECT 383.6000 71.6000 384.4000 72.4000 ;
	    RECT 385.2000 71.6000 386.0000 72.4000 ;
	    RECT 383.7000 68.4000 384.3000 71.6000 ;
	    RECT 385.3000 70.4000 385.9000 71.6000 ;
	    RECT 385.2000 69.6000 386.0000 70.4000 ;
	    RECT 388.4000 70.3000 389.2000 70.4000 ;
	    RECT 388.4000 69.7000 390.7000 70.3000 ;
	    RECT 388.4000 69.6000 389.2000 69.7000 ;
	    RECT 390.1000 68.4000 390.7000 69.7000 ;
	    RECT 393.2000 69.6000 394.0000 70.4000 ;
	    RECT 383.6000 67.6000 384.4000 68.4000 ;
	    RECT 388.4000 67.6000 389.2000 68.4000 ;
	    RECT 390.0000 67.6000 390.8000 68.4000 ;
	    RECT 375.6000 53.6000 376.4000 54.4000 ;
	    RECT 377.2000 53.6000 378.0000 54.4000 ;
	    RECT 374.0000 31.6000 374.8000 32.4000 ;
	    RECT 364.4000 29.6000 365.2000 30.4000 ;
	    RECT 366.0000 29.6000 366.8000 30.4000 ;
	    RECT 369.2000 29.6000 370.0000 30.4000 ;
	    RECT 367.6000 27.6000 368.4000 28.4000 ;
	    RECT 369.2000 27.6000 370.0000 28.4000 ;
	    RECT 367.7000 24.4000 368.3000 27.6000 ;
	    RECT 374.1000 26.4000 374.7000 31.6000 ;
	    RECT 375.7000 28.4000 376.3000 53.6000 ;
	    RECT 378.8000 51.6000 379.6000 52.6000 ;
	    RECT 380.4000 46.2000 381.2000 57.8000 ;
	    RECT 382.0000 53.6000 382.8000 54.4000 ;
	    RECT 382.1000 46.4000 382.7000 53.6000 ;
	    RECT 383.6000 50.2000 384.4000 55.8000 ;
	    RECT 385.2000 53.6000 386.0000 54.4000 ;
	    RECT 388.5000 54.3000 389.1000 67.6000 ;
	    RECT 390.1000 60.4000 390.7000 67.6000 ;
	    RECT 390.0000 59.6000 390.8000 60.4000 ;
	    RECT 394.8000 59.6000 395.6000 60.4000 ;
	    RECT 390.0000 54.3000 390.8000 54.4000 ;
	    RECT 388.5000 53.7000 390.8000 54.3000 ;
	    RECT 390.0000 53.6000 390.8000 53.7000 ;
	    RECT 391.6000 53.6000 392.4000 54.4000 ;
	    RECT 385.3000 52.4000 385.9000 53.6000 ;
	    RECT 385.2000 51.6000 386.0000 52.4000 ;
	    RECT 388.4000 51.6000 389.2000 52.4000 ;
	    RECT 385.2000 49.6000 386.0000 50.4000 ;
	    RECT 385.3000 48.4000 385.9000 49.6000 ;
	    RECT 385.2000 47.6000 386.0000 48.4000 ;
	    RECT 382.0000 45.6000 382.8000 46.4000 ;
	    RECT 385.2000 45.6000 386.0000 46.4000 ;
	    RECT 382.0000 37.6000 382.8000 38.4000 ;
	    RECT 385.3000 34.4000 385.9000 45.6000 ;
	    RECT 385.2000 33.6000 386.0000 34.4000 ;
	    RECT 378.8000 29.6000 379.6000 30.4000 ;
	    RECT 375.6000 27.6000 376.4000 28.4000 ;
	    RECT 377.2000 27.6000 378.0000 28.4000 ;
	    RECT 380.4000 27.6000 381.2000 28.4000 ;
	    RECT 374.0000 25.6000 374.8000 26.4000 ;
	    RECT 366.0000 23.6000 366.8000 24.4000 ;
	    RECT 367.6000 23.6000 368.4000 24.4000 ;
	    RECT 359.6000 19.6000 360.4000 20.4000 ;
	    RECT 353.2000 17.6000 354.0000 18.4000 ;
	    RECT 366.1000 16.4000 366.7000 23.6000 ;
	    RECT 369.2000 17.6000 370.0000 18.4000 ;
	    RECT 369.3000 16.4000 369.9000 17.6000 ;
	    RECT 366.0000 15.6000 366.8000 16.4000 ;
	    RECT 369.2000 15.6000 370.0000 16.4000 ;
	    RECT 366.1000 12.4000 366.7000 15.6000 ;
	    RECT 319.6000 11.6000 320.4000 12.4000 ;
	    RECT 322.8000 11.6000 323.6000 12.4000 ;
	    RECT 327.6000 11.6000 328.4000 12.4000 ;
	    RECT 330.8000 11.6000 331.6000 12.4000 ;
	    RECT 332.4000 11.6000 333.2000 12.4000 ;
	    RECT 338.8000 11.6000 339.6000 12.4000 ;
	    RECT 342.0000 11.6000 342.8000 12.4000 ;
	    RECT 343.6000 11.6000 344.4000 12.4000 ;
	    RECT 350.0000 11.6000 350.8000 12.4000 ;
	    RECT 356.4000 11.6000 357.2000 12.4000 ;
	    RECT 358.0000 11.6000 358.8000 12.4000 ;
	    RECT 361.2000 11.6000 362.0000 12.4000 ;
	    RECT 366.0000 11.6000 366.8000 12.4000 ;
	    RECT 322.9000 10.4000 323.5000 11.6000 ;
	    RECT 322.8000 9.6000 323.6000 10.4000 ;
	    RECT 316.4000 7.6000 317.2000 8.4000 ;
	    RECT 332.5000 2.4000 333.1000 11.6000 ;
	    RECT 338.9000 6.4000 339.5000 11.6000 ;
	    RECT 356.5000 8.4000 357.1000 11.6000 ;
	    RECT 361.3000 10.4000 361.9000 11.6000 ;
	    RECT 361.2000 9.6000 362.0000 10.4000 ;
	    RECT 356.4000 7.6000 357.2000 8.4000 ;
	    RECT 338.8000 5.6000 339.6000 6.4000 ;
	    RECT 362.8000 5.6000 363.6000 6.4000 ;
	    RECT 374.0000 6.2000 374.8000 17.8000 ;
	    RECT 377.3000 12.4000 377.9000 27.6000 ;
	    RECT 380.5000 14.4000 381.1000 27.6000 ;
	    RECT 385.3000 20.4000 385.9000 33.6000 ;
	    RECT 386.8000 24.2000 387.6000 35.8000 ;
	    RECT 388.5000 30.4000 389.1000 51.6000 ;
	    RECT 391.7000 38.4000 392.3000 53.6000 ;
	    RECT 394.9000 52.4000 395.5000 59.6000 ;
	    RECT 396.5000 54.4000 397.1000 89.7000 ;
	    RECT 402.8000 86.2000 403.6000 97.8000 ;
	    RECT 404.4000 93.6000 405.2000 94.4000 ;
	    RECT 406.0000 90.2000 406.8000 95.8000 ;
	    RECT 407.7000 86.4000 408.3000 107.6000 ;
	    RECT 415.6000 104.2000 416.4000 115.8000 ;
	    RECT 422.0000 111.6000 422.8000 112.4000 ;
	    RECT 422.1000 110.4000 422.7000 111.6000 ;
	    RECT 422.0000 109.6000 422.8000 110.4000 ;
	    RECT 423.6000 105.6000 424.4000 106.4000 ;
	    RECT 414.0000 99.6000 414.8000 100.4000 ;
	    RECT 414.1000 98.4000 414.7000 99.6000 ;
	    RECT 414.0000 97.6000 414.8000 98.4000 ;
	    RECT 407.6000 85.6000 408.4000 86.4000 ;
	    RECT 418.8000 86.2000 419.6000 97.8000 ;
	    RECT 423.7000 94.4000 424.3000 105.6000 ;
	    RECT 425.2000 104.2000 426.0000 115.8000 ;
	    RECT 433.3000 112.4000 433.9000 139.6000 ;
	    RECT 434.8000 135.6000 435.6000 136.4000 ;
	    RECT 434.9000 134.4000 435.5000 135.6000 ;
	    RECT 434.8000 133.6000 435.6000 134.4000 ;
	    RECT 442.8000 133.6000 443.6000 134.4000 ;
	    RECT 434.8000 131.6000 435.6000 132.4000 ;
	    RECT 439.6000 131.6000 440.4000 132.4000 ;
	    RECT 439.7000 130.4000 440.3000 131.6000 ;
	    RECT 439.6000 129.6000 440.4000 130.4000 ;
	    RECT 442.9000 118.4000 443.5000 133.6000 ;
	    RECT 444.5000 132.4000 445.1000 139.6000 ;
	    RECT 449.2000 133.6000 450.0000 134.4000 ;
	    RECT 449.3000 132.4000 449.9000 133.6000 ;
	    RECT 444.4000 131.6000 445.2000 132.4000 ;
	    RECT 449.2000 131.6000 450.0000 132.4000 ;
	    RECT 444.5000 130.4000 445.1000 131.6000 ;
	    RECT 444.4000 129.6000 445.2000 130.4000 ;
	    RECT 449.2000 129.6000 450.0000 130.4000 ;
	    RECT 442.8000 117.6000 443.6000 118.4000 ;
	    RECT 428.4000 106.2000 429.2000 111.8000 ;
	    RECT 433.2000 111.6000 434.0000 112.4000 ;
	    RECT 430.0000 107.6000 430.8000 108.4000 ;
	    RECT 430.1000 100.4000 430.7000 107.6000 ;
	    RECT 433.2000 103.6000 434.0000 104.4000 ;
	    RECT 434.8000 103.6000 435.6000 104.4000 ;
	    RECT 439.6000 104.2000 440.4000 115.8000 ;
	    RECT 430.0000 99.6000 430.8000 100.4000 ;
	    RECT 423.6000 93.6000 424.4000 94.4000 ;
	    RECT 426.8000 91.6000 427.6000 92.6000 ;
	    RECT 428.4000 86.2000 429.2000 97.8000 ;
	    RECT 430.0000 93.6000 430.8000 94.4000 ;
	    RECT 431.6000 90.2000 432.4000 95.8000 ;
	    RECT 433.3000 90.4000 433.9000 103.6000 ;
	    RECT 439.6000 97.6000 440.4000 98.4000 ;
	    RECT 439.7000 96.4000 440.3000 97.6000 ;
	    RECT 439.6000 95.6000 440.4000 96.4000 ;
	    RECT 438.0000 94.3000 438.8000 94.4000 ;
	    RECT 436.5000 93.7000 438.8000 94.3000 ;
	    RECT 434.8000 91.6000 435.6000 92.4000 ;
	    RECT 433.2000 89.6000 434.0000 90.4000 ;
	    RECT 430.0000 85.6000 430.8000 86.4000 ;
	    RECT 399.6000 64.2000 400.4000 75.8000 ;
	    RECT 407.6000 71.6000 408.4000 72.4000 ;
	    RECT 407.7000 70.2000 408.3000 71.6000 ;
	    RECT 407.6000 69.4000 408.4000 70.2000 ;
	    RECT 409.2000 64.2000 410.0000 75.8000 ;
	    RECT 414.0000 73.6000 414.8000 74.4000 ;
	    RECT 410.8000 67.6000 411.6000 68.4000 ;
	    RECT 410.9000 60.4000 411.5000 67.6000 ;
	    RECT 412.4000 66.2000 413.2000 71.8000 ;
	    RECT 414.1000 68.4000 414.7000 73.6000 ;
	    RECT 423.6000 71.6000 424.4000 72.4000 ;
	    RECT 425.2000 71.6000 426.0000 72.4000 ;
	    RECT 423.7000 70.4000 424.3000 71.6000 ;
	    RECT 423.6000 69.6000 424.4000 70.4000 ;
	    RECT 425.3000 68.4000 425.9000 71.6000 ;
	    RECT 428.4000 69.6000 429.2000 70.4000 ;
	    RECT 430.1000 68.4000 430.7000 85.6000 ;
	    RECT 436.5000 78.4000 437.1000 93.7000 ;
	    RECT 438.0000 93.6000 438.8000 93.7000 ;
	    RECT 438.0000 91.6000 438.8000 92.4000 ;
	    RECT 439.6000 83.6000 440.4000 84.4000 ;
	    RECT 436.4000 77.6000 437.2000 78.4000 ;
	    RECT 414.0000 67.6000 414.8000 68.4000 ;
	    RECT 425.2000 67.6000 426.0000 68.4000 ;
	    RECT 430.0000 67.6000 430.8000 68.4000 ;
	    RECT 430.1000 62.4000 430.7000 67.6000 ;
	    RECT 433.2000 63.6000 434.0000 64.4000 ;
	    RECT 430.0000 61.6000 430.8000 62.4000 ;
	    RECT 433.3000 60.4000 433.9000 63.6000 ;
	    RECT 410.8000 59.6000 411.6000 60.4000 ;
	    RECT 425.2000 59.6000 426.0000 60.4000 ;
	    RECT 433.2000 59.6000 434.0000 60.4000 ;
	    RECT 409.2000 57.6000 410.0000 58.4000 ;
	    RECT 409.3000 56.4000 409.9000 57.6000 ;
	    RECT 409.2000 55.6000 410.0000 56.4000 ;
	    RECT 396.4000 53.6000 397.2000 54.4000 ;
	    RECT 409.3000 52.4000 409.9000 55.6000 ;
	    RECT 394.8000 51.6000 395.6000 52.4000 ;
	    RECT 409.2000 51.6000 410.0000 52.4000 ;
	    RECT 394.9000 50.4000 395.5000 51.6000 ;
	    RECT 393.2000 49.6000 394.0000 50.4000 ;
	    RECT 394.8000 49.6000 395.6000 50.4000 ;
	    RECT 401.2000 49.6000 402.0000 50.4000 ;
	    RECT 391.6000 37.6000 392.4000 38.4000 ;
	    RECT 394.9000 32.4000 395.5000 49.6000 ;
	    RECT 414.0000 46.2000 414.8000 57.8000 ;
	    RECT 422.0000 55.6000 422.8000 56.4000 ;
	    RECT 422.1000 52.6000 422.7000 55.6000 ;
	    RECT 422.0000 51.8000 422.8000 52.6000 ;
	    RECT 422.1000 51.7000 422.7000 51.8000 ;
	    RECT 423.6000 46.2000 424.4000 57.8000 ;
	    RECT 425.3000 54.4000 425.9000 59.6000 ;
	    RECT 436.5000 56.4000 437.1000 77.6000 ;
	    RECT 438.0000 57.6000 438.8000 58.4000 ;
	    RECT 425.2000 53.6000 426.0000 54.4000 ;
	    RECT 398.0000 43.6000 398.8000 44.4000 ;
	    RECT 394.8000 31.6000 395.6000 32.4000 ;
	    RECT 388.4000 29.6000 389.2000 30.4000 ;
	    RECT 394.8000 29.4000 395.6000 30.4000 ;
	    RECT 396.4000 24.2000 397.2000 35.8000 ;
	    RECT 398.1000 30.4000 398.7000 43.6000 ;
	    RECT 401.2000 39.6000 402.0000 40.4000 ;
	    RECT 401.3000 38.4000 401.9000 39.6000 ;
	    RECT 401.2000 37.6000 402.0000 38.4000 ;
	    RECT 418.8000 37.6000 419.6000 38.4000 ;
	    RECT 398.0000 29.6000 398.8000 30.4000 ;
	    RECT 398.0000 27.6000 398.8000 28.4000 ;
	    RECT 385.2000 19.6000 386.0000 20.4000 ;
	    RECT 380.4000 13.6000 381.2000 14.4000 ;
	    RECT 377.2000 11.6000 378.0000 12.4000 ;
	    RECT 383.6000 6.2000 384.4000 17.8000 ;
	    RECT 385.3000 14.4000 385.9000 19.6000 ;
	    RECT 385.2000 13.6000 386.0000 14.4000 ;
	    RECT 386.8000 10.2000 387.6000 15.8000 ;
	    RECT 388.4000 9.6000 389.2000 10.4000 ;
	    RECT 388.5000 8.4000 389.1000 9.6000 ;
	    RECT 388.4000 7.6000 389.2000 8.4000 ;
	    RECT 393.2000 6.2000 394.0000 17.8000 ;
	    RECT 398.1000 14.4000 398.7000 27.6000 ;
	    RECT 399.6000 26.2000 400.4000 31.8000 ;
	    RECT 401.3000 28.4000 401.9000 37.6000 ;
	    RECT 415.6000 35.6000 416.4000 36.4000 ;
	    RECT 415.7000 32.4000 416.3000 35.6000 ;
	    RECT 404.4000 31.6000 405.2000 32.4000 ;
	    RECT 415.6000 31.6000 416.4000 32.4000 ;
	    RECT 415.7000 30.4000 416.3000 31.6000 ;
	    RECT 414.0000 29.6000 414.8000 30.4000 ;
	    RECT 415.6000 29.6000 416.4000 30.4000 ;
	    RECT 401.2000 27.6000 402.0000 28.4000 ;
	    RECT 417.2000 27.6000 418.0000 28.4000 ;
	    RECT 417.3000 24.4000 417.9000 27.6000 ;
	    RECT 417.2000 23.6000 418.0000 24.4000 ;
	    RECT 423.6000 24.2000 424.4000 35.8000 ;
	    RECT 425.3000 30.4000 425.9000 53.6000 ;
	    RECT 426.8000 50.2000 427.6000 55.8000 ;
	    RECT 433.2000 55.6000 434.0000 56.4000 ;
	    RECT 436.4000 55.6000 437.2000 56.4000 ;
	    RECT 438.1000 54.4000 438.7000 57.6000 ;
	    RECT 428.4000 53.6000 429.2000 54.4000 ;
	    RECT 438.0000 53.6000 438.8000 54.4000 ;
	    RECT 428.5000 52.4000 429.1000 53.6000 ;
	    RECT 439.7000 52.4000 440.3000 83.6000 ;
	    RECT 442.9000 56.3000 443.5000 117.6000 ;
	    RECT 447.6000 109.4000 448.4000 110.4000 ;
	    RECT 447.6000 105.6000 448.4000 106.4000 ;
	    RECT 444.4000 86.2000 445.2000 97.8000 ;
	    RECT 447.7000 94.4000 448.3000 105.6000 ;
	    RECT 449.2000 104.2000 450.0000 115.8000 ;
	    RECT 450.9000 98.4000 451.5000 143.6000 ;
	    RECT 452.4000 133.6000 453.2000 134.4000 ;
	    RECT 452.5000 128.4000 453.1000 133.6000 ;
	    RECT 457.2000 129.6000 458.0000 130.4000 ;
	    RECT 452.4000 127.6000 453.2000 128.4000 ;
	    RECT 452.5000 126.4000 453.1000 127.6000 ;
	    RECT 452.4000 125.6000 453.2000 126.4000 ;
	    RECT 457.3000 112.4000 457.9000 129.6000 ;
	    RECT 458.8000 126.2000 459.6000 137.8000 ;
	    RECT 452.4000 106.2000 453.2000 111.8000 ;
	    RECT 457.2000 111.6000 458.0000 112.4000 ;
	    RECT 457.2000 109.6000 458.0000 110.4000 ;
	    RECT 457.3000 108.4000 457.9000 109.6000 ;
	    RECT 454.0000 107.6000 454.8000 108.4000 ;
	    RECT 457.2000 107.6000 458.0000 108.4000 ;
	    RECT 454.1000 104.4000 454.7000 107.6000 ;
	    RECT 460.5000 106.4000 461.1000 163.6000 ;
	    RECT 462.1000 114.4000 462.7000 167.6000 ;
	    RECT 478.0000 163.6000 478.8000 164.4000 ;
	    RECT 484.4000 163.6000 485.2000 164.4000 ;
	    RECT 463.6000 144.2000 464.4000 155.8000 ;
	    RECT 471.6000 149.4000 472.4000 150.4000 ;
	    RECT 470.0000 147.6000 470.8000 148.4000 ;
	    RECT 463.6000 131.6000 464.4000 132.4000 ;
	    RECT 468.4000 126.2000 469.2000 137.8000 ;
	    RECT 470.1000 134.4000 470.7000 147.6000 ;
	    RECT 473.2000 144.2000 474.0000 155.8000 ;
	    RECT 478.1000 152.4000 478.7000 163.6000 ;
	    RECT 476.4000 146.2000 477.2000 151.8000 ;
	    RECT 478.0000 151.6000 478.8000 152.4000 ;
	    RECT 478.0000 149.6000 478.8000 150.4000 ;
	    RECT 481.2000 149.6000 482.0000 150.4000 ;
	    RECT 473.2000 137.6000 474.0000 138.4000 ;
	    RECT 470.0000 133.6000 470.8000 134.4000 ;
	    RECT 470.1000 132.4000 470.7000 133.6000 ;
	    RECT 470.0000 131.6000 470.8000 132.4000 ;
	    RECT 471.6000 130.2000 472.4000 135.8000 ;
	    RECT 478.0000 126.2000 478.8000 137.8000 ;
	    RECT 465.2000 117.6000 466.0000 118.4000 ;
	    RECT 471.6000 115.6000 472.4000 116.4000 ;
	    RECT 471.7000 114.4000 472.3000 115.6000 ;
	    RECT 462.0000 113.6000 462.8000 114.4000 ;
	    RECT 471.6000 113.6000 472.4000 114.4000 ;
	    RECT 471.7000 112.4000 472.3000 113.6000 ;
	    RECT 462.0000 111.6000 462.8000 112.4000 ;
	    RECT 471.6000 111.6000 472.4000 112.4000 ;
	    RECT 462.1000 110.4000 462.7000 111.6000 ;
	    RECT 462.0000 109.6000 462.8000 110.4000 ;
	    RECT 460.4000 105.6000 461.2000 106.4000 ;
	    RECT 454.0000 103.6000 454.8000 104.4000 ;
	    RECT 460.4000 103.6000 461.2000 104.4000 ;
	    RECT 450.8000 97.6000 451.6000 98.4000 ;
	    RECT 447.6000 93.6000 448.4000 94.4000 ;
	    RECT 452.4000 93.6000 453.2000 94.4000 ;
	    RECT 452.5000 92.6000 453.1000 93.6000 ;
	    RECT 452.4000 91.8000 453.2000 92.6000 ;
	    RECT 454.0000 86.2000 454.8000 97.8000 ;
	    RECT 455.6000 93.6000 456.4000 94.4000 ;
	    RECT 455.7000 80.4000 456.3000 93.6000 ;
	    RECT 457.2000 90.2000 458.0000 95.8000 ;
	    RECT 458.8000 95.6000 459.6000 96.4000 ;
	    RECT 460.5000 88.4000 461.1000 103.6000 ;
	    RECT 462.1000 92.4000 462.7000 109.6000 ;
	    RECT 463.6000 107.6000 464.4000 108.4000 ;
	    RECT 463.7000 100.4000 464.3000 107.6000 ;
	    RECT 468.4000 103.6000 469.2000 104.4000 ;
	    RECT 476.4000 104.2000 477.2000 115.8000 ;
	    RECT 484.5000 114.4000 485.1000 163.6000 ;
	    RECT 486.1000 158.4000 486.7000 167.6000 ;
	    RECT 486.0000 157.6000 486.8000 158.4000 ;
	    RECT 487.7000 148.4000 488.3000 167.6000 ;
	    RECT 489.3000 150.4000 489.9000 169.6000 ;
	    RECT 490.8000 166.2000 491.6000 177.8000 ;
	    RECT 494.1000 158.4000 494.7000 213.7000 ;
	    RECT 498.8000 206.2000 499.6000 217.8000 ;
	    RECT 500.4000 213.6000 501.2000 214.4000 ;
	    RECT 500.5000 212.4000 501.1000 213.6000 ;
	    RECT 500.4000 211.6000 501.2000 212.4000 ;
	    RECT 497.2000 185.6000 498.0000 186.4000 ;
	    RECT 495.6000 183.6000 496.4000 184.4000 ;
	    RECT 494.0000 157.6000 494.8000 158.4000 ;
	    RECT 489.2000 149.6000 490.0000 150.4000 ;
	    RECT 492.4000 149.6000 493.2000 150.4000 ;
	    RECT 487.6000 147.6000 488.4000 148.4000 ;
	    RECT 486.0000 145.6000 486.8000 146.4000 ;
	    RECT 486.1000 144.4000 486.7000 145.6000 ;
	    RECT 486.0000 143.6000 486.8000 144.4000 ;
	    RECT 487.7000 140.4000 488.3000 147.6000 ;
	    RECT 487.6000 139.6000 488.4000 140.4000 ;
	    RECT 486.0000 133.6000 486.8000 134.4000 ;
	    RECT 486.1000 132.6000 486.7000 133.6000 ;
	    RECT 486.0000 131.8000 486.8000 132.6000 ;
	    RECT 487.6000 126.2000 488.4000 137.8000 ;
	    RECT 492.4000 137.6000 493.2000 138.4000 ;
	    RECT 492.5000 136.4000 493.1000 137.6000 ;
	    RECT 489.2000 133.6000 490.0000 134.4000 ;
	    RECT 489.3000 132.4000 489.9000 133.6000 ;
	    RECT 489.2000 131.6000 490.0000 132.4000 ;
	    RECT 490.8000 130.2000 491.6000 135.8000 ;
	    RECT 492.4000 135.6000 493.2000 136.4000 ;
	    RECT 495.7000 132.4000 496.3000 183.6000 ;
	    RECT 497.3000 174.4000 497.9000 185.6000 ;
	    RECT 498.8000 184.2000 499.6000 195.8000 ;
	    RECT 500.5000 188.4000 501.1000 211.6000 ;
	    RECT 500.4000 187.6000 501.2000 188.4000 ;
	    RECT 502.0000 186.2000 502.8000 191.8000 ;
	    RECT 503.7000 178.3000 504.3000 237.6000 ;
	    RECT 508.4000 224.2000 509.2000 235.8000 ;
	    RECT 505.2000 211.6000 506.0000 212.4000 ;
	    RECT 508.4000 206.2000 509.2000 217.8000 ;
	    RECT 510.1000 204.3000 510.7000 251.6000 ;
	    RECT 511.7000 232.3000 512.3000 307.6000 ;
	    RECT 513.2000 255.6000 514.0000 256.4000 ;
	    RECT 513.2000 233.6000 514.0000 234.4000 ;
	    RECT 511.7000 231.7000 513.9000 232.3000 ;
	    RECT 511.6000 210.2000 512.4000 215.8000 ;
	    RECT 508.5000 203.7000 510.7000 204.3000 ;
	    RECT 505.2000 193.6000 506.0000 194.4000 ;
	    RECT 508.5000 194.3000 509.1000 203.7000 ;
	    RECT 510.0000 195.6000 510.8000 196.4000 ;
	    RECT 508.5000 193.7000 510.7000 194.3000 ;
	    RECT 506.8000 189.6000 507.6000 190.4000 ;
	    RECT 506.9000 188.4000 507.5000 189.6000 ;
	    RECT 506.8000 187.6000 507.6000 188.4000 ;
	    RECT 506.8000 183.6000 507.6000 184.4000 ;
	    RECT 497.2000 173.6000 498.0000 174.4000 ;
	    RECT 498.8000 173.6000 499.6000 174.4000 ;
	    RECT 497.3000 154.4000 497.9000 173.6000 ;
	    RECT 498.9000 172.6000 499.5000 173.6000 ;
	    RECT 498.8000 171.8000 499.6000 172.6000 ;
	    RECT 500.4000 166.2000 501.2000 177.8000 ;
	    RECT 502.1000 177.7000 504.3000 178.3000 ;
	    RECT 497.2000 153.6000 498.0000 154.4000 ;
	    RECT 497.2000 149.6000 498.0000 150.4000 ;
	    RECT 495.6000 131.6000 496.4000 132.4000 ;
	    RECT 484.4000 113.6000 485.2000 114.4000 ;
	    RECT 484.4000 109.4000 485.2000 110.4000 ;
	    RECT 484.4000 105.6000 485.2000 106.4000 ;
	    RECT 463.6000 99.6000 464.4000 100.4000 ;
	    RECT 468.4000 97.6000 469.2000 98.4000 ;
	    RECT 468.5000 94.4000 469.1000 97.6000 ;
	    RECT 465.2000 93.6000 466.0000 94.4000 ;
	    RECT 468.4000 93.6000 469.2000 94.4000 ;
	    RECT 462.0000 91.6000 462.8000 92.4000 ;
	    RECT 463.6000 91.6000 464.4000 92.4000 ;
	    RECT 468.5000 90.4000 469.1000 93.6000 ;
	    RECT 466.8000 89.6000 467.6000 90.4000 ;
	    RECT 468.4000 89.6000 469.2000 90.4000 ;
	    RECT 466.9000 88.4000 467.5000 89.6000 ;
	    RECT 460.4000 87.6000 461.2000 88.4000 ;
	    RECT 466.8000 87.6000 467.6000 88.4000 ;
	    RECT 462.0000 85.6000 462.8000 86.4000 ;
	    RECT 473.2000 86.2000 474.0000 97.8000 ;
	    RECT 481.2000 95.6000 482.0000 96.4000 ;
	    RECT 481.3000 92.6000 481.9000 95.6000 ;
	    RECT 474.8000 91.6000 475.6000 92.4000 ;
	    RECT 478.0000 91.6000 478.8000 92.4000 ;
	    RECT 481.2000 91.8000 482.0000 92.6000 ;
	    RECT 474.9000 86.4000 475.5000 91.6000 ;
	    RECT 474.8000 85.6000 475.6000 86.4000 ;
	    RECT 462.1000 80.4000 462.7000 85.6000 ;
	    RECT 455.6000 79.6000 456.4000 80.4000 ;
	    RECT 462.0000 79.6000 462.8000 80.4000 ;
	    RECT 455.6000 73.6000 456.4000 74.4000 ;
	    RECT 454.0000 71.6000 454.8000 72.4000 ;
	    RECT 450.8000 69.6000 451.6000 70.4000 ;
	    RECT 450.9000 68.4000 451.5000 69.6000 ;
	    RECT 450.8000 67.6000 451.6000 68.4000 ;
	    RECT 446.0000 65.6000 446.8000 66.4000 ;
	    RECT 446.1000 64.4000 446.7000 65.6000 ;
	    RECT 446.0000 63.6000 446.8000 64.4000 ;
	    RECT 454.0000 63.6000 454.8000 64.4000 ;
	    RECT 460.4000 64.2000 461.2000 75.8000 ;
	    RECT 462.1000 70.4000 462.7000 79.6000 ;
	    RECT 468.4000 71.6000 469.2000 72.4000 ;
	    RECT 462.0000 69.6000 462.8000 70.4000 ;
	    RECT 468.5000 70.2000 469.1000 71.6000 ;
	    RECT 444.4000 58.3000 445.2000 58.4000 ;
	    RECT 446.1000 58.3000 446.7000 63.6000 ;
	    RECT 444.4000 57.7000 446.7000 58.3000 ;
	    RECT 444.4000 57.6000 445.2000 57.7000 ;
	    RECT 442.9000 55.7000 445.1000 56.3000 ;
	    RECT 442.8000 53.6000 443.6000 54.4000 ;
	    RECT 442.9000 52.4000 443.5000 53.6000 ;
	    RECT 428.4000 51.6000 429.2000 52.4000 ;
	    RECT 431.6000 51.6000 432.4000 52.4000 ;
	    RECT 436.4000 51.6000 437.2000 52.4000 ;
	    RECT 439.6000 51.6000 440.4000 52.4000 ;
	    RECT 442.8000 51.6000 443.6000 52.4000 ;
	    RECT 431.7000 50.4000 432.3000 51.6000 ;
	    RECT 431.6000 49.6000 432.4000 50.4000 ;
	    RECT 425.2000 29.6000 426.0000 30.4000 ;
	    RECT 426.8000 29.6000 427.6000 30.4000 ;
	    RECT 425.3000 28.4000 425.9000 29.6000 ;
	    RECT 425.2000 27.6000 426.0000 28.4000 ;
	    RECT 433.2000 24.2000 434.0000 35.8000 ;
	    RECT 434.8000 27.6000 435.6000 28.4000 ;
	    RECT 423.6000 19.6000 424.4000 20.4000 ;
	    RECT 401.2000 15.6000 402.0000 16.4000 ;
	    RECT 398.0000 13.6000 398.8000 14.4000 ;
	    RECT 401.3000 12.6000 401.9000 15.6000 ;
	    RECT 401.2000 11.8000 402.0000 12.6000 ;
	    RECT 401.3000 11.7000 401.9000 11.8000 ;
	    RECT 402.8000 6.2000 403.6000 17.8000 ;
	    RECT 406.0000 10.2000 406.8000 15.8000 ;
	    RECT 418.8000 15.6000 419.6000 16.4000 ;
	    RECT 423.7000 14.4000 424.3000 19.6000 ;
	    RECT 414.0000 13.6000 414.8000 14.4000 ;
	    RECT 423.6000 13.6000 424.4000 14.4000 ;
	    RECT 425.2000 13.6000 426.0000 14.4000 ;
	    RECT 414.1000 10.4000 414.7000 13.6000 ;
	    RECT 417.2000 11.6000 418.0000 12.4000 ;
	    RECT 422.0000 11.6000 422.8000 12.4000 ;
	    RECT 417.3000 10.4000 417.9000 11.6000 ;
	    RECT 414.0000 9.6000 414.8000 10.4000 ;
	    RECT 417.2000 9.6000 418.0000 10.4000 ;
	    RECT 425.3000 8.4000 425.9000 13.6000 ;
	    RECT 425.2000 7.6000 426.0000 8.4000 ;
	    RECT 430.0000 6.2000 430.8000 17.8000 ;
	    RECT 434.9000 14.4000 435.5000 27.6000 ;
	    RECT 436.4000 26.2000 437.2000 31.8000 ;
	    RECT 438.0000 25.6000 438.8000 26.4000 ;
	    RECT 438.1000 24.4000 438.7000 25.6000 ;
	    RECT 438.0000 23.6000 438.8000 24.4000 ;
	    RECT 442.8000 24.2000 443.6000 35.8000 ;
	    RECT 444.5000 24.4000 445.1000 55.7000 ;
	    RECT 446.0000 51.6000 446.8000 52.4000 ;
	    RECT 444.4000 23.6000 445.2000 24.4000 ;
	    RECT 438.1000 22.4000 438.7000 23.6000 ;
	    RECT 438.0000 21.6000 438.8000 22.4000 ;
	    RECT 434.8000 13.6000 435.6000 14.4000 ;
	    RECT 438.0000 11.8000 438.8000 12.6000 ;
	    RECT 438.1000 10.4000 438.7000 11.8000 ;
	    RECT 438.0000 9.6000 438.8000 10.4000 ;
	    RECT 439.6000 6.2000 440.4000 17.8000 ;
	    RECT 442.8000 10.2000 443.6000 15.8000 ;
	    RECT 444.5000 14.4000 445.1000 23.6000 ;
	    RECT 444.4000 13.6000 445.2000 14.4000 ;
	    RECT 446.1000 12.4000 446.7000 51.6000 ;
	    RECT 449.2000 46.2000 450.0000 57.8000 ;
	    RECT 454.1000 52.4000 454.7000 63.6000 ;
	    RECT 462.1000 62.3000 462.7000 69.6000 ;
	    RECT 468.4000 69.4000 469.2000 70.2000 ;
	    RECT 470.0000 64.2000 470.8000 75.8000 ;
	    RECT 474.8000 73.6000 475.6000 74.4000 ;
	    RECT 473.2000 66.2000 474.0000 71.8000 ;
	    RECT 474.9000 66.4000 475.5000 73.6000 ;
	    RECT 478.1000 70.4000 478.7000 91.6000 ;
	    RECT 482.8000 86.2000 483.6000 97.8000 ;
	    RECT 484.5000 94.4000 485.1000 105.6000 ;
	    RECT 486.0000 104.2000 486.8000 115.8000 ;
	    RECT 495.7000 114.3000 496.3000 131.6000 ;
	    RECT 494.1000 113.7000 496.3000 114.3000 ;
	    RECT 489.2000 106.2000 490.0000 111.8000 ;
	    RECT 490.8000 111.6000 491.6000 112.4000 ;
	    RECT 490.9000 106.4000 491.5000 111.6000 ;
	    RECT 494.1000 110.4000 494.7000 113.7000 ;
	    RECT 495.6000 111.6000 496.4000 112.4000 ;
	    RECT 495.7000 110.4000 496.3000 111.6000 ;
	    RECT 494.0000 109.6000 494.8000 110.4000 ;
	    RECT 495.6000 109.6000 496.4000 110.4000 ;
	    RECT 490.8000 105.6000 491.6000 106.4000 ;
	    RECT 494.1000 98.3000 494.7000 109.6000 ;
	    RECT 497.3000 100.3000 497.9000 149.6000 ;
	    RECT 498.8000 144.2000 499.6000 155.8000 ;
	    RECT 502.1000 136.4000 502.7000 177.7000 ;
	    RECT 503.6000 170.2000 504.4000 175.8000 ;
	    RECT 505.2000 175.6000 506.0000 176.4000 ;
	    RECT 505.3000 172.4000 505.9000 175.6000 ;
	    RECT 506.9000 172.4000 507.5000 183.6000 ;
	    RECT 510.1000 172.4000 510.7000 193.7000 ;
	    RECT 513.3000 190.4000 513.9000 231.7000 ;
	    RECT 513.2000 189.6000 514.0000 190.4000 ;
	    RECT 511.6000 173.6000 512.4000 174.4000 ;
	    RECT 505.2000 171.6000 506.0000 172.4000 ;
	    RECT 506.8000 171.6000 507.6000 172.4000 ;
	    RECT 510.0000 171.6000 510.8000 172.4000 ;
	    RECT 513.2000 171.6000 514.0000 172.4000 ;
	    RECT 503.6000 149.6000 504.4000 150.4000 ;
	    RECT 502.0000 135.6000 502.8000 136.4000 ;
	    RECT 498.8000 133.6000 499.6000 134.4000 ;
	    RECT 502.0000 133.6000 502.8000 134.4000 ;
	    RECT 503.7000 132.4000 504.3000 149.6000 ;
	    RECT 506.8000 149.4000 507.6000 150.2000 ;
	    RECT 505.2000 147.6000 506.0000 148.4000 ;
	    RECT 505.3000 132.4000 505.9000 147.6000 ;
	    RECT 506.9000 138.4000 507.5000 149.4000 ;
	    RECT 508.4000 144.2000 509.2000 155.8000 ;
	    RECT 510.1000 150.4000 510.7000 171.6000 ;
	    RECT 513.3000 170.4000 513.9000 171.6000 ;
	    RECT 513.2000 169.6000 514.0000 170.4000 ;
	    RECT 510.0000 149.6000 510.8000 150.4000 ;
	    RECT 511.6000 146.2000 512.4000 151.8000 ;
	    RECT 511.6000 139.6000 512.4000 140.4000 ;
	    RECT 506.8000 137.6000 507.6000 138.4000 ;
	    RECT 503.6000 131.6000 504.4000 132.4000 ;
	    RECT 505.2000 131.6000 506.0000 132.4000 ;
	    RECT 510.0000 131.6000 510.8000 132.4000 ;
	    RECT 500.4000 130.3000 501.2000 130.4000 ;
	    RECT 500.4000 129.7000 502.7000 130.3000 ;
	    RECT 500.4000 129.6000 501.2000 129.7000 ;
	    RECT 502.1000 118.4000 502.7000 129.7000 ;
	    RECT 498.8000 117.6000 499.6000 118.4000 ;
	    RECT 502.0000 117.6000 502.8000 118.4000 ;
	    RECT 498.9000 112.4000 499.5000 117.6000 ;
	    RECT 502.0000 113.6000 502.8000 114.4000 ;
	    RECT 503.6000 113.6000 504.4000 114.4000 ;
	    RECT 498.8000 111.6000 499.6000 112.4000 ;
	    RECT 502.1000 110.4000 502.7000 113.6000 ;
	    RECT 498.8000 109.6000 499.6000 110.4000 ;
	    RECT 502.0000 109.6000 502.8000 110.4000 ;
	    RECT 492.5000 97.7000 494.7000 98.3000 ;
	    RECT 495.7000 99.7000 497.9000 100.3000 ;
	    RECT 484.4000 93.6000 485.2000 94.4000 ;
	    RECT 486.0000 90.2000 486.8000 95.8000 ;
	    RECT 487.6000 95.6000 488.4000 96.4000 ;
	    RECT 492.5000 92.4000 493.1000 97.7000 ;
	    RECT 494.0000 95.6000 494.8000 96.4000 ;
	    RECT 494.1000 94.4000 494.7000 95.6000 ;
	    RECT 494.0000 93.6000 494.8000 94.4000 ;
	    RECT 492.4000 91.6000 493.2000 92.4000 ;
	    RECT 487.6000 89.6000 488.4000 90.4000 ;
	    RECT 486.0000 79.6000 486.8000 80.4000 ;
	    RECT 486.1000 74.4000 486.7000 79.6000 ;
	    RECT 487.7000 78.4000 488.3000 89.6000 ;
	    RECT 487.6000 77.6000 488.4000 78.4000 ;
	    RECT 482.8000 73.6000 483.6000 74.4000 ;
	    RECT 486.0000 73.6000 486.8000 74.4000 ;
	    RECT 482.9000 72.4000 483.5000 73.6000 ;
	    RECT 479.6000 71.6000 480.4000 72.4000 ;
	    RECT 482.8000 71.6000 483.6000 72.4000 ;
	    RECT 478.0000 69.6000 478.8000 70.4000 ;
	    RECT 474.8000 65.6000 475.6000 66.4000 ;
	    RECT 460.5000 61.7000 462.7000 62.3000 ;
	    RECT 450.8000 51.6000 451.6000 52.4000 ;
	    RECT 454.0000 51.6000 454.8000 52.4000 ;
	    RECT 449.2000 31.6000 450.0000 32.4000 ;
	    RECT 449.3000 30.4000 449.9000 31.6000 ;
	    RECT 449.2000 29.6000 450.0000 30.4000 ;
	    RECT 450.9000 28.4000 451.5000 51.6000 ;
	    RECT 458.8000 46.2000 459.6000 57.8000 ;
	    RECT 460.5000 54.4000 461.1000 61.7000 ;
	    RECT 463.6000 61.6000 464.4000 62.4000 ;
	    RECT 463.7000 58.4000 464.3000 61.6000 ;
	    RECT 463.6000 57.6000 464.4000 58.4000 ;
	    RECT 482.8000 57.6000 483.6000 58.4000 ;
	    RECT 460.4000 53.6000 461.2000 54.4000 ;
	    RECT 462.0000 50.2000 462.8000 55.8000 ;
	    RECT 473.2000 55.6000 474.0000 56.4000 ;
	    RECT 470.0000 51.6000 470.8000 52.4000 ;
	    RECT 478.0000 51.6000 478.8000 52.4000 ;
	    RECT 486.1000 48.4000 486.7000 73.6000 ;
	    RECT 487.6000 71.6000 488.4000 72.4000 ;
	    RECT 487.7000 70.4000 488.3000 71.6000 ;
	    RECT 495.7000 70.4000 496.3000 99.7000 ;
	    RECT 498.9000 92.4000 499.5000 109.6000 ;
	    RECT 505.3000 94.4000 505.9000 131.6000 ;
	    RECT 506.8000 129.6000 507.6000 130.4000 ;
	    RECT 506.9000 128.4000 507.5000 129.6000 ;
	    RECT 511.7000 128.4000 512.3000 139.6000 ;
	    RECT 506.8000 127.6000 507.6000 128.4000 ;
	    RECT 510.0000 127.6000 510.8000 128.4000 ;
	    RECT 511.6000 127.6000 512.4000 128.4000 ;
	    RECT 510.1000 126.4000 510.7000 127.6000 ;
	    RECT 510.0000 125.6000 510.8000 126.4000 ;
	    RECT 508.4000 117.6000 509.2000 118.4000 ;
	    RECT 510.0000 114.3000 510.8000 114.4000 ;
	    RECT 511.7000 114.3000 512.3000 127.6000 ;
	    RECT 510.0000 113.7000 512.3000 114.3000 ;
	    RECT 510.0000 113.6000 510.8000 113.7000 ;
	    RECT 506.8000 109.6000 507.6000 110.4000 ;
	    RECT 508.4000 109.6000 509.2000 110.4000 ;
	    RECT 502.0000 93.6000 502.8000 94.4000 ;
	    RECT 505.2000 93.6000 506.0000 94.4000 ;
	    RECT 498.8000 91.6000 499.6000 92.4000 ;
	    RECT 498.8000 87.6000 499.6000 88.4000 ;
	    RECT 500.4000 87.6000 501.2000 88.4000 ;
	    RECT 498.9000 86.4000 499.5000 87.6000 ;
	    RECT 498.8000 85.6000 499.6000 86.4000 ;
	    RECT 500.5000 80.4000 501.1000 87.6000 ;
	    RECT 500.4000 79.6000 501.2000 80.4000 ;
	    RECT 502.1000 78.4000 502.7000 93.6000 ;
	    RECT 506.9000 92.4000 507.5000 109.6000 ;
	    RECT 506.8000 91.6000 507.6000 92.4000 ;
	    RECT 505.2000 87.6000 506.0000 88.4000 ;
	    RECT 503.6000 83.6000 504.4000 84.4000 ;
	    RECT 502.0000 77.6000 502.8000 78.4000 ;
	    RECT 498.8000 75.6000 499.6000 76.4000 ;
	    RECT 498.9000 72.4000 499.5000 75.6000 ;
	    RECT 503.7000 74.4000 504.3000 83.6000 ;
	    RECT 505.3000 80.4000 505.9000 87.6000 ;
	    RECT 505.2000 79.6000 506.0000 80.4000 ;
	    RECT 503.6000 73.6000 504.4000 74.4000 ;
	    RECT 506.9000 72.4000 507.5000 91.6000 ;
	    RECT 498.8000 71.6000 499.6000 72.4000 ;
	    RECT 506.8000 71.6000 507.6000 72.4000 ;
	    RECT 487.6000 69.6000 488.4000 70.4000 ;
	    RECT 495.6000 69.6000 496.4000 70.4000 ;
	    RECT 495.7000 68.4000 496.3000 69.6000 ;
	    RECT 495.6000 67.6000 496.4000 68.4000 ;
	    RECT 490.8000 65.6000 491.6000 66.4000 ;
	    RECT 490.9000 60.4000 491.5000 65.6000 ;
	    RECT 490.8000 59.6000 491.6000 60.4000 ;
	    RECT 490.9000 58.3000 491.5000 59.6000 ;
	    RECT 492.4000 58.3000 493.2000 58.4000 ;
	    RECT 490.9000 57.7000 493.2000 58.3000 ;
	    RECT 492.4000 57.6000 493.2000 57.7000 ;
	    RECT 489.2000 51.6000 490.0000 52.4000 ;
	    RECT 468.4000 47.6000 469.2000 48.4000 ;
	    RECT 479.6000 47.6000 480.4000 48.4000 ;
	    RECT 486.0000 48.3000 486.8000 48.4000 ;
	    RECT 487.6000 48.3000 488.4000 48.4000 ;
	    RECT 486.0000 47.7000 488.4000 48.3000 ;
	    RECT 486.0000 47.6000 486.8000 47.7000 ;
	    RECT 487.6000 47.6000 488.4000 47.7000 ;
	    RECT 463.6000 43.6000 464.4000 44.4000 ;
	    RECT 470.0000 43.6000 470.8000 44.4000 ;
	    RECT 478.0000 43.6000 478.8000 44.4000 ;
	    RECT 489.2000 43.6000 490.0000 44.4000 ;
	    RECT 450.8000 27.6000 451.6000 28.4000 ;
	    RECT 452.4000 24.2000 453.2000 35.8000 ;
	    RECT 457.2000 35.6000 458.0000 36.4000 ;
	    RECT 457.3000 32.4000 457.9000 35.6000 ;
	    RECT 454.0000 27.6000 454.8000 28.4000 ;
	    RECT 455.6000 26.2000 456.4000 31.8000 ;
	    RECT 457.2000 31.6000 458.0000 32.4000 ;
	    RECT 455.6000 19.6000 456.4000 20.4000 ;
	    RECT 455.7000 14.4000 456.3000 19.6000 ;
	    RECT 454.0000 13.6000 454.8000 14.4000 ;
	    RECT 455.6000 13.6000 456.4000 14.4000 ;
	    RECT 457.3000 12.4000 457.9000 31.6000 ;
	    RECT 460.4000 27.6000 461.2000 28.4000 ;
	    RECT 458.8000 23.6000 459.6000 24.4000 ;
	    RECT 460.5000 24.3000 461.1000 27.6000 ;
	    RECT 462.0000 25.6000 462.8000 26.4000 ;
	    RECT 460.5000 23.7000 462.7000 24.3000 ;
	    RECT 446.0000 11.6000 446.8000 12.4000 ;
	    RECT 447.6000 11.6000 448.4000 12.4000 ;
	    RECT 450.8000 11.6000 451.6000 12.4000 ;
	    RECT 457.2000 11.6000 458.0000 12.4000 ;
	    RECT 447.7000 10.4000 448.3000 11.6000 ;
	    RECT 450.9000 10.4000 451.5000 11.6000 ;
	    RECT 447.6000 9.6000 448.4000 10.4000 ;
	    RECT 450.8000 9.6000 451.6000 10.4000 ;
	    RECT 458.9000 10.3000 459.5000 23.6000 ;
	    RECT 462.1000 18.4000 462.7000 23.7000 ;
	    RECT 463.7000 20.4000 464.3000 43.6000 ;
	    RECT 470.1000 32.4000 470.7000 43.6000 ;
	    RECT 476.4000 37.6000 477.2000 38.4000 ;
	    RECT 466.8000 31.6000 467.6000 32.4000 ;
	    RECT 470.0000 31.6000 470.8000 32.4000 ;
	    RECT 476.5000 30.4000 477.1000 37.6000 ;
	    RECT 478.1000 32.3000 478.7000 43.6000 ;
	    RECT 486.0000 37.6000 486.8000 38.4000 ;
	    RECT 481.2000 33.6000 482.0000 34.4000 ;
	    RECT 479.6000 32.3000 480.4000 32.4000 ;
	    RECT 478.1000 31.7000 480.4000 32.3000 ;
	    RECT 479.6000 31.6000 480.4000 31.7000 ;
	    RECT 466.8000 29.6000 467.6000 30.4000 ;
	    RECT 476.4000 29.6000 477.2000 30.4000 ;
	    RECT 468.4000 27.6000 469.2000 28.4000 ;
	    RECT 463.6000 19.6000 464.4000 20.4000 ;
	    RECT 462.0000 17.6000 462.8000 18.4000 ;
	    RECT 460.4000 13.6000 461.2000 14.4000 ;
	    RECT 460.4000 10.3000 461.2000 10.4000 ;
	    RECT 458.9000 9.7000 461.2000 10.3000 ;
	    RECT 460.4000 9.6000 461.2000 9.7000 ;
	    RECT 466.8000 6.2000 467.6000 17.8000 ;
	    RECT 468.5000 14.4000 469.1000 27.6000 ;
	    RECT 481.3000 26.4000 481.9000 33.6000 ;
	    RECT 486.1000 30.4000 486.7000 37.6000 ;
	    RECT 489.3000 32.4000 489.9000 43.6000 ;
	    RECT 495.7000 38.4000 496.3000 67.6000 ;
	    RECT 498.8000 63.6000 499.6000 64.4000 ;
	    RECT 497.2000 46.2000 498.0000 57.8000 ;
	    RECT 498.9000 52.3000 499.5000 63.6000 ;
	    RECT 502.0000 53.6000 502.8000 54.4000 ;
	    RECT 500.4000 52.3000 501.2000 52.4000 ;
	    RECT 498.9000 51.7000 501.2000 52.3000 ;
	    RECT 500.4000 51.6000 501.2000 51.7000 ;
	    RECT 495.6000 37.6000 496.4000 38.4000 ;
	    RECT 490.8000 33.6000 491.6000 34.4000 ;
	    RECT 489.2000 31.6000 490.0000 32.4000 ;
	    RECT 486.0000 29.6000 486.8000 30.4000 ;
	    RECT 489.2000 29.6000 490.0000 30.4000 ;
	    RECT 471.6000 25.6000 472.4000 26.4000 ;
	    RECT 481.2000 25.6000 482.0000 26.4000 ;
	    RECT 471.7000 18.4000 472.3000 25.6000 ;
	    RECT 479.6000 23.6000 480.4000 24.4000 ;
	    RECT 495.6000 24.2000 496.4000 35.8000 ;
	    RECT 500.4000 29.6000 501.2000 30.4000 ;
	    RECT 502.1000 28.4000 502.7000 53.6000 ;
	    RECT 506.8000 46.2000 507.6000 57.8000 ;
	    RECT 510.0000 50.2000 510.8000 55.8000 ;
	    RECT 497.2000 27.6000 498.0000 28.4000 ;
	    RECT 502.0000 27.6000 502.8000 28.4000 ;
	    RECT 479.7000 20.4000 480.3000 23.6000 ;
	    RECT 479.6000 19.6000 480.4000 20.4000 ;
	    RECT 492.4000 19.6000 493.2000 20.4000 ;
	    RECT 471.6000 17.6000 472.4000 18.4000 ;
	    RECT 468.4000 13.6000 469.2000 14.4000 ;
	    RECT 470.0000 13.6000 470.8000 14.4000 ;
	    RECT 470.1000 12.4000 470.7000 13.6000 ;
	    RECT 470.0000 11.6000 470.8000 12.4000 ;
	    RECT 476.4000 6.2000 477.2000 17.8000 ;
	    RECT 481.2000 17.6000 482.0000 18.4000 ;
	    RECT 478.0000 13.6000 478.8000 14.4000 ;
	    RECT 479.6000 10.2000 480.4000 15.8000 ;
	    RECT 486.0000 6.2000 486.8000 17.8000 ;
	    RECT 487.6000 13.6000 488.4000 14.4000 ;
	    RECT 492.5000 12.4000 493.1000 19.6000 ;
	    RECT 492.4000 11.6000 493.2000 12.4000 ;
	    RECT 495.6000 6.2000 496.4000 17.8000 ;
	    RECT 497.3000 14.4000 497.9000 27.6000 ;
	    RECT 502.1000 18.4000 502.7000 27.6000 ;
	    RECT 505.2000 24.2000 506.0000 35.8000 ;
	    RECT 508.4000 26.2000 509.2000 31.8000 ;
	    RECT 502.0000 17.6000 502.8000 18.4000 ;
	    RECT 497.2000 13.6000 498.0000 14.4000 ;
	    RECT 498.8000 10.2000 499.6000 15.8000 ;
	    RECT 338.8000 3.6000 339.6000 4.4000 ;
	    RECT 462.0000 3.6000 462.8000 4.4000 ;
	    RECT 276.4000 1.6000 277.2000 2.4000 ;
	    RECT 332.4000 1.6000 333.2000 2.4000 ;
         LAYER metal3 ;
	    RECT 130.8000 338.3000 131.6000 338.4000 ;
	    RECT 150.0000 338.3000 150.8000 338.4000 ;
	    RECT 151.6000 338.3000 152.4000 338.4000 ;
	    RECT 130.8000 337.7000 152.4000 338.3000 ;
	    RECT 130.8000 337.6000 131.6000 337.7000 ;
	    RECT 150.0000 337.6000 150.8000 337.7000 ;
	    RECT 151.6000 337.6000 152.4000 337.7000 ;
	    RECT 263.6000 338.3000 264.4000 338.4000 ;
	    RECT 292.4000 338.3000 293.2000 338.4000 ;
	    RECT 430.0000 338.3000 430.8000 338.4000 ;
	    RECT 439.6000 338.3000 440.4000 338.4000 ;
	    RECT 263.6000 337.7000 440.4000 338.3000 ;
	    RECT 263.6000 337.6000 264.4000 337.7000 ;
	    RECT 292.4000 337.6000 293.2000 337.7000 ;
	    RECT 430.0000 337.6000 430.8000 337.7000 ;
	    RECT 439.6000 337.6000 440.4000 337.7000 ;
	    RECT 14.0000 336.3000 14.8000 336.4000 ;
	    RECT 36.4000 336.3000 37.2000 336.4000 ;
	    RECT 164.4000 336.3000 165.2000 336.4000 ;
	    RECT 193.2000 336.3000 194.0000 336.4000 ;
	    RECT 14.0000 335.7000 37.2000 336.3000 ;
	    RECT 14.0000 335.6000 14.8000 335.7000 ;
	    RECT 36.4000 335.6000 37.2000 335.7000 ;
	    RECT 159.7000 335.7000 194.0000 336.3000 ;
	    RECT 159.7000 334.4000 160.3000 335.7000 ;
	    RECT 164.4000 335.6000 165.2000 335.7000 ;
	    RECT 193.2000 335.6000 194.0000 335.7000 ;
	    RECT 242.8000 336.3000 243.6000 336.4000 ;
	    RECT 262.0000 336.3000 262.8000 336.4000 ;
	    RECT 242.8000 335.7000 262.8000 336.3000 ;
	    RECT 242.8000 335.6000 243.6000 335.7000 ;
	    RECT 262.0000 335.6000 262.8000 335.7000 ;
	    RECT 263.6000 336.3000 264.4000 336.4000 ;
	    RECT 279.6000 336.3000 280.4000 336.4000 ;
	    RECT 263.6000 335.7000 280.4000 336.3000 ;
	    RECT 263.6000 335.6000 264.4000 335.7000 ;
	    RECT 279.6000 335.6000 280.4000 335.7000 ;
	    RECT 284.4000 336.3000 285.2000 336.4000 ;
	    RECT 294.0000 336.3000 294.8000 336.4000 ;
	    RECT 335.6000 336.3000 336.4000 336.4000 ;
	    RECT 346.8000 336.3000 347.6000 336.4000 ;
	    RECT 284.4000 335.7000 347.6000 336.3000 ;
	    RECT 284.4000 335.6000 285.2000 335.7000 ;
	    RECT 294.0000 335.6000 294.8000 335.7000 ;
	    RECT 335.6000 335.6000 336.4000 335.7000 ;
	    RECT 346.8000 335.6000 347.6000 335.7000 ;
	    RECT 34.8000 334.3000 35.6000 334.4000 ;
	    RECT 47.6000 334.3000 48.4000 334.4000 ;
	    RECT 34.8000 333.7000 48.4000 334.3000 ;
	    RECT 34.8000 333.6000 35.6000 333.7000 ;
	    RECT 47.6000 333.6000 48.4000 333.7000 ;
	    RECT 66.8000 334.3000 67.6000 334.4000 ;
	    RECT 73.2000 334.3000 74.0000 334.4000 ;
	    RECT 66.8000 333.7000 74.0000 334.3000 ;
	    RECT 66.8000 333.6000 67.6000 333.7000 ;
	    RECT 73.2000 333.6000 74.0000 333.7000 ;
	    RECT 106.8000 334.3000 107.6000 334.4000 ;
	    RECT 122.8000 334.3000 123.6000 334.4000 ;
	    RECT 106.8000 333.7000 123.6000 334.3000 ;
	    RECT 106.8000 333.6000 107.6000 333.7000 ;
	    RECT 122.8000 333.6000 123.6000 333.7000 ;
	    RECT 129.2000 334.3000 130.0000 334.4000 ;
	    RECT 159.6000 334.3000 160.4000 334.4000 ;
	    RECT 129.2000 333.7000 160.4000 334.3000 ;
	    RECT 129.2000 333.6000 130.0000 333.7000 ;
	    RECT 159.6000 333.6000 160.4000 333.7000 ;
	    RECT 183.6000 334.3000 184.4000 334.4000 ;
	    RECT 217.2000 334.3000 218.0000 334.4000 ;
	    RECT 183.6000 333.7000 218.0000 334.3000 ;
	    RECT 183.6000 333.6000 184.4000 333.7000 ;
	    RECT 217.2000 333.6000 218.0000 333.7000 ;
	    RECT 218.8000 334.3000 219.6000 334.4000 ;
	    RECT 222.0000 334.3000 222.8000 334.4000 ;
	    RECT 218.8000 333.7000 222.8000 334.3000 ;
	    RECT 218.8000 333.6000 219.6000 333.7000 ;
	    RECT 222.0000 333.6000 222.8000 333.7000 ;
	    RECT 255.6000 334.3000 256.4000 334.4000 ;
	    RECT 274.8000 334.3000 275.6000 334.4000 ;
	    RECT 255.6000 333.7000 275.6000 334.3000 ;
	    RECT 255.6000 333.6000 256.4000 333.7000 ;
	    RECT 274.8000 333.6000 275.6000 333.7000 ;
	    RECT 278.0000 334.3000 278.8000 334.4000 ;
	    RECT 289.2000 334.3000 290.0000 334.4000 ;
	    RECT 298.8000 334.3000 299.6000 334.4000 ;
	    RECT 278.0000 333.7000 299.6000 334.3000 ;
	    RECT 278.0000 333.6000 278.8000 333.7000 ;
	    RECT 289.2000 333.6000 290.0000 333.7000 ;
	    RECT 298.8000 333.6000 299.6000 333.7000 ;
	    RECT 303.6000 334.3000 304.4000 334.4000 ;
	    RECT 313.2000 334.3000 314.0000 334.4000 ;
	    RECT 303.6000 333.7000 314.0000 334.3000 ;
	    RECT 303.6000 333.6000 304.4000 333.7000 ;
	    RECT 313.2000 333.6000 314.0000 333.7000 ;
	    RECT 332.4000 334.3000 333.2000 334.4000 ;
	    RECT 362.8000 334.3000 363.6000 334.4000 ;
	    RECT 378.8000 334.3000 379.6000 334.4000 ;
	    RECT 332.4000 333.7000 379.6000 334.3000 ;
	    RECT 332.4000 333.6000 333.2000 333.7000 ;
	    RECT 362.8000 333.6000 363.6000 333.7000 ;
	    RECT 378.8000 333.6000 379.6000 333.7000 ;
	    RECT 438.0000 334.3000 438.8000 334.4000 ;
	    RECT 450.8000 334.3000 451.6000 334.4000 ;
	    RECT 438.0000 333.7000 451.6000 334.3000 ;
	    RECT 438.0000 333.6000 438.8000 333.7000 ;
	    RECT 450.8000 333.6000 451.6000 333.7000 ;
	    RECT 462.0000 334.3000 462.8000 334.4000 ;
	    RECT 503.6000 334.3000 504.4000 334.4000 ;
	    RECT 462.0000 333.7000 504.4000 334.3000 ;
	    RECT 462.0000 333.6000 462.8000 333.7000 ;
	    RECT 503.6000 333.6000 504.4000 333.7000 ;
	    RECT 1.2000 332.3000 2.0000 332.4000 ;
	    RECT 23.6000 332.3000 24.4000 332.4000 ;
	    RECT 30.0000 332.3000 30.8000 332.4000 ;
	    RECT 1.2000 331.7000 30.8000 332.3000 ;
	    RECT 1.2000 331.6000 2.0000 331.7000 ;
	    RECT 23.6000 331.6000 24.4000 331.7000 ;
	    RECT 30.0000 331.6000 30.8000 331.7000 ;
	    RECT 34.8000 332.3000 35.6000 332.4000 ;
	    RECT 49.2000 332.3000 50.0000 332.4000 ;
	    RECT 34.8000 331.7000 50.0000 332.3000 ;
	    RECT 34.8000 331.6000 35.6000 331.7000 ;
	    RECT 49.2000 331.6000 50.0000 331.7000 ;
	    RECT 52.4000 332.3000 53.2000 332.4000 ;
	    RECT 73.2000 332.3000 74.0000 332.4000 ;
	    RECT 52.4000 331.7000 74.0000 332.3000 ;
	    RECT 52.4000 331.6000 53.2000 331.7000 ;
	    RECT 73.2000 331.6000 74.0000 331.7000 ;
	    RECT 122.8000 332.3000 123.6000 332.4000 ;
	    RECT 127.6000 332.3000 128.4000 332.4000 ;
	    RECT 129.2000 332.3000 130.0000 332.4000 ;
	    RECT 122.8000 331.7000 130.0000 332.3000 ;
	    RECT 122.8000 331.6000 123.6000 331.7000 ;
	    RECT 127.6000 331.6000 128.4000 331.7000 ;
	    RECT 129.2000 331.6000 130.0000 331.7000 ;
	    RECT 143.6000 332.3000 144.4000 332.4000 ;
	    RECT 153.2000 332.3000 154.0000 332.4000 ;
	    RECT 143.6000 331.7000 154.0000 332.3000 ;
	    RECT 143.6000 331.6000 144.4000 331.7000 ;
	    RECT 153.2000 331.6000 154.0000 331.7000 ;
	    RECT 174.0000 332.3000 174.8000 332.4000 ;
	    RECT 186.8000 332.3000 187.6000 332.4000 ;
	    RECT 174.0000 331.7000 187.6000 332.3000 ;
	    RECT 174.0000 331.6000 174.8000 331.7000 ;
	    RECT 186.8000 331.6000 187.6000 331.7000 ;
	    RECT 190.0000 332.3000 190.8000 332.4000 ;
	    RECT 225.2000 332.3000 226.0000 332.4000 ;
	    RECT 190.0000 331.7000 226.0000 332.3000 ;
	    RECT 190.0000 331.6000 190.8000 331.7000 ;
	    RECT 225.2000 331.6000 226.0000 331.7000 ;
	    RECT 234.8000 332.3000 235.6000 332.4000 ;
	    RECT 241.2000 332.3000 242.0000 332.4000 ;
	    RECT 249.2000 332.3000 250.0000 332.4000 ;
	    RECT 263.6000 332.3000 264.4000 332.4000 ;
	    RECT 234.8000 331.7000 250.0000 332.3000 ;
	    RECT 234.8000 331.6000 235.6000 331.7000 ;
	    RECT 241.2000 331.6000 242.0000 331.7000 ;
	    RECT 249.2000 331.6000 250.0000 331.7000 ;
	    RECT 250.9000 331.7000 264.4000 332.3000 ;
	    RECT 33.2000 330.3000 34.0000 330.4000 ;
	    RECT 36.4000 330.3000 37.2000 330.4000 ;
	    RECT 33.2000 329.7000 37.2000 330.3000 ;
	    RECT 33.2000 329.6000 34.0000 329.7000 ;
	    RECT 36.4000 329.6000 37.2000 329.7000 ;
	    RECT 46.0000 330.3000 46.8000 330.4000 ;
	    RECT 52.4000 330.3000 53.2000 330.4000 ;
	    RECT 46.0000 329.7000 53.2000 330.3000 ;
	    RECT 46.0000 329.6000 46.8000 329.7000 ;
	    RECT 52.4000 329.6000 53.2000 329.7000 ;
	    RECT 100.4000 330.3000 101.2000 330.4000 ;
	    RECT 137.2000 330.3000 138.0000 330.4000 ;
	    RECT 156.4000 330.3000 157.2000 330.4000 ;
	    RECT 100.4000 329.7000 157.2000 330.3000 ;
	    RECT 100.4000 329.6000 101.2000 329.7000 ;
	    RECT 137.2000 329.6000 138.0000 329.7000 ;
	    RECT 156.4000 329.6000 157.2000 329.7000 ;
	    RECT 183.6000 330.3000 184.4000 330.4000 ;
	    RECT 186.8000 330.3000 187.6000 330.4000 ;
	    RECT 183.6000 329.7000 187.6000 330.3000 ;
	    RECT 183.6000 329.6000 184.4000 329.7000 ;
	    RECT 186.8000 329.6000 187.6000 329.7000 ;
	    RECT 207.6000 330.3000 208.4000 330.4000 ;
	    RECT 234.8000 330.3000 235.6000 330.4000 ;
	    RECT 207.6000 329.7000 235.6000 330.3000 ;
	    RECT 207.6000 329.6000 208.4000 329.7000 ;
	    RECT 234.8000 329.6000 235.6000 329.7000 ;
	    RECT 242.8000 330.3000 243.6000 330.4000 ;
	    RECT 250.9000 330.3000 251.5000 331.7000 ;
	    RECT 263.6000 331.6000 264.4000 331.7000 ;
	    RECT 273.2000 331.6000 274.0000 332.4000 ;
	    RECT 279.6000 332.3000 280.4000 332.4000 ;
	    RECT 286.0000 332.3000 286.8000 332.4000 ;
	    RECT 279.6000 331.7000 286.8000 332.3000 ;
	    RECT 279.6000 331.6000 280.4000 331.7000 ;
	    RECT 286.0000 331.6000 286.8000 331.7000 ;
	    RECT 295.6000 332.3000 296.4000 332.4000 ;
	    RECT 305.2000 332.3000 306.0000 332.4000 ;
	    RECT 295.6000 331.7000 306.0000 332.3000 ;
	    RECT 295.6000 331.6000 296.4000 331.7000 ;
	    RECT 305.2000 331.6000 306.0000 331.7000 ;
	    RECT 338.8000 332.3000 339.6000 332.4000 ;
	    RECT 343.6000 332.3000 344.4000 332.4000 ;
	    RECT 338.8000 331.7000 344.4000 332.3000 ;
	    RECT 338.8000 331.6000 339.6000 331.7000 ;
	    RECT 343.6000 331.6000 344.4000 331.7000 ;
	    RECT 345.2000 332.3000 346.0000 332.4000 ;
	    RECT 366.0000 332.3000 366.8000 332.4000 ;
	    RECT 345.2000 331.7000 366.8000 332.3000 ;
	    RECT 345.2000 331.6000 346.0000 331.7000 ;
	    RECT 366.0000 331.6000 366.8000 331.7000 ;
	    RECT 391.6000 332.3000 392.4000 332.4000 ;
	    RECT 393.2000 332.3000 394.0000 332.4000 ;
	    RECT 391.6000 331.7000 394.0000 332.3000 ;
	    RECT 391.6000 331.6000 392.4000 331.7000 ;
	    RECT 393.2000 331.6000 394.0000 331.7000 ;
	    RECT 418.8000 332.3000 419.6000 332.4000 ;
	    RECT 425.2000 332.3000 426.0000 332.4000 ;
	    RECT 462.0000 332.3000 462.8000 332.4000 ;
	    RECT 418.8000 331.7000 462.8000 332.3000 ;
	    RECT 418.8000 331.6000 419.6000 331.7000 ;
	    RECT 425.2000 331.6000 426.0000 331.7000 ;
	    RECT 462.0000 331.6000 462.8000 331.7000 ;
	    RECT 473.2000 332.3000 474.0000 332.4000 ;
	    RECT 490.8000 332.3000 491.6000 332.4000 ;
	    RECT 473.2000 331.7000 491.6000 332.3000 ;
	    RECT 473.2000 331.6000 474.0000 331.7000 ;
	    RECT 490.8000 331.6000 491.6000 331.7000 ;
	    RECT 242.8000 329.7000 251.5000 330.3000 ;
	    RECT 286.1000 330.3000 286.7000 331.6000 ;
	    RECT 297.2000 330.3000 298.0000 330.4000 ;
	    RECT 286.1000 329.7000 298.0000 330.3000 ;
	    RECT 242.8000 329.6000 243.6000 329.7000 ;
	    RECT 297.2000 329.6000 298.0000 329.7000 ;
	    RECT 298.8000 330.3000 299.6000 330.4000 ;
	    RECT 382.0000 330.3000 382.8000 330.4000 ;
	    RECT 393.2000 330.3000 394.0000 330.4000 ;
	    RECT 298.8000 329.7000 369.9000 330.3000 ;
	    RECT 298.8000 329.6000 299.6000 329.7000 ;
	    RECT 369.3000 328.4000 369.9000 329.7000 ;
	    RECT 382.0000 329.7000 394.0000 330.3000 ;
	    RECT 382.0000 329.6000 382.8000 329.7000 ;
	    RECT 393.2000 329.6000 394.0000 329.7000 ;
	    RECT 396.4000 330.3000 397.2000 330.4000 ;
	    RECT 415.6000 330.3000 416.4000 330.4000 ;
	    RECT 396.4000 329.7000 416.4000 330.3000 ;
	    RECT 396.4000 329.6000 397.2000 329.7000 ;
	    RECT 415.6000 329.6000 416.4000 329.7000 ;
	    RECT 430.0000 330.3000 430.8000 330.4000 ;
	    RECT 438.0000 330.3000 438.8000 330.4000 ;
	    RECT 430.0000 329.7000 438.8000 330.3000 ;
	    RECT 430.0000 329.6000 430.8000 329.7000 ;
	    RECT 438.0000 329.6000 438.8000 329.7000 ;
	    RECT 458.8000 330.3000 459.6000 330.4000 ;
	    RECT 471.6000 330.3000 472.4000 330.4000 ;
	    RECT 458.8000 329.7000 472.4000 330.3000 ;
	    RECT 458.8000 329.6000 459.6000 329.7000 ;
	    RECT 471.6000 329.6000 472.4000 329.7000 ;
	    RECT 39.6000 328.3000 40.4000 328.4000 ;
	    RECT 65.2000 328.3000 66.0000 328.4000 ;
	    RECT 39.6000 327.7000 66.0000 328.3000 ;
	    RECT 39.6000 327.6000 40.4000 327.7000 ;
	    RECT 65.2000 327.6000 66.0000 327.7000 ;
	    RECT 119.6000 328.3000 120.4000 328.4000 ;
	    RECT 129.2000 328.3000 130.0000 328.4000 ;
	    RECT 119.6000 327.7000 130.0000 328.3000 ;
	    RECT 119.6000 327.6000 120.4000 327.7000 ;
	    RECT 129.2000 327.6000 130.0000 327.7000 ;
	    RECT 161.2000 328.3000 162.0000 328.4000 ;
	    RECT 180.4000 328.3000 181.2000 328.4000 ;
	    RECT 161.2000 327.7000 181.2000 328.3000 ;
	    RECT 161.2000 327.6000 162.0000 327.7000 ;
	    RECT 180.4000 327.6000 181.2000 327.7000 ;
	    RECT 202.8000 328.3000 203.6000 328.4000 ;
	    RECT 212.4000 328.3000 213.2000 328.4000 ;
	    RECT 202.8000 327.7000 213.2000 328.3000 ;
	    RECT 202.8000 327.6000 203.6000 327.7000 ;
	    RECT 212.4000 327.6000 213.2000 327.7000 ;
	    RECT 214.0000 328.3000 214.8000 328.4000 ;
	    RECT 220.4000 328.3000 221.2000 328.4000 ;
	    RECT 233.2000 328.3000 234.0000 328.4000 ;
	    RECT 214.0000 327.7000 234.0000 328.3000 ;
	    RECT 214.0000 327.6000 214.8000 327.7000 ;
	    RECT 220.4000 327.6000 221.2000 327.7000 ;
	    RECT 233.2000 327.6000 234.0000 327.7000 ;
	    RECT 262.0000 328.3000 262.8000 328.4000 ;
	    RECT 274.8000 328.3000 275.6000 328.4000 ;
	    RECT 262.0000 327.7000 275.6000 328.3000 ;
	    RECT 262.0000 327.6000 262.8000 327.7000 ;
	    RECT 274.8000 327.6000 275.6000 327.7000 ;
	    RECT 298.8000 328.3000 299.6000 328.4000 ;
	    RECT 308.4000 328.3000 309.2000 328.4000 ;
	    RECT 316.4000 328.3000 317.2000 328.4000 ;
	    RECT 334.0000 328.3000 334.8000 328.4000 ;
	    RECT 298.8000 327.7000 334.8000 328.3000 ;
	    RECT 298.8000 327.6000 299.6000 327.7000 ;
	    RECT 308.4000 327.6000 309.2000 327.7000 ;
	    RECT 316.4000 327.6000 317.2000 327.7000 ;
	    RECT 334.0000 327.6000 334.8000 327.7000 ;
	    RECT 343.6000 328.3000 344.4000 328.4000 ;
	    RECT 358.0000 328.3000 358.8000 328.4000 ;
	    RECT 343.6000 327.7000 358.8000 328.3000 ;
	    RECT 343.6000 327.6000 344.4000 327.7000 ;
	    RECT 358.0000 327.6000 358.8000 327.7000 ;
	    RECT 369.2000 328.3000 370.0000 328.4000 ;
	    RECT 388.4000 328.3000 389.2000 328.4000 ;
	    RECT 369.2000 327.7000 389.2000 328.3000 ;
	    RECT 369.2000 327.6000 370.0000 327.7000 ;
	    RECT 388.4000 327.6000 389.2000 327.7000 ;
	    RECT 398.0000 328.3000 398.8000 328.4000 ;
	    RECT 401.2000 328.3000 402.0000 328.4000 ;
	    RECT 414.0000 328.3000 414.8000 328.4000 ;
	    RECT 417.2000 328.3000 418.0000 328.4000 ;
	    RECT 426.8000 328.3000 427.6000 328.4000 ;
	    RECT 398.0000 327.7000 427.6000 328.3000 ;
	    RECT 398.0000 327.6000 398.8000 327.7000 ;
	    RECT 401.2000 327.6000 402.0000 327.7000 ;
	    RECT 414.0000 327.6000 414.8000 327.7000 ;
	    RECT 417.2000 327.6000 418.0000 327.7000 ;
	    RECT 426.8000 327.6000 427.6000 327.7000 ;
	    RECT 468.4000 328.3000 469.2000 328.4000 ;
	    RECT 508.4000 328.3000 509.2000 328.4000 ;
	    RECT 468.4000 327.7000 509.2000 328.3000 ;
	    RECT 468.4000 327.6000 469.2000 327.7000 ;
	    RECT 508.4000 327.6000 509.2000 327.7000 ;
	    RECT 36.4000 326.3000 37.2000 326.4000 ;
	    RECT 60.4000 326.3000 61.2000 326.4000 ;
	    RECT 86.0000 326.3000 86.8000 326.4000 ;
	    RECT 100.4000 326.3000 101.2000 326.4000 ;
	    RECT 36.4000 325.7000 101.2000 326.3000 ;
	    RECT 36.4000 325.6000 37.2000 325.7000 ;
	    RECT 60.4000 325.6000 61.2000 325.7000 ;
	    RECT 86.0000 325.6000 86.8000 325.7000 ;
	    RECT 100.4000 325.6000 101.2000 325.7000 ;
	    RECT 118.0000 326.3000 118.8000 326.4000 ;
	    RECT 338.8000 326.3000 339.6000 326.4000 ;
	    RECT 118.0000 325.7000 339.6000 326.3000 ;
	    RECT 118.0000 325.6000 118.8000 325.7000 ;
	    RECT 338.8000 325.6000 339.6000 325.7000 ;
	    RECT 396.4000 326.3000 397.2000 326.4000 ;
	    RECT 399.6000 326.3000 400.4000 326.4000 ;
	    RECT 412.4000 326.3000 413.2000 326.4000 ;
	    RECT 466.8000 326.3000 467.6000 326.4000 ;
	    RECT 498.8000 326.3000 499.6000 326.4000 ;
	    RECT 396.4000 325.7000 499.6000 326.3000 ;
	    RECT 396.4000 325.6000 397.2000 325.7000 ;
	    RECT 399.6000 325.6000 400.4000 325.7000 ;
	    RECT 412.4000 325.6000 413.2000 325.7000 ;
	    RECT 466.8000 325.6000 467.6000 325.7000 ;
	    RECT 498.8000 325.6000 499.6000 325.7000 ;
	    RECT 41.2000 324.3000 42.0000 324.4000 ;
	    RECT 58.8000 324.3000 59.6000 324.4000 ;
	    RECT 41.2000 323.7000 59.6000 324.3000 ;
	    RECT 41.2000 323.6000 42.0000 323.7000 ;
	    RECT 58.8000 323.6000 59.6000 323.7000 ;
	    RECT 71.6000 324.3000 72.4000 324.4000 ;
	    RECT 78.0000 324.3000 78.8000 324.4000 ;
	    RECT 71.6000 323.7000 78.8000 324.3000 ;
	    RECT 71.6000 323.6000 72.4000 323.7000 ;
	    RECT 78.0000 323.6000 78.8000 323.7000 ;
	    RECT 94.0000 324.3000 94.8000 324.4000 ;
	    RECT 116.4000 324.3000 117.2000 324.4000 ;
	    RECT 94.0000 323.7000 117.2000 324.3000 ;
	    RECT 94.0000 323.6000 94.8000 323.7000 ;
	    RECT 116.4000 323.6000 117.2000 323.7000 ;
	    RECT 185.2000 324.3000 186.0000 324.4000 ;
	    RECT 215.6000 324.3000 216.4000 324.4000 ;
	    RECT 218.8000 324.3000 219.6000 324.4000 ;
	    RECT 185.2000 323.7000 219.6000 324.3000 ;
	    RECT 185.2000 323.6000 186.0000 323.7000 ;
	    RECT 215.6000 323.6000 216.4000 323.7000 ;
	    RECT 218.8000 323.6000 219.6000 323.7000 ;
	    RECT 228.4000 324.3000 229.2000 324.4000 ;
	    RECT 244.4000 324.3000 245.2000 324.4000 ;
	    RECT 289.2000 324.3000 290.0000 324.4000 ;
	    RECT 228.4000 323.7000 243.5000 324.3000 ;
	    RECT 228.4000 323.6000 229.2000 323.7000 ;
	    RECT 153.2000 322.3000 154.0000 322.4000 ;
	    RECT 158.0000 322.3000 158.8000 322.4000 ;
	    RECT 194.8000 322.3000 195.6000 322.4000 ;
	    RECT 153.2000 321.7000 195.6000 322.3000 ;
	    RECT 153.2000 321.6000 154.0000 321.7000 ;
	    RECT 158.0000 321.6000 158.8000 321.7000 ;
	    RECT 194.8000 321.6000 195.6000 321.7000 ;
	    RECT 201.2000 322.3000 202.0000 322.4000 ;
	    RECT 210.8000 322.3000 211.6000 322.4000 ;
	    RECT 228.4000 322.3000 229.2000 322.4000 ;
	    RECT 241.2000 322.3000 242.0000 322.4000 ;
	    RECT 201.2000 321.7000 229.2000 322.3000 ;
	    RECT 201.2000 321.6000 202.0000 321.7000 ;
	    RECT 210.8000 321.6000 211.6000 321.7000 ;
	    RECT 228.4000 321.6000 229.2000 321.7000 ;
	    RECT 238.1000 321.7000 242.0000 322.3000 ;
	    RECT 242.9000 322.3000 243.5000 323.7000 ;
	    RECT 244.4000 323.7000 290.0000 324.3000 ;
	    RECT 244.4000 323.6000 245.2000 323.7000 ;
	    RECT 289.2000 323.6000 290.0000 323.7000 ;
	    RECT 302.0000 324.3000 302.8000 324.4000 ;
	    RECT 310.0000 324.3000 310.8000 324.4000 ;
	    RECT 479.6000 324.3000 480.4000 324.4000 ;
	    RECT 302.0000 323.7000 480.4000 324.3000 ;
	    RECT 302.0000 323.6000 302.8000 323.7000 ;
	    RECT 310.0000 323.6000 310.8000 323.7000 ;
	    RECT 479.6000 323.6000 480.4000 323.7000 ;
	    RECT 399.6000 322.3000 400.4000 322.4000 ;
	    RECT 242.9000 321.7000 400.4000 322.3000 ;
	    RECT 180.4000 320.3000 181.2000 320.4000 ;
	    RECT 215.6000 320.3000 216.4000 320.4000 ;
	    RECT 238.1000 320.3000 238.7000 321.7000 ;
	    RECT 241.2000 321.6000 242.0000 321.7000 ;
	    RECT 399.6000 321.6000 400.4000 321.7000 ;
	    RECT 431.6000 322.3000 432.4000 322.4000 ;
	    RECT 434.8000 322.3000 435.6000 322.4000 ;
	    RECT 466.8000 322.3000 467.6000 322.4000 ;
	    RECT 474.8000 322.3000 475.6000 322.4000 ;
	    RECT 431.6000 321.7000 475.6000 322.3000 ;
	    RECT 431.6000 321.6000 432.4000 321.7000 ;
	    RECT 434.8000 321.6000 435.6000 321.7000 ;
	    RECT 466.8000 321.6000 467.6000 321.7000 ;
	    RECT 474.8000 321.6000 475.6000 321.7000 ;
	    RECT 180.4000 319.7000 238.7000 320.3000 ;
	    RECT 252.4000 320.3000 253.2000 320.4000 ;
	    RECT 268.4000 320.3000 269.2000 320.4000 ;
	    RECT 252.4000 319.7000 269.2000 320.3000 ;
	    RECT 180.4000 319.6000 181.2000 319.7000 ;
	    RECT 215.6000 319.6000 216.4000 319.7000 ;
	    RECT 252.4000 319.6000 253.2000 319.7000 ;
	    RECT 268.4000 319.6000 269.2000 319.7000 ;
	    RECT 276.4000 320.3000 277.2000 320.4000 ;
	    RECT 399.6000 320.3000 400.4000 320.4000 ;
	    RECT 276.4000 319.7000 400.4000 320.3000 ;
	    RECT 276.4000 319.6000 277.2000 319.7000 ;
	    RECT 399.6000 319.6000 400.4000 319.7000 ;
	    RECT 71.6000 318.3000 72.4000 318.4000 ;
	    RECT 81.2000 318.3000 82.0000 318.4000 ;
	    RECT 71.6000 317.7000 82.0000 318.3000 ;
	    RECT 71.6000 317.6000 72.4000 317.7000 ;
	    RECT 81.2000 317.6000 82.0000 317.7000 ;
	    RECT 82.8000 318.3000 83.6000 318.4000 ;
	    RECT 122.8000 318.3000 123.6000 318.4000 ;
	    RECT 82.8000 317.7000 123.6000 318.3000 ;
	    RECT 82.8000 317.6000 83.6000 317.7000 ;
	    RECT 122.8000 317.6000 123.6000 317.7000 ;
	    RECT 191.6000 318.3000 192.4000 318.4000 ;
	    RECT 204.4000 318.3000 205.2000 318.4000 ;
	    RECT 220.4000 318.3000 221.2000 318.4000 ;
	    RECT 191.6000 317.7000 221.2000 318.3000 ;
	    RECT 191.6000 317.6000 192.4000 317.7000 ;
	    RECT 204.4000 317.6000 205.2000 317.7000 ;
	    RECT 220.4000 317.6000 221.2000 317.7000 ;
	    RECT 226.8000 318.3000 227.6000 318.4000 ;
	    RECT 292.4000 318.3000 293.2000 318.4000 ;
	    RECT 332.4000 318.3000 333.2000 318.4000 ;
	    RECT 226.8000 317.7000 333.2000 318.3000 ;
	    RECT 226.8000 317.6000 227.6000 317.7000 ;
	    RECT 292.4000 317.6000 293.2000 317.7000 ;
	    RECT 332.4000 317.6000 333.2000 317.7000 ;
	    RECT 38.0000 316.3000 38.8000 316.4000 ;
	    RECT 54.0000 316.3000 54.8000 316.4000 ;
	    RECT 38.0000 315.7000 54.8000 316.3000 ;
	    RECT 38.0000 315.6000 38.8000 315.7000 ;
	    RECT 54.0000 315.6000 54.8000 315.7000 ;
	    RECT 66.8000 316.3000 67.6000 316.4000 ;
	    RECT 130.8000 316.3000 131.6000 316.4000 ;
	    RECT 434.8000 316.3000 435.6000 316.4000 ;
	    RECT 66.8000 315.7000 83.5000 316.3000 ;
	    RECT 66.8000 315.6000 67.6000 315.7000 ;
	    RECT 9.2000 314.3000 10.0000 314.4000 ;
	    RECT 25.2000 314.3000 26.0000 314.4000 ;
	    RECT 44.4000 314.3000 45.2000 314.4000 ;
	    RECT 9.2000 313.7000 45.2000 314.3000 ;
	    RECT 9.2000 313.6000 10.0000 313.7000 ;
	    RECT 25.2000 313.6000 26.0000 313.7000 ;
	    RECT 44.4000 313.6000 45.2000 313.7000 ;
	    RECT 55.6000 314.3000 56.4000 314.4000 ;
	    RECT 81.2000 314.3000 82.0000 314.4000 ;
	    RECT 55.6000 313.7000 82.0000 314.3000 ;
	    RECT 82.9000 314.3000 83.5000 315.7000 ;
	    RECT 130.8000 315.7000 435.6000 316.3000 ;
	    RECT 130.8000 315.6000 131.6000 315.7000 ;
	    RECT 434.8000 315.6000 435.6000 315.7000 ;
	    RECT 172.4000 314.3000 173.2000 314.4000 ;
	    RECT 82.9000 313.7000 173.2000 314.3000 ;
	    RECT 55.6000 313.6000 56.4000 313.7000 ;
	    RECT 81.2000 313.6000 82.0000 313.7000 ;
	    RECT 172.4000 313.6000 173.2000 313.7000 ;
	    RECT 182.0000 314.3000 182.8000 314.4000 ;
	    RECT 223.6000 314.3000 224.4000 314.4000 ;
	    RECT 182.0000 313.7000 224.4000 314.3000 ;
	    RECT 182.0000 313.6000 182.8000 313.7000 ;
	    RECT 223.6000 313.6000 224.4000 313.7000 ;
	    RECT 233.2000 314.3000 234.0000 314.4000 ;
	    RECT 266.8000 314.3000 267.6000 314.4000 ;
	    RECT 233.2000 313.7000 267.6000 314.3000 ;
	    RECT 233.2000 313.6000 234.0000 313.7000 ;
	    RECT 266.8000 313.6000 267.6000 313.7000 ;
	    RECT 268.4000 314.3000 269.2000 314.4000 ;
	    RECT 279.6000 314.3000 280.4000 314.4000 ;
	    RECT 268.4000 313.7000 280.4000 314.3000 ;
	    RECT 268.4000 313.6000 269.2000 313.7000 ;
	    RECT 279.6000 313.6000 280.4000 313.7000 ;
	    RECT 282.8000 314.3000 283.6000 314.4000 ;
	    RECT 303.6000 314.3000 304.4000 314.4000 ;
	    RECT 322.8000 314.3000 323.6000 314.4000 ;
	    RECT 282.8000 313.7000 323.6000 314.3000 ;
	    RECT 282.8000 313.6000 283.6000 313.7000 ;
	    RECT 303.6000 313.6000 304.4000 313.7000 ;
	    RECT 322.8000 313.6000 323.6000 313.7000 ;
	    RECT 329.2000 314.3000 330.0000 314.4000 ;
	    RECT 340.4000 314.3000 341.2000 314.4000 ;
	    RECT 329.2000 313.7000 341.2000 314.3000 ;
	    RECT 329.2000 313.6000 330.0000 313.7000 ;
	    RECT 340.4000 313.6000 341.2000 313.7000 ;
	    RECT 343.6000 314.3000 344.4000 314.4000 ;
	    RECT 372.4000 314.3000 373.2000 314.4000 ;
	    RECT 374.0000 314.3000 374.8000 314.4000 ;
	    RECT 399.6000 314.3000 400.4000 314.4000 ;
	    RECT 415.6000 314.3000 416.4000 314.4000 ;
	    RECT 343.6000 313.7000 416.4000 314.3000 ;
	    RECT 343.6000 313.6000 344.4000 313.7000 ;
	    RECT 372.4000 313.6000 373.2000 313.7000 ;
	    RECT 374.0000 313.6000 374.8000 313.7000 ;
	    RECT 399.6000 313.6000 400.4000 313.7000 ;
	    RECT 415.6000 313.6000 416.4000 313.7000 ;
	    RECT 47.6000 312.3000 48.4000 312.4000 ;
	    RECT 50.8000 312.3000 51.6000 312.4000 ;
	    RECT 47.6000 311.7000 51.6000 312.3000 ;
	    RECT 47.6000 311.6000 48.4000 311.7000 ;
	    RECT 50.8000 311.6000 51.6000 311.7000 ;
	    RECT 63.6000 312.3000 64.4000 312.4000 ;
	    RECT 78.0000 312.3000 78.8000 312.4000 ;
	    RECT 63.6000 311.7000 78.8000 312.3000 ;
	    RECT 63.6000 311.6000 64.4000 311.7000 ;
	    RECT 78.0000 311.6000 78.8000 311.7000 ;
	    RECT 90.8000 312.3000 91.6000 312.4000 ;
	    RECT 114.8000 312.3000 115.6000 312.4000 ;
	    RECT 90.8000 311.7000 115.6000 312.3000 ;
	    RECT 90.8000 311.6000 91.6000 311.7000 ;
	    RECT 114.8000 311.6000 115.6000 311.7000 ;
	    RECT 116.4000 312.3000 117.2000 312.4000 ;
	    RECT 138.8000 312.3000 139.6000 312.4000 ;
	    RECT 116.4000 311.7000 139.6000 312.3000 ;
	    RECT 116.4000 311.6000 117.2000 311.7000 ;
	    RECT 138.8000 311.6000 139.6000 311.7000 ;
	    RECT 148.4000 312.3000 149.2000 312.4000 ;
	    RECT 198.0000 312.3000 198.8000 312.4000 ;
	    RECT 148.4000 311.7000 198.8000 312.3000 ;
	    RECT 148.4000 311.6000 149.2000 311.7000 ;
	    RECT 198.0000 311.6000 198.8000 311.7000 ;
	    RECT 199.6000 312.3000 200.4000 312.4000 ;
	    RECT 207.6000 312.3000 208.4000 312.4000 ;
	    RECT 199.6000 311.7000 208.4000 312.3000 ;
	    RECT 199.6000 311.6000 200.4000 311.7000 ;
	    RECT 207.6000 311.6000 208.4000 311.7000 ;
	    RECT 214.0000 312.3000 214.8000 312.4000 ;
	    RECT 234.8000 312.3000 235.6000 312.4000 ;
	    RECT 214.0000 311.7000 235.6000 312.3000 ;
	    RECT 214.0000 311.6000 214.8000 311.7000 ;
	    RECT 234.8000 311.6000 235.6000 311.7000 ;
	    RECT 236.4000 312.3000 237.2000 312.4000 ;
	    RECT 260.4000 312.3000 261.2000 312.4000 ;
	    RECT 236.4000 311.7000 261.2000 312.3000 ;
	    RECT 236.4000 311.6000 237.2000 311.7000 ;
	    RECT 260.4000 311.6000 261.2000 311.7000 ;
	    RECT 263.6000 312.3000 264.4000 312.4000 ;
	    RECT 292.4000 312.3000 293.2000 312.4000 ;
	    RECT 263.6000 311.7000 293.2000 312.3000 ;
	    RECT 263.6000 311.6000 264.4000 311.7000 ;
	    RECT 292.4000 311.6000 293.2000 311.7000 ;
	    RECT 295.6000 312.3000 296.4000 312.4000 ;
	    RECT 300.4000 312.3000 301.2000 312.4000 ;
	    RECT 295.6000 311.7000 301.2000 312.3000 ;
	    RECT 295.6000 311.6000 296.4000 311.7000 ;
	    RECT 300.4000 311.6000 301.2000 311.7000 ;
	    RECT 313.2000 312.3000 314.0000 312.4000 ;
	    RECT 407.6000 312.3000 408.4000 312.4000 ;
	    RECT 428.4000 312.3000 429.2000 312.4000 ;
	    RECT 313.2000 311.7000 429.2000 312.3000 ;
	    RECT 313.2000 311.6000 314.0000 311.7000 ;
	    RECT 407.6000 311.6000 408.4000 311.7000 ;
	    RECT 428.4000 311.6000 429.2000 311.7000 ;
	    RECT 470.0000 312.3000 470.8000 312.4000 ;
	    RECT 478.0000 312.3000 478.8000 312.4000 ;
	    RECT 470.0000 311.7000 478.8000 312.3000 ;
	    RECT 470.0000 311.6000 470.8000 311.7000 ;
	    RECT 478.0000 311.6000 478.8000 311.7000 ;
	    RECT 34.8000 310.3000 35.6000 310.4000 ;
	    RECT 47.6000 310.3000 48.4000 310.4000 ;
	    RECT 34.8000 309.7000 48.4000 310.3000 ;
	    RECT 34.8000 309.6000 35.6000 309.7000 ;
	    RECT 47.6000 309.6000 48.4000 309.7000 ;
	    RECT 54.0000 310.3000 54.8000 310.4000 ;
	    RECT 65.2000 310.3000 66.0000 310.4000 ;
	    RECT 54.0000 309.7000 66.0000 310.3000 ;
	    RECT 54.0000 309.6000 54.8000 309.7000 ;
	    RECT 65.2000 309.6000 66.0000 309.7000 ;
	    RECT 113.2000 310.3000 114.0000 310.4000 ;
	    RECT 118.0000 310.3000 118.8000 310.4000 ;
	    RECT 119.6000 310.3000 120.4000 310.4000 ;
	    RECT 113.2000 309.7000 120.4000 310.3000 ;
	    RECT 113.2000 309.6000 114.0000 309.7000 ;
	    RECT 118.0000 309.6000 118.8000 309.7000 ;
	    RECT 119.6000 309.6000 120.4000 309.7000 ;
	    RECT 126.0000 310.3000 126.8000 310.4000 ;
	    RECT 146.8000 310.3000 147.6000 310.4000 ;
	    RECT 126.0000 309.7000 147.6000 310.3000 ;
	    RECT 126.0000 309.6000 126.8000 309.7000 ;
	    RECT 146.8000 309.6000 147.6000 309.7000 ;
	    RECT 161.2000 310.3000 162.0000 310.4000 ;
	    RECT 170.8000 310.3000 171.6000 310.4000 ;
	    RECT 175.6000 310.3000 176.4000 310.4000 ;
	    RECT 161.2000 309.7000 176.4000 310.3000 ;
	    RECT 161.2000 309.6000 162.0000 309.7000 ;
	    RECT 170.8000 309.6000 171.6000 309.7000 ;
	    RECT 175.6000 309.6000 176.4000 309.7000 ;
	    RECT 194.8000 310.3000 195.6000 310.4000 ;
	    RECT 199.6000 310.3000 200.4000 310.4000 ;
	    RECT 194.8000 309.7000 200.4000 310.3000 ;
	    RECT 194.8000 309.6000 195.6000 309.7000 ;
	    RECT 199.6000 309.6000 200.4000 309.7000 ;
	    RECT 204.4000 310.3000 205.2000 310.4000 ;
	    RECT 206.0000 310.3000 206.8000 310.4000 ;
	    RECT 204.4000 309.7000 206.8000 310.3000 ;
	    RECT 204.4000 309.6000 205.2000 309.7000 ;
	    RECT 206.0000 309.6000 206.8000 309.7000 ;
	    RECT 223.6000 310.3000 224.4000 310.4000 ;
	    RECT 273.2000 310.3000 274.0000 310.4000 ;
	    RECT 223.6000 309.7000 274.0000 310.3000 ;
	    RECT 223.6000 309.6000 224.4000 309.7000 ;
	    RECT 273.2000 309.6000 274.0000 309.7000 ;
	    RECT 276.4000 310.3000 277.2000 310.4000 ;
	    RECT 290.8000 310.3000 291.6000 310.4000 ;
	    RECT 276.4000 309.7000 291.6000 310.3000 ;
	    RECT 276.4000 309.6000 277.2000 309.7000 ;
	    RECT 290.8000 309.6000 291.6000 309.7000 ;
	    RECT 298.8000 309.6000 299.6000 310.4000 ;
	    RECT 316.4000 310.3000 317.2000 310.4000 ;
	    RECT 326.0000 310.3000 326.8000 310.4000 ;
	    RECT 330.8000 310.3000 331.6000 310.4000 ;
	    RECT 337.2000 310.3000 338.0000 310.4000 ;
	    RECT 342.0000 310.3000 342.8000 310.4000 ;
	    RECT 316.4000 309.7000 325.1000 310.3000 ;
	    RECT 316.4000 309.6000 317.2000 309.7000 ;
	    RECT 116.4000 308.3000 117.2000 308.4000 ;
	    RECT 94.1000 307.7000 117.2000 308.3000 ;
	    RECT 74.8000 306.3000 75.6000 306.4000 ;
	    RECT 94.1000 306.3000 94.7000 307.7000 ;
	    RECT 116.4000 307.6000 117.2000 307.7000 ;
	    RECT 121.2000 308.3000 122.0000 308.4000 ;
	    RECT 129.2000 308.3000 130.0000 308.4000 ;
	    RECT 121.2000 307.7000 130.0000 308.3000 ;
	    RECT 121.2000 307.6000 122.0000 307.7000 ;
	    RECT 129.2000 307.6000 130.0000 307.7000 ;
	    RECT 148.4000 308.3000 149.2000 308.4000 ;
	    RECT 159.6000 308.3000 160.4000 308.4000 ;
	    RECT 148.4000 307.7000 160.4000 308.3000 ;
	    RECT 148.4000 307.6000 149.2000 307.7000 ;
	    RECT 159.6000 307.6000 160.4000 307.7000 ;
	    RECT 202.8000 308.3000 203.6000 308.4000 ;
	    RECT 204.4000 308.3000 205.2000 308.4000 ;
	    RECT 202.8000 307.7000 205.2000 308.3000 ;
	    RECT 202.8000 307.6000 203.6000 307.7000 ;
	    RECT 204.4000 307.6000 205.2000 307.7000 ;
	    RECT 209.2000 308.3000 210.0000 308.4000 ;
	    RECT 225.2000 308.3000 226.0000 308.4000 ;
	    RECT 209.2000 307.7000 226.0000 308.3000 ;
	    RECT 209.2000 307.6000 210.0000 307.7000 ;
	    RECT 225.2000 307.6000 226.0000 307.7000 ;
	    RECT 228.4000 308.3000 229.2000 308.4000 ;
	    RECT 244.4000 308.3000 245.2000 308.4000 ;
	    RECT 228.4000 307.7000 245.2000 308.3000 ;
	    RECT 228.4000 307.6000 229.2000 307.7000 ;
	    RECT 244.4000 307.6000 245.2000 307.7000 ;
	    RECT 247.6000 308.3000 248.4000 308.4000 ;
	    RECT 273.2000 308.3000 274.0000 308.4000 ;
	    RECT 247.6000 307.7000 274.0000 308.3000 ;
	    RECT 247.6000 307.6000 248.4000 307.7000 ;
	    RECT 273.2000 307.6000 274.0000 307.7000 ;
	    RECT 278.0000 308.3000 278.8000 308.4000 ;
	    RECT 282.8000 308.3000 283.6000 308.4000 ;
	    RECT 278.0000 307.7000 283.6000 308.3000 ;
	    RECT 278.0000 307.6000 278.8000 307.7000 ;
	    RECT 282.8000 307.6000 283.6000 307.7000 ;
	    RECT 292.4000 308.3000 293.2000 308.4000 ;
	    RECT 298.8000 308.3000 299.6000 308.4000 ;
	    RECT 313.2000 308.3000 314.0000 308.4000 ;
	    RECT 292.4000 307.7000 299.6000 308.3000 ;
	    RECT 292.4000 307.6000 293.2000 307.7000 ;
	    RECT 298.8000 307.6000 299.6000 307.7000 ;
	    RECT 300.5000 307.7000 314.0000 308.3000 ;
	    RECT 324.5000 308.3000 325.1000 309.7000 ;
	    RECT 326.0000 309.7000 342.8000 310.3000 ;
	    RECT 326.0000 309.6000 326.8000 309.7000 ;
	    RECT 330.8000 309.6000 331.6000 309.7000 ;
	    RECT 337.2000 309.6000 338.0000 309.7000 ;
	    RECT 342.0000 309.6000 342.8000 309.7000 ;
	    RECT 367.6000 310.3000 368.4000 310.4000 ;
	    RECT 372.4000 310.3000 373.2000 310.4000 ;
	    RECT 367.6000 309.7000 373.2000 310.3000 ;
	    RECT 367.6000 309.6000 368.4000 309.7000 ;
	    RECT 372.4000 309.6000 373.2000 309.7000 ;
	    RECT 388.4000 310.3000 389.2000 310.4000 ;
	    RECT 402.8000 310.3000 403.6000 310.4000 ;
	    RECT 388.4000 309.7000 403.6000 310.3000 ;
	    RECT 388.4000 309.6000 389.2000 309.7000 ;
	    RECT 402.8000 309.6000 403.6000 309.7000 ;
	    RECT 430.0000 310.3000 430.8000 310.4000 ;
	    RECT 446.0000 310.3000 446.8000 310.4000 ;
	    RECT 430.0000 309.7000 446.8000 310.3000 ;
	    RECT 430.0000 309.6000 430.8000 309.7000 ;
	    RECT 446.0000 309.6000 446.8000 309.7000 ;
	    RECT 471.6000 310.3000 472.4000 310.4000 ;
	    RECT 478.0000 310.3000 478.8000 310.4000 ;
	    RECT 471.6000 309.7000 478.8000 310.3000 ;
	    RECT 471.6000 309.6000 472.4000 309.7000 ;
	    RECT 478.0000 309.6000 478.8000 309.7000 ;
	    RECT 482.8000 310.3000 483.6000 310.4000 ;
	    RECT 495.6000 310.3000 496.4000 310.4000 ;
	    RECT 513.2000 310.3000 514.0000 310.4000 ;
	    RECT 482.8000 309.7000 514.0000 310.3000 ;
	    RECT 482.8000 309.6000 483.6000 309.7000 ;
	    RECT 495.6000 309.6000 496.4000 309.7000 ;
	    RECT 513.2000 309.6000 514.0000 309.7000 ;
	    RECT 327.6000 308.3000 328.4000 308.4000 ;
	    RECT 324.5000 307.7000 328.4000 308.3000 ;
	    RECT 74.8000 305.7000 94.7000 306.3000 ;
	    RECT 100.4000 306.3000 101.2000 306.4000 ;
	    RECT 132.4000 306.3000 133.2000 306.4000 ;
	    RECT 100.4000 305.7000 133.2000 306.3000 ;
	    RECT 74.8000 305.6000 75.6000 305.7000 ;
	    RECT 100.4000 305.6000 101.2000 305.7000 ;
	    RECT 132.4000 305.6000 133.2000 305.7000 ;
	    RECT 142.0000 306.3000 142.8000 306.4000 ;
	    RECT 169.2000 306.3000 170.0000 306.4000 ;
	    RECT 188.4000 306.3000 189.2000 306.4000 ;
	    RECT 142.0000 305.7000 189.2000 306.3000 ;
	    RECT 142.0000 305.6000 142.8000 305.7000 ;
	    RECT 169.2000 305.6000 170.0000 305.7000 ;
	    RECT 188.4000 305.6000 189.2000 305.7000 ;
	    RECT 190.0000 306.3000 190.8000 306.4000 ;
	    RECT 222.0000 306.3000 222.8000 306.4000 ;
	    RECT 263.6000 306.3000 264.4000 306.4000 ;
	    RECT 300.5000 306.3000 301.1000 307.7000 ;
	    RECT 313.2000 307.6000 314.0000 307.7000 ;
	    RECT 327.6000 307.6000 328.4000 307.7000 ;
	    RECT 332.4000 308.3000 333.2000 308.4000 ;
	    RECT 345.2000 308.3000 346.0000 308.4000 ;
	    RECT 332.4000 307.7000 346.0000 308.3000 ;
	    RECT 332.4000 307.6000 333.2000 307.7000 ;
	    RECT 345.2000 307.6000 346.0000 307.7000 ;
	    RECT 358.0000 308.3000 358.8000 308.4000 ;
	    RECT 367.6000 308.3000 368.4000 308.4000 ;
	    RECT 358.0000 307.7000 368.4000 308.3000 ;
	    RECT 358.0000 307.6000 358.8000 307.7000 ;
	    RECT 367.6000 307.6000 368.4000 307.7000 ;
	    RECT 452.4000 308.3000 453.2000 308.4000 ;
	    RECT 465.2000 308.3000 466.0000 308.4000 ;
	    RECT 452.4000 307.7000 466.0000 308.3000 ;
	    RECT 452.4000 307.6000 453.2000 307.7000 ;
	    RECT 465.2000 307.6000 466.0000 307.7000 ;
	    RECT 505.2000 308.3000 506.0000 308.4000 ;
	    RECT 506.8000 308.3000 507.6000 308.4000 ;
	    RECT 511.6000 308.3000 512.4000 308.4000 ;
	    RECT 505.2000 307.7000 512.4000 308.3000 ;
	    RECT 505.2000 307.6000 506.0000 307.7000 ;
	    RECT 506.8000 307.6000 507.6000 307.7000 ;
	    RECT 511.6000 307.6000 512.4000 307.7000 ;
	    RECT 190.0000 305.7000 222.8000 306.3000 ;
	    RECT 190.0000 305.6000 190.8000 305.7000 ;
	    RECT 222.0000 305.6000 222.8000 305.7000 ;
	    RECT 223.7000 305.7000 264.4000 306.3000 ;
	    RECT 70.0000 304.3000 70.8000 304.4000 ;
	    RECT 79.6000 304.3000 80.4000 304.4000 ;
	    RECT 70.0000 303.7000 80.4000 304.3000 ;
	    RECT 70.0000 303.6000 70.8000 303.7000 ;
	    RECT 79.6000 303.6000 80.4000 303.7000 ;
	    RECT 103.6000 304.3000 104.4000 304.4000 ;
	    RECT 137.2000 304.3000 138.0000 304.4000 ;
	    RECT 103.6000 303.7000 138.0000 304.3000 ;
	    RECT 103.6000 303.6000 104.4000 303.7000 ;
	    RECT 137.2000 303.6000 138.0000 303.7000 ;
	    RECT 138.8000 304.3000 139.6000 304.4000 ;
	    RECT 223.7000 304.3000 224.3000 305.7000 ;
	    RECT 263.6000 305.6000 264.4000 305.7000 ;
	    RECT 265.3000 305.7000 301.1000 306.3000 ;
	    RECT 306.8000 306.3000 307.6000 306.4000 ;
	    RECT 314.8000 306.3000 315.6000 306.4000 ;
	    RECT 306.8000 305.7000 315.6000 306.3000 ;
	    RECT 138.8000 303.7000 224.3000 304.3000 ;
	    RECT 225.2000 304.3000 226.0000 304.4000 ;
	    RECT 249.2000 304.3000 250.0000 304.4000 ;
	    RECT 225.2000 303.7000 250.0000 304.3000 ;
	    RECT 138.8000 303.6000 139.6000 303.7000 ;
	    RECT 225.2000 303.6000 226.0000 303.7000 ;
	    RECT 249.2000 303.6000 250.0000 303.7000 ;
	    RECT 263.6000 304.3000 264.4000 304.4000 ;
	    RECT 265.3000 304.3000 265.9000 305.7000 ;
	    RECT 306.8000 305.6000 307.6000 305.7000 ;
	    RECT 314.8000 305.6000 315.6000 305.7000 ;
	    RECT 457.2000 306.3000 458.0000 306.4000 ;
	    RECT 462.0000 306.3000 462.8000 306.4000 ;
	    RECT 457.2000 305.7000 462.8000 306.3000 ;
	    RECT 457.2000 305.6000 458.0000 305.7000 ;
	    RECT 462.0000 305.6000 462.8000 305.7000 ;
	    RECT 263.6000 303.7000 265.9000 304.3000 ;
	    RECT 268.4000 304.3000 269.2000 304.4000 ;
	    RECT 327.6000 304.3000 328.4000 304.4000 ;
	    RECT 268.4000 303.7000 328.4000 304.3000 ;
	    RECT 263.6000 303.6000 264.4000 303.7000 ;
	    RECT 268.4000 303.6000 269.2000 303.7000 ;
	    RECT 327.6000 303.6000 328.4000 303.7000 ;
	    RECT 332.4000 304.3000 333.2000 304.4000 ;
	    RECT 342.0000 304.3000 342.8000 304.4000 ;
	    RECT 345.2000 304.3000 346.0000 304.4000 ;
	    RECT 364.4000 304.3000 365.2000 304.4000 ;
	    RECT 332.4000 303.7000 365.2000 304.3000 ;
	    RECT 332.4000 303.6000 333.2000 303.7000 ;
	    RECT 342.0000 303.6000 342.8000 303.7000 ;
	    RECT 345.2000 303.6000 346.0000 303.7000 ;
	    RECT 364.4000 303.6000 365.2000 303.7000 ;
	    RECT 458.8000 304.3000 459.6000 304.4000 ;
	    RECT 486.0000 304.3000 486.8000 304.4000 ;
	    RECT 458.8000 303.7000 486.8000 304.3000 ;
	    RECT 458.8000 303.6000 459.6000 303.7000 ;
	    RECT 486.0000 303.6000 486.8000 303.7000 ;
	    RECT 60.4000 302.3000 61.2000 302.4000 ;
	    RECT 242.8000 302.3000 243.6000 302.4000 ;
	    RECT 60.4000 301.7000 243.6000 302.3000 ;
	    RECT 60.4000 301.6000 61.2000 301.7000 ;
	    RECT 242.8000 301.6000 243.6000 301.7000 ;
	    RECT 244.4000 302.3000 245.2000 302.4000 ;
	    RECT 252.4000 302.3000 253.2000 302.4000 ;
	    RECT 244.4000 301.7000 253.2000 302.3000 ;
	    RECT 244.4000 301.6000 245.2000 301.7000 ;
	    RECT 252.4000 301.6000 253.2000 301.7000 ;
	    RECT 271.6000 302.3000 272.4000 302.4000 ;
	    RECT 289.2000 302.3000 290.0000 302.4000 ;
	    RECT 334.0000 302.3000 334.8000 302.4000 ;
	    RECT 271.6000 301.7000 334.8000 302.3000 ;
	    RECT 271.6000 301.6000 272.4000 301.7000 ;
	    RECT 289.2000 301.6000 290.0000 301.7000 ;
	    RECT 334.0000 301.6000 334.8000 301.7000 ;
	    RECT 337.2000 302.3000 338.0000 302.4000 ;
	    RECT 346.8000 302.3000 347.6000 302.4000 ;
	    RECT 458.9000 302.3000 459.5000 303.6000 ;
	    RECT 337.2000 301.7000 459.5000 302.3000 ;
	    RECT 337.2000 301.6000 338.0000 301.7000 ;
	    RECT 346.8000 301.6000 347.6000 301.7000 ;
	    RECT 1.2000 300.3000 2.0000 300.4000 ;
	    RECT 4.4000 300.3000 5.2000 300.4000 ;
	    RECT 1.2000 299.7000 5.2000 300.3000 ;
	    RECT 1.2000 299.6000 2.0000 299.7000 ;
	    RECT 4.4000 299.6000 5.2000 299.7000 ;
	    RECT 84.4000 300.3000 85.2000 300.4000 ;
	    RECT 118.0000 300.3000 118.8000 300.4000 ;
	    RECT 150.0000 300.3000 150.8000 300.4000 ;
	    RECT 170.8000 300.3000 171.6000 300.4000 ;
	    RECT 84.4000 299.7000 117.1000 300.3000 ;
	    RECT 84.4000 299.6000 85.2000 299.7000 ;
	    RECT 26.8000 298.3000 27.6000 298.4000 ;
	    RECT 39.6000 298.3000 40.4000 298.4000 ;
	    RECT 26.8000 297.7000 40.4000 298.3000 ;
	    RECT 116.5000 298.3000 117.1000 299.7000 ;
	    RECT 118.0000 299.7000 171.6000 300.3000 ;
	    RECT 118.0000 299.6000 118.8000 299.7000 ;
	    RECT 150.0000 299.6000 150.8000 299.7000 ;
	    RECT 170.8000 299.6000 171.6000 299.7000 ;
	    RECT 172.4000 300.3000 173.2000 300.4000 ;
	    RECT 247.6000 300.3000 248.4000 300.4000 ;
	    RECT 172.4000 299.7000 248.4000 300.3000 ;
	    RECT 172.4000 299.6000 173.2000 299.7000 ;
	    RECT 247.6000 299.6000 248.4000 299.7000 ;
	    RECT 270.0000 300.3000 270.8000 300.4000 ;
	    RECT 302.0000 300.3000 302.8000 300.4000 ;
	    RECT 350.0000 300.3000 350.8000 300.4000 ;
	    RECT 369.2000 300.3000 370.0000 300.4000 ;
	    RECT 270.0000 299.7000 370.0000 300.3000 ;
	    RECT 270.0000 299.6000 270.8000 299.7000 ;
	    RECT 302.0000 299.6000 302.8000 299.7000 ;
	    RECT 350.0000 299.6000 350.8000 299.7000 ;
	    RECT 369.2000 299.6000 370.0000 299.7000 ;
	    RECT 417.2000 300.3000 418.0000 300.4000 ;
	    RECT 458.8000 300.3000 459.6000 300.4000 ;
	    RECT 417.2000 299.7000 459.6000 300.3000 ;
	    RECT 417.2000 299.6000 418.0000 299.7000 ;
	    RECT 458.8000 299.6000 459.6000 299.7000 ;
	    RECT 119.6000 298.3000 120.4000 298.4000 ;
	    RECT 116.5000 297.7000 120.4000 298.3000 ;
	    RECT 26.8000 297.6000 27.6000 297.7000 ;
	    RECT 39.6000 297.6000 40.4000 297.7000 ;
	    RECT 119.6000 297.6000 120.4000 297.7000 ;
	    RECT 122.8000 298.3000 123.6000 298.4000 ;
	    RECT 138.8000 298.3000 139.6000 298.4000 ;
	    RECT 122.8000 297.7000 139.6000 298.3000 ;
	    RECT 122.8000 297.6000 123.6000 297.7000 ;
	    RECT 138.8000 297.6000 139.6000 297.7000 ;
	    RECT 140.4000 298.3000 141.2000 298.4000 ;
	    RECT 146.8000 298.3000 147.6000 298.4000 ;
	    RECT 140.4000 297.7000 147.6000 298.3000 ;
	    RECT 140.4000 297.6000 141.2000 297.7000 ;
	    RECT 146.8000 297.6000 147.6000 297.7000 ;
	    RECT 151.6000 298.3000 152.4000 298.4000 ;
	    RECT 158.0000 298.3000 158.8000 298.4000 ;
	    RECT 151.6000 297.7000 158.8000 298.3000 ;
	    RECT 151.6000 297.6000 152.4000 297.7000 ;
	    RECT 158.0000 297.6000 158.8000 297.7000 ;
	    RECT 162.8000 298.3000 163.6000 298.4000 ;
	    RECT 169.2000 298.3000 170.0000 298.4000 ;
	    RECT 162.8000 297.7000 170.0000 298.3000 ;
	    RECT 162.8000 297.6000 163.6000 297.7000 ;
	    RECT 169.2000 297.6000 170.0000 297.7000 ;
	    RECT 170.8000 298.3000 171.6000 298.4000 ;
	    RECT 198.0000 298.3000 198.8000 298.4000 ;
	    RECT 206.0000 298.3000 206.8000 298.4000 ;
	    RECT 170.8000 297.7000 198.8000 298.3000 ;
	    RECT 170.8000 297.6000 171.6000 297.7000 ;
	    RECT 198.0000 297.6000 198.8000 297.7000 ;
	    RECT 199.7000 297.7000 206.8000 298.3000 ;
	    RECT 58.8000 296.3000 59.6000 296.4000 ;
	    RECT 62.0000 296.3000 62.8000 296.4000 ;
	    RECT 70.0000 296.3000 70.8000 296.4000 ;
	    RECT 58.8000 295.7000 70.8000 296.3000 ;
	    RECT 58.8000 295.6000 59.6000 295.7000 ;
	    RECT 62.0000 295.6000 62.8000 295.7000 ;
	    RECT 70.0000 295.6000 70.8000 295.7000 ;
	    RECT 71.6000 296.3000 72.4000 296.4000 ;
	    RECT 94.0000 296.3000 94.8000 296.4000 ;
	    RECT 124.4000 296.3000 125.2000 296.4000 ;
	    RECT 135.6000 296.3000 136.4000 296.4000 ;
	    RECT 153.2000 296.3000 154.0000 296.4000 ;
	    RECT 177.2000 296.3000 178.0000 296.4000 ;
	    RECT 71.6000 295.7000 89.9000 296.3000 ;
	    RECT 71.6000 295.6000 72.4000 295.7000 ;
	    RECT 62.0000 294.3000 62.8000 294.4000 ;
	    RECT 68.4000 294.3000 69.2000 294.4000 ;
	    RECT 73.2000 294.3000 74.0000 294.4000 ;
	    RECT 62.0000 293.7000 74.0000 294.3000 ;
	    RECT 62.0000 293.6000 62.8000 293.7000 ;
	    RECT 68.4000 293.6000 69.2000 293.7000 ;
	    RECT 73.2000 293.6000 74.0000 293.7000 ;
	    RECT 74.8000 294.3000 75.6000 294.4000 ;
	    RECT 86.0000 294.3000 86.8000 294.4000 ;
	    RECT 87.6000 294.3000 88.4000 294.4000 ;
	    RECT 74.8000 293.7000 88.4000 294.3000 ;
	    RECT 89.3000 294.3000 89.9000 295.7000 ;
	    RECT 94.0000 295.7000 105.9000 296.3000 ;
	    RECT 94.0000 295.6000 94.8000 295.7000 ;
	    RECT 95.6000 294.3000 96.4000 294.4000 ;
	    RECT 89.3000 293.7000 96.4000 294.3000 ;
	    RECT 74.8000 293.6000 75.6000 293.7000 ;
	    RECT 86.0000 293.6000 86.8000 293.7000 ;
	    RECT 87.6000 293.6000 88.4000 293.7000 ;
	    RECT 95.6000 293.6000 96.4000 293.7000 ;
	    RECT 97.2000 294.3000 98.0000 294.4000 ;
	    RECT 103.6000 294.3000 104.4000 294.4000 ;
	    RECT 97.2000 293.7000 104.4000 294.3000 ;
	    RECT 105.3000 294.3000 105.9000 295.7000 ;
	    RECT 124.4000 295.7000 178.0000 296.3000 ;
	    RECT 124.4000 295.6000 125.2000 295.7000 ;
	    RECT 135.6000 295.6000 136.4000 295.7000 ;
	    RECT 153.2000 295.6000 154.0000 295.7000 ;
	    RECT 177.2000 295.6000 178.0000 295.7000 ;
	    RECT 194.8000 296.3000 195.6000 296.4000 ;
	    RECT 199.7000 296.3000 200.3000 297.7000 ;
	    RECT 206.0000 297.6000 206.8000 297.7000 ;
	    RECT 207.6000 298.3000 208.4000 298.4000 ;
	    RECT 217.2000 298.3000 218.0000 298.4000 ;
	    RECT 225.2000 298.3000 226.0000 298.4000 ;
	    RECT 207.6000 297.7000 213.1000 298.3000 ;
	    RECT 207.6000 297.6000 208.4000 297.7000 ;
	    RECT 194.8000 295.7000 200.3000 296.3000 ;
	    RECT 201.2000 296.3000 202.0000 296.4000 ;
	    RECT 210.8000 296.3000 211.6000 296.4000 ;
	    RECT 201.2000 295.7000 211.6000 296.3000 ;
	    RECT 212.5000 296.3000 213.1000 297.7000 ;
	    RECT 217.2000 297.7000 226.0000 298.3000 ;
	    RECT 217.2000 297.6000 218.0000 297.7000 ;
	    RECT 225.2000 297.6000 226.0000 297.7000 ;
	    RECT 228.4000 298.3000 229.2000 298.4000 ;
	    RECT 250.8000 298.3000 251.6000 298.4000 ;
	    RECT 375.6000 298.3000 376.4000 298.4000 ;
	    RECT 417.2000 298.3000 418.0000 298.4000 ;
	    RECT 228.4000 297.7000 418.0000 298.3000 ;
	    RECT 228.4000 297.6000 229.2000 297.7000 ;
	    RECT 250.8000 297.6000 251.6000 297.7000 ;
	    RECT 375.6000 297.6000 376.4000 297.7000 ;
	    RECT 417.2000 297.6000 418.0000 297.7000 ;
	    RECT 430.0000 298.3000 430.8000 298.4000 ;
	    RECT 462.0000 298.3000 462.8000 298.4000 ;
	    RECT 471.6000 298.3000 472.4000 298.4000 ;
	    RECT 430.0000 297.7000 472.4000 298.3000 ;
	    RECT 430.0000 297.6000 430.8000 297.7000 ;
	    RECT 462.0000 297.6000 462.8000 297.7000 ;
	    RECT 471.6000 297.6000 472.4000 297.7000 ;
	    RECT 484.4000 298.3000 485.2000 298.4000 ;
	    RECT 489.2000 298.3000 490.0000 298.4000 ;
	    RECT 484.4000 297.7000 490.0000 298.3000 ;
	    RECT 484.4000 297.6000 485.2000 297.7000 ;
	    RECT 489.2000 297.6000 490.0000 297.7000 ;
	    RECT 263.6000 296.3000 264.4000 296.4000 ;
	    RECT 212.5000 295.7000 264.4000 296.3000 ;
	    RECT 194.8000 295.6000 195.6000 295.7000 ;
	    RECT 201.2000 295.6000 202.0000 295.7000 ;
	    RECT 210.8000 295.6000 211.6000 295.7000 ;
	    RECT 263.6000 295.6000 264.4000 295.7000 ;
	    RECT 266.8000 296.3000 267.6000 296.4000 ;
	    RECT 270.0000 296.3000 270.8000 296.4000 ;
	    RECT 266.8000 295.7000 270.8000 296.3000 ;
	    RECT 266.8000 295.6000 267.6000 295.7000 ;
	    RECT 270.0000 295.6000 270.8000 295.7000 ;
	    RECT 271.6000 296.3000 272.4000 296.4000 ;
	    RECT 282.8000 296.3000 283.6000 296.4000 ;
	    RECT 271.6000 295.7000 283.6000 296.3000 ;
	    RECT 271.6000 295.6000 272.4000 295.7000 ;
	    RECT 282.8000 295.6000 283.6000 295.7000 ;
	    RECT 290.8000 296.3000 291.6000 296.4000 ;
	    RECT 308.4000 296.3000 309.2000 296.4000 ;
	    RECT 290.8000 295.7000 309.2000 296.3000 ;
	    RECT 290.8000 295.6000 291.6000 295.7000 ;
	    RECT 308.4000 295.6000 309.2000 295.7000 ;
	    RECT 321.2000 296.3000 322.0000 296.4000 ;
	    RECT 329.2000 296.3000 330.0000 296.4000 ;
	    RECT 321.2000 295.7000 330.0000 296.3000 ;
	    RECT 321.2000 295.6000 322.0000 295.7000 ;
	    RECT 329.2000 295.6000 330.0000 295.7000 ;
	    RECT 362.8000 296.3000 363.6000 296.4000 ;
	    RECT 366.0000 296.3000 366.8000 296.4000 ;
	    RECT 378.8000 296.3000 379.6000 296.4000 ;
	    RECT 434.8000 296.3000 435.6000 296.4000 ;
	    RECT 362.8000 295.7000 379.6000 296.3000 ;
	    RECT 362.8000 295.6000 363.6000 295.7000 ;
	    RECT 366.0000 295.6000 366.8000 295.7000 ;
	    RECT 378.8000 295.6000 379.6000 295.7000 ;
	    RECT 414.1000 295.7000 435.6000 296.3000 ;
	    RECT 126.0000 294.3000 126.8000 294.4000 ;
	    RECT 105.3000 293.7000 126.8000 294.3000 ;
	    RECT 97.2000 293.6000 98.0000 293.7000 ;
	    RECT 103.6000 293.6000 104.4000 293.7000 ;
	    RECT 126.0000 293.6000 126.8000 293.7000 ;
	    RECT 134.0000 294.3000 134.8000 294.4000 ;
	    RECT 162.8000 294.3000 163.6000 294.4000 ;
	    RECT 134.0000 293.7000 163.6000 294.3000 ;
	    RECT 134.0000 293.6000 134.8000 293.7000 ;
	    RECT 162.8000 293.6000 163.6000 293.7000 ;
	    RECT 164.4000 293.6000 165.2000 294.4000 ;
	    RECT 169.2000 294.3000 170.0000 294.4000 ;
	    RECT 175.6000 294.3000 176.4000 294.4000 ;
	    RECT 186.8000 294.3000 187.6000 294.4000 ;
	    RECT 169.2000 293.7000 187.6000 294.3000 ;
	    RECT 169.2000 293.6000 170.0000 293.7000 ;
	    RECT 175.6000 293.6000 176.4000 293.7000 ;
	    RECT 186.8000 293.6000 187.6000 293.7000 ;
	    RECT 198.0000 294.3000 198.8000 294.4000 ;
	    RECT 202.8000 294.3000 203.6000 294.4000 ;
	    RECT 198.0000 293.7000 203.6000 294.3000 ;
	    RECT 198.0000 293.6000 198.8000 293.7000 ;
	    RECT 202.8000 293.6000 203.6000 293.7000 ;
	    RECT 204.4000 294.3000 205.2000 294.4000 ;
	    RECT 209.2000 294.3000 210.0000 294.4000 ;
	    RECT 204.4000 293.7000 210.0000 294.3000 ;
	    RECT 204.4000 293.6000 205.2000 293.7000 ;
	    RECT 209.2000 293.6000 210.0000 293.7000 ;
	    RECT 210.8000 294.3000 211.6000 294.4000 ;
	    RECT 215.6000 294.3000 216.4000 294.4000 ;
	    RECT 210.8000 293.7000 216.4000 294.3000 ;
	    RECT 210.8000 293.6000 211.6000 293.7000 ;
	    RECT 215.6000 293.6000 216.4000 293.7000 ;
	    RECT 222.0000 294.3000 222.8000 294.4000 ;
	    RECT 223.6000 294.3000 224.4000 294.4000 ;
	    RECT 222.0000 293.7000 224.4000 294.3000 ;
	    RECT 222.0000 293.6000 222.8000 293.7000 ;
	    RECT 223.6000 293.6000 224.4000 293.7000 ;
	    RECT 225.2000 294.3000 226.0000 294.4000 ;
	    RECT 233.2000 294.3000 234.0000 294.4000 ;
	    RECT 225.2000 293.7000 234.0000 294.3000 ;
	    RECT 225.2000 293.6000 226.0000 293.7000 ;
	    RECT 233.2000 293.6000 234.0000 293.7000 ;
	    RECT 238.0000 294.3000 238.8000 294.4000 ;
	    RECT 244.4000 294.3000 245.2000 294.4000 ;
	    RECT 238.0000 293.7000 245.2000 294.3000 ;
	    RECT 238.0000 293.6000 238.8000 293.7000 ;
	    RECT 244.4000 293.6000 245.2000 293.7000 ;
	    RECT 246.0000 294.3000 246.8000 294.4000 ;
	    RECT 260.4000 294.3000 261.2000 294.4000 ;
	    RECT 265.2000 294.3000 266.0000 294.4000 ;
	    RECT 297.2000 294.3000 298.0000 294.4000 ;
	    RECT 324.4000 294.3000 325.2000 294.4000 ;
	    RECT 246.0000 293.7000 325.2000 294.3000 ;
	    RECT 246.0000 293.6000 246.8000 293.7000 ;
	    RECT 260.4000 293.6000 261.2000 293.7000 ;
	    RECT 265.2000 293.6000 266.0000 293.7000 ;
	    RECT 297.2000 293.6000 298.0000 293.7000 ;
	    RECT 324.4000 293.6000 325.2000 293.7000 ;
	    RECT 329.2000 294.3000 330.0000 294.4000 ;
	    RECT 414.1000 294.3000 414.7000 295.7000 ;
	    RECT 434.8000 295.6000 435.6000 295.7000 ;
	    RECT 487.6000 295.6000 488.4000 296.4000 ;
	    RECT 490.8000 296.3000 491.6000 296.4000 ;
	    RECT 500.4000 296.3000 501.2000 296.4000 ;
	    RECT 490.8000 295.7000 501.2000 296.3000 ;
	    RECT 490.8000 295.6000 491.6000 295.7000 ;
	    RECT 500.4000 295.6000 501.2000 295.7000 ;
	    RECT 329.2000 293.7000 414.7000 294.3000 ;
	    RECT 415.6000 294.3000 416.4000 294.4000 ;
	    RECT 425.2000 294.3000 426.0000 294.4000 ;
	    RECT 455.6000 294.3000 456.4000 294.4000 ;
	    RECT 415.6000 293.7000 456.4000 294.3000 ;
	    RECT 329.2000 293.6000 330.0000 293.7000 ;
	    RECT 415.6000 293.6000 416.4000 293.7000 ;
	    RECT 425.2000 293.6000 426.0000 293.7000 ;
	    RECT 455.6000 293.6000 456.4000 293.7000 ;
	    RECT 470.0000 294.3000 470.8000 294.4000 ;
	    RECT 482.8000 294.3000 483.6000 294.4000 ;
	    RECT 470.0000 293.7000 483.6000 294.3000 ;
	    RECT 470.0000 293.6000 470.8000 293.7000 ;
	    RECT 482.8000 293.6000 483.6000 293.7000 ;
	    RECT 487.6000 294.3000 488.4000 294.4000 ;
	    RECT 492.4000 294.3000 493.2000 294.4000 ;
	    RECT 487.6000 293.7000 493.2000 294.3000 ;
	    RECT 487.6000 293.6000 488.4000 293.7000 ;
	    RECT 492.4000 293.6000 493.2000 293.7000 ;
	    RECT 12.4000 292.3000 13.2000 292.4000 ;
	    RECT 26.8000 292.3000 27.6000 292.4000 ;
	    RECT 46.0000 292.3000 46.8000 292.4000 ;
	    RECT 12.4000 291.7000 46.8000 292.3000 ;
	    RECT 12.4000 291.6000 13.2000 291.7000 ;
	    RECT 26.8000 291.6000 27.6000 291.7000 ;
	    RECT 46.0000 291.6000 46.8000 291.7000 ;
	    RECT 78.0000 292.3000 78.8000 292.4000 ;
	    RECT 82.8000 292.3000 83.6000 292.4000 ;
	    RECT 84.4000 292.3000 85.2000 292.4000 ;
	    RECT 78.0000 291.7000 85.2000 292.3000 ;
	    RECT 78.0000 291.6000 78.8000 291.7000 ;
	    RECT 82.8000 291.6000 83.6000 291.7000 ;
	    RECT 84.4000 291.6000 85.2000 291.7000 ;
	    RECT 90.8000 292.3000 91.6000 292.4000 ;
	    RECT 98.8000 292.3000 99.6000 292.4000 ;
	    RECT 90.8000 291.7000 99.6000 292.3000 ;
	    RECT 90.8000 291.6000 91.6000 291.7000 ;
	    RECT 98.8000 291.6000 99.6000 291.7000 ;
	    RECT 102.0000 292.3000 102.8000 292.4000 ;
	    RECT 116.4000 292.3000 117.2000 292.4000 ;
	    RECT 122.8000 292.3000 123.6000 292.4000 ;
	    RECT 102.0000 291.7000 123.6000 292.3000 ;
	    RECT 102.0000 291.6000 102.8000 291.7000 ;
	    RECT 116.4000 291.6000 117.2000 291.7000 ;
	    RECT 122.8000 291.6000 123.6000 291.7000 ;
	    RECT 126.0000 292.3000 126.8000 292.4000 ;
	    RECT 132.4000 292.3000 133.2000 292.4000 ;
	    RECT 143.6000 292.3000 144.4000 292.4000 ;
	    RECT 126.0000 291.7000 144.4000 292.3000 ;
	    RECT 126.0000 291.6000 126.8000 291.7000 ;
	    RECT 132.4000 291.6000 133.2000 291.7000 ;
	    RECT 143.6000 291.6000 144.4000 291.7000 ;
	    RECT 151.6000 292.3000 152.4000 292.4000 ;
	    RECT 154.8000 292.3000 155.6000 292.4000 ;
	    RECT 151.6000 291.7000 155.6000 292.3000 ;
	    RECT 151.6000 291.6000 152.4000 291.7000 ;
	    RECT 154.8000 291.6000 155.6000 291.7000 ;
	    RECT 164.4000 292.3000 165.2000 292.4000 ;
	    RECT 222.0000 292.3000 222.8000 292.4000 ;
	    RECT 164.4000 291.7000 222.8000 292.3000 ;
	    RECT 164.4000 291.6000 165.2000 291.7000 ;
	    RECT 222.0000 291.6000 222.8000 291.7000 ;
	    RECT 231.6000 292.3000 232.4000 292.4000 ;
	    RECT 244.4000 292.3000 245.2000 292.4000 ;
	    RECT 279.6000 292.3000 280.4000 292.4000 ;
	    RECT 303.6000 292.3000 304.4000 292.4000 ;
	    RECT 322.8000 292.3000 323.6000 292.4000 ;
	    RECT 340.4000 292.3000 341.2000 292.4000 ;
	    RECT 231.6000 291.7000 341.2000 292.3000 ;
	    RECT 231.6000 291.6000 232.4000 291.7000 ;
	    RECT 244.4000 291.6000 245.2000 291.7000 ;
	    RECT 279.6000 291.6000 280.4000 291.7000 ;
	    RECT 303.6000 291.6000 304.4000 291.7000 ;
	    RECT 322.8000 291.6000 323.6000 291.7000 ;
	    RECT 340.4000 291.6000 341.2000 291.7000 ;
	    RECT 361.2000 292.3000 362.0000 292.4000 ;
	    RECT 375.6000 292.3000 376.4000 292.4000 ;
	    RECT 361.2000 291.7000 376.4000 292.3000 ;
	    RECT 361.2000 291.6000 362.0000 291.7000 ;
	    RECT 375.6000 291.6000 376.4000 291.7000 ;
	    RECT 434.8000 292.3000 435.6000 292.4000 ;
	    RECT 444.4000 292.3000 445.2000 292.4000 ;
	    RECT 434.8000 291.7000 445.2000 292.3000 ;
	    RECT 434.8000 291.6000 435.6000 291.7000 ;
	    RECT 444.4000 291.6000 445.2000 291.7000 ;
	    RECT 457.2000 292.3000 458.0000 292.4000 ;
	    RECT 492.4000 292.3000 493.2000 292.4000 ;
	    RECT 457.2000 291.7000 493.2000 292.3000 ;
	    RECT 457.2000 291.6000 458.0000 291.7000 ;
	    RECT 492.4000 291.6000 493.2000 291.7000 ;
	    RECT 86.0000 290.3000 86.8000 290.4000 ;
	    RECT 97.2000 290.3000 98.0000 290.4000 ;
	    RECT 100.4000 290.3000 101.2000 290.4000 ;
	    RECT 86.0000 289.7000 101.2000 290.3000 ;
	    RECT 86.0000 289.6000 86.8000 289.7000 ;
	    RECT 97.2000 289.6000 98.0000 289.7000 ;
	    RECT 100.4000 289.6000 101.2000 289.7000 ;
	    RECT 150.0000 290.3000 150.8000 290.4000 ;
	    RECT 161.2000 290.3000 162.0000 290.4000 ;
	    RECT 150.0000 289.7000 162.0000 290.3000 ;
	    RECT 150.0000 289.6000 150.8000 289.7000 ;
	    RECT 161.2000 289.6000 162.0000 289.7000 ;
	    RECT 162.8000 290.3000 163.6000 290.4000 ;
	    RECT 164.4000 290.3000 165.2000 290.4000 ;
	    RECT 162.8000 289.7000 165.2000 290.3000 ;
	    RECT 162.8000 289.6000 163.6000 289.7000 ;
	    RECT 164.4000 289.6000 165.2000 289.7000 ;
	    RECT 166.0000 290.3000 166.8000 290.4000 ;
	    RECT 170.8000 290.3000 171.6000 290.4000 ;
	    RECT 166.0000 289.7000 171.6000 290.3000 ;
	    RECT 166.0000 289.6000 166.8000 289.7000 ;
	    RECT 170.8000 289.6000 171.6000 289.7000 ;
	    RECT 234.8000 290.3000 235.6000 290.4000 ;
	    RECT 244.4000 290.3000 245.2000 290.4000 ;
	    RECT 234.8000 289.7000 245.2000 290.3000 ;
	    RECT 234.8000 289.6000 235.6000 289.7000 ;
	    RECT 244.4000 289.6000 245.2000 289.7000 ;
	    RECT 266.8000 290.3000 267.6000 290.4000 ;
	    RECT 281.2000 290.3000 282.0000 290.4000 ;
	    RECT 266.8000 289.7000 282.0000 290.3000 ;
	    RECT 266.8000 289.6000 267.6000 289.7000 ;
	    RECT 281.2000 289.6000 282.0000 289.7000 ;
	    RECT 289.2000 289.6000 290.0000 290.4000 ;
	    RECT 297.2000 290.3000 298.0000 290.4000 ;
	    RECT 305.2000 290.3000 306.0000 290.4000 ;
	    RECT 297.2000 289.7000 306.0000 290.3000 ;
	    RECT 297.2000 289.6000 298.0000 289.7000 ;
	    RECT 305.2000 289.6000 306.0000 289.7000 ;
	    RECT 306.8000 290.3000 307.6000 290.4000 ;
	    RECT 318.0000 290.3000 318.8000 290.4000 ;
	    RECT 306.8000 289.7000 318.8000 290.3000 ;
	    RECT 306.8000 289.6000 307.6000 289.7000 ;
	    RECT 318.0000 289.6000 318.8000 289.7000 ;
	    RECT 322.8000 290.3000 323.6000 290.4000 ;
	    RECT 335.6000 290.3000 336.4000 290.4000 ;
	    RECT 322.8000 289.7000 336.4000 290.3000 ;
	    RECT 322.8000 289.6000 323.6000 289.7000 ;
	    RECT 335.6000 289.6000 336.4000 289.7000 ;
	    RECT 372.4000 290.3000 373.2000 290.4000 ;
	    RECT 378.8000 290.3000 379.6000 290.4000 ;
	    RECT 372.4000 289.7000 379.6000 290.3000 ;
	    RECT 372.4000 289.6000 373.2000 289.7000 ;
	    RECT 378.8000 289.6000 379.6000 289.7000 ;
	    RECT 426.8000 290.3000 427.6000 290.4000 ;
	    RECT 431.6000 290.3000 432.4000 290.4000 ;
	    RECT 426.8000 289.7000 432.4000 290.3000 ;
	    RECT 426.8000 289.6000 427.6000 289.7000 ;
	    RECT 431.6000 289.6000 432.4000 289.7000 ;
	    RECT 505.2000 290.3000 506.0000 290.4000 ;
	    RECT 510.0000 290.3000 510.8000 290.4000 ;
	    RECT 505.2000 289.7000 510.8000 290.3000 ;
	    RECT 505.2000 289.6000 506.0000 289.7000 ;
	    RECT 510.0000 289.6000 510.8000 289.7000 ;
	    RECT 63.6000 288.3000 64.4000 288.4000 ;
	    RECT 76.4000 288.3000 77.2000 288.4000 ;
	    RECT 63.6000 287.7000 77.2000 288.3000 ;
	    RECT 63.6000 287.6000 64.4000 287.7000 ;
	    RECT 76.4000 287.6000 77.2000 287.7000 ;
	    RECT 97.2000 288.3000 98.0000 288.4000 ;
	    RECT 129.2000 288.3000 130.0000 288.4000 ;
	    RECT 202.8000 288.3000 203.6000 288.4000 ;
	    RECT 207.6000 288.3000 208.4000 288.4000 ;
	    RECT 97.2000 287.7000 208.4000 288.3000 ;
	    RECT 97.2000 287.6000 98.0000 287.7000 ;
	    RECT 129.2000 287.6000 130.0000 287.7000 ;
	    RECT 202.8000 287.6000 203.6000 287.7000 ;
	    RECT 207.6000 287.6000 208.4000 287.7000 ;
	    RECT 209.2000 288.3000 210.0000 288.4000 ;
	    RECT 276.4000 288.3000 277.2000 288.4000 ;
	    RECT 209.2000 287.7000 277.2000 288.3000 ;
	    RECT 209.2000 287.6000 210.0000 287.7000 ;
	    RECT 276.4000 287.6000 277.2000 287.7000 ;
	    RECT 279.6000 288.3000 280.4000 288.4000 ;
	    RECT 287.6000 288.3000 288.4000 288.4000 ;
	    RECT 279.6000 287.7000 288.4000 288.3000 ;
	    RECT 289.3000 288.3000 289.9000 289.6000 ;
	    RECT 407.6000 288.3000 408.4000 288.4000 ;
	    RECT 289.3000 287.7000 408.4000 288.3000 ;
	    RECT 279.6000 287.6000 280.4000 287.7000 ;
	    RECT 287.6000 287.6000 288.4000 287.7000 ;
	    RECT 407.6000 287.6000 408.4000 287.7000 ;
	    RECT 420.4000 288.3000 421.2000 288.4000 ;
	    RECT 430.0000 288.3000 430.8000 288.4000 ;
	    RECT 420.4000 287.7000 430.8000 288.3000 ;
	    RECT 420.4000 287.6000 421.2000 287.7000 ;
	    RECT 430.0000 287.6000 430.8000 287.7000 ;
	    RECT 462.0000 288.3000 462.8000 288.4000 ;
	    RECT 470.0000 288.3000 470.8000 288.4000 ;
	    RECT 462.0000 287.7000 470.8000 288.3000 ;
	    RECT 462.0000 287.6000 462.8000 287.7000 ;
	    RECT 470.0000 287.6000 470.8000 287.7000 ;
	    RECT 87.6000 286.3000 88.4000 286.4000 ;
	    RECT 113.2000 286.3000 114.0000 286.4000 ;
	    RECT 87.6000 285.7000 114.0000 286.3000 ;
	    RECT 87.6000 285.6000 88.4000 285.7000 ;
	    RECT 113.2000 285.6000 114.0000 285.7000 ;
	    RECT 114.8000 286.3000 115.6000 286.4000 ;
	    RECT 166.0000 286.3000 166.8000 286.4000 ;
	    RECT 114.8000 285.7000 166.8000 286.3000 ;
	    RECT 114.8000 285.6000 115.6000 285.7000 ;
	    RECT 166.0000 285.6000 166.8000 285.7000 ;
	    RECT 170.8000 286.3000 171.6000 286.4000 ;
	    RECT 174.0000 286.3000 174.8000 286.4000 ;
	    RECT 214.0000 286.3000 214.8000 286.4000 ;
	    RECT 170.8000 285.7000 214.8000 286.3000 ;
	    RECT 170.8000 285.6000 171.6000 285.7000 ;
	    RECT 174.0000 285.6000 174.8000 285.7000 ;
	    RECT 214.0000 285.6000 214.8000 285.7000 ;
	    RECT 217.2000 286.3000 218.0000 286.4000 ;
	    RECT 218.8000 286.3000 219.6000 286.4000 ;
	    RECT 217.2000 285.7000 219.6000 286.3000 ;
	    RECT 217.2000 285.6000 218.0000 285.7000 ;
	    RECT 218.8000 285.6000 219.6000 285.7000 ;
	    RECT 220.4000 286.3000 221.2000 286.4000 ;
	    RECT 250.8000 286.3000 251.6000 286.4000 ;
	    RECT 220.4000 285.7000 251.6000 286.3000 ;
	    RECT 220.4000 285.6000 221.2000 285.7000 ;
	    RECT 250.8000 285.6000 251.6000 285.7000 ;
	    RECT 257.2000 286.3000 258.0000 286.4000 ;
	    RECT 263.6000 286.3000 264.4000 286.4000 ;
	    RECT 268.4000 286.3000 269.2000 286.4000 ;
	    RECT 257.2000 285.7000 269.2000 286.3000 ;
	    RECT 257.2000 285.6000 258.0000 285.7000 ;
	    RECT 263.6000 285.6000 264.4000 285.7000 ;
	    RECT 268.4000 285.6000 269.2000 285.7000 ;
	    RECT 278.0000 286.3000 278.8000 286.4000 ;
	    RECT 284.4000 286.3000 285.2000 286.4000 ;
	    RECT 286.0000 286.3000 286.8000 286.4000 ;
	    RECT 294.0000 286.3000 294.8000 286.4000 ;
	    RECT 298.8000 286.3000 299.6000 286.4000 ;
	    RECT 306.8000 286.3000 307.6000 286.4000 ;
	    RECT 278.0000 285.7000 307.6000 286.3000 ;
	    RECT 278.0000 285.6000 278.8000 285.7000 ;
	    RECT 284.4000 285.6000 285.2000 285.7000 ;
	    RECT 286.0000 285.6000 286.8000 285.7000 ;
	    RECT 294.0000 285.6000 294.8000 285.7000 ;
	    RECT 298.8000 285.6000 299.6000 285.7000 ;
	    RECT 306.8000 285.6000 307.6000 285.7000 ;
	    RECT 308.4000 286.3000 309.2000 286.4000 ;
	    RECT 327.6000 286.3000 328.4000 286.4000 ;
	    RECT 308.4000 285.7000 328.4000 286.3000 ;
	    RECT 308.4000 285.6000 309.2000 285.7000 ;
	    RECT 327.6000 285.6000 328.4000 285.7000 ;
	    RECT 334.0000 286.3000 334.8000 286.4000 ;
	    RECT 338.8000 286.3000 339.6000 286.4000 ;
	    RECT 334.0000 285.7000 339.6000 286.3000 ;
	    RECT 334.0000 285.6000 334.8000 285.7000 ;
	    RECT 338.8000 285.6000 339.6000 285.7000 ;
	    RECT 342.0000 286.3000 342.8000 286.4000 ;
	    RECT 380.4000 286.3000 381.2000 286.4000 ;
	    RECT 342.0000 285.7000 381.2000 286.3000 ;
	    RECT 342.0000 285.6000 342.8000 285.7000 ;
	    RECT 380.4000 285.6000 381.2000 285.7000 ;
	    RECT 394.8000 286.3000 395.6000 286.4000 ;
	    RECT 418.8000 286.3000 419.6000 286.4000 ;
	    RECT 434.8000 286.3000 435.6000 286.4000 ;
	    RECT 394.8000 285.7000 435.6000 286.3000 ;
	    RECT 394.8000 285.6000 395.6000 285.7000 ;
	    RECT 418.8000 285.6000 419.6000 285.7000 ;
	    RECT 434.8000 285.6000 435.6000 285.7000 ;
	    RECT 470.0000 286.3000 470.8000 286.4000 ;
	    RECT 494.0000 286.3000 494.8000 286.4000 ;
	    RECT 497.2000 286.3000 498.0000 286.4000 ;
	    RECT 470.0000 285.7000 498.0000 286.3000 ;
	    RECT 470.0000 285.6000 470.8000 285.7000 ;
	    RECT 494.0000 285.6000 494.8000 285.7000 ;
	    RECT 497.2000 285.6000 498.0000 285.7000 ;
	    RECT 506.8000 286.3000 507.6000 286.4000 ;
	    RECT 508.4000 286.3000 509.2000 286.4000 ;
	    RECT 506.8000 285.7000 509.2000 286.3000 ;
	    RECT 506.8000 285.6000 507.6000 285.7000 ;
	    RECT 508.4000 285.6000 509.2000 285.7000 ;
	    RECT 73.2000 284.3000 74.0000 284.4000 ;
	    RECT 138.8000 284.3000 139.6000 284.4000 ;
	    RECT 206.0000 284.3000 206.8000 284.4000 ;
	    RECT 73.2000 283.7000 112.3000 284.3000 ;
	    RECT 73.2000 283.6000 74.0000 283.7000 ;
	    RECT 33.2000 282.3000 34.0000 282.4000 ;
	    RECT 65.2000 282.3000 66.0000 282.4000 ;
	    RECT 33.2000 281.7000 66.0000 282.3000 ;
	    RECT 33.2000 281.6000 34.0000 281.7000 ;
	    RECT 65.2000 281.6000 66.0000 281.7000 ;
	    RECT 89.2000 282.3000 90.0000 282.4000 ;
	    RECT 102.0000 282.3000 102.8000 282.4000 ;
	    RECT 89.2000 281.7000 102.8000 282.3000 ;
	    RECT 111.7000 282.3000 112.3000 283.7000 ;
	    RECT 138.8000 283.7000 206.8000 284.3000 ;
	    RECT 138.8000 283.6000 139.6000 283.7000 ;
	    RECT 206.0000 283.6000 206.8000 283.7000 ;
	    RECT 207.6000 284.3000 208.4000 284.4000 ;
	    RECT 273.2000 284.3000 274.0000 284.4000 ;
	    RECT 207.6000 283.7000 274.0000 284.3000 ;
	    RECT 207.6000 283.6000 208.4000 283.7000 ;
	    RECT 273.2000 283.6000 274.0000 283.7000 ;
	    RECT 276.4000 284.3000 277.2000 284.4000 ;
	    RECT 295.6000 284.3000 296.4000 284.4000 ;
	    RECT 276.4000 283.7000 296.4000 284.3000 ;
	    RECT 276.4000 283.6000 277.2000 283.7000 ;
	    RECT 295.6000 283.6000 296.4000 283.7000 ;
	    RECT 297.2000 284.3000 298.0000 284.4000 ;
	    RECT 300.4000 284.3000 301.2000 284.4000 ;
	    RECT 297.2000 283.7000 301.2000 284.3000 ;
	    RECT 297.2000 283.6000 298.0000 283.7000 ;
	    RECT 300.4000 283.6000 301.2000 283.7000 ;
	    RECT 302.0000 284.3000 302.8000 284.4000 ;
	    RECT 310.0000 284.3000 310.8000 284.4000 ;
	    RECT 302.0000 283.7000 310.8000 284.3000 ;
	    RECT 302.0000 283.6000 302.8000 283.7000 ;
	    RECT 310.0000 283.6000 310.8000 283.7000 ;
	    RECT 313.2000 284.3000 314.0000 284.4000 ;
	    RECT 327.6000 284.3000 328.4000 284.4000 ;
	    RECT 313.2000 283.7000 328.4000 284.3000 ;
	    RECT 313.2000 283.6000 314.0000 283.7000 ;
	    RECT 327.6000 283.6000 328.4000 283.7000 ;
	    RECT 334.0000 284.3000 334.8000 284.4000 ;
	    RECT 351.6000 284.3000 352.4000 284.4000 ;
	    RECT 334.0000 283.7000 352.4000 284.3000 ;
	    RECT 334.0000 283.6000 334.8000 283.7000 ;
	    RECT 351.6000 283.6000 352.4000 283.7000 ;
	    RECT 361.2000 284.3000 362.0000 284.4000 ;
	    RECT 406.0000 284.3000 406.8000 284.4000 ;
	    RECT 361.2000 283.7000 406.8000 284.3000 ;
	    RECT 361.2000 283.6000 362.0000 283.7000 ;
	    RECT 406.0000 283.6000 406.8000 283.7000 ;
	    RECT 407.6000 284.3000 408.4000 284.4000 ;
	    RECT 415.6000 284.3000 416.4000 284.4000 ;
	    RECT 422.0000 284.3000 422.8000 284.4000 ;
	    RECT 407.6000 283.7000 422.8000 284.3000 ;
	    RECT 407.6000 283.6000 408.4000 283.7000 ;
	    RECT 415.6000 283.6000 416.4000 283.7000 ;
	    RECT 422.0000 283.6000 422.8000 283.7000 ;
	    RECT 198.0000 282.3000 198.8000 282.4000 ;
	    RECT 111.7000 281.7000 198.8000 282.3000 ;
	    RECT 89.2000 281.6000 90.0000 281.7000 ;
	    RECT 102.0000 281.6000 102.8000 281.7000 ;
	    RECT 198.0000 281.6000 198.8000 281.7000 ;
	    RECT 199.6000 282.3000 200.4000 282.4000 ;
	    RECT 206.0000 282.3000 206.8000 282.4000 ;
	    RECT 199.6000 281.7000 206.8000 282.3000 ;
	    RECT 199.6000 281.6000 200.4000 281.7000 ;
	    RECT 206.0000 281.6000 206.8000 281.7000 ;
	    RECT 214.0000 282.3000 214.8000 282.4000 ;
	    RECT 356.4000 282.3000 357.2000 282.4000 ;
	    RECT 214.0000 281.7000 357.2000 282.3000 ;
	    RECT 214.0000 281.6000 214.8000 281.7000 ;
	    RECT 356.4000 281.6000 357.2000 281.7000 ;
	    RECT 358.0000 282.3000 358.8000 282.4000 ;
	    RECT 383.6000 282.3000 384.4000 282.4000 ;
	    RECT 391.6000 282.3000 392.4000 282.4000 ;
	    RECT 358.0000 281.7000 392.4000 282.3000 ;
	    RECT 358.0000 281.6000 358.8000 281.7000 ;
	    RECT 383.6000 281.6000 384.4000 281.7000 ;
	    RECT 391.6000 281.6000 392.4000 281.7000 ;
	    RECT 92.4000 280.3000 93.2000 280.4000 ;
	    RECT 100.4000 280.3000 101.2000 280.4000 ;
	    RECT 92.4000 279.7000 101.2000 280.3000 ;
	    RECT 92.4000 279.6000 93.2000 279.7000 ;
	    RECT 100.4000 279.6000 101.2000 279.7000 ;
	    RECT 111.6000 280.3000 112.4000 280.4000 ;
	    RECT 129.2000 280.3000 130.0000 280.4000 ;
	    RECT 111.6000 279.7000 130.0000 280.3000 ;
	    RECT 111.6000 279.6000 112.4000 279.7000 ;
	    RECT 129.2000 279.6000 130.0000 279.7000 ;
	    RECT 132.4000 280.3000 133.2000 280.4000 ;
	    RECT 150.0000 280.3000 150.8000 280.4000 ;
	    RECT 132.4000 279.7000 150.8000 280.3000 ;
	    RECT 132.4000 279.6000 133.2000 279.7000 ;
	    RECT 150.0000 279.6000 150.8000 279.7000 ;
	    RECT 170.8000 280.3000 171.6000 280.4000 ;
	    RECT 190.0000 280.3000 190.8000 280.4000 ;
	    RECT 170.8000 279.7000 190.8000 280.3000 ;
	    RECT 170.8000 279.6000 171.6000 279.7000 ;
	    RECT 190.0000 279.6000 190.8000 279.7000 ;
	    RECT 193.2000 280.3000 194.0000 280.4000 ;
	    RECT 199.6000 280.3000 200.4000 280.4000 ;
	    RECT 225.2000 280.3000 226.0000 280.4000 ;
	    RECT 193.2000 279.7000 226.0000 280.3000 ;
	    RECT 193.2000 279.6000 194.0000 279.7000 ;
	    RECT 199.6000 279.6000 200.4000 279.7000 ;
	    RECT 225.2000 279.6000 226.0000 279.7000 ;
	    RECT 231.6000 280.3000 232.4000 280.4000 ;
	    RECT 246.0000 280.3000 246.8000 280.4000 ;
	    RECT 231.6000 279.7000 246.8000 280.3000 ;
	    RECT 231.6000 279.6000 232.4000 279.7000 ;
	    RECT 246.0000 279.6000 246.8000 279.7000 ;
	    RECT 249.2000 280.3000 250.0000 280.4000 ;
	    RECT 249.2000 279.7000 360.3000 280.3000 ;
	    RECT 249.2000 279.6000 250.0000 279.7000 ;
	    RECT 20.4000 278.3000 21.2000 278.4000 ;
	    RECT 55.6000 278.3000 56.4000 278.4000 ;
	    RECT 20.4000 277.7000 56.4000 278.3000 ;
	    RECT 20.4000 277.6000 21.2000 277.7000 ;
	    RECT 55.6000 277.6000 56.4000 277.7000 ;
	    RECT 86.0000 278.3000 86.8000 278.4000 ;
	    RECT 114.8000 278.3000 115.6000 278.4000 ;
	    RECT 86.0000 277.7000 115.6000 278.3000 ;
	    RECT 86.0000 277.6000 86.8000 277.7000 ;
	    RECT 114.8000 277.6000 115.6000 277.7000 ;
	    RECT 126.0000 278.3000 126.8000 278.4000 ;
	    RECT 127.6000 278.3000 128.4000 278.4000 ;
	    RECT 145.2000 278.3000 146.0000 278.4000 ;
	    RECT 158.0000 278.3000 158.8000 278.4000 ;
	    RECT 186.8000 278.3000 187.6000 278.4000 ;
	    RECT 210.8000 278.3000 211.6000 278.4000 ;
	    RECT 126.0000 277.7000 184.3000 278.3000 ;
	    RECT 126.0000 277.6000 126.8000 277.7000 ;
	    RECT 127.6000 277.6000 128.4000 277.7000 ;
	    RECT 145.2000 277.6000 146.0000 277.7000 ;
	    RECT 158.0000 277.6000 158.8000 277.7000 ;
	    RECT 183.7000 276.4000 184.3000 277.7000 ;
	    RECT 186.8000 277.7000 211.6000 278.3000 ;
	    RECT 186.8000 277.6000 187.6000 277.7000 ;
	    RECT 210.8000 277.6000 211.6000 277.7000 ;
	    RECT 212.4000 278.3000 213.2000 278.4000 ;
	    RECT 226.8000 278.3000 227.6000 278.4000 ;
	    RECT 212.4000 277.7000 227.6000 278.3000 ;
	    RECT 212.4000 277.6000 213.2000 277.7000 ;
	    RECT 226.8000 277.6000 227.6000 277.7000 ;
	    RECT 239.6000 278.3000 240.4000 278.4000 ;
	    RECT 249.2000 278.3000 250.0000 278.4000 ;
	    RECT 239.6000 277.7000 250.0000 278.3000 ;
	    RECT 239.6000 277.6000 240.4000 277.7000 ;
	    RECT 249.2000 277.6000 250.0000 277.7000 ;
	    RECT 250.8000 278.3000 251.6000 278.4000 ;
	    RECT 308.4000 278.3000 309.2000 278.4000 ;
	    RECT 250.8000 277.7000 309.2000 278.3000 ;
	    RECT 250.8000 277.6000 251.6000 277.7000 ;
	    RECT 308.4000 277.6000 309.2000 277.7000 ;
	    RECT 311.6000 278.3000 312.4000 278.4000 ;
	    RECT 316.4000 278.3000 317.2000 278.4000 ;
	    RECT 358.0000 278.3000 358.8000 278.4000 ;
	    RECT 311.6000 277.7000 358.8000 278.3000 ;
	    RECT 359.7000 278.3000 360.3000 279.7000 ;
	    RECT 471.6000 278.3000 472.4000 278.4000 ;
	    RECT 359.7000 277.7000 472.4000 278.3000 ;
	    RECT 311.6000 277.6000 312.4000 277.7000 ;
	    RECT 316.4000 277.6000 317.2000 277.7000 ;
	    RECT 358.0000 277.6000 358.8000 277.7000 ;
	    RECT 471.6000 277.6000 472.4000 277.7000 ;
	    RECT 478.0000 278.3000 478.8000 278.4000 ;
	    RECT 492.4000 278.3000 493.2000 278.4000 ;
	    RECT 478.0000 277.7000 493.2000 278.3000 ;
	    RECT 478.0000 277.6000 478.8000 277.7000 ;
	    RECT 492.4000 277.6000 493.2000 277.7000 ;
	    RECT 47.6000 276.3000 48.4000 276.4000 ;
	    RECT 70.0000 276.3000 70.8000 276.4000 ;
	    RECT 47.6000 275.7000 70.8000 276.3000 ;
	    RECT 47.6000 275.6000 48.4000 275.7000 ;
	    RECT 70.0000 275.6000 70.8000 275.7000 ;
	    RECT 73.2000 276.3000 74.0000 276.4000 ;
	    RECT 84.4000 276.3000 85.2000 276.4000 ;
	    RECT 148.4000 276.3000 149.2000 276.4000 ;
	    RECT 73.2000 275.7000 81.9000 276.3000 ;
	    RECT 73.2000 275.6000 74.0000 275.7000 ;
	    RECT 14.0000 274.3000 14.8000 274.4000 ;
	    RECT 58.8000 274.3000 59.6000 274.4000 ;
	    RECT 14.0000 273.7000 59.6000 274.3000 ;
	    RECT 14.0000 273.6000 14.8000 273.7000 ;
	    RECT 58.8000 273.6000 59.6000 273.7000 ;
	    RECT 66.8000 274.3000 67.6000 274.4000 ;
	    RECT 79.6000 274.3000 80.4000 274.4000 ;
	    RECT 66.8000 273.7000 80.4000 274.3000 ;
	    RECT 81.3000 274.3000 81.9000 275.7000 ;
	    RECT 84.4000 275.7000 149.2000 276.3000 ;
	    RECT 84.4000 275.6000 85.2000 275.7000 ;
	    RECT 148.4000 275.6000 149.2000 275.7000 ;
	    RECT 150.0000 276.3000 150.8000 276.4000 ;
	    RECT 182.0000 276.3000 182.8000 276.4000 ;
	    RECT 150.0000 275.7000 182.8000 276.3000 ;
	    RECT 150.0000 275.6000 150.8000 275.7000 ;
	    RECT 182.0000 275.6000 182.8000 275.7000 ;
	    RECT 183.6000 276.3000 184.4000 276.4000 ;
	    RECT 209.2000 276.3000 210.0000 276.4000 ;
	    RECT 222.0000 276.3000 222.8000 276.4000 ;
	    RECT 242.8000 276.3000 243.6000 276.4000 ;
	    RECT 265.2000 276.3000 266.0000 276.4000 ;
	    RECT 279.6000 276.3000 280.4000 276.4000 ;
	    RECT 183.6000 275.7000 243.6000 276.3000 ;
	    RECT 183.6000 275.6000 184.4000 275.7000 ;
	    RECT 209.2000 275.6000 210.0000 275.7000 ;
	    RECT 222.0000 275.6000 222.8000 275.7000 ;
	    RECT 242.8000 275.6000 243.6000 275.7000 ;
	    RECT 244.5000 275.7000 266.0000 276.3000 ;
	    RECT 87.6000 274.3000 88.4000 274.4000 ;
	    RECT 81.3000 273.7000 88.4000 274.3000 ;
	    RECT 66.8000 273.6000 67.6000 273.7000 ;
	    RECT 79.6000 273.6000 80.4000 273.7000 ;
	    RECT 87.6000 273.6000 88.4000 273.7000 ;
	    RECT 90.8000 274.3000 91.6000 274.4000 ;
	    RECT 114.8000 274.3000 115.6000 274.4000 ;
	    RECT 121.2000 274.3000 122.0000 274.4000 ;
	    RECT 145.2000 274.3000 146.0000 274.4000 ;
	    RECT 185.2000 274.3000 186.0000 274.4000 ;
	    RECT 90.8000 273.7000 186.0000 274.3000 ;
	    RECT 90.8000 273.6000 91.6000 273.7000 ;
	    RECT 114.8000 273.6000 115.6000 273.7000 ;
	    RECT 121.2000 273.6000 122.0000 273.7000 ;
	    RECT 145.2000 273.6000 146.0000 273.7000 ;
	    RECT 185.2000 273.6000 186.0000 273.7000 ;
	    RECT 186.8000 274.3000 187.6000 274.4000 ;
	    RECT 196.4000 274.3000 197.2000 274.4000 ;
	    RECT 186.8000 273.7000 197.2000 274.3000 ;
	    RECT 186.8000 273.6000 187.6000 273.7000 ;
	    RECT 196.4000 273.6000 197.2000 273.7000 ;
	    RECT 198.0000 274.3000 198.8000 274.4000 ;
	    RECT 220.4000 274.3000 221.2000 274.4000 ;
	    RECT 198.0000 273.7000 221.2000 274.3000 ;
	    RECT 198.0000 273.6000 198.8000 273.7000 ;
	    RECT 220.4000 273.6000 221.2000 273.7000 ;
	    RECT 228.4000 274.3000 229.2000 274.4000 ;
	    RECT 244.5000 274.3000 245.1000 275.7000 ;
	    RECT 265.2000 275.6000 266.0000 275.7000 ;
	    RECT 266.9000 275.7000 280.4000 276.3000 ;
	    RECT 228.4000 273.7000 245.1000 274.3000 ;
	    RECT 250.8000 274.3000 251.6000 274.4000 ;
	    RECT 266.9000 274.3000 267.5000 275.7000 ;
	    RECT 279.6000 275.6000 280.4000 275.7000 ;
	    RECT 284.4000 276.3000 285.2000 276.4000 ;
	    RECT 378.8000 276.3000 379.6000 276.4000 ;
	    RECT 390.0000 276.3000 390.8000 276.4000 ;
	    RECT 420.4000 276.3000 421.2000 276.4000 ;
	    RECT 426.8000 276.3000 427.6000 276.4000 ;
	    RECT 284.4000 275.7000 377.9000 276.3000 ;
	    RECT 284.4000 275.6000 285.2000 275.7000 ;
	    RECT 250.8000 273.7000 267.5000 274.3000 ;
	    RECT 276.4000 274.3000 277.2000 274.4000 ;
	    RECT 290.8000 274.3000 291.6000 274.4000 ;
	    RECT 276.4000 273.7000 291.6000 274.3000 ;
	    RECT 228.4000 273.6000 229.2000 273.7000 ;
	    RECT 250.8000 273.6000 251.6000 273.7000 ;
	    RECT 276.4000 273.6000 277.2000 273.7000 ;
	    RECT 290.8000 273.6000 291.6000 273.7000 ;
	    RECT 298.8000 274.3000 299.6000 274.4000 ;
	    RECT 302.0000 274.3000 302.8000 274.4000 ;
	    RECT 298.8000 273.7000 302.8000 274.3000 ;
	    RECT 298.8000 273.6000 299.6000 273.7000 ;
	    RECT 302.0000 273.6000 302.8000 273.7000 ;
	    RECT 305.2000 274.3000 306.0000 274.4000 ;
	    RECT 308.4000 274.3000 309.2000 274.4000 ;
	    RECT 305.2000 273.7000 309.2000 274.3000 ;
	    RECT 305.2000 273.6000 306.0000 273.7000 ;
	    RECT 308.4000 273.6000 309.2000 273.7000 ;
	    RECT 310.0000 274.3000 310.8000 274.4000 ;
	    RECT 319.6000 274.3000 320.4000 274.4000 ;
	    RECT 310.0000 273.7000 320.4000 274.3000 ;
	    RECT 310.0000 273.6000 310.8000 273.7000 ;
	    RECT 319.6000 273.6000 320.4000 273.7000 ;
	    RECT 330.8000 274.3000 331.6000 274.4000 ;
	    RECT 340.4000 274.3000 341.2000 274.4000 ;
	    RECT 375.6000 274.3000 376.4000 274.4000 ;
	    RECT 330.8000 273.7000 376.4000 274.3000 ;
	    RECT 377.3000 274.3000 377.9000 275.7000 ;
	    RECT 378.8000 275.7000 427.6000 276.3000 ;
	    RECT 378.8000 275.6000 379.6000 275.7000 ;
	    RECT 390.0000 275.6000 390.8000 275.7000 ;
	    RECT 420.4000 275.6000 421.2000 275.7000 ;
	    RECT 426.8000 275.6000 427.6000 275.7000 ;
	    RECT 484.4000 276.3000 485.2000 276.4000 ;
	    RECT 487.6000 276.3000 488.4000 276.4000 ;
	    RECT 484.4000 275.7000 488.4000 276.3000 ;
	    RECT 484.4000 275.6000 485.2000 275.7000 ;
	    RECT 487.6000 275.6000 488.4000 275.7000 ;
	    RECT 393.2000 274.3000 394.0000 274.4000 ;
	    RECT 417.2000 274.3000 418.0000 274.4000 ;
	    RECT 377.3000 273.7000 418.0000 274.3000 ;
	    RECT 330.8000 273.6000 331.6000 273.7000 ;
	    RECT 340.4000 273.6000 341.2000 273.7000 ;
	    RECT 375.6000 273.6000 376.4000 273.7000 ;
	    RECT 393.2000 273.6000 394.0000 273.7000 ;
	    RECT 417.2000 273.6000 418.0000 273.7000 ;
	    RECT 454.0000 274.3000 454.8000 274.4000 ;
	    RECT 457.2000 274.3000 458.0000 274.4000 ;
	    RECT 454.0000 273.7000 458.0000 274.3000 ;
	    RECT 454.0000 273.6000 454.8000 273.7000 ;
	    RECT 457.2000 273.6000 458.0000 273.7000 ;
	    RECT 458.8000 274.3000 459.6000 274.4000 ;
	    RECT 462.0000 274.3000 462.8000 274.4000 ;
	    RECT 458.8000 273.7000 462.8000 274.3000 ;
	    RECT 458.8000 273.6000 459.6000 273.7000 ;
	    RECT 462.0000 273.6000 462.8000 273.7000 ;
	    RECT 471.6000 274.3000 472.4000 274.4000 ;
	    RECT 490.8000 274.3000 491.6000 274.4000 ;
	    RECT 471.6000 273.7000 491.6000 274.3000 ;
	    RECT 471.6000 273.6000 472.4000 273.7000 ;
	    RECT 490.8000 273.6000 491.6000 273.7000 ;
	    RECT 4.4000 272.3000 5.2000 272.4000 ;
	    RECT 17.2000 272.3000 18.0000 272.4000 ;
	    RECT 4.4000 271.7000 18.0000 272.3000 ;
	    RECT 4.4000 271.6000 5.2000 271.7000 ;
	    RECT 17.2000 271.6000 18.0000 271.7000 ;
	    RECT 54.0000 272.3000 54.8000 272.4000 ;
	    RECT 63.6000 272.3000 64.4000 272.4000 ;
	    RECT 54.0000 271.7000 64.4000 272.3000 ;
	    RECT 54.0000 271.6000 54.8000 271.7000 ;
	    RECT 63.6000 271.6000 64.4000 271.7000 ;
	    RECT 76.4000 272.3000 77.2000 272.4000 ;
	    RECT 82.8000 272.3000 83.6000 272.4000 ;
	    RECT 89.2000 272.3000 90.0000 272.4000 ;
	    RECT 76.4000 271.7000 90.0000 272.3000 ;
	    RECT 76.4000 271.6000 77.2000 271.7000 ;
	    RECT 82.8000 271.6000 83.6000 271.7000 ;
	    RECT 89.2000 271.6000 90.0000 271.7000 ;
	    RECT 90.8000 272.3000 91.6000 272.4000 ;
	    RECT 142.0000 272.3000 142.8000 272.4000 ;
	    RECT 90.8000 271.7000 142.8000 272.3000 ;
	    RECT 90.8000 271.6000 91.6000 271.7000 ;
	    RECT 142.0000 271.6000 142.8000 271.7000 ;
	    RECT 143.6000 272.3000 144.4000 272.4000 ;
	    RECT 146.8000 272.3000 147.6000 272.4000 ;
	    RECT 143.6000 271.7000 147.6000 272.3000 ;
	    RECT 143.6000 271.6000 144.4000 271.7000 ;
	    RECT 146.8000 271.6000 147.6000 271.7000 ;
	    RECT 148.4000 272.3000 149.2000 272.4000 ;
	    RECT 180.4000 272.3000 181.2000 272.4000 ;
	    RECT 148.4000 271.7000 181.2000 272.3000 ;
	    RECT 148.4000 271.6000 149.2000 271.7000 ;
	    RECT 180.4000 271.6000 181.2000 271.7000 ;
	    RECT 186.8000 272.3000 187.6000 272.4000 ;
	    RECT 193.2000 272.3000 194.0000 272.4000 ;
	    RECT 186.8000 271.7000 194.0000 272.3000 ;
	    RECT 186.8000 271.6000 187.6000 271.7000 ;
	    RECT 193.2000 271.6000 194.0000 271.7000 ;
	    RECT 194.8000 272.3000 195.6000 272.4000 ;
	    RECT 215.6000 272.3000 216.4000 272.4000 ;
	    RECT 194.8000 271.7000 216.4000 272.3000 ;
	    RECT 194.8000 271.6000 195.6000 271.7000 ;
	    RECT 215.6000 271.6000 216.4000 271.7000 ;
	    RECT 223.6000 272.3000 224.4000 272.4000 ;
	    RECT 233.2000 272.3000 234.0000 272.4000 ;
	    RECT 223.6000 271.7000 234.0000 272.3000 ;
	    RECT 223.6000 271.6000 224.4000 271.7000 ;
	    RECT 233.2000 271.6000 234.0000 271.7000 ;
	    RECT 234.8000 272.3000 235.6000 272.4000 ;
	    RECT 238.0000 272.3000 238.8000 272.4000 ;
	    RECT 234.8000 271.7000 238.8000 272.3000 ;
	    RECT 234.8000 271.6000 235.6000 271.7000 ;
	    RECT 238.0000 271.6000 238.8000 271.7000 ;
	    RECT 250.8000 272.3000 251.6000 272.4000 ;
	    RECT 284.4000 272.3000 285.2000 272.4000 ;
	    RECT 250.8000 271.7000 285.2000 272.3000 ;
	    RECT 250.8000 271.6000 251.6000 271.7000 ;
	    RECT 284.4000 271.6000 285.2000 271.7000 ;
	    RECT 286.0000 272.3000 286.8000 272.4000 ;
	    RECT 290.8000 272.3000 291.6000 272.4000 ;
	    RECT 286.0000 271.7000 291.6000 272.3000 ;
	    RECT 286.0000 271.6000 286.8000 271.7000 ;
	    RECT 290.8000 271.6000 291.6000 271.7000 ;
	    RECT 292.4000 271.6000 293.2000 272.4000 ;
	    RECT 295.6000 272.3000 296.4000 272.4000 ;
	    RECT 313.2000 272.3000 314.0000 272.4000 ;
	    RECT 295.6000 271.7000 314.0000 272.3000 ;
	    RECT 295.6000 271.6000 296.4000 271.7000 ;
	    RECT 313.2000 271.6000 314.0000 271.7000 ;
	    RECT 318.0000 272.3000 318.8000 272.4000 ;
	    RECT 326.0000 272.3000 326.8000 272.4000 ;
	    RECT 318.0000 271.7000 326.8000 272.3000 ;
	    RECT 318.0000 271.6000 318.8000 271.7000 ;
	    RECT 326.0000 271.6000 326.8000 271.7000 ;
	    RECT 327.6000 272.3000 328.4000 272.4000 ;
	    RECT 343.6000 272.3000 344.4000 272.4000 ;
	    RECT 327.6000 271.7000 344.4000 272.3000 ;
	    RECT 327.6000 271.6000 328.4000 271.7000 ;
	    RECT 343.6000 271.6000 344.4000 271.7000 ;
	    RECT 345.2000 272.3000 346.0000 272.4000 ;
	    RECT 359.6000 272.3000 360.4000 272.4000 ;
	    RECT 345.2000 271.7000 360.4000 272.3000 ;
	    RECT 345.2000 271.6000 346.0000 271.7000 ;
	    RECT 359.6000 271.6000 360.4000 271.7000 ;
	    RECT 374.0000 272.3000 374.8000 272.4000 ;
	    RECT 402.8000 272.3000 403.6000 272.4000 ;
	    RECT 414.0000 272.3000 414.8000 272.4000 ;
	    RECT 374.0000 271.7000 414.8000 272.3000 ;
	    RECT 374.0000 271.6000 374.8000 271.7000 ;
	    RECT 402.8000 271.6000 403.6000 271.7000 ;
	    RECT 414.0000 271.6000 414.8000 271.7000 ;
	    RECT 417.2000 272.3000 418.0000 272.4000 ;
	    RECT 422.0000 272.3000 422.8000 272.4000 ;
	    RECT 417.2000 271.7000 422.8000 272.3000 ;
	    RECT 417.2000 271.6000 418.0000 271.7000 ;
	    RECT 422.0000 271.6000 422.8000 271.7000 ;
	    RECT 457.2000 272.3000 458.0000 272.4000 ;
	    RECT 474.8000 272.3000 475.6000 272.4000 ;
	    RECT 510.0000 272.3000 510.8000 272.4000 ;
	    RECT 457.2000 271.7000 510.8000 272.3000 ;
	    RECT 457.2000 271.6000 458.0000 271.7000 ;
	    RECT 474.8000 271.6000 475.6000 271.7000 ;
	    RECT 510.0000 271.6000 510.8000 271.7000 ;
	    RECT 17.2000 270.3000 18.0000 270.4000 ;
	    RECT 38.0000 270.3000 38.8000 270.4000 ;
	    RECT 17.2000 269.7000 38.8000 270.3000 ;
	    RECT 17.2000 269.6000 18.0000 269.7000 ;
	    RECT 38.0000 269.6000 38.8000 269.7000 ;
	    RECT 52.4000 270.3000 53.2000 270.4000 ;
	    RECT 71.6000 270.3000 72.4000 270.4000 ;
	    RECT 52.4000 269.7000 72.4000 270.3000 ;
	    RECT 52.4000 269.6000 53.2000 269.7000 ;
	    RECT 71.6000 269.6000 72.4000 269.7000 ;
	    RECT 74.8000 270.3000 75.6000 270.4000 ;
	    RECT 78.0000 270.3000 78.8000 270.4000 ;
	    RECT 74.8000 269.7000 78.8000 270.3000 ;
	    RECT 74.8000 269.6000 75.6000 269.7000 ;
	    RECT 78.0000 269.6000 78.8000 269.7000 ;
	    RECT 81.2000 270.3000 82.0000 270.4000 ;
	    RECT 100.4000 270.3000 101.2000 270.4000 ;
	    RECT 81.2000 269.7000 101.2000 270.3000 ;
	    RECT 81.2000 269.6000 82.0000 269.7000 ;
	    RECT 100.4000 269.6000 101.2000 269.7000 ;
	    RECT 103.6000 270.3000 104.4000 270.4000 ;
	    RECT 146.8000 270.3000 147.6000 270.4000 ;
	    RECT 103.6000 269.7000 147.6000 270.3000 ;
	    RECT 103.6000 269.6000 104.4000 269.7000 ;
	    RECT 146.8000 269.6000 147.6000 269.7000 ;
	    RECT 161.2000 270.3000 162.0000 270.4000 ;
	    RECT 186.8000 270.3000 187.6000 270.4000 ;
	    RECT 161.2000 269.7000 187.6000 270.3000 ;
	    RECT 161.2000 269.6000 162.0000 269.7000 ;
	    RECT 186.8000 269.6000 187.6000 269.7000 ;
	    RECT 190.0000 270.3000 190.8000 270.4000 ;
	    RECT 196.4000 270.3000 197.2000 270.4000 ;
	    RECT 190.0000 269.7000 197.2000 270.3000 ;
	    RECT 190.0000 269.6000 190.8000 269.7000 ;
	    RECT 196.4000 269.6000 197.2000 269.7000 ;
	    RECT 198.0000 270.3000 198.8000 270.4000 ;
	    RECT 206.0000 270.3000 206.8000 270.4000 ;
	    RECT 212.4000 270.3000 213.2000 270.4000 ;
	    RECT 198.0000 269.7000 213.2000 270.3000 ;
	    RECT 198.0000 269.6000 198.8000 269.7000 ;
	    RECT 206.0000 269.6000 206.8000 269.7000 ;
	    RECT 212.4000 269.6000 213.2000 269.7000 ;
	    RECT 215.6000 270.3000 216.4000 270.4000 ;
	    RECT 225.2000 270.3000 226.0000 270.4000 ;
	    RECT 215.6000 269.7000 226.0000 270.3000 ;
	    RECT 215.6000 269.6000 216.4000 269.7000 ;
	    RECT 225.2000 269.6000 226.0000 269.7000 ;
	    RECT 228.4000 270.3000 229.2000 270.4000 ;
	    RECT 244.4000 270.3000 245.2000 270.4000 ;
	    RECT 270.0000 270.3000 270.8000 270.4000 ;
	    RECT 286.0000 270.3000 286.8000 270.4000 ;
	    RECT 314.8000 270.3000 315.6000 270.4000 ;
	    RECT 319.6000 270.3000 320.4000 270.4000 ;
	    RECT 338.8000 270.3000 339.6000 270.4000 ;
	    RECT 228.4000 269.7000 339.6000 270.3000 ;
	    RECT 228.4000 269.6000 229.2000 269.7000 ;
	    RECT 244.4000 269.6000 245.2000 269.7000 ;
	    RECT 270.0000 269.6000 270.8000 269.7000 ;
	    RECT 286.0000 269.6000 286.8000 269.7000 ;
	    RECT 314.8000 269.6000 315.6000 269.7000 ;
	    RECT 319.6000 269.6000 320.4000 269.7000 ;
	    RECT 338.8000 269.6000 339.6000 269.7000 ;
	    RECT 353.2000 269.6000 354.0000 270.4000 ;
	    RECT 354.8000 270.3000 355.6000 270.4000 ;
	    RECT 364.4000 270.3000 365.2000 270.4000 ;
	    RECT 354.8000 269.7000 365.2000 270.3000 ;
	    RECT 354.8000 269.6000 355.6000 269.7000 ;
	    RECT 364.4000 269.6000 365.2000 269.7000 ;
	    RECT 372.4000 270.3000 373.2000 270.4000 ;
	    RECT 374.0000 270.3000 374.8000 270.4000 ;
	    RECT 372.4000 269.7000 374.8000 270.3000 ;
	    RECT 372.4000 269.6000 373.2000 269.7000 ;
	    RECT 374.0000 269.6000 374.8000 269.7000 ;
	    RECT 380.4000 270.3000 381.2000 270.4000 ;
	    RECT 396.4000 270.3000 397.2000 270.4000 ;
	    RECT 380.4000 269.7000 397.2000 270.3000 ;
	    RECT 380.4000 269.6000 381.2000 269.7000 ;
	    RECT 396.4000 269.6000 397.2000 269.7000 ;
	    RECT 404.4000 270.3000 405.2000 270.4000 ;
	    RECT 422.0000 270.3000 422.8000 270.4000 ;
	    RECT 404.4000 269.7000 422.8000 270.3000 ;
	    RECT 404.4000 269.6000 405.2000 269.7000 ;
	    RECT 422.0000 269.6000 422.8000 269.7000 ;
	    RECT 450.8000 270.3000 451.6000 270.4000 ;
	    RECT 495.6000 270.3000 496.4000 270.4000 ;
	    RECT 450.8000 269.7000 496.4000 270.3000 ;
	    RECT 450.8000 269.6000 451.6000 269.7000 ;
	    RECT 495.6000 269.6000 496.4000 269.7000 ;
	    RECT 497.2000 270.3000 498.0000 270.4000 ;
	    RECT 500.4000 270.3000 501.2000 270.4000 ;
	    RECT 497.2000 269.7000 501.2000 270.3000 ;
	    RECT 497.2000 269.6000 498.0000 269.7000 ;
	    RECT 500.4000 269.6000 501.2000 269.7000 ;
	    RECT 4.4000 268.3000 5.2000 268.4000 ;
	    RECT 20.4000 268.3000 21.2000 268.4000 ;
	    RECT 4.4000 267.7000 21.2000 268.3000 ;
	    RECT 4.4000 267.6000 5.2000 267.7000 ;
	    RECT 20.4000 267.6000 21.2000 267.7000 ;
	    RECT 31.6000 268.3000 32.4000 268.4000 ;
	    RECT 38.0000 268.3000 38.8000 268.4000 ;
	    RECT 31.6000 267.7000 38.8000 268.3000 ;
	    RECT 31.6000 267.6000 32.4000 267.7000 ;
	    RECT 38.0000 267.6000 38.8000 267.7000 ;
	    RECT 42.8000 268.3000 43.6000 268.4000 ;
	    RECT 60.4000 268.3000 61.2000 268.4000 ;
	    RECT 79.6000 268.3000 80.4000 268.4000 ;
	    RECT 42.8000 267.7000 51.5000 268.3000 ;
	    RECT 42.8000 267.6000 43.6000 267.7000 ;
	    RECT 10.8000 266.3000 11.6000 266.4000 ;
	    RECT 49.2000 266.3000 50.0000 266.4000 ;
	    RECT 10.8000 265.7000 50.0000 266.3000 ;
	    RECT 50.9000 266.3000 51.5000 267.7000 ;
	    RECT 60.4000 267.7000 80.4000 268.3000 ;
	    RECT 60.4000 267.6000 61.2000 267.7000 ;
	    RECT 79.6000 267.6000 80.4000 267.7000 ;
	    RECT 81.2000 268.3000 82.0000 268.4000 ;
	    RECT 87.6000 268.3000 88.4000 268.4000 ;
	    RECT 92.4000 268.3000 93.2000 268.4000 ;
	    RECT 81.2000 267.7000 93.2000 268.3000 ;
	    RECT 81.2000 267.6000 82.0000 267.7000 ;
	    RECT 87.6000 267.6000 88.4000 267.7000 ;
	    RECT 92.4000 267.6000 93.2000 267.7000 ;
	    RECT 100.4000 268.3000 101.2000 268.4000 ;
	    RECT 111.6000 268.3000 112.4000 268.4000 ;
	    RECT 100.4000 267.7000 112.4000 268.3000 ;
	    RECT 100.4000 267.6000 101.2000 267.7000 ;
	    RECT 111.6000 267.6000 112.4000 267.7000 ;
	    RECT 121.2000 268.3000 122.0000 268.4000 ;
	    RECT 122.8000 268.3000 123.6000 268.4000 ;
	    RECT 124.4000 268.3000 125.2000 268.4000 ;
	    RECT 121.2000 267.7000 125.2000 268.3000 ;
	    RECT 121.2000 267.6000 122.0000 267.7000 ;
	    RECT 122.8000 267.6000 123.6000 267.7000 ;
	    RECT 124.4000 267.6000 125.2000 267.7000 ;
	    RECT 129.2000 268.3000 130.0000 268.4000 ;
	    RECT 150.0000 268.3000 150.8000 268.4000 ;
	    RECT 129.2000 267.7000 150.8000 268.3000 ;
	    RECT 129.2000 267.6000 130.0000 267.7000 ;
	    RECT 150.0000 267.6000 150.8000 267.7000 ;
	    RECT 290.8000 268.3000 291.6000 268.4000 ;
	    RECT 300.4000 268.3000 301.2000 268.4000 ;
	    RECT 321.2000 268.3000 322.0000 268.4000 ;
	    RECT 367.6000 268.3000 368.4000 268.4000 ;
	    RECT 372.4000 268.3000 373.2000 268.4000 ;
	    RECT 290.8000 267.7000 373.2000 268.3000 ;
	    RECT 290.8000 267.6000 291.6000 267.7000 ;
	    RECT 300.4000 267.6000 301.2000 267.7000 ;
	    RECT 321.2000 267.6000 322.0000 267.7000 ;
	    RECT 367.6000 267.6000 368.4000 267.7000 ;
	    RECT 372.4000 267.6000 373.2000 267.7000 ;
	    RECT 478.0000 268.3000 478.8000 268.4000 ;
	    RECT 503.6000 268.3000 504.4000 268.4000 ;
	    RECT 478.0000 267.7000 504.4000 268.3000 ;
	    RECT 478.0000 267.6000 478.8000 267.7000 ;
	    RECT 503.6000 267.6000 504.4000 267.7000 ;
	    RECT 103.6000 266.3000 104.4000 266.4000 ;
	    RECT 50.9000 265.7000 104.4000 266.3000 ;
	    RECT 10.8000 265.6000 11.6000 265.7000 ;
	    RECT 49.2000 265.6000 50.0000 265.7000 ;
	    RECT 103.6000 265.6000 104.4000 265.7000 ;
	    RECT 119.6000 266.3000 120.4000 266.4000 ;
	    RECT 129.2000 266.3000 130.0000 266.4000 ;
	    RECT 119.6000 265.7000 130.0000 266.3000 ;
	    RECT 119.6000 265.6000 120.4000 265.7000 ;
	    RECT 129.2000 265.6000 130.0000 265.7000 ;
	    RECT 130.8000 266.3000 131.6000 266.4000 ;
	    RECT 134.0000 266.3000 134.8000 266.4000 ;
	    RECT 130.8000 265.7000 134.8000 266.3000 ;
	    RECT 130.8000 265.6000 131.6000 265.7000 ;
	    RECT 134.0000 265.6000 134.8000 265.7000 ;
	    RECT 135.6000 266.3000 136.4000 266.4000 ;
	    RECT 140.4000 266.3000 141.2000 266.4000 ;
	    RECT 142.0000 266.3000 142.8000 266.4000 ;
	    RECT 135.6000 265.7000 142.8000 266.3000 ;
	    RECT 135.6000 265.6000 136.4000 265.7000 ;
	    RECT 140.4000 265.6000 141.2000 265.7000 ;
	    RECT 142.0000 265.6000 142.8000 265.7000 ;
	    RECT 182.0000 266.3000 182.8000 266.4000 ;
	    RECT 183.6000 266.3000 184.4000 266.4000 ;
	    RECT 182.0000 265.7000 184.4000 266.3000 ;
	    RECT 182.0000 265.6000 182.8000 265.7000 ;
	    RECT 183.6000 265.6000 184.4000 265.7000 ;
	    RECT 185.2000 266.3000 186.0000 266.4000 ;
	    RECT 188.4000 266.3000 189.2000 266.4000 ;
	    RECT 185.2000 265.7000 189.2000 266.3000 ;
	    RECT 185.2000 265.6000 186.0000 265.7000 ;
	    RECT 188.4000 265.6000 189.2000 265.7000 ;
	    RECT 191.6000 266.3000 192.4000 266.4000 ;
	    RECT 198.0000 266.3000 198.8000 266.4000 ;
	    RECT 191.6000 265.7000 198.8000 266.3000 ;
	    RECT 191.6000 265.6000 192.4000 265.7000 ;
	    RECT 198.0000 265.6000 198.8000 265.7000 ;
	    RECT 202.8000 265.6000 203.6000 266.4000 ;
	    RECT 210.8000 266.3000 211.6000 266.4000 ;
	    RECT 214.0000 266.3000 214.8000 266.4000 ;
	    RECT 210.8000 265.7000 214.8000 266.3000 ;
	    RECT 210.8000 265.6000 211.6000 265.7000 ;
	    RECT 214.0000 265.6000 214.8000 265.7000 ;
	    RECT 215.6000 266.3000 216.4000 266.4000 ;
	    RECT 234.8000 266.3000 235.6000 266.4000 ;
	    RECT 215.6000 265.7000 235.6000 266.3000 ;
	    RECT 215.6000 265.6000 216.4000 265.7000 ;
	    RECT 234.8000 265.6000 235.6000 265.7000 ;
	    RECT 236.4000 266.3000 237.2000 266.4000 ;
	    RECT 244.4000 266.3000 245.2000 266.4000 ;
	    RECT 303.6000 266.3000 304.4000 266.4000 ;
	    RECT 236.4000 265.7000 304.4000 266.3000 ;
	    RECT 236.4000 265.6000 237.2000 265.7000 ;
	    RECT 244.4000 265.6000 245.2000 265.7000 ;
	    RECT 303.6000 265.6000 304.4000 265.7000 ;
	    RECT 305.2000 265.6000 306.0000 266.4000 ;
	    RECT 306.8000 266.3000 307.6000 266.4000 ;
	    RECT 324.4000 266.3000 325.2000 266.4000 ;
	    RECT 306.8000 265.7000 325.2000 266.3000 ;
	    RECT 306.8000 265.6000 307.6000 265.7000 ;
	    RECT 324.4000 265.6000 325.2000 265.7000 ;
	    RECT 351.6000 266.3000 352.4000 266.4000 ;
	    RECT 356.4000 266.3000 357.2000 266.4000 ;
	    RECT 374.0000 266.3000 374.8000 266.4000 ;
	    RECT 399.6000 266.3000 400.4000 266.4000 ;
	    RECT 351.6000 265.7000 373.1000 266.3000 ;
	    RECT 351.6000 265.6000 352.4000 265.7000 ;
	    RECT 356.4000 265.6000 357.2000 265.7000 ;
	    RECT 6.0000 264.3000 6.8000 264.4000 ;
	    RECT 57.2000 264.3000 58.0000 264.4000 ;
	    RECT 6.0000 263.7000 58.0000 264.3000 ;
	    RECT 6.0000 263.6000 6.8000 263.7000 ;
	    RECT 57.2000 263.6000 58.0000 263.7000 ;
	    RECT 68.4000 264.3000 69.2000 264.4000 ;
	    RECT 137.2000 264.3000 138.0000 264.4000 ;
	    RECT 68.4000 263.7000 138.0000 264.3000 ;
	    RECT 142.1000 264.3000 142.7000 265.6000 ;
	    RECT 204.4000 264.3000 205.2000 264.4000 ;
	    RECT 206.0000 264.3000 206.8000 264.4000 ;
	    RECT 142.1000 263.7000 206.8000 264.3000 ;
	    RECT 68.4000 263.6000 69.2000 263.7000 ;
	    RECT 137.2000 263.6000 138.0000 263.7000 ;
	    RECT 204.4000 263.6000 205.2000 263.7000 ;
	    RECT 206.0000 263.6000 206.8000 263.7000 ;
	    RECT 209.2000 264.3000 210.0000 264.4000 ;
	    RECT 236.4000 264.3000 237.2000 264.4000 ;
	    RECT 209.2000 263.7000 237.2000 264.3000 ;
	    RECT 209.2000 263.6000 210.0000 263.7000 ;
	    RECT 236.4000 263.6000 237.2000 263.7000 ;
	    RECT 250.8000 264.3000 251.6000 264.4000 ;
	    RECT 262.0000 264.3000 262.8000 264.4000 ;
	    RECT 297.2000 264.3000 298.0000 264.4000 ;
	    RECT 298.8000 264.3000 299.6000 264.4000 ;
	    RECT 313.2000 264.3000 314.0000 264.4000 ;
	    RECT 250.8000 263.7000 314.0000 264.3000 ;
	    RECT 250.8000 263.6000 251.6000 263.7000 ;
	    RECT 262.0000 263.6000 262.8000 263.7000 ;
	    RECT 297.2000 263.6000 298.0000 263.7000 ;
	    RECT 298.8000 263.6000 299.6000 263.7000 ;
	    RECT 313.2000 263.6000 314.0000 263.7000 ;
	    RECT 314.8000 264.3000 315.6000 264.4000 ;
	    RECT 330.8000 264.3000 331.6000 264.4000 ;
	    RECT 354.8000 264.3000 355.6000 264.4000 ;
	    RECT 314.8000 263.7000 355.6000 264.3000 ;
	    RECT 314.8000 263.6000 315.6000 263.7000 ;
	    RECT 330.8000 263.6000 331.6000 263.7000 ;
	    RECT 354.8000 263.6000 355.6000 263.7000 ;
	    RECT 356.4000 264.3000 357.2000 264.4000 ;
	    RECT 358.0000 264.3000 358.8000 264.4000 ;
	    RECT 356.4000 263.7000 358.8000 264.3000 ;
	    RECT 372.5000 264.3000 373.1000 265.7000 ;
	    RECT 374.0000 265.7000 400.4000 266.3000 ;
	    RECT 374.0000 265.6000 374.8000 265.7000 ;
	    RECT 399.6000 265.6000 400.4000 265.7000 ;
	    RECT 484.4000 266.3000 485.2000 266.4000 ;
	    RECT 497.2000 266.3000 498.0000 266.4000 ;
	    RECT 484.4000 265.7000 498.0000 266.3000 ;
	    RECT 484.4000 265.6000 485.2000 265.7000 ;
	    RECT 497.2000 265.6000 498.0000 265.7000 ;
	    RECT 426.8000 264.3000 427.6000 264.4000 ;
	    RECT 433.2000 264.3000 434.0000 264.4000 ;
	    RECT 372.5000 263.7000 434.0000 264.3000 ;
	    RECT 356.4000 263.6000 357.2000 263.7000 ;
	    RECT 358.0000 263.6000 358.8000 263.7000 ;
	    RECT 426.8000 263.6000 427.6000 263.7000 ;
	    RECT 433.2000 263.6000 434.0000 263.7000 ;
	    RECT 439.6000 264.3000 440.4000 264.4000 ;
	    RECT 454.0000 264.3000 454.8000 264.4000 ;
	    RECT 439.6000 263.7000 454.8000 264.3000 ;
	    RECT 439.6000 263.6000 440.4000 263.7000 ;
	    RECT 454.0000 263.6000 454.8000 263.7000 ;
	    RECT 41.2000 262.3000 42.0000 262.4000 ;
	    RECT 57.2000 262.3000 58.0000 262.4000 ;
	    RECT 41.2000 261.7000 58.0000 262.3000 ;
	    RECT 41.2000 261.6000 42.0000 261.7000 ;
	    RECT 57.2000 261.6000 58.0000 261.7000 ;
	    RECT 60.4000 262.3000 61.2000 262.4000 ;
	    RECT 126.0000 262.3000 126.8000 262.4000 ;
	    RECT 60.4000 261.7000 126.8000 262.3000 ;
	    RECT 60.4000 261.6000 61.2000 261.7000 ;
	    RECT 126.0000 261.6000 126.8000 261.7000 ;
	    RECT 132.4000 262.3000 133.2000 262.4000 ;
	    RECT 135.6000 262.3000 136.4000 262.4000 ;
	    RECT 148.4000 262.3000 149.2000 262.4000 ;
	    RECT 175.6000 262.3000 176.4000 262.4000 ;
	    RECT 177.2000 262.3000 178.0000 262.4000 ;
	    RECT 194.8000 262.3000 195.6000 262.4000 ;
	    RECT 132.4000 261.7000 195.6000 262.3000 ;
	    RECT 132.4000 261.6000 133.2000 261.7000 ;
	    RECT 135.6000 261.6000 136.4000 261.7000 ;
	    RECT 148.4000 261.6000 149.2000 261.7000 ;
	    RECT 175.6000 261.6000 176.4000 261.7000 ;
	    RECT 177.2000 261.6000 178.0000 261.7000 ;
	    RECT 194.8000 261.6000 195.6000 261.7000 ;
	    RECT 209.2000 262.3000 210.0000 262.4000 ;
	    RECT 218.8000 262.3000 219.6000 262.4000 ;
	    RECT 209.2000 261.7000 219.6000 262.3000 ;
	    RECT 209.2000 261.6000 210.0000 261.7000 ;
	    RECT 218.8000 261.6000 219.6000 261.7000 ;
	    RECT 263.6000 262.3000 264.4000 262.4000 ;
	    RECT 266.8000 262.3000 267.6000 262.4000 ;
	    RECT 350.0000 262.3000 350.8000 262.4000 ;
	    RECT 263.6000 261.7000 350.8000 262.3000 ;
	    RECT 263.6000 261.6000 264.4000 261.7000 ;
	    RECT 266.8000 261.6000 267.6000 261.7000 ;
	    RECT 350.0000 261.6000 350.8000 261.7000 ;
	    RECT 353.2000 262.3000 354.0000 262.4000 ;
	    RECT 385.2000 262.3000 386.0000 262.4000 ;
	    RECT 388.4000 262.3000 389.2000 262.4000 ;
	    RECT 425.2000 262.3000 426.0000 262.4000 ;
	    RECT 431.6000 262.3000 432.4000 262.4000 ;
	    RECT 449.2000 262.3000 450.0000 262.4000 ;
	    RECT 353.2000 261.7000 450.0000 262.3000 ;
	    RECT 353.2000 261.6000 354.0000 261.7000 ;
	    RECT 385.2000 261.6000 386.0000 261.7000 ;
	    RECT 388.4000 261.6000 389.2000 261.7000 ;
	    RECT 425.2000 261.6000 426.0000 261.7000 ;
	    RECT 431.6000 261.6000 432.4000 261.7000 ;
	    RECT 449.2000 261.6000 450.0000 261.7000 ;
	    RECT 44.4000 260.3000 45.2000 260.4000 ;
	    RECT 47.6000 260.3000 48.4000 260.4000 ;
	    RECT 44.4000 259.7000 48.4000 260.3000 ;
	    RECT 44.4000 259.6000 45.2000 259.7000 ;
	    RECT 47.6000 259.6000 48.4000 259.7000 ;
	    RECT 58.8000 260.3000 59.6000 260.4000 ;
	    RECT 62.0000 260.3000 62.8000 260.4000 ;
	    RECT 63.6000 260.3000 64.4000 260.4000 ;
	    RECT 129.2000 260.3000 130.0000 260.4000 ;
	    RECT 58.8000 259.7000 64.4000 260.3000 ;
	    RECT 58.8000 259.6000 59.6000 259.7000 ;
	    RECT 62.0000 259.6000 62.8000 259.7000 ;
	    RECT 63.6000 259.6000 64.4000 259.7000 ;
	    RECT 65.3000 259.7000 130.0000 260.3000 ;
	    RECT 62.0000 258.3000 62.8000 258.4000 ;
	    RECT 65.3000 258.3000 65.9000 259.7000 ;
	    RECT 129.2000 259.6000 130.0000 259.7000 ;
	    RECT 132.4000 260.3000 133.2000 260.4000 ;
	    RECT 140.4000 260.3000 141.2000 260.4000 ;
	    RECT 204.4000 260.3000 205.2000 260.4000 ;
	    RECT 239.6000 260.3000 240.4000 260.4000 ;
	    RECT 250.8000 260.3000 251.6000 260.4000 ;
	    RECT 132.4000 259.7000 201.9000 260.3000 ;
	    RECT 132.4000 259.6000 133.2000 259.7000 ;
	    RECT 140.4000 259.6000 141.2000 259.7000 ;
	    RECT 124.4000 258.3000 125.2000 258.4000 ;
	    RECT 62.0000 257.7000 65.9000 258.3000 ;
	    RECT 100.5000 257.7000 125.2000 258.3000 ;
	    RECT 62.0000 257.6000 62.8000 257.7000 ;
	    RECT 100.5000 256.4000 101.1000 257.7000 ;
	    RECT 124.4000 257.6000 125.2000 257.7000 ;
	    RECT 126.0000 258.3000 126.8000 258.4000 ;
	    RECT 164.4000 258.3000 165.2000 258.4000 ;
	    RECT 126.0000 257.7000 165.2000 258.3000 ;
	    RECT 126.0000 257.6000 126.8000 257.7000 ;
	    RECT 164.4000 257.6000 165.2000 257.7000 ;
	    RECT 172.4000 258.3000 173.2000 258.4000 ;
	    RECT 177.2000 258.3000 178.0000 258.4000 ;
	    RECT 193.2000 258.3000 194.0000 258.4000 ;
	    RECT 199.6000 258.3000 200.4000 258.4000 ;
	    RECT 172.4000 257.7000 200.4000 258.3000 ;
	    RECT 201.3000 258.3000 201.9000 259.7000 ;
	    RECT 204.4000 259.7000 235.5000 260.3000 ;
	    RECT 204.4000 259.6000 205.2000 259.7000 ;
	    RECT 234.9000 258.4000 235.5000 259.7000 ;
	    RECT 239.6000 259.7000 251.6000 260.3000 ;
	    RECT 239.6000 259.6000 240.4000 259.7000 ;
	    RECT 250.8000 259.6000 251.6000 259.7000 ;
	    RECT 266.8000 260.3000 267.6000 260.4000 ;
	    RECT 276.4000 260.3000 277.2000 260.4000 ;
	    RECT 266.8000 259.7000 277.2000 260.3000 ;
	    RECT 266.8000 259.6000 267.6000 259.7000 ;
	    RECT 276.4000 259.6000 277.2000 259.7000 ;
	    RECT 302.0000 259.6000 302.8000 260.4000 ;
	    RECT 303.6000 260.3000 304.4000 260.4000 ;
	    RECT 374.0000 260.3000 374.8000 260.4000 ;
	    RECT 303.6000 259.7000 374.8000 260.3000 ;
	    RECT 303.6000 259.6000 304.4000 259.7000 ;
	    RECT 374.0000 259.6000 374.8000 259.7000 ;
	    RECT 378.8000 260.3000 379.6000 260.4000 ;
	    RECT 382.0000 260.3000 382.8000 260.4000 ;
	    RECT 378.8000 259.7000 382.8000 260.3000 ;
	    RECT 378.8000 259.6000 379.6000 259.7000 ;
	    RECT 382.0000 259.6000 382.8000 259.7000 ;
	    RECT 452.4000 260.3000 453.2000 260.4000 ;
	    RECT 465.2000 260.3000 466.0000 260.4000 ;
	    RECT 452.4000 259.7000 466.0000 260.3000 ;
	    RECT 452.4000 259.6000 453.2000 259.7000 ;
	    RECT 465.2000 259.6000 466.0000 259.7000 ;
	    RECT 476.4000 260.3000 477.2000 260.4000 ;
	    RECT 479.6000 260.3000 480.4000 260.4000 ;
	    RECT 486.0000 260.3000 486.8000 260.4000 ;
	    RECT 476.4000 259.7000 486.8000 260.3000 ;
	    RECT 476.4000 259.6000 477.2000 259.7000 ;
	    RECT 479.6000 259.6000 480.4000 259.7000 ;
	    RECT 486.0000 259.6000 486.8000 259.7000 ;
	    RECT 502.0000 260.3000 502.8000 260.4000 ;
	    RECT 503.6000 260.3000 504.4000 260.4000 ;
	    RECT 502.0000 259.7000 504.4000 260.3000 ;
	    RECT 502.0000 259.6000 502.8000 259.7000 ;
	    RECT 503.6000 259.6000 504.4000 259.7000 ;
	    RECT 207.6000 258.3000 208.4000 258.4000 ;
	    RECT 201.3000 257.7000 208.4000 258.3000 ;
	    RECT 172.4000 257.6000 173.2000 257.7000 ;
	    RECT 177.2000 257.6000 178.0000 257.7000 ;
	    RECT 193.2000 257.6000 194.0000 257.7000 ;
	    RECT 199.6000 257.6000 200.4000 257.7000 ;
	    RECT 207.6000 257.6000 208.4000 257.7000 ;
	    RECT 210.8000 258.3000 211.6000 258.4000 ;
	    RECT 215.6000 258.3000 216.4000 258.4000 ;
	    RECT 210.8000 257.7000 216.4000 258.3000 ;
	    RECT 210.8000 257.6000 211.6000 257.7000 ;
	    RECT 215.6000 257.6000 216.4000 257.7000 ;
	    RECT 217.2000 257.6000 218.0000 258.4000 ;
	    RECT 220.4000 258.3000 221.2000 258.4000 ;
	    RECT 231.6000 258.3000 232.4000 258.4000 ;
	    RECT 220.4000 257.7000 232.4000 258.3000 ;
	    RECT 220.4000 257.6000 221.2000 257.7000 ;
	    RECT 231.6000 257.6000 232.4000 257.7000 ;
	    RECT 234.8000 258.3000 235.6000 258.4000 ;
	    RECT 430.0000 258.3000 430.8000 258.4000 ;
	    RECT 234.8000 257.7000 430.8000 258.3000 ;
	    RECT 234.8000 257.6000 235.6000 257.7000 ;
	    RECT 430.0000 257.6000 430.8000 257.7000 ;
	    RECT 450.8000 258.3000 451.6000 258.4000 ;
	    RECT 470.0000 258.3000 470.8000 258.4000 ;
	    RECT 450.8000 257.7000 470.8000 258.3000 ;
	    RECT 450.8000 257.6000 451.6000 257.7000 ;
	    RECT 470.0000 257.6000 470.8000 257.7000 ;
	    RECT 490.8000 258.3000 491.6000 258.4000 ;
	    RECT 505.2000 258.3000 506.0000 258.4000 ;
	    RECT 490.8000 257.7000 506.0000 258.3000 ;
	    RECT 490.8000 257.6000 491.6000 257.7000 ;
	    RECT 505.2000 257.6000 506.0000 257.7000 ;
	    RECT 33.2000 256.3000 34.0000 256.4000 ;
	    RECT 71.6000 256.3000 72.4000 256.4000 ;
	    RECT 73.2000 256.3000 74.0000 256.4000 ;
	    RECT 33.2000 255.7000 38.7000 256.3000 ;
	    RECT 33.2000 255.6000 34.0000 255.7000 ;
	    RECT 26.8000 254.3000 27.6000 254.4000 ;
	    RECT 31.6000 254.3000 32.4000 254.4000 ;
	    RECT 36.4000 254.3000 37.2000 254.4000 ;
	    RECT 26.8000 253.7000 37.2000 254.3000 ;
	    RECT 38.1000 254.3000 38.7000 255.7000 ;
	    RECT 71.6000 255.7000 74.0000 256.3000 ;
	    RECT 71.6000 255.6000 72.4000 255.7000 ;
	    RECT 73.2000 255.6000 74.0000 255.7000 ;
	    RECT 74.8000 256.3000 75.6000 256.4000 ;
	    RECT 76.4000 256.3000 77.2000 256.4000 ;
	    RECT 74.8000 255.7000 77.2000 256.3000 ;
	    RECT 74.8000 255.6000 75.6000 255.7000 ;
	    RECT 76.4000 255.6000 77.2000 255.7000 ;
	    RECT 87.6000 256.3000 88.4000 256.4000 ;
	    RECT 100.4000 256.3000 101.2000 256.4000 ;
	    RECT 87.6000 255.7000 101.2000 256.3000 ;
	    RECT 87.6000 255.6000 88.4000 255.7000 ;
	    RECT 100.4000 255.6000 101.2000 255.7000 ;
	    RECT 158.0000 256.3000 158.8000 256.4000 ;
	    RECT 161.2000 256.3000 162.0000 256.4000 ;
	    RECT 158.0000 255.7000 162.0000 256.3000 ;
	    RECT 158.0000 255.6000 158.8000 255.7000 ;
	    RECT 161.2000 255.6000 162.0000 255.7000 ;
	    RECT 170.8000 256.3000 171.6000 256.4000 ;
	    RECT 183.6000 256.3000 184.4000 256.4000 ;
	    RECT 196.4000 256.3000 197.2000 256.4000 ;
	    RECT 170.8000 255.7000 197.2000 256.3000 ;
	    RECT 170.8000 255.6000 171.6000 255.7000 ;
	    RECT 183.6000 255.6000 184.4000 255.7000 ;
	    RECT 196.4000 255.6000 197.2000 255.7000 ;
	    RECT 198.0000 256.3000 198.8000 256.4000 ;
	    RECT 217.3000 256.3000 217.9000 257.6000 ;
	    RECT 198.0000 255.7000 217.9000 256.3000 ;
	    RECT 218.8000 256.3000 219.6000 256.4000 ;
	    RECT 238.0000 256.3000 238.8000 256.4000 ;
	    RECT 258.8000 256.3000 259.6000 256.4000 ;
	    RECT 218.8000 255.7000 237.1000 256.3000 ;
	    RECT 198.0000 255.6000 198.8000 255.7000 ;
	    RECT 218.8000 255.6000 219.6000 255.7000 ;
	    RECT 50.8000 254.3000 51.6000 254.4000 ;
	    RECT 38.1000 253.7000 51.6000 254.3000 ;
	    RECT 26.8000 253.6000 27.6000 253.7000 ;
	    RECT 31.6000 253.6000 32.4000 253.7000 ;
	    RECT 36.4000 253.6000 37.2000 253.7000 ;
	    RECT 50.8000 253.6000 51.6000 253.7000 ;
	    RECT 55.6000 254.3000 56.4000 254.4000 ;
	    RECT 63.6000 254.3000 64.4000 254.4000 ;
	    RECT 55.6000 253.7000 64.4000 254.3000 ;
	    RECT 55.6000 253.6000 56.4000 253.7000 ;
	    RECT 63.6000 253.6000 64.4000 253.7000 ;
	    RECT 76.4000 254.3000 77.2000 254.4000 ;
	    RECT 90.8000 254.3000 91.6000 254.4000 ;
	    RECT 76.4000 253.7000 91.6000 254.3000 ;
	    RECT 76.4000 253.6000 77.2000 253.7000 ;
	    RECT 90.8000 253.6000 91.6000 253.7000 ;
	    RECT 113.2000 254.3000 114.0000 254.4000 ;
	    RECT 116.4000 254.3000 117.2000 254.4000 ;
	    RECT 113.2000 253.7000 117.2000 254.3000 ;
	    RECT 113.2000 253.6000 114.0000 253.7000 ;
	    RECT 116.4000 253.6000 117.2000 253.7000 ;
	    RECT 122.8000 254.3000 123.6000 254.4000 ;
	    RECT 138.8000 254.3000 139.6000 254.4000 ;
	    RECT 167.6000 254.3000 168.4000 254.4000 ;
	    RECT 122.8000 253.7000 139.6000 254.3000 ;
	    RECT 122.8000 253.6000 123.6000 253.7000 ;
	    RECT 138.8000 253.6000 139.6000 253.7000 ;
	    RECT 142.1000 253.7000 168.4000 254.3000 ;
	    RECT 142.1000 252.4000 142.7000 253.7000 ;
	    RECT 167.6000 253.6000 168.4000 253.7000 ;
	    RECT 182.0000 254.3000 182.8000 254.4000 ;
	    RECT 190.0000 254.3000 190.8000 254.4000 ;
	    RECT 214.0000 254.3000 214.8000 254.4000 ;
	    RECT 233.2000 254.3000 234.0000 254.4000 ;
	    RECT 234.8000 254.3000 235.6000 254.4000 ;
	    RECT 182.0000 253.7000 235.6000 254.3000 ;
	    RECT 236.5000 254.3000 237.1000 255.7000 ;
	    RECT 238.0000 255.7000 259.6000 256.3000 ;
	    RECT 238.0000 255.6000 238.8000 255.7000 ;
	    RECT 258.8000 255.6000 259.6000 255.7000 ;
	    RECT 260.4000 256.3000 261.2000 256.4000 ;
	    RECT 270.0000 256.3000 270.8000 256.4000 ;
	    RECT 260.4000 255.7000 270.8000 256.3000 ;
	    RECT 260.4000 255.6000 261.2000 255.7000 ;
	    RECT 270.0000 255.6000 270.8000 255.7000 ;
	    RECT 271.6000 256.3000 272.4000 256.4000 ;
	    RECT 386.8000 256.3000 387.6000 256.4000 ;
	    RECT 404.4000 256.3000 405.2000 256.4000 ;
	    RECT 271.6000 255.7000 365.1000 256.3000 ;
	    RECT 271.6000 255.6000 272.4000 255.7000 ;
	    RECT 313.2000 254.3000 314.0000 254.4000 ;
	    RECT 332.4000 254.3000 333.2000 254.4000 ;
	    RECT 236.5000 253.7000 333.2000 254.3000 ;
	    RECT 182.0000 253.6000 182.8000 253.7000 ;
	    RECT 190.0000 253.6000 190.8000 253.7000 ;
	    RECT 214.0000 253.6000 214.8000 253.7000 ;
	    RECT 233.2000 253.6000 234.0000 253.7000 ;
	    RECT 234.8000 253.6000 235.6000 253.7000 ;
	    RECT 313.2000 253.6000 314.0000 253.7000 ;
	    RECT 332.4000 253.6000 333.2000 253.7000 ;
	    RECT 348.4000 254.3000 349.2000 254.4000 ;
	    RECT 361.2000 254.3000 362.0000 254.4000 ;
	    RECT 362.8000 254.3000 363.6000 254.4000 ;
	    RECT 348.4000 253.7000 363.6000 254.3000 ;
	    RECT 364.5000 254.3000 365.1000 255.7000 ;
	    RECT 386.8000 255.7000 405.2000 256.3000 ;
	    RECT 386.8000 255.6000 387.6000 255.7000 ;
	    RECT 404.4000 255.6000 405.2000 255.7000 ;
	    RECT 409.2000 256.3000 410.0000 256.4000 ;
	    RECT 420.4000 256.3000 421.2000 256.4000 ;
	    RECT 409.2000 255.7000 421.2000 256.3000 ;
	    RECT 409.2000 255.6000 410.0000 255.7000 ;
	    RECT 420.4000 255.6000 421.2000 255.7000 ;
	    RECT 428.4000 256.3000 429.2000 256.4000 ;
	    RECT 447.6000 256.3000 448.4000 256.4000 ;
	    RECT 428.4000 255.7000 448.4000 256.3000 ;
	    RECT 428.4000 255.6000 429.2000 255.7000 ;
	    RECT 447.6000 255.6000 448.4000 255.7000 ;
	    RECT 463.6000 256.3000 464.4000 256.4000 ;
	    RECT 476.4000 256.3000 477.2000 256.4000 ;
	    RECT 463.6000 255.7000 477.2000 256.3000 ;
	    RECT 463.6000 255.6000 464.4000 255.7000 ;
	    RECT 476.4000 255.6000 477.2000 255.7000 ;
	    RECT 479.6000 256.3000 480.4000 256.4000 ;
	    RECT 513.2000 256.3000 514.0000 256.4000 ;
	    RECT 479.6000 255.7000 514.0000 256.3000 ;
	    RECT 479.6000 255.6000 480.4000 255.7000 ;
	    RECT 513.2000 255.6000 514.0000 255.7000 ;
	    RECT 479.7000 254.3000 480.3000 255.6000 ;
	    RECT 364.5000 253.7000 480.3000 254.3000 ;
	    RECT 481.2000 254.3000 482.0000 254.4000 ;
	    RECT 502.0000 254.3000 502.8000 254.4000 ;
	    RECT 506.8000 254.3000 507.6000 254.4000 ;
	    RECT 481.2000 253.7000 507.6000 254.3000 ;
	    RECT 348.4000 253.6000 349.2000 253.7000 ;
	    RECT 361.2000 253.6000 362.0000 253.7000 ;
	    RECT 362.8000 253.6000 363.6000 253.7000 ;
	    RECT 481.2000 253.6000 482.0000 253.7000 ;
	    RECT 502.0000 253.6000 502.8000 253.7000 ;
	    RECT 506.8000 253.6000 507.6000 253.7000 ;
	    RECT 23.6000 252.3000 24.4000 252.4000 ;
	    RECT 30.0000 252.3000 30.8000 252.4000 ;
	    RECT 23.6000 251.7000 30.8000 252.3000 ;
	    RECT 23.6000 251.6000 24.4000 251.7000 ;
	    RECT 30.0000 251.6000 30.8000 251.7000 ;
	    RECT 34.8000 252.3000 35.6000 252.4000 ;
	    RECT 62.0000 252.3000 62.8000 252.4000 ;
	    RECT 34.8000 251.7000 62.8000 252.3000 ;
	    RECT 34.8000 251.6000 35.6000 251.7000 ;
	    RECT 62.0000 251.6000 62.8000 251.7000 ;
	    RECT 90.8000 252.3000 91.6000 252.4000 ;
	    RECT 95.6000 252.3000 96.4000 252.4000 ;
	    RECT 97.2000 252.3000 98.0000 252.4000 ;
	    RECT 90.8000 251.7000 98.0000 252.3000 ;
	    RECT 90.8000 251.6000 91.6000 251.7000 ;
	    RECT 95.6000 251.6000 96.4000 251.7000 ;
	    RECT 97.2000 251.6000 98.0000 251.7000 ;
	    RECT 113.2000 252.3000 114.0000 252.4000 ;
	    RECT 129.2000 252.3000 130.0000 252.4000 ;
	    RECT 142.0000 252.3000 142.8000 252.4000 ;
	    RECT 113.2000 251.7000 142.8000 252.3000 ;
	    RECT 113.2000 251.6000 114.0000 251.7000 ;
	    RECT 129.2000 251.6000 130.0000 251.7000 ;
	    RECT 142.0000 251.6000 142.8000 251.7000 ;
	    RECT 154.8000 252.3000 155.6000 252.4000 ;
	    RECT 166.0000 252.3000 166.8000 252.4000 ;
	    RECT 154.8000 251.7000 166.8000 252.3000 ;
	    RECT 154.8000 251.6000 155.6000 251.7000 ;
	    RECT 166.0000 251.6000 166.8000 251.7000 ;
	    RECT 186.8000 252.3000 187.6000 252.4000 ;
	    RECT 196.4000 252.3000 197.2000 252.4000 ;
	    RECT 198.0000 252.3000 198.8000 252.4000 ;
	    RECT 186.8000 251.7000 195.5000 252.3000 ;
	    RECT 186.8000 251.6000 187.6000 251.7000 ;
	    RECT 50.8000 250.3000 51.6000 250.4000 ;
	    RECT 55.6000 250.3000 56.4000 250.4000 ;
	    RECT 50.8000 249.7000 56.4000 250.3000 ;
	    RECT 50.8000 249.6000 51.6000 249.7000 ;
	    RECT 55.6000 249.6000 56.4000 249.7000 ;
	    RECT 66.8000 250.3000 67.6000 250.4000 ;
	    RECT 111.6000 250.3000 112.4000 250.4000 ;
	    RECT 66.8000 249.7000 112.4000 250.3000 ;
	    RECT 66.8000 249.6000 67.6000 249.7000 ;
	    RECT 111.6000 249.6000 112.4000 249.7000 ;
	    RECT 119.6000 250.3000 120.4000 250.4000 ;
	    RECT 134.0000 250.3000 134.8000 250.4000 ;
	    RECT 140.4000 250.3000 141.2000 250.4000 ;
	    RECT 119.6000 249.7000 134.8000 250.3000 ;
	    RECT 119.6000 249.6000 120.4000 249.7000 ;
	    RECT 134.0000 249.6000 134.8000 249.7000 ;
	    RECT 135.7000 249.7000 141.2000 250.3000 ;
	    RECT 54.0000 248.3000 54.8000 248.4000 ;
	    RECT 116.4000 248.3000 117.2000 248.4000 ;
	    RECT 54.0000 247.7000 117.2000 248.3000 ;
	    RECT 54.0000 247.6000 54.8000 247.7000 ;
	    RECT 116.4000 247.6000 117.2000 247.7000 ;
	    RECT 121.2000 248.3000 122.0000 248.4000 ;
	    RECT 135.7000 248.3000 136.3000 249.7000 ;
	    RECT 140.4000 249.6000 141.2000 249.7000 ;
	    RECT 148.4000 250.3000 149.2000 250.4000 ;
	    RECT 150.0000 250.3000 150.8000 250.4000 ;
	    RECT 148.4000 249.7000 150.8000 250.3000 ;
	    RECT 148.4000 249.6000 149.2000 249.7000 ;
	    RECT 150.0000 249.6000 150.8000 249.7000 ;
	    RECT 161.2000 250.3000 162.0000 250.4000 ;
	    RECT 162.8000 250.3000 163.6000 250.4000 ;
	    RECT 161.2000 249.7000 163.6000 250.3000 ;
	    RECT 161.2000 249.6000 162.0000 249.7000 ;
	    RECT 162.8000 249.6000 163.6000 249.7000 ;
	    RECT 164.4000 250.3000 165.2000 250.4000 ;
	    RECT 190.0000 250.3000 190.8000 250.4000 ;
	    RECT 193.2000 250.3000 194.0000 250.4000 ;
	    RECT 164.4000 249.7000 189.1000 250.3000 ;
	    RECT 164.4000 249.6000 165.2000 249.7000 ;
	    RECT 121.2000 247.7000 136.3000 248.3000 ;
	    RECT 137.2000 248.3000 138.0000 248.4000 ;
	    RECT 150.0000 248.3000 150.8000 248.4000 ;
	    RECT 164.4000 248.3000 165.2000 248.4000 ;
	    RECT 186.8000 248.3000 187.6000 248.4000 ;
	    RECT 137.2000 247.7000 187.6000 248.3000 ;
	    RECT 188.5000 248.3000 189.1000 249.7000 ;
	    RECT 190.0000 249.7000 194.0000 250.3000 ;
	    RECT 194.9000 250.3000 195.5000 251.7000 ;
	    RECT 196.4000 251.7000 198.8000 252.3000 ;
	    RECT 196.4000 251.6000 197.2000 251.7000 ;
	    RECT 198.0000 251.6000 198.8000 251.7000 ;
	    RECT 212.4000 252.3000 213.2000 252.4000 ;
	    RECT 225.2000 252.3000 226.0000 252.4000 ;
	    RECT 212.4000 251.7000 226.0000 252.3000 ;
	    RECT 212.4000 251.6000 213.2000 251.7000 ;
	    RECT 225.2000 251.6000 226.0000 251.7000 ;
	    RECT 230.0000 252.3000 230.8000 252.4000 ;
	    RECT 255.6000 252.3000 256.4000 252.4000 ;
	    RECT 230.0000 251.7000 256.4000 252.3000 ;
	    RECT 230.0000 251.6000 230.8000 251.7000 ;
	    RECT 255.6000 251.6000 256.4000 251.7000 ;
	    RECT 257.2000 252.3000 258.0000 252.4000 ;
	    RECT 266.8000 252.3000 267.6000 252.4000 ;
	    RECT 257.2000 251.7000 267.6000 252.3000 ;
	    RECT 257.2000 251.6000 258.0000 251.7000 ;
	    RECT 266.8000 251.6000 267.6000 251.7000 ;
	    RECT 268.4000 252.3000 269.2000 252.4000 ;
	    RECT 271.6000 252.3000 272.4000 252.4000 ;
	    RECT 268.4000 251.7000 272.4000 252.3000 ;
	    RECT 268.4000 251.6000 269.2000 251.7000 ;
	    RECT 271.6000 251.6000 272.4000 251.7000 ;
	    RECT 273.2000 252.3000 274.0000 252.4000 ;
	    RECT 279.6000 252.3000 280.4000 252.4000 ;
	    RECT 292.4000 252.3000 293.2000 252.4000 ;
	    RECT 273.2000 251.7000 293.2000 252.3000 ;
	    RECT 273.2000 251.6000 274.0000 251.7000 ;
	    RECT 279.6000 251.6000 280.4000 251.7000 ;
	    RECT 292.4000 251.6000 293.2000 251.7000 ;
	    RECT 295.6000 252.3000 296.4000 252.4000 ;
	    RECT 300.4000 252.3000 301.2000 252.4000 ;
	    RECT 295.6000 251.7000 301.2000 252.3000 ;
	    RECT 295.6000 251.6000 296.4000 251.7000 ;
	    RECT 300.4000 251.6000 301.2000 251.7000 ;
	    RECT 326.0000 252.3000 326.8000 252.4000 ;
	    RECT 337.2000 252.3000 338.0000 252.4000 ;
	    RECT 326.0000 251.7000 338.0000 252.3000 ;
	    RECT 326.0000 251.6000 326.8000 251.7000 ;
	    RECT 337.2000 251.6000 338.0000 251.7000 ;
	    RECT 343.6000 251.6000 344.4000 252.4000 ;
	    RECT 350.0000 252.3000 350.8000 252.4000 ;
	    RECT 450.8000 252.3000 451.6000 252.4000 ;
	    RECT 350.0000 251.7000 451.6000 252.3000 ;
	    RECT 350.0000 251.6000 350.8000 251.7000 ;
	    RECT 450.8000 251.6000 451.6000 251.7000 ;
	    RECT 454.0000 252.3000 454.8000 252.4000 ;
	    RECT 466.8000 252.3000 467.6000 252.4000 ;
	    RECT 474.8000 252.3000 475.6000 252.4000 ;
	    RECT 510.0000 252.3000 510.8000 252.4000 ;
	    RECT 454.0000 251.7000 510.8000 252.3000 ;
	    RECT 454.0000 251.6000 454.8000 251.7000 ;
	    RECT 466.8000 251.6000 467.6000 251.7000 ;
	    RECT 474.8000 251.6000 475.6000 251.7000 ;
	    RECT 510.0000 251.6000 510.8000 251.7000 ;
	    RECT 196.4000 250.3000 197.2000 250.4000 ;
	    RECT 194.9000 249.7000 197.2000 250.3000 ;
	    RECT 190.0000 249.6000 190.8000 249.7000 ;
	    RECT 193.2000 249.6000 194.0000 249.7000 ;
	    RECT 196.4000 249.6000 197.2000 249.7000 ;
	    RECT 206.0000 250.3000 206.8000 250.4000 ;
	    RECT 218.8000 250.3000 219.6000 250.4000 ;
	    RECT 220.4000 250.3000 221.2000 250.4000 ;
	    RECT 206.0000 249.7000 221.2000 250.3000 ;
	    RECT 206.0000 249.6000 206.8000 249.7000 ;
	    RECT 218.8000 249.6000 219.6000 249.7000 ;
	    RECT 220.4000 249.6000 221.2000 249.7000 ;
	    RECT 226.8000 250.3000 227.6000 250.4000 ;
	    RECT 249.2000 250.3000 250.0000 250.4000 ;
	    RECT 266.8000 250.3000 267.6000 250.4000 ;
	    RECT 226.8000 249.7000 245.1000 250.3000 ;
	    RECT 226.8000 249.6000 227.6000 249.7000 ;
	    RECT 244.5000 248.4000 245.1000 249.7000 ;
	    RECT 249.2000 249.7000 267.6000 250.3000 ;
	    RECT 249.2000 249.6000 250.0000 249.7000 ;
	    RECT 266.8000 249.6000 267.6000 249.7000 ;
	    RECT 270.0000 250.3000 270.8000 250.4000 ;
	    RECT 305.2000 250.3000 306.0000 250.4000 ;
	    RECT 270.0000 249.7000 306.0000 250.3000 ;
	    RECT 270.0000 249.6000 270.8000 249.7000 ;
	    RECT 305.2000 249.6000 306.0000 249.7000 ;
	    RECT 335.6000 250.3000 336.4000 250.4000 ;
	    RECT 340.4000 250.3000 341.2000 250.4000 ;
	    RECT 335.6000 249.7000 341.2000 250.3000 ;
	    RECT 335.6000 249.6000 336.4000 249.7000 ;
	    RECT 340.4000 249.6000 341.2000 249.7000 ;
	    RECT 346.8000 250.3000 347.6000 250.4000 ;
	    RECT 353.2000 250.3000 354.0000 250.4000 ;
	    RECT 346.8000 249.7000 354.0000 250.3000 ;
	    RECT 346.8000 249.6000 347.6000 249.7000 ;
	    RECT 353.2000 249.6000 354.0000 249.7000 ;
	    RECT 356.4000 250.3000 357.2000 250.4000 ;
	    RECT 361.2000 250.3000 362.0000 250.4000 ;
	    RECT 356.4000 249.7000 362.0000 250.3000 ;
	    RECT 356.4000 249.6000 357.2000 249.7000 ;
	    RECT 361.2000 249.6000 362.0000 249.7000 ;
	    RECT 370.8000 250.3000 371.6000 250.4000 ;
	    RECT 383.6000 250.3000 384.4000 250.4000 ;
	    RECT 370.8000 249.7000 384.4000 250.3000 ;
	    RECT 370.8000 249.6000 371.6000 249.7000 ;
	    RECT 383.6000 249.6000 384.4000 249.7000 ;
	    RECT 406.0000 250.3000 406.8000 250.4000 ;
	    RECT 418.8000 250.3000 419.6000 250.4000 ;
	    RECT 406.0000 249.7000 419.6000 250.3000 ;
	    RECT 406.0000 249.6000 406.8000 249.7000 ;
	    RECT 418.8000 249.6000 419.6000 249.7000 ;
	    RECT 420.4000 250.3000 421.2000 250.4000 ;
	    RECT 430.0000 250.3000 430.8000 250.4000 ;
	    RECT 441.2000 250.3000 442.0000 250.4000 ;
	    RECT 457.2000 250.3000 458.0000 250.4000 ;
	    RECT 420.4000 249.7000 458.0000 250.3000 ;
	    RECT 420.4000 249.6000 421.2000 249.7000 ;
	    RECT 430.0000 249.6000 430.8000 249.7000 ;
	    RECT 441.2000 249.6000 442.0000 249.7000 ;
	    RECT 457.2000 249.6000 458.0000 249.7000 ;
	    RECT 463.6000 250.3000 464.4000 250.4000 ;
	    RECT 474.8000 250.3000 475.6000 250.4000 ;
	    RECT 463.6000 249.7000 475.6000 250.3000 ;
	    RECT 463.6000 249.6000 464.4000 249.7000 ;
	    RECT 474.8000 249.6000 475.6000 249.7000 ;
	    RECT 506.8000 249.6000 507.6000 250.4000 ;
	    RECT 225.2000 248.3000 226.0000 248.4000 ;
	    RECT 188.5000 247.7000 226.0000 248.3000 ;
	    RECT 121.2000 247.6000 122.0000 247.7000 ;
	    RECT 137.2000 247.6000 138.0000 247.7000 ;
	    RECT 150.0000 247.6000 150.8000 247.7000 ;
	    RECT 164.4000 247.6000 165.2000 247.7000 ;
	    RECT 186.8000 247.6000 187.6000 247.7000 ;
	    RECT 225.2000 247.6000 226.0000 247.7000 ;
	    RECT 226.8000 248.3000 227.6000 248.4000 ;
	    RECT 238.0000 248.3000 238.8000 248.4000 ;
	    RECT 226.8000 247.7000 238.8000 248.3000 ;
	    RECT 226.8000 247.6000 227.6000 247.7000 ;
	    RECT 238.0000 247.6000 238.8000 247.7000 ;
	    RECT 239.6000 248.3000 240.4000 248.4000 ;
	    RECT 242.8000 248.3000 243.6000 248.4000 ;
	    RECT 239.6000 247.7000 243.6000 248.3000 ;
	    RECT 239.6000 247.6000 240.4000 247.7000 ;
	    RECT 242.8000 247.6000 243.6000 247.7000 ;
	    RECT 244.4000 247.6000 245.2000 248.4000 ;
	    RECT 246.0000 248.3000 246.8000 248.4000 ;
	    RECT 257.2000 248.3000 258.0000 248.4000 ;
	    RECT 246.0000 247.7000 258.0000 248.3000 ;
	    RECT 246.0000 247.6000 246.8000 247.7000 ;
	    RECT 257.2000 247.6000 258.0000 247.7000 ;
	    RECT 258.8000 248.3000 259.6000 248.4000 ;
	    RECT 265.2000 248.3000 266.0000 248.4000 ;
	    RECT 284.4000 248.3000 285.2000 248.4000 ;
	    RECT 258.8000 247.7000 285.2000 248.3000 ;
	    RECT 258.8000 247.6000 259.6000 247.7000 ;
	    RECT 265.2000 247.6000 266.0000 247.7000 ;
	    RECT 284.4000 247.6000 285.2000 247.7000 ;
	    RECT 286.0000 248.3000 286.8000 248.4000 ;
	    RECT 294.0000 248.3000 294.8000 248.4000 ;
	    RECT 286.0000 247.7000 294.8000 248.3000 ;
	    RECT 286.0000 247.6000 286.8000 247.7000 ;
	    RECT 294.0000 247.6000 294.8000 247.7000 ;
	    RECT 12.4000 246.3000 13.2000 246.4000 ;
	    RECT 30.0000 246.3000 30.8000 246.4000 ;
	    RECT 12.4000 245.7000 30.8000 246.3000 ;
	    RECT 12.4000 245.6000 13.2000 245.7000 ;
	    RECT 30.0000 245.6000 30.8000 245.7000 ;
	    RECT 113.2000 246.3000 114.0000 246.4000 ;
	    RECT 169.2000 246.3000 170.0000 246.4000 ;
	    RECT 172.4000 246.3000 173.2000 246.4000 ;
	    RECT 190.0000 246.3000 190.8000 246.4000 ;
	    RECT 113.2000 245.7000 190.8000 246.3000 ;
	    RECT 113.2000 245.6000 114.0000 245.7000 ;
	    RECT 169.2000 245.6000 170.0000 245.7000 ;
	    RECT 172.4000 245.6000 173.2000 245.7000 ;
	    RECT 190.0000 245.6000 190.8000 245.7000 ;
	    RECT 196.4000 246.3000 197.2000 246.4000 ;
	    RECT 199.6000 246.3000 200.4000 246.4000 ;
	    RECT 196.4000 245.7000 200.4000 246.3000 ;
	    RECT 196.4000 245.6000 197.2000 245.7000 ;
	    RECT 199.6000 245.6000 200.4000 245.7000 ;
	    RECT 202.8000 246.3000 203.6000 246.4000 ;
	    RECT 428.4000 246.3000 429.2000 246.4000 ;
	    RECT 202.8000 245.7000 429.2000 246.3000 ;
	    RECT 202.8000 245.6000 203.6000 245.7000 ;
	    RECT 428.4000 245.6000 429.2000 245.7000 ;
	    RECT 502.0000 246.3000 502.8000 246.4000 ;
	    RECT 505.2000 246.3000 506.0000 246.4000 ;
	    RECT 502.0000 245.7000 506.0000 246.3000 ;
	    RECT 502.0000 245.6000 502.8000 245.7000 ;
	    RECT 505.2000 245.6000 506.0000 245.7000 ;
	    RECT 10.8000 244.3000 11.6000 244.4000 ;
	    RECT 15.6000 244.3000 16.4000 244.4000 ;
	    RECT 10.8000 243.7000 16.4000 244.3000 ;
	    RECT 10.8000 243.6000 11.6000 243.7000 ;
	    RECT 15.6000 243.6000 16.4000 243.7000 ;
	    RECT 86.0000 244.3000 86.8000 244.4000 ;
	    RECT 153.2000 244.3000 154.0000 244.4000 ;
	    RECT 86.0000 243.7000 154.0000 244.3000 ;
	    RECT 86.0000 243.6000 86.8000 243.7000 ;
	    RECT 153.2000 243.6000 154.0000 243.7000 ;
	    RECT 164.4000 244.3000 165.2000 244.4000 ;
	    RECT 177.2000 244.3000 178.0000 244.4000 ;
	    RECT 182.0000 244.3000 182.8000 244.4000 ;
	    RECT 164.4000 243.7000 182.8000 244.3000 ;
	    RECT 164.4000 243.6000 165.2000 243.7000 ;
	    RECT 177.2000 243.6000 178.0000 243.7000 ;
	    RECT 182.0000 243.6000 182.8000 243.7000 ;
	    RECT 186.8000 244.3000 187.6000 244.4000 ;
	    RECT 201.2000 244.3000 202.0000 244.4000 ;
	    RECT 186.8000 243.7000 202.0000 244.3000 ;
	    RECT 186.8000 243.6000 187.6000 243.7000 ;
	    RECT 201.2000 243.6000 202.0000 243.7000 ;
	    RECT 218.8000 244.3000 219.6000 244.4000 ;
	    RECT 222.0000 244.3000 222.8000 244.4000 ;
	    RECT 218.8000 243.7000 222.8000 244.3000 ;
	    RECT 218.8000 243.6000 219.6000 243.7000 ;
	    RECT 222.0000 243.6000 222.8000 243.7000 ;
	    RECT 223.6000 244.3000 224.4000 244.4000 ;
	    RECT 231.6000 244.3000 232.4000 244.4000 ;
	    RECT 223.6000 243.7000 232.4000 244.3000 ;
	    RECT 223.6000 243.6000 224.4000 243.7000 ;
	    RECT 231.6000 243.6000 232.4000 243.7000 ;
	    RECT 244.4000 244.3000 245.2000 244.4000 ;
	    RECT 249.2000 244.3000 250.0000 244.4000 ;
	    RECT 244.4000 243.7000 250.0000 244.3000 ;
	    RECT 244.4000 243.6000 245.2000 243.7000 ;
	    RECT 249.2000 243.6000 250.0000 243.7000 ;
	    RECT 252.4000 244.3000 253.2000 244.4000 ;
	    RECT 263.6000 244.3000 264.4000 244.4000 ;
	    RECT 252.4000 243.7000 264.4000 244.3000 ;
	    RECT 252.4000 243.6000 253.2000 243.7000 ;
	    RECT 263.6000 243.6000 264.4000 243.7000 ;
	    RECT 265.2000 244.3000 266.0000 244.4000 ;
	    RECT 271.6000 244.3000 272.4000 244.4000 ;
	    RECT 265.2000 243.7000 272.4000 244.3000 ;
	    RECT 265.2000 243.6000 266.0000 243.7000 ;
	    RECT 271.6000 243.6000 272.4000 243.7000 ;
	    RECT 276.4000 244.3000 277.2000 244.4000 ;
	    RECT 310.0000 244.3000 310.8000 244.4000 ;
	    RECT 276.4000 243.7000 310.8000 244.3000 ;
	    RECT 276.4000 243.6000 277.2000 243.7000 ;
	    RECT 310.0000 243.6000 310.8000 243.7000 ;
	    RECT 346.8000 244.3000 347.6000 244.4000 ;
	    RECT 380.4000 244.3000 381.2000 244.4000 ;
	    RECT 346.8000 243.7000 381.2000 244.3000 ;
	    RECT 346.8000 243.6000 347.6000 243.7000 ;
	    RECT 380.4000 243.6000 381.2000 243.7000 ;
	    RECT 390.0000 244.3000 390.8000 244.4000 ;
	    RECT 433.2000 244.3000 434.0000 244.4000 ;
	    RECT 390.0000 243.7000 434.0000 244.3000 ;
	    RECT 390.0000 243.6000 390.8000 243.7000 ;
	    RECT 433.2000 243.6000 434.0000 243.7000 ;
	    RECT 442.8000 244.3000 443.6000 244.4000 ;
	    RECT 481.2000 244.3000 482.0000 244.4000 ;
	    RECT 442.8000 243.7000 482.0000 244.3000 ;
	    RECT 442.8000 243.6000 443.6000 243.7000 ;
	    RECT 481.2000 243.6000 482.0000 243.7000 ;
	    RECT 487.6000 244.3000 488.4000 244.4000 ;
	    RECT 490.8000 244.3000 491.6000 244.4000 ;
	    RECT 487.6000 243.7000 491.6000 244.3000 ;
	    RECT 487.6000 243.6000 488.4000 243.7000 ;
	    RECT 490.8000 243.6000 491.6000 243.7000 ;
	    RECT 130.8000 242.3000 131.6000 242.4000 ;
	    RECT 137.2000 242.3000 138.0000 242.4000 ;
	    RECT 130.8000 241.7000 138.0000 242.3000 ;
	    RECT 130.8000 241.6000 131.6000 241.7000 ;
	    RECT 137.2000 241.6000 138.0000 241.7000 ;
	    RECT 145.2000 241.6000 146.0000 242.4000 ;
	    RECT 158.0000 242.3000 158.8000 242.4000 ;
	    RECT 202.8000 242.3000 203.6000 242.4000 ;
	    RECT 158.0000 241.7000 203.6000 242.3000 ;
	    RECT 158.0000 241.6000 158.8000 241.7000 ;
	    RECT 202.8000 241.6000 203.6000 241.7000 ;
	    RECT 206.0000 242.3000 206.8000 242.4000 ;
	    RECT 231.6000 242.3000 232.4000 242.4000 ;
	    RECT 206.0000 241.7000 232.4000 242.3000 ;
	    RECT 206.0000 241.6000 206.8000 241.7000 ;
	    RECT 231.6000 241.6000 232.4000 241.7000 ;
	    RECT 284.4000 242.3000 285.2000 242.4000 ;
	    RECT 302.0000 242.3000 302.8000 242.4000 ;
	    RECT 284.4000 241.7000 302.8000 242.3000 ;
	    RECT 284.4000 241.6000 285.2000 241.7000 ;
	    RECT 302.0000 241.6000 302.8000 241.7000 ;
	    RECT 305.2000 242.3000 306.0000 242.4000 ;
	    RECT 382.0000 242.3000 382.8000 242.4000 ;
	    RECT 305.2000 241.7000 382.8000 242.3000 ;
	    RECT 305.2000 241.6000 306.0000 241.7000 ;
	    RECT 382.0000 241.6000 382.8000 241.7000 ;
	    RECT 412.4000 242.3000 413.2000 242.4000 ;
	    RECT 425.2000 242.3000 426.0000 242.4000 ;
	    RECT 412.4000 241.7000 426.0000 242.3000 ;
	    RECT 412.4000 241.6000 413.2000 241.7000 ;
	    RECT 425.2000 241.6000 426.0000 241.7000 ;
	    RECT 111.6000 240.3000 112.4000 240.4000 ;
	    RECT 209.2000 240.3000 210.0000 240.4000 ;
	    RECT 111.6000 239.7000 210.0000 240.3000 ;
	    RECT 111.6000 239.6000 112.4000 239.7000 ;
	    RECT 209.2000 239.6000 210.0000 239.7000 ;
	    RECT 222.0000 240.3000 222.8000 240.4000 ;
	    RECT 289.2000 240.3000 290.0000 240.4000 ;
	    RECT 342.0000 240.3000 342.8000 240.4000 ;
	    RECT 346.8000 240.3000 347.6000 240.4000 ;
	    RECT 222.0000 239.7000 347.6000 240.3000 ;
	    RECT 222.0000 239.6000 222.8000 239.7000 ;
	    RECT 289.2000 239.6000 290.0000 239.7000 ;
	    RECT 342.0000 239.6000 342.8000 239.7000 ;
	    RECT 346.8000 239.6000 347.6000 239.7000 ;
	    RECT 356.4000 240.3000 357.2000 240.4000 ;
	    RECT 382.0000 240.3000 382.8000 240.4000 ;
	    RECT 356.4000 239.7000 382.8000 240.3000 ;
	    RECT 356.4000 239.6000 357.2000 239.7000 ;
	    RECT 382.0000 239.6000 382.8000 239.7000 ;
	    RECT 98.8000 238.3000 99.6000 238.4000 ;
	    RECT 161.2000 238.3000 162.0000 238.4000 ;
	    RECT 303.6000 238.3000 304.4000 238.4000 ;
	    RECT 345.2000 238.3000 346.0000 238.4000 ;
	    RECT 412.4000 238.3000 413.2000 238.4000 ;
	    RECT 98.8000 237.7000 413.2000 238.3000 ;
	    RECT 98.8000 237.6000 99.6000 237.7000 ;
	    RECT 161.2000 237.6000 162.0000 237.7000 ;
	    RECT 303.6000 237.6000 304.4000 237.7000 ;
	    RECT 345.2000 237.6000 346.0000 237.7000 ;
	    RECT 412.4000 237.6000 413.2000 237.7000 ;
	    RECT 414.0000 238.3000 414.8000 238.4000 ;
	    RECT 494.0000 238.3000 494.8000 238.4000 ;
	    RECT 414.0000 237.7000 494.8000 238.3000 ;
	    RECT 414.0000 237.6000 414.8000 237.7000 ;
	    RECT 494.0000 237.6000 494.8000 237.7000 ;
	    RECT 503.6000 238.3000 504.4000 238.4000 ;
	    RECT 508.4000 238.3000 509.2000 238.4000 ;
	    RECT 503.6000 237.7000 509.2000 238.3000 ;
	    RECT 503.6000 237.6000 504.4000 237.7000 ;
	    RECT 508.4000 237.6000 509.2000 237.7000 ;
	    RECT 10.8000 236.3000 11.6000 236.4000 ;
	    RECT 47.6000 236.3000 48.4000 236.4000 ;
	    RECT 62.0000 236.3000 62.8000 236.4000 ;
	    RECT 10.8000 235.7000 62.8000 236.3000 ;
	    RECT 10.8000 235.6000 11.6000 235.7000 ;
	    RECT 47.6000 235.6000 48.4000 235.7000 ;
	    RECT 62.0000 235.6000 62.8000 235.7000 ;
	    RECT 135.6000 236.3000 136.4000 236.4000 ;
	    RECT 193.2000 236.3000 194.0000 236.4000 ;
	    RECT 135.6000 235.7000 194.0000 236.3000 ;
	    RECT 135.6000 235.6000 136.4000 235.7000 ;
	    RECT 193.2000 235.6000 194.0000 235.7000 ;
	    RECT 194.8000 236.3000 195.6000 236.4000 ;
	    RECT 215.6000 236.3000 216.4000 236.4000 ;
	    RECT 194.8000 235.7000 216.4000 236.3000 ;
	    RECT 194.8000 235.6000 195.6000 235.7000 ;
	    RECT 215.6000 235.6000 216.4000 235.7000 ;
	    RECT 217.2000 236.3000 218.0000 236.4000 ;
	    RECT 234.8000 236.3000 235.6000 236.4000 ;
	    RECT 217.2000 235.7000 235.6000 236.3000 ;
	    RECT 217.2000 235.6000 218.0000 235.7000 ;
	    RECT 234.8000 235.6000 235.6000 235.7000 ;
	    RECT 238.0000 236.3000 238.8000 236.4000 ;
	    RECT 249.2000 236.3000 250.0000 236.4000 ;
	    RECT 250.8000 236.3000 251.6000 236.4000 ;
	    RECT 458.8000 236.3000 459.6000 236.4000 ;
	    RECT 238.0000 235.7000 251.6000 236.3000 ;
	    RECT 238.0000 235.6000 238.8000 235.7000 ;
	    RECT 249.2000 235.6000 250.0000 235.7000 ;
	    RECT 250.8000 235.6000 251.6000 235.7000 ;
	    RECT 252.5000 235.7000 459.6000 236.3000 ;
	    RECT 18.8000 234.3000 19.6000 234.4000 ;
	    RECT 49.2000 234.3000 50.0000 234.4000 ;
	    RECT 18.8000 233.7000 50.0000 234.3000 ;
	    RECT 18.8000 233.6000 19.6000 233.7000 ;
	    RECT 49.2000 233.6000 50.0000 233.7000 ;
	    RECT 60.4000 234.3000 61.2000 234.4000 ;
	    RECT 151.6000 234.3000 152.4000 234.4000 ;
	    RECT 252.5000 234.3000 253.1000 235.7000 ;
	    RECT 458.8000 235.6000 459.6000 235.7000 ;
	    RECT 489.2000 236.3000 490.0000 236.4000 ;
	    RECT 495.6000 236.3000 496.4000 236.4000 ;
	    RECT 489.2000 235.7000 496.4000 236.3000 ;
	    RECT 489.2000 235.6000 490.0000 235.7000 ;
	    RECT 495.6000 235.6000 496.4000 235.7000 ;
	    RECT 60.4000 233.7000 139.5000 234.3000 ;
	    RECT 60.4000 233.6000 61.2000 233.7000 ;
	    RECT 4.4000 232.3000 5.2000 232.4000 ;
	    RECT 22.0000 232.3000 22.8000 232.4000 ;
	    RECT 4.4000 231.7000 22.8000 232.3000 ;
	    RECT 4.4000 231.6000 5.2000 231.7000 ;
	    RECT 22.0000 231.6000 22.8000 231.7000 ;
	    RECT 36.4000 232.3000 37.2000 232.4000 ;
	    RECT 46.0000 232.3000 46.8000 232.4000 ;
	    RECT 36.4000 231.7000 46.8000 232.3000 ;
	    RECT 36.4000 231.6000 37.2000 231.7000 ;
	    RECT 46.0000 231.6000 46.8000 231.7000 ;
	    RECT 90.8000 232.3000 91.6000 232.4000 ;
	    RECT 122.8000 232.3000 123.6000 232.4000 ;
	    RECT 90.8000 231.7000 123.6000 232.3000 ;
	    RECT 90.8000 231.6000 91.6000 231.7000 ;
	    RECT 122.8000 231.6000 123.6000 231.7000 ;
	    RECT 124.4000 232.3000 125.2000 232.4000 ;
	    RECT 137.2000 232.3000 138.0000 232.4000 ;
	    RECT 124.4000 231.7000 138.0000 232.3000 ;
	    RECT 138.9000 232.3000 139.5000 233.7000 ;
	    RECT 151.6000 233.7000 253.1000 234.3000 ;
	    RECT 254.0000 234.3000 254.8000 234.4000 ;
	    RECT 276.4000 234.3000 277.2000 234.4000 ;
	    RECT 254.0000 233.7000 277.2000 234.3000 ;
	    RECT 151.6000 233.6000 152.4000 233.7000 ;
	    RECT 254.0000 233.6000 254.8000 233.7000 ;
	    RECT 276.4000 233.6000 277.2000 233.7000 ;
	    RECT 282.8000 234.3000 283.6000 234.4000 ;
	    RECT 305.2000 234.3000 306.0000 234.4000 ;
	    RECT 282.8000 233.7000 306.0000 234.3000 ;
	    RECT 282.8000 233.6000 283.6000 233.7000 ;
	    RECT 305.2000 233.6000 306.0000 233.7000 ;
	    RECT 308.4000 234.3000 309.2000 234.4000 ;
	    RECT 318.0000 234.3000 318.8000 234.4000 ;
	    RECT 414.0000 234.3000 414.8000 234.4000 ;
	    RECT 308.4000 233.7000 414.8000 234.3000 ;
	    RECT 308.4000 233.6000 309.2000 233.7000 ;
	    RECT 318.0000 233.6000 318.8000 233.7000 ;
	    RECT 414.0000 233.6000 414.8000 233.7000 ;
	    RECT 436.4000 234.3000 437.2000 234.4000 ;
	    RECT 441.2000 234.3000 442.0000 234.4000 ;
	    RECT 481.2000 234.3000 482.0000 234.4000 ;
	    RECT 436.4000 233.7000 482.0000 234.3000 ;
	    RECT 436.4000 233.6000 437.2000 233.7000 ;
	    RECT 441.2000 233.6000 442.0000 233.7000 ;
	    RECT 481.2000 233.6000 482.0000 233.7000 ;
	    RECT 494.0000 234.3000 494.8000 234.4000 ;
	    RECT 513.2000 234.3000 514.0000 234.4000 ;
	    RECT 494.0000 233.7000 514.0000 234.3000 ;
	    RECT 494.0000 233.6000 494.8000 233.7000 ;
	    RECT 513.2000 233.6000 514.0000 233.7000 ;
	    RECT 194.8000 232.3000 195.6000 232.4000 ;
	    RECT 250.8000 232.3000 251.6000 232.4000 ;
	    RECT 138.9000 231.7000 195.6000 232.3000 ;
	    RECT 124.4000 231.6000 125.2000 231.7000 ;
	    RECT 137.2000 231.6000 138.0000 231.7000 ;
	    RECT 194.8000 231.6000 195.6000 231.7000 ;
	    RECT 212.5000 231.7000 251.6000 232.3000 ;
	    RECT 212.5000 230.4000 213.1000 231.7000 ;
	    RECT 250.8000 231.6000 251.6000 231.7000 ;
	    RECT 254.0000 232.3000 254.8000 232.4000 ;
	    RECT 266.8000 232.3000 267.6000 232.4000 ;
	    RECT 268.4000 232.3000 269.2000 232.4000 ;
	    RECT 274.8000 232.3000 275.6000 232.4000 ;
	    RECT 254.0000 231.7000 265.9000 232.3000 ;
	    RECT 254.0000 231.6000 254.8000 231.7000 ;
	    RECT 12.4000 230.3000 13.2000 230.4000 ;
	    RECT 14.0000 230.3000 14.8000 230.4000 ;
	    RECT 18.8000 230.3000 19.6000 230.4000 ;
	    RECT 12.4000 229.7000 19.6000 230.3000 ;
	    RECT 12.4000 229.6000 13.2000 229.7000 ;
	    RECT 14.0000 229.6000 14.8000 229.7000 ;
	    RECT 18.8000 229.6000 19.6000 229.7000 ;
	    RECT 31.6000 230.3000 32.4000 230.4000 ;
	    RECT 68.4000 230.3000 69.2000 230.4000 ;
	    RECT 31.6000 229.7000 69.2000 230.3000 ;
	    RECT 31.6000 229.6000 32.4000 229.7000 ;
	    RECT 68.4000 229.6000 69.2000 229.7000 ;
	    RECT 74.8000 230.3000 75.6000 230.4000 ;
	    RECT 82.8000 230.3000 83.6000 230.4000 ;
	    RECT 74.8000 229.7000 83.6000 230.3000 ;
	    RECT 74.8000 229.6000 75.6000 229.7000 ;
	    RECT 82.8000 229.6000 83.6000 229.7000 ;
	    RECT 95.6000 230.3000 96.4000 230.4000 ;
	    RECT 111.6000 230.3000 112.4000 230.4000 ;
	    RECT 95.6000 229.7000 112.4000 230.3000 ;
	    RECT 95.6000 229.6000 96.4000 229.7000 ;
	    RECT 111.6000 229.6000 112.4000 229.7000 ;
	    RECT 126.0000 230.3000 126.8000 230.4000 ;
	    RECT 134.0000 230.3000 134.8000 230.4000 ;
	    RECT 126.0000 229.7000 134.8000 230.3000 ;
	    RECT 126.0000 229.6000 126.8000 229.7000 ;
	    RECT 134.0000 229.6000 134.8000 229.7000 ;
	    RECT 135.6000 230.3000 136.4000 230.4000 ;
	    RECT 142.0000 230.3000 142.8000 230.4000 ;
	    RECT 148.4000 230.3000 149.2000 230.4000 ;
	    RECT 135.6000 229.7000 149.2000 230.3000 ;
	    RECT 135.6000 229.6000 136.4000 229.7000 ;
	    RECT 142.0000 229.6000 142.8000 229.7000 ;
	    RECT 148.4000 229.6000 149.2000 229.7000 ;
	    RECT 159.6000 230.3000 160.4000 230.4000 ;
	    RECT 167.6000 230.3000 168.4000 230.4000 ;
	    RECT 159.6000 229.7000 168.4000 230.3000 ;
	    RECT 159.6000 229.6000 160.4000 229.7000 ;
	    RECT 167.6000 229.6000 168.4000 229.7000 ;
	    RECT 177.2000 229.6000 178.0000 230.4000 ;
	    RECT 178.8000 230.3000 179.6000 230.4000 ;
	    RECT 196.4000 230.3000 197.2000 230.4000 ;
	    RECT 178.8000 229.7000 197.2000 230.3000 ;
	    RECT 178.8000 229.6000 179.6000 229.7000 ;
	    RECT 196.4000 229.6000 197.2000 229.7000 ;
	    RECT 202.8000 230.3000 203.6000 230.4000 ;
	    RECT 210.8000 230.3000 211.6000 230.4000 ;
	    RECT 202.8000 229.7000 211.6000 230.3000 ;
	    RECT 202.8000 229.6000 203.6000 229.7000 ;
	    RECT 210.8000 229.6000 211.6000 229.7000 ;
	    RECT 212.4000 229.6000 213.2000 230.4000 ;
	    RECT 215.6000 230.3000 216.4000 230.4000 ;
	    RECT 218.8000 230.3000 219.6000 230.4000 ;
	    RECT 215.6000 229.7000 219.6000 230.3000 ;
	    RECT 215.6000 229.6000 216.4000 229.7000 ;
	    RECT 218.8000 229.6000 219.6000 229.7000 ;
	    RECT 220.4000 230.3000 221.2000 230.4000 ;
	    RECT 223.6000 230.3000 224.4000 230.4000 ;
	    RECT 228.4000 230.3000 229.2000 230.4000 ;
	    RECT 220.4000 229.7000 229.2000 230.3000 ;
	    RECT 220.4000 229.6000 221.2000 229.7000 ;
	    RECT 223.6000 229.6000 224.4000 229.7000 ;
	    RECT 228.4000 229.6000 229.2000 229.7000 ;
	    RECT 236.4000 230.3000 237.2000 230.4000 ;
	    RECT 263.6000 230.3000 264.4000 230.4000 ;
	    RECT 236.4000 229.7000 264.4000 230.3000 ;
	    RECT 265.3000 230.3000 265.9000 231.7000 ;
	    RECT 266.8000 231.7000 269.2000 232.3000 ;
	    RECT 266.8000 231.6000 267.6000 231.7000 ;
	    RECT 268.4000 231.6000 269.2000 231.7000 ;
	    RECT 270.1000 231.7000 275.6000 232.3000 ;
	    RECT 270.1000 230.3000 270.7000 231.7000 ;
	    RECT 274.8000 231.6000 275.6000 231.7000 ;
	    RECT 281.2000 232.3000 282.0000 232.4000 ;
	    RECT 282.8000 232.3000 283.6000 232.4000 ;
	    RECT 281.2000 231.7000 283.6000 232.3000 ;
	    RECT 281.2000 231.6000 282.0000 231.7000 ;
	    RECT 282.8000 231.6000 283.6000 231.7000 ;
	    RECT 284.4000 232.3000 285.2000 232.4000 ;
	    RECT 292.4000 232.3000 293.2000 232.4000 ;
	    RECT 284.4000 231.7000 293.2000 232.3000 ;
	    RECT 284.4000 231.6000 285.2000 231.7000 ;
	    RECT 292.4000 231.6000 293.2000 231.7000 ;
	    RECT 298.8000 232.3000 299.6000 232.4000 ;
	    RECT 366.0000 232.3000 366.8000 232.4000 ;
	    RECT 298.8000 231.7000 366.8000 232.3000 ;
	    RECT 298.8000 231.6000 299.6000 231.7000 ;
	    RECT 366.0000 231.6000 366.8000 231.7000 ;
	    RECT 375.6000 232.3000 376.4000 232.4000 ;
	    RECT 386.8000 232.3000 387.6000 232.4000 ;
	    RECT 375.6000 231.7000 387.6000 232.3000 ;
	    RECT 375.6000 231.6000 376.4000 231.7000 ;
	    RECT 386.8000 231.6000 387.6000 231.7000 ;
	    RECT 399.6000 232.3000 400.4000 232.4000 ;
	    RECT 402.8000 232.3000 403.6000 232.4000 ;
	    RECT 404.4000 232.3000 405.2000 232.4000 ;
	    RECT 399.6000 231.7000 405.2000 232.3000 ;
	    RECT 399.6000 231.6000 400.4000 231.7000 ;
	    RECT 402.8000 231.6000 403.6000 231.7000 ;
	    RECT 404.4000 231.6000 405.2000 231.7000 ;
	    RECT 449.2000 232.3000 450.0000 232.4000 ;
	    RECT 452.4000 232.3000 453.2000 232.4000 ;
	    RECT 449.2000 231.7000 453.2000 232.3000 ;
	    RECT 449.2000 231.6000 450.0000 231.7000 ;
	    RECT 452.4000 231.6000 453.2000 231.7000 ;
	    RECT 482.8000 232.3000 483.6000 232.4000 ;
	    RECT 486.0000 232.3000 486.8000 232.4000 ;
	    RECT 482.8000 231.7000 486.8000 232.3000 ;
	    RECT 482.8000 231.6000 483.6000 231.7000 ;
	    RECT 486.0000 231.6000 486.8000 231.7000 ;
	    RECT 265.3000 229.7000 270.7000 230.3000 ;
	    RECT 271.6000 230.3000 272.4000 230.4000 ;
	    RECT 279.6000 230.3000 280.4000 230.4000 ;
	    RECT 324.4000 230.3000 325.2000 230.4000 ;
	    RECT 271.6000 229.7000 280.4000 230.3000 ;
	    RECT 236.4000 229.6000 237.2000 229.7000 ;
	    RECT 263.6000 229.6000 264.4000 229.7000 ;
	    RECT 271.6000 229.6000 272.4000 229.7000 ;
	    RECT 279.6000 229.6000 280.4000 229.7000 ;
	    RECT 281.3000 229.7000 325.2000 230.3000 ;
	    RECT 10.8000 228.3000 11.6000 228.4000 ;
	    RECT 17.2000 228.3000 18.0000 228.4000 ;
	    RECT 42.8000 228.3000 43.6000 228.4000 ;
	    RECT 10.8000 227.7000 43.6000 228.3000 ;
	    RECT 10.8000 227.6000 11.6000 227.7000 ;
	    RECT 17.2000 227.6000 18.0000 227.7000 ;
	    RECT 42.8000 227.6000 43.6000 227.7000 ;
	    RECT 47.6000 228.3000 48.4000 228.4000 ;
	    RECT 81.2000 228.3000 82.0000 228.4000 ;
	    RECT 47.6000 227.7000 82.0000 228.3000 ;
	    RECT 47.6000 227.6000 48.4000 227.7000 ;
	    RECT 81.2000 227.6000 82.0000 227.7000 ;
	    RECT 92.4000 228.3000 93.2000 228.4000 ;
	    RECT 94.0000 228.3000 94.8000 228.4000 ;
	    RECT 92.4000 227.7000 94.8000 228.3000 ;
	    RECT 92.4000 227.6000 93.2000 227.7000 ;
	    RECT 94.0000 227.6000 94.8000 227.7000 ;
	    RECT 114.8000 228.3000 115.6000 228.4000 ;
	    RECT 166.0000 228.3000 166.8000 228.4000 ;
	    RECT 114.8000 227.7000 166.8000 228.3000 ;
	    RECT 114.8000 227.6000 115.6000 227.7000 ;
	    RECT 166.0000 227.6000 166.8000 227.7000 ;
	    RECT 170.8000 228.3000 171.6000 228.4000 ;
	    RECT 175.6000 228.3000 176.4000 228.4000 ;
	    RECT 170.8000 227.7000 176.4000 228.3000 ;
	    RECT 170.8000 227.6000 171.6000 227.7000 ;
	    RECT 175.6000 227.6000 176.4000 227.7000 ;
	    RECT 177.2000 228.3000 178.0000 228.4000 ;
	    RECT 186.8000 228.3000 187.6000 228.4000 ;
	    RECT 177.2000 227.7000 187.6000 228.3000 ;
	    RECT 177.2000 227.6000 178.0000 227.7000 ;
	    RECT 186.8000 227.6000 187.6000 227.7000 ;
	    RECT 190.0000 228.3000 190.8000 228.4000 ;
	    RECT 201.2000 228.3000 202.0000 228.4000 ;
	    RECT 190.0000 227.7000 202.0000 228.3000 ;
	    RECT 190.0000 227.6000 190.8000 227.7000 ;
	    RECT 201.2000 227.6000 202.0000 227.7000 ;
	    RECT 206.0000 228.3000 206.8000 228.4000 ;
	    RECT 214.0000 228.3000 214.8000 228.4000 ;
	    RECT 206.0000 227.7000 214.8000 228.3000 ;
	    RECT 218.9000 228.3000 219.5000 229.6000 ;
	    RECT 281.3000 228.4000 281.9000 229.7000 ;
	    RECT 324.4000 229.6000 325.2000 229.7000 ;
	    RECT 337.2000 230.3000 338.0000 230.4000 ;
	    RECT 348.4000 230.3000 349.2000 230.4000 ;
	    RECT 337.2000 229.7000 349.2000 230.3000 ;
	    RECT 337.2000 229.6000 338.0000 229.7000 ;
	    RECT 348.4000 229.6000 349.2000 229.7000 ;
	    RECT 386.8000 230.3000 387.6000 230.4000 ;
	    RECT 391.6000 230.3000 392.4000 230.4000 ;
	    RECT 386.8000 229.7000 392.4000 230.3000 ;
	    RECT 386.8000 229.6000 387.6000 229.7000 ;
	    RECT 391.6000 229.6000 392.4000 229.7000 ;
	    RECT 402.8000 230.3000 403.6000 230.4000 ;
	    RECT 425.2000 230.3000 426.0000 230.4000 ;
	    RECT 402.8000 229.7000 426.0000 230.3000 ;
	    RECT 402.8000 229.6000 403.6000 229.7000 ;
	    RECT 425.2000 229.6000 426.0000 229.7000 ;
	    RECT 441.2000 230.3000 442.0000 230.4000 ;
	    RECT 450.8000 230.3000 451.6000 230.4000 ;
	    RECT 441.2000 229.7000 451.6000 230.3000 ;
	    RECT 441.2000 229.6000 442.0000 229.7000 ;
	    RECT 450.8000 229.6000 451.6000 229.7000 ;
	    RECT 474.8000 230.3000 475.6000 230.4000 ;
	    RECT 482.8000 230.3000 483.6000 230.4000 ;
	    RECT 474.8000 229.7000 483.6000 230.3000 ;
	    RECT 474.8000 229.6000 475.6000 229.7000 ;
	    RECT 482.8000 229.6000 483.6000 229.7000 ;
	    RECT 486.0000 230.3000 486.8000 230.4000 ;
	    RECT 500.4000 230.3000 501.2000 230.4000 ;
	    RECT 486.0000 229.7000 501.2000 230.3000 ;
	    RECT 486.0000 229.6000 486.8000 229.7000 ;
	    RECT 500.4000 229.6000 501.2000 229.7000 ;
	    RECT 226.8000 228.3000 227.6000 228.4000 ;
	    RECT 230.0000 228.3000 230.8000 228.4000 ;
	    RECT 249.2000 228.3000 250.0000 228.4000 ;
	    RECT 218.9000 227.7000 227.6000 228.3000 ;
	    RECT 206.0000 227.6000 206.8000 227.7000 ;
	    RECT 214.0000 227.6000 214.8000 227.7000 ;
	    RECT 226.8000 227.6000 227.6000 227.7000 ;
	    RECT 228.5000 227.7000 230.8000 228.3000 ;
	    RECT 68.4000 226.3000 69.2000 226.4000 ;
	    RECT 74.8000 226.3000 75.6000 226.4000 ;
	    RECT 87.6000 226.3000 88.4000 226.4000 ;
	    RECT 68.4000 225.7000 88.4000 226.3000 ;
	    RECT 68.4000 225.6000 69.2000 225.7000 ;
	    RECT 74.8000 225.6000 75.6000 225.7000 ;
	    RECT 87.6000 225.6000 88.4000 225.7000 ;
	    RECT 92.4000 226.3000 93.2000 226.4000 ;
	    RECT 124.4000 226.3000 125.2000 226.4000 ;
	    RECT 92.4000 225.7000 125.2000 226.3000 ;
	    RECT 92.4000 225.6000 93.2000 225.7000 ;
	    RECT 124.4000 225.6000 125.2000 225.7000 ;
	    RECT 142.0000 226.3000 142.8000 226.4000 ;
	    RECT 151.6000 226.3000 152.4000 226.4000 ;
	    RECT 142.0000 225.7000 152.4000 226.3000 ;
	    RECT 142.0000 225.6000 142.8000 225.7000 ;
	    RECT 151.6000 225.6000 152.4000 225.7000 ;
	    RECT 166.0000 226.3000 166.8000 226.4000 ;
	    RECT 178.8000 226.3000 179.6000 226.4000 ;
	    RECT 166.0000 225.7000 179.6000 226.3000 ;
	    RECT 166.0000 225.6000 166.8000 225.7000 ;
	    RECT 178.8000 225.6000 179.6000 225.7000 ;
	    RECT 190.0000 226.3000 190.8000 226.4000 ;
	    RECT 196.4000 226.3000 197.2000 226.4000 ;
	    RECT 190.0000 225.7000 197.2000 226.3000 ;
	    RECT 190.0000 225.6000 190.8000 225.7000 ;
	    RECT 196.4000 225.6000 197.2000 225.7000 ;
	    RECT 198.0000 226.3000 198.8000 226.4000 ;
	    RECT 202.8000 226.3000 203.6000 226.4000 ;
	    RECT 228.5000 226.3000 229.1000 227.7000 ;
	    RECT 230.0000 227.6000 230.8000 227.7000 ;
	    RECT 231.7000 227.7000 250.0000 228.3000 ;
	    RECT 198.0000 225.7000 229.1000 226.3000 ;
	    RECT 230.0000 226.3000 230.8000 226.4000 ;
	    RECT 231.7000 226.3000 232.3000 227.7000 ;
	    RECT 249.2000 227.6000 250.0000 227.7000 ;
	    RECT 260.4000 228.3000 261.2000 228.4000 ;
	    RECT 266.8000 228.3000 267.6000 228.4000 ;
	    RECT 260.4000 227.7000 267.6000 228.3000 ;
	    RECT 260.4000 227.6000 261.2000 227.7000 ;
	    RECT 266.8000 227.6000 267.6000 227.7000 ;
	    RECT 274.8000 228.3000 275.6000 228.4000 ;
	    RECT 276.4000 228.3000 277.2000 228.4000 ;
	    RECT 274.8000 227.7000 277.2000 228.3000 ;
	    RECT 274.8000 227.6000 275.6000 227.7000 ;
	    RECT 276.4000 227.6000 277.2000 227.7000 ;
	    RECT 281.2000 227.6000 282.0000 228.4000 ;
	    RECT 282.8000 228.3000 283.6000 228.4000 ;
	    RECT 302.0000 228.3000 302.8000 228.4000 ;
	    RECT 282.8000 227.7000 302.8000 228.3000 ;
	    RECT 282.8000 227.6000 283.6000 227.7000 ;
	    RECT 302.0000 227.6000 302.8000 227.7000 ;
	    RECT 303.6000 228.3000 304.4000 228.4000 ;
	    RECT 313.2000 228.3000 314.0000 228.4000 ;
	    RECT 396.4000 228.3000 397.2000 228.4000 ;
	    RECT 303.6000 227.7000 397.2000 228.3000 ;
	    RECT 303.6000 227.6000 304.4000 227.7000 ;
	    RECT 313.2000 227.6000 314.0000 227.7000 ;
	    RECT 396.4000 227.6000 397.2000 227.7000 ;
	    RECT 436.4000 228.3000 437.2000 228.4000 ;
	    RECT 474.9000 228.3000 475.5000 229.6000 ;
	    RECT 436.4000 227.7000 475.5000 228.3000 ;
	    RECT 476.4000 228.3000 477.2000 228.4000 ;
	    RECT 497.2000 228.3000 498.0000 228.4000 ;
	    RECT 476.4000 227.7000 498.0000 228.3000 ;
	    RECT 436.4000 227.6000 437.2000 227.7000 ;
	    RECT 476.4000 227.6000 477.2000 227.7000 ;
	    RECT 497.2000 227.6000 498.0000 227.7000 ;
	    RECT 230.0000 225.7000 232.3000 226.3000 ;
	    RECT 198.0000 225.6000 198.8000 225.7000 ;
	    RECT 202.8000 225.6000 203.6000 225.7000 ;
	    RECT 230.0000 225.6000 230.8000 225.7000 ;
	    RECT 234.8000 225.6000 235.6000 226.4000 ;
	    RECT 244.4000 226.3000 245.2000 226.4000 ;
	    RECT 247.6000 226.3000 248.4000 226.4000 ;
	    RECT 244.4000 225.7000 248.4000 226.3000 ;
	    RECT 244.4000 225.6000 245.2000 225.7000 ;
	    RECT 247.6000 225.6000 248.4000 225.7000 ;
	    RECT 249.2000 226.3000 250.0000 226.4000 ;
	    RECT 254.0000 226.3000 254.8000 226.4000 ;
	    RECT 249.2000 225.7000 254.8000 226.3000 ;
	    RECT 249.2000 225.6000 250.0000 225.7000 ;
	    RECT 254.0000 225.6000 254.8000 225.7000 ;
	    RECT 265.2000 226.3000 266.0000 226.4000 ;
	    RECT 274.8000 226.3000 275.6000 226.4000 ;
	    RECT 265.2000 225.7000 275.6000 226.3000 ;
	    RECT 265.2000 225.6000 266.0000 225.7000 ;
	    RECT 274.8000 225.6000 275.6000 225.7000 ;
	    RECT 278.0000 226.3000 278.8000 226.4000 ;
	    RECT 294.0000 226.3000 294.8000 226.4000 ;
	    RECT 326.0000 226.3000 326.8000 226.4000 ;
	    RECT 351.6000 226.3000 352.4000 226.4000 ;
	    RECT 278.0000 225.7000 352.4000 226.3000 ;
	    RECT 278.0000 225.6000 278.8000 225.7000 ;
	    RECT 294.0000 225.6000 294.8000 225.7000 ;
	    RECT 326.0000 225.6000 326.8000 225.7000 ;
	    RECT 351.6000 225.6000 352.4000 225.7000 ;
	    RECT 396.4000 226.3000 397.2000 226.4000 ;
	    RECT 414.0000 226.3000 414.8000 226.4000 ;
	    RECT 396.4000 225.7000 414.8000 226.3000 ;
	    RECT 396.4000 225.6000 397.2000 225.7000 ;
	    RECT 414.0000 225.6000 414.8000 225.7000 ;
	    RECT 450.8000 226.3000 451.6000 226.4000 ;
	    RECT 471.6000 226.3000 472.4000 226.4000 ;
	    RECT 450.8000 225.7000 472.4000 226.3000 ;
	    RECT 450.8000 225.6000 451.6000 225.7000 ;
	    RECT 471.6000 225.6000 472.4000 225.7000 ;
	    RECT 62.0000 224.3000 62.8000 224.4000 ;
	    RECT 167.6000 224.3000 168.4000 224.4000 ;
	    RECT 62.0000 223.7000 168.4000 224.3000 ;
	    RECT 62.0000 223.6000 62.8000 223.7000 ;
	    RECT 167.6000 223.6000 168.4000 223.7000 ;
	    RECT 177.2000 224.3000 178.0000 224.4000 ;
	    RECT 225.2000 224.3000 226.0000 224.4000 ;
	    RECT 177.2000 223.7000 226.0000 224.3000 ;
	    RECT 177.2000 223.6000 178.0000 223.7000 ;
	    RECT 225.2000 223.6000 226.0000 223.7000 ;
	    RECT 231.6000 224.3000 232.4000 224.4000 ;
	    RECT 246.0000 224.3000 246.8000 224.4000 ;
	    RECT 231.6000 223.7000 246.8000 224.3000 ;
	    RECT 231.6000 223.6000 232.4000 223.7000 ;
	    RECT 246.0000 223.6000 246.8000 223.7000 ;
	    RECT 250.8000 224.3000 251.6000 224.4000 ;
	    RECT 270.0000 224.3000 270.8000 224.4000 ;
	    RECT 250.8000 223.7000 270.8000 224.3000 ;
	    RECT 250.8000 223.6000 251.6000 223.7000 ;
	    RECT 270.0000 223.6000 270.8000 223.7000 ;
	    RECT 286.0000 223.6000 286.8000 224.4000 ;
	    RECT 287.6000 224.3000 288.4000 224.4000 ;
	    RECT 314.8000 224.3000 315.6000 224.4000 ;
	    RECT 287.6000 223.7000 315.6000 224.3000 ;
	    RECT 287.6000 223.6000 288.4000 223.7000 ;
	    RECT 314.8000 223.6000 315.6000 223.7000 ;
	    RECT 316.4000 224.3000 317.2000 224.4000 ;
	    RECT 322.8000 224.3000 323.6000 224.4000 ;
	    RECT 362.8000 224.3000 363.6000 224.4000 ;
	    RECT 382.0000 224.3000 382.8000 224.4000 ;
	    RECT 316.4000 223.7000 382.8000 224.3000 ;
	    RECT 316.4000 223.6000 317.2000 223.7000 ;
	    RECT 322.8000 223.6000 323.6000 223.7000 ;
	    RECT 362.8000 223.6000 363.6000 223.7000 ;
	    RECT 382.0000 223.6000 382.8000 223.7000 ;
	    RECT 396.4000 224.3000 397.2000 224.4000 ;
	    RECT 439.6000 224.3000 440.4000 224.4000 ;
	    RECT 396.4000 223.7000 440.4000 224.3000 ;
	    RECT 396.4000 223.6000 397.2000 223.7000 ;
	    RECT 439.6000 223.6000 440.4000 223.7000 ;
	    RECT 490.8000 224.3000 491.6000 224.4000 ;
	    RECT 494.0000 224.3000 494.8000 224.4000 ;
	    RECT 490.8000 223.7000 494.8000 224.3000 ;
	    RECT 490.8000 223.6000 491.6000 223.7000 ;
	    RECT 494.0000 223.6000 494.8000 223.7000 ;
	    RECT 84.4000 222.3000 85.2000 222.4000 ;
	    RECT 97.2000 222.3000 98.0000 222.4000 ;
	    RECT 154.8000 222.3000 155.6000 222.4000 ;
	    RECT 215.6000 222.3000 216.4000 222.4000 ;
	    RECT 220.4000 222.3000 221.2000 222.4000 ;
	    RECT 239.6000 222.3000 240.4000 222.4000 ;
	    RECT 84.4000 221.7000 240.4000 222.3000 ;
	    RECT 84.4000 221.6000 85.2000 221.7000 ;
	    RECT 97.2000 221.6000 98.0000 221.7000 ;
	    RECT 154.8000 221.6000 155.6000 221.7000 ;
	    RECT 215.6000 221.6000 216.4000 221.7000 ;
	    RECT 220.4000 221.6000 221.2000 221.7000 ;
	    RECT 239.6000 221.6000 240.4000 221.7000 ;
	    RECT 242.8000 222.3000 243.6000 222.4000 ;
	    RECT 252.4000 222.3000 253.2000 222.4000 ;
	    RECT 242.8000 221.7000 253.2000 222.3000 ;
	    RECT 242.8000 221.6000 243.6000 221.7000 ;
	    RECT 252.4000 221.6000 253.2000 221.7000 ;
	    RECT 262.0000 222.3000 262.8000 222.4000 ;
	    RECT 282.8000 222.3000 283.6000 222.4000 ;
	    RECT 262.0000 221.7000 283.6000 222.3000 ;
	    RECT 262.0000 221.6000 262.8000 221.7000 ;
	    RECT 282.8000 221.6000 283.6000 221.7000 ;
	    RECT 287.6000 222.3000 288.4000 222.4000 ;
	    RECT 289.2000 222.3000 290.0000 222.4000 ;
	    RECT 287.6000 221.7000 290.0000 222.3000 ;
	    RECT 287.6000 221.6000 288.4000 221.7000 ;
	    RECT 289.2000 221.6000 290.0000 221.7000 ;
	    RECT 290.8000 222.3000 291.6000 222.4000 ;
	    RECT 350.0000 222.3000 350.8000 222.4000 ;
	    RECT 290.8000 221.7000 350.8000 222.3000 ;
	    RECT 290.8000 221.6000 291.6000 221.7000 ;
	    RECT 350.0000 221.6000 350.8000 221.7000 ;
	    RECT 361.2000 222.3000 362.0000 222.4000 ;
	    RECT 490.9000 222.3000 491.5000 223.6000 ;
	    RECT 361.2000 221.7000 491.5000 222.3000 ;
	    RECT 361.2000 221.6000 362.0000 221.7000 ;
	    RECT 119.6000 220.3000 120.4000 220.4000 ;
	    RECT 146.8000 220.3000 147.6000 220.4000 ;
	    RECT 119.6000 219.7000 147.6000 220.3000 ;
	    RECT 119.6000 219.6000 120.4000 219.7000 ;
	    RECT 146.8000 219.6000 147.6000 219.7000 ;
	    RECT 151.6000 219.6000 152.4000 220.4000 ;
	    RECT 178.8000 220.3000 179.6000 220.4000 ;
	    RECT 185.2000 220.3000 186.0000 220.4000 ;
	    RECT 178.8000 219.7000 186.0000 220.3000 ;
	    RECT 178.8000 219.6000 179.6000 219.7000 ;
	    RECT 185.2000 219.6000 186.0000 219.7000 ;
	    RECT 186.8000 219.6000 187.6000 220.4000 ;
	    RECT 188.4000 220.3000 189.2000 220.4000 ;
	    RECT 209.2000 220.3000 210.0000 220.4000 ;
	    RECT 188.4000 219.7000 210.0000 220.3000 ;
	    RECT 188.4000 219.6000 189.2000 219.7000 ;
	    RECT 209.2000 219.6000 210.0000 219.7000 ;
	    RECT 212.4000 220.3000 213.2000 220.4000 ;
	    RECT 217.2000 220.3000 218.0000 220.4000 ;
	    RECT 212.4000 219.7000 218.0000 220.3000 ;
	    RECT 212.4000 219.6000 213.2000 219.7000 ;
	    RECT 217.2000 219.6000 218.0000 219.7000 ;
	    RECT 218.8000 220.3000 219.6000 220.4000 ;
	    RECT 222.0000 220.3000 222.8000 220.4000 ;
	    RECT 231.6000 220.3000 232.4000 220.4000 ;
	    RECT 218.8000 219.7000 222.8000 220.3000 ;
	    RECT 218.8000 219.6000 219.6000 219.7000 ;
	    RECT 222.0000 219.6000 222.8000 219.7000 ;
	    RECT 223.7000 219.7000 232.4000 220.3000 ;
	    RECT 90.8000 218.3000 91.6000 218.4000 ;
	    RECT 97.2000 218.3000 98.0000 218.4000 ;
	    RECT 159.6000 218.3000 160.4000 218.4000 ;
	    RECT 162.8000 218.3000 163.6000 218.4000 ;
	    RECT 90.8000 217.7000 163.6000 218.3000 ;
	    RECT 90.8000 217.6000 91.6000 217.7000 ;
	    RECT 97.2000 217.6000 98.0000 217.7000 ;
	    RECT 159.6000 217.6000 160.4000 217.7000 ;
	    RECT 162.8000 217.6000 163.6000 217.7000 ;
	    RECT 164.4000 218.3000 165.2000 218.4000 ;
	    RECT 207.6000 218.3000 208.4000 218.4000 ;
	    RECT 164.4000 217.7000 208.4000 218.3000 ;
	    RECT 164.4000 217.6000 165.2000 217.7000 ;
	    RECT 207.6000 217.6000 208.4000 217.7000 ;
	    RECT 209.2000 218.3000 210.0000 218.4000 ;
	    RECT 223.7000 218.3000 224.3000 219.7000 ;
	    RECT 231.6000 219.6000 232.4000 219.7000 ;
	    RECT 233.2000 220.3000 234.0000 220.4000 ;
	    RECT 241.2000 220.3000 242.0000 220.4000 ;
	    RECT 233.2000 219.7000 242.0000 220.3000 ;
	    RECT 233.2000 219.6000 234.0000 219.7000 ;
	    RECT 241.2000 219.6000 242.0000 219.7000 ;
	    RECT 244.4000 220.3000 245.2000 220.4000 ;
	    RECT 247.6000 220.3000 248.4000 220.4000 ;
	    RECT 249.2000 220.3000 250.0000 220.4000 ;
	    RECT 244.4000 219.7000 250.0000 220.3000 ;
	    RECT 244.4000 219.6000 245.2000 219.7000 ;
	    RECT 247.6000 219.6000 248.4000 219.7000 ;
	    RECT 249.2000 219.6000 250.0000 219.7000 ;
	    RECT 263.6000 220.3000 264.4000 220.4000 ;
	    RECT 289.2000 220.3000 290.0000 220.4000 ;
	    RECT 263.6000 219.7000 290.0000 220.3000 ;
	    RECT 263.6000 219.6000 264.4000 219.7000 ;
	    RECT 289.2000 219.6000 290.0000 219.7000 ;
	    RECT 308.4000 220.3000 309.2000 220.4000 ;
	    RECT 334.0000 220.3000 334.8000 220.4000 ;
	    RECT 359.6000 220.3000 360.4000 220.4000 ;
	    RECT 308.4000 219.7000 360.4000 220.3000 ;
	    RECT 308.4000 219.6000 309.2000 219.7000 ;
	    RECT 334.0000 219.6000 334.8000 219.7000 ;
	    RECT 359.6000 219.6000 360.4000 219.7000 ;
	    RECT 364.4000 220.3000 365.2000 220.4000 ;
	    RECT 383.6000 220.3000 384.4000 220.4000 ;
	    RECT 492.4000 220.3000 493.2000 220.4000 ;
	    RECT 364.4000 219.7000 384.4000 220.3000 ;
	    RECT 364.4000 219.6000 365.2000 219.7000 ;
	    RECT 383.6000 219.6000 384.4000 219.7000 ;
	    RECT 385.3000 219.7000 493.2000 220.3000 ;
	    RECT 209.2000 217.7000 224.3000 218.3000 ;
	    RECT 225.2000 218.3000 226.0000 218.4000 ;
	    RECT 385.3000 218.3000 385.9000 219.7000 ;
	    RECT 492.4000 219.6000 493.2000 219.7000 ;
	    RECT 225.2000 217.7000 385.9000 218.3000 ;
	    RECT 399.6000 218.3000 400.4000 218.4000 ;
	    RECT 417.2000 218.3000 418.0000 218.4000 ;
	    RECT 399.6000 217.7000 418.0000 218.3000 ;
	    RECT 209.2000 217.6000 210.0000 217.7000 ;
	    RECT 225.2000 217.6000 226.0000 217.7000 ;
	    RECT 399.6000 217.6000 400.4000 217.7000 ;
	    RECT 417.2000 217.6000 418.0000 217.7000 ;
	    RECT 39.6000 216.3000 40.4000 216.4000 ;
	    RECT 47.6000 216.3000 48.4000 216.4000 ;
	    RECT 39.6000 215.7000 48.4000 216.3000 ;
	    RECT 39.6000 215.6000 40.4000 215.7000 ;
	    RECT 47.6000 215.6000 48.4000 215.7000 ;
	    RECT 52.4000 216.3000 53.2000 216.4000 ;
	    RECT 62.0000 216.3000 62.8000 216.4000 ;
	    RECT 52.4000 215.7000 62.8000 216.3000 ;
	    RECT 52.4000 215.6000 53.2000 215.7000 ;
	    RECT 62.0000 215.6000 62.8000 215.7000 ;
	    RECT 105.2000 216.3000 106.0000 216.4000 ;
	    RECT 119.6000 216.3000 120.4000 216.4000 ;
	    RECT 105.2000 215.7000 120.4000 216.3000 ;
	    RECT 105.2000 215.6000 106.0000 215.7000 ;
	    RECT 119.6000 215.6000 120.4000 215.7000 ;
	    RECT 154.8000 216.3000 155.6000 216.4000 ;
	    RECT 183.6000 216.3000 184.4000 216.4000 ;
	    RECT 154.8000 215.7000 184.4000 216.3000 ;
	    RECT 154.8000 215.6000 155.6000 215.7000 ;
	    RECT 183.6000 215.6000 184.4000 215.7000 ;
	    RECT 185.2000 216.3000 186.0000 216.4000 ;
	    RECT 190.0000 216.3000 190.8000 216.4000 ;
	    RECT 185.2000 215.7000 190.8000 216.3000 ;
	    RECT 185.2000 215.6000 186.0000 215.7000 ;
	    RECT 190.0000 215.6000 190.8000 215.7000 ;
	    RECT 193.2000 216.3000 194.0000 216.4000 ;
	    RECT 202.8000 216.3000 203.6000 216.4000 ;
	    RECT 193.2000 215.7000 203.6000 216.3000 ;
	    RECT 193.2000 215.6000 194.0000 215.7000 ;
	    RECT 202.8000 215.6000 203.6000 215.7000 ;
	    RECT 206.0000 216.3000 206.8000 216.4000 ;
	    RECT 207.6000 216.3000 208.4000 216.4000 ;
	    RECT 206.0000 215.7000 208.4000 216.3000 ;
	    RECT 206.0000 215.6000 206.8000 215.7000 ;
	    RECT 207.6000 215.6000 208.4000 215.7000 ;
	    RECT 228.4000 215.6000 229.2000 216.4000 ;
	    RECT 238.0000 216.3000 238.8000 216.4000 ;
	    RECT 230.1000 215.7000 238.8000 216.3000 ;
	    RECT 41.2000 214.3000 42.0000 214.4000 ;
	    RECT 57.2000 214.3000 58.0000 214.4000 ;
	    RECT 41.2000 213.7000 58.0000 214.3000 ;
	    RECT 41.2000 213.6000 42.0000 213.7000 ;
	    RECT 57.2000 213.6000 58.0000 213.7000 ;
	    RECT 62.0000 213.6000 62.8000 214.4000 ;
	    RECT 81.2000 214.3000 82.0000 214.4000 ;
	    RECT 100.4000 214.3000 101.2000 214.4000 ;
	    RECT 81.2000 213.7000 101.2000 214.3000 ;
	    RECT 81.2000 213.6000 82.0000 213.7000 ;
	    RECT 100.4000 213.6000 101.2000 213.7000 ;
	    RECT 111.6000 214.3000 112.4000 214.4000 ;
	    RECT 130.8000 214.3000 131.6000 214.4000 ;
	    RECT 156.4000 214.3000 157.2000 214.4000 ;
	    RECT 169.2000 214.3000 170.0000 214.4000 ;
	    RECT 111.6000 213.7000 170.0000 214.3000 ;
	    RECT 111.6000 213.6000 112.4000 213.7000 ;
	    RECT 130.8000 213.6000 131.6000 213.7000 ;
	    RECT 156.4000 213.6000 157.2000 213.7000 ;
	    RECT 169.2000 213.6000 170.0000 213.7000 ;
	    RECT 174.0000 214.3000 174.8000 214.4000 ;
	    RECT 199.6000 214.3000 200.4000 214.4000 ;
	    RECT 174.0000 213.7000 200.4000 214.3000 ;
	    RECT 174.0000 213.6000 174.8000 213.7000 ;
	    RECT 199.6000 213.6000 200.4000 213.7000 ;
	    RECT 206.0000 214.3000 206.8000 214.4000 ;
	    RECT 222.0000 214.3000 222.8000 214.4000 ;
	    RECT 206.0000 213.7000 222.8000 214.3000 ;
	    RECT 206.0000 213.6000 206.8000 213.7000 ;
	    RECT 222.0000 213.6000 222.8000 213.7000 ;
	    RECT 225.2000 214.3000 226.0000 214.4000 ;
	    RECT 230.1000 214.3000 230.7000 215.7000 ;
	    RECT 238.0000 215.6000 238.8000 215.7000 ;
	    RECT 249.2000 216.3000 250.0000 216.4000 ;
	    RECT 265.2000 216.3000 266.0000 216.4000 ;
	    RECT 278.0000 216.3000 278.8000 216.4000 ;
	    RECT 289.2000 216.3000 290.0000 216.4000 ;
	    RECT 308.4000 216.3000 309.2000 216.4000 ;
	    RECT 249.2000 215.7000 290.0000 216.3000 ;
	    RECT 249.2000 215.6000 250.0000 215.7000 ;
	    RECT 265.2000 215.6000 266.0000 215.7000 ;
	    RECT 278.0000 215.6000 278.8000 215.7000 ;
	    RECT 289.2000 215.6000 290.0000 215.7000 ;
	    RECT 295.7000 215.7000 309.2000 216.3000 ;
	    RECT 225.2000 213.7000 230.7000 214.3000 ;
	    RECT 234.8000 214.3000 235.6000 214.4000 ;
	    RECT 250.8000 214.3000 251.6000 214.4000 ;
	    RECT 234.8000 213.7000 251.6000 214.3000 ;
	    RECT 225.2000 213.6000 226.0000 213.7000 ;
	    RECT 234.8000 213.6000 235.6000 213.7000 ;
	    RECT 250.8000 213.6000 251.6000 213.7000 ;
	    RECT 252.4000 214.3000 253.2000 214.4000 ;
	    RECT 266.8000 214.3000 267.6000 214.4000 ;
	    RECT 271.6000 214.3000 272.4000 214.4000 ;
	    RECT 281.2000 214.3000 282.0000 214.4000 ;
	    RECT 252.4000 213.7000 265.9000 214.3000 ;
	    RECT 252.4000 213.6000 253.2000 213.7000 ;
	    RECT 4.4000 212.3000 5.2000 212.4000 ;
	    RECT 15.6000 212.3000 16.4000 212.4000 ;
	    RECT 4.4000 211.7000 16.4000 212.3000 ;
	    RECT 4.4000 211.6000 5.2000 211.7000 ;
	    RECT 15.6000 211.6000 16.4000 211.7000 ;
	    RECT 30.0000 212.3000 30.8000 212.4000 ;
	    RECT 36.4000 212.3000 37.2000 212.4000 ;
	    RECT 30.0000 211.7000 37.2000 212.3000 ;
	    RECT 30.0000 211.6000 30.8000 211.7000 ;
	    RECT 36.4000 211.6000 37.2000 211.7000 ;
	    RECT 41.2000 212.3000 42.0000 212.4000 ;
	    RECT 71.6000 212.3000 72.4000 212.4000 ;
	    RECT 41.2000 211.7000 72.4000 212.3000 ;
	    RECT 41.2000 211.6000 42.0000 211.7000 ;
	    RECT 71.6000 211.6000 72.4000 211.7000 ;
	    RECT 92.4000 212.3000 93.2000 212.4000 ;
	    RECT 94.0000 212.3000 94.8000 212.4000 ;
	    RECT 92.4000 211.7000 94.8000 212.3000 ;
	    RECT 92.4000 211.6000 93.2000 211.7000 ;
	    RECT 94.0000 211.6000 94.8000 211.7000 ;
	    RECT 121.2000 212.3000 122.0000 212.4000 ;
	    RECT 126.0000 212.3000 126.8000 212.4000 ;
	    RECT 135.6000 212.3000 136.4000 212.4000 ;
	    RECT 121.2000 211.7000 136.4000 212.3000 ;
	    RECT 121.2000 211.6000 122.0000 211.7000 ;
	    RECT 126.0000 211.6000 126.8000 211.7000 ;
	    RECT 135.6000 211.6000 136.4000 211.7000 ;
	    RECT 154.8000 212.3000 155.6000 212.4000 ;
	    RECT 158.0000 212.3000 158.8000 212.4000 ;
	    RECT 154.8000 211.7000 158.8000 212.3000 ;
	    RECT 154.8000 211.6000 155.6000 211.7000 ;
	    RECT 158.0000 211.6000 158.8000 211.7000 ;
	    RECT 218.8000 212.3000 219.6000 212.4000 ;
	    RECT 228.4000 212.3000 229.2000 212.4000 ;
	    RECT 218.8000 211.7000 229.2000 212.3000 ;
	    RECT 218.8000 211.6000 219.6000 211.7000 ;
	    RECT 228.4000 211.6000 229.2000 211.7000 ;
	    RECT 231.6000 212.3000 232.4000 212.4000 ;
	    RECT 263.6000 212.3000 264.4000 212.4000 ;
	    RECT 231.6000 211.7000 264.4000 212.3000 ;
	    RECT 265.3000 212.3000 265.9000 213.7000 ;
	    RECT 266.8000 213.7000 282.0000 214.3000 ;
	    RECT 266.8000 213.6000 267.6000 213.7000 ;
	    RECT 271.6000 213.6000 272.4000 213.7000 ;
	    RECT 281.2000 213.6000 282.0000 213.7000 ;
	    RECT 282.8000 214.3000 283.6000 214.4000 ;
	    RECT 295.7000 214.3000 296.3000 215.7000 ;
	    RECT 308.4000 215.6000 309.2000 215.7000 ;
	    RECT 310.0000 216.3000 310.8000 216.4000 ;
	    RECT 319.6000 216.3000 320.4000 216.4000 ;
	    RECT 364.4000 216.3000 365.2000 216.4000 ;
	    RECT 310.0000 215.7000 365.2000 216.3000 ;
	    RECT 310.0000 215.6000 310.8000 215.7000 ;
	    RECT 319.6000 215.6000 320.4000 215.7000 ;
	    RECT 364.4000 215.6000 365.2000 215.7000 ;
	    RECT 366.0000 216.3000 366.8000 216.4000 ;
	    RECT 393.2000 216.3000 394.0000 216.4000 ;
	    RECT 436.4000 216.3000 437.2000 216.4000 ;
	    RECT 366.0000 215.7000 437.2000 216.3000 ;
	    RECT 366.0000 215.6000 366.8000 215.7000 ;
	    RECT 393.2000 215.6000 394.0000 215.7000 ;
	    RECT 436.4000 215.6000 437.2000 215.7000 ;
	    RECT 441.2000 216.3000 442.0000 216.4000 ;
	    RECT 458.8000 216.3000 459.6000 216.4000 ;
	    RECT 484.4000 216.3000 485.2000 216.4000 ;
	    RECT 441.2000 215.7000 485.2000 216.3000 ;
	    RECT 441.2000 215.6000 442.0000 215.7000 ;
	    RECT 458.8000 215.6000 459.6000 215.7000 ;
	    RECT 484.4000 215.6000 485.2000 215.7000 ;
	    RECT 282.8000 213.7000 296.3000 214.3000 ;
	    RECT 305.2000 214.3000 306.0000 214.4000 ;
	    RECT 338.8000 214.3000 339.6000 214.4000 ;
	    RECT 305.2000 213.7000 339.6000 214.3000 ;
	    RECT 282.8000 213.6000 283.6000 213.7000 ;
	    RECT 305.2000 213.6000 306.0000 213.7000 ;
	    RECT 338.8000 213.6000 339.6000 213.7000 ;
	    RECT 346.8000 213.6000 347.6000 214.4000 ;
	    RECT 350.0000 214.3000 350.8000 214.4000 ;
	    RECT 412.4000 214.3000 413.2000 214.4000 ;
	    RECT 350.0000 213.7000 413.2000 214.3000 ;
	    RECT 350.0000 213.6000 350.8000 213.7000 ;
	    RECT 412.4000 213.6000 413.2000 213.7000 ;
	    RECT 414.0000 214.3000 414.8000 214.4000 ;
	    RECT 415.6000 214.3000 416.4000 214.4000 ;
	    RECT 414.0000 213.7000 416.4000 214.3000 ;
	    RECT 414.0000 213.6000 414.8000 213.7000 ;
	    RECT 415.6000 213.6000 416.4000 213.7000 ;
	    RECT 442.8000 214.3000 443.6000 214.4000 ;
	    RECT 447.6000 214.3000 448.4000 214.4000 ;
	    RECT 442.8000 213.7000 448.4000 214.3000 ;
	    RECT 442.8000 213.6000 443.6000 213.7000 ;
	    RECT 447.6000 213.6000 448.4000 213.7000 ;
	    RECT 449.2000 214.3000 450.0000 214.4000 ;
	    RECT 450.8000 214.3000 451.6000 214.4000 ;
	    RECT 449.2000 213.7000 451.6000 214.3000 ;
	    RECT 449.2000 213.6000 450.0000 213.7000 ;
	    RECT 450.8000 213.6000 451.6000 213.7000 ;
	    RECT 474.8000 214.3000 475.6000 214.4000 ;
	    RECT 500.4000 214.3000 501.2000 214.4000 ;
	    RECT 474.8000 213.7000 501.2000 214.3000 ;
	    RECT 474.8000 213.6000 475.6000 213.7000 ;
	    RECT 500.4000 213.6000 501.2000 213.7000 ;
	    RECT 270.0000 212.3000 270.8000 212.4000 ;
	    RECT 265.3000 211.7000 270.8000 212.3000 ;
	    RECT 231.6000 211.6000 232.4000 211.7000 ;
	    RECT 263.6000 211.6000 264.4000 211.7000 ;
	    RECT 270.0000 211.6000 270.8000 211.7000 ;
	    RECT 273.2000 212.3000 274.0000 212.4000 ;
	    RECT 386.8000 212.3000 387.6000 212.4000 ;
	    RECT 481.2000 212.3000 482.0000 212.4000 ;
	    RECT 489.2000 212.3000 490.0000 212.4000 ;
	    RECT 273.2000 211.7000 490.0000 212.3000 ;
	    RECT 273.2000 211.6000 274.0000 211.7000 ;
	    RECT 386.8000 211.6000 387.6000 211.7000 ;
	    RECT 481.2000 211.6000 482.0000 211.7000 ;
	    RECT 489.2000 211.6000 490.0000 211.7000 ;
	    RECT 492.4000 212.3000 493.2000 212.4000 ;
	    RECT 505.2000 212.3000 506.0000 212.4000 ;
	    RECT 492.4000 211.7000 506.0000 212.3000 ;
	    RECT 492.4000 211.6000 493.2000 211.7000 ;
	    RECT 505.2000 211.6000 506.0000 211.7000 ;
	    RECT 14.0000 210.3000 14.8000 210.4000 ;
	    RECT 36.4000 210.3000 37.2000 210.4000 ;
	    RECT 14.0000 209.7000 37.2000 210.3000 ;
	    RECT 14.0000 209.6000 14.8000 209.7000 ;
	    RECT 36.4000 209.6000 37.2000 209.7000 ;
	    RECT 100.4000 210.3000 101.2000 210.4000 ;
	    RECT 105.2000 210.3000 106.0000 210.4000 ;
	    RECT 100.4000 209.7000 106.0000 210.3000 ;
	    RECT 100.4000 209.6000 101.2000 209.7000 ;
	    RECT 105.2000 209.6000 106.0000 209.7000 ;
	    RECT 114.8000 210.3000 115.6000 210.4000 ;
	    RECT 122.8000 210.3000 123.6000 210.4000 ;
	    RECT 114.8000 209.7000 123.6000 210.3000 ;
	    RECT 114.8000 209.6000 115.6000 209.7000 ;
	    RECT 122.8000 209.6000 123.6000 209.7000 ;
	    RECT 137.2000 210.3000 138.0000 210.4000 ;
	    RECT 148.4000 210.3000 149.2000 210.4000 ;
	    RECT 137.2000 209.7000 149.2000 210.3000 ;
	    RECT 137.2000 209.6000 138.0000 209.7000 ;
	    RECT 148.4000 209.6000 149.2000 209.7000 ;
	    RECT 154.8000 210.3000 155.6000 210.4000 ;
	    RECT 162.8000 210.3000 163.6000 210.4000 ;
	    RECT 154.8000 209.7000 163.6000 210.3000 ;
	    RECT 154.8000 209.6000 155.6000 209.7000 ;
	    RECT 162.8000 209.6000 163.6000 209.7000 ;
	    RECT 182.0000 210.3000 182.8000 210.4000 ;
	    RECT 199.6000 210.3000 200.4000 210.4000 ;
	    RECT 238.0000 210.3000 238.8000 210.4000 ;
	    RECT 182.0000 209.7000 238.8000 210.3000 ;
	    RECT 182.0000 209.6000 182.8000 209.7000 ;
	    RECT 199.6000 209.6000 200.4000 209.7000 ;
	    RECT 238.0000 209.6000 238.8000 209.7000 ;
	    RECT 244.4000 210.3000 245.2000 210.4000 ;
	    RECT 284.4000 210.3000 285.2000 210.4000 ;
	    RECT 244.4000 209.7000 285.2000 210.3000 ;
	    RECT 244.4000 209.6000 245.2000 209.7000 ;
	    RECT 284.4000 209.6000 285.2000 209.7000 ;
	    RECT 286.0000 210.3000 286.8000 210.4000 ;
	    RECT 300.4000 210.3000 301.2000 210.4000 ;
	    RECT 286.0000 209.7000 301.2000 210.3000 ;
	    RECT 286.0000 209.6000 286.8000 209.7000 ;
	    RECT 300.4000 209.6000 301.2000 209.7000 ;
	    RECT 302.0000 210.3000 302.8000 210.4000 ;
	    RECT 310.0000 210.3000 310.8000 210.4000 ;
	    RECT 311.6000 210.3000 312.4000 210.4000 ;
	    RECT 318.0000 210.3000 318.8000 210.4000 ;
	    RECT 302.0000 209.7000 318.8000 210.3000 ;
	    RECT 302.0000 209.6000 302.8000 209.7000 ;
	    RECT 310.0000 209.6000 310.8000 209.7000 ;
	    RECT 311.6000 209.6000 312.4000 209.7000 ;
	    RECT 318.0000 209.6000 318.8000 209.7000 ;
	    RECT 340.4000 210.3000 341.2000 210.4000 ;
	    RECT 348.4000 210.3000 349.2000 210.4000 ;
	    RECT 340.4000 209.7000 349.2000 210.3000 ;
	    RECT 340.4000 209.6000 341.2000 209.7000 ;
	    RECT 348.4000 209.6000 349.2000 209.7000 ;
	    RECT 377.2000 210.3000 378.0000 210.4000 ;
	    RECT 388.4000 210.3000 389.2000 210.4000 ;
	    RECT 377.2000 209.7000 389.2000 210.3000 ;
	    RECT 377.2000 209.6000 378.0000 209.7000 ;
	    RECT 388.4000 209.6000 389.2000 209.7000 ;
	    RECT 394.8000 210.3000 395.6000 210.4000 ;
	    RECT 396.4000 210.3000 397.2000 210.4000 ;
	    RECT 394.8000 209.7000 397.2000 210.3000 ;
	    RECT 394.8000 209.6000 395.6000 209.7000 ;
	    RECT 396.4000 209.6000 397.2000 209.7000 ;
	    RECT 414.0000 210.3000 414.8000 210.4000 ;
	    RECT 428.4000 210.3000 429.2000 210.4000 ;
	    RECT 414.0000 209.7000 429.2000 210.3000 ;
	    RECT 414.0000 209.6000 414.8000 209.7000 ;
	    RECT 428.4000 209.6000 429.2000 209.7000 ;
	    RECT 471.6000 210.3000 472.4000 210.4000 ;
	    RECT 479.6000 210.3000 480.4000 210.4000 ;
	    RECT 471.6000 209.7000 480.4000 210.3000 ;
	    RECT 471.6000 209.6000 472.4000 209.7000 ;
	    RECT 479.6000 209.6000 480.4000 209.7000 ;
	    RECT 50.8000 208.3000 51.6000 208.4000 ;
	    RECT 118.0000 208.3000 118.8000 208.4000 ;
	    RECT 50.8000 207.7000 118.8000 208.3000 ;
	    RECT 50.8000 207.6000 51.6000 207.7000 ;
	    RECT 118.0000 207.6000 118.8000 207.7000 ;
	    RECT 146.8000 208.3000 147.6000 208.4000 ;
	    RECT 158.0000 208.3000 158.8000 208.4000 ;
	    RECT 183.6000 208.3000 184.4000 208.4000 ;
	    RECT 146.8000 207.7000 184.4000 208.3000 ;
	    RECT 146.8000 207.6000 147.6000 207.7000 ;
	    RECT 158.0000 207.6000 158.8000 207.7000 ;
	    RECT 183.6000 207.6000 184.4000 207.7000 ;
	    RECT 185.2000 208.3000 186.0000 208.4000 ;
	    RECT 188.4000 208.3000 189.2000 208.4000 ;
	    RECT 185.2000 207.7000 189.2000 208.3000 ;
	    RECT 185.2000 207.6000 186.0000 207.7000 ;
	    RECT 188.4000 207.6000 189.2000 207.7000 ;
	    RECT 233.2000 208.3000 234.0000 208.4000 ;
	    RECT 241.2000 208.3000 242.0000 208.4000 ;
	    RECT 233.2000 207.7000 242.0000 208.3000 ;
	    RECT 233.2000 207.6000 234.0000 207.7000 ;
	    RECT 241.2000 207.6000 242.0000 207.7000 ;
	    RECT 242.8000 208.3000 243.6000 208.4000 ;
	    RECT 247.6000 208.3000 248.4000 208.4000 ;
	    RECT 242.8000 207.7000 248.4000 208.3000 ;
	    RECT 242.8000 207.6000 243.6000 207.7000 ;
	    RECT 247.6000 207.6000 248.4000 207.7000 ;
	    RECT 249.2000 208.3000 250.0000 208.4000 ;
	    RECT 270.0000 208.3000 270.8000 208.4000 ;
	    RECT 321.2000 208.3000 322.0000 208.4000 ;
	    RECT 249.2000 207.7000 269.1000 208.3000 ;
	    RECT 249.2000 207.6000 250.0000 207.7000 ;
	    RECT 62.0000 206.3000 62.8000 206.4000 ;
	    RECT 164.4000 206.3000 165.2000 206.4000 ;
	    RECT 62.0000 205.7000 165.2000 206.3000 ;
	    RECT 62.0000 205.6000 62.8000 205.7000 ;
	    RECT 164.4000 205.6000 165.2000 205.7000 ;
	    RECT 174.0000 206.3000 174.8000 206.4000 ;
	    RECT 220.4000 206.3000 221.2000 206.4000 ;
	    RECT 174.0000 205.7000 221.2000 206.3000 ;
	    RECT 174.0000 205.6000 174.8000 205.7000 ;
	    RECT 220.4000 205.6000 221.2000 205.7000 ;
	    RECT 228.4000 206.3000 229.2000 206.4000 ;
	    RECT 230.0000 206.3000 230.8000 206.4000 ;
	    RECT 228.4000 205.7000 230.8000 206.3000 ;
	    RECT 228.4000 205.6000 229.2000 205.7000 ;
	    RECT 230.0000 205.6000 230.8000 205.7000 ;
	    RECT 231.6000 206.3000 232.4000 206.4000 ;
	    RECT 266.8000 206.3000 267.6000 206.4000 ;
	    RECT 231.6000 205.7000 267.6000 206.3000 ;
	    RECT 268.5000 206.3000 269.1000 207.7000 ;
	    RECT 270.0000 207.7000 322.0000 208.3000 ;
	    RECT 270.0000 207.6000 270.8000 207.7000 ;
	    RECT 321.2000 207.6000 322.0000 207.7000 ;
	    RECT 338.8000 208.3000 339.6000 208.4000 ;
	    RECT 418.8000 208.3000 419.6000 208.4000 ;
	    RECT 430.0000 208.3000 430.8000 208.4000 ;
	    RECT 338.8000 207.7000 430.8000 208.3000 ;
	    RECT 338.8000 207.6000 339.6000 207.7000 ;
	    RECT 418.8000 207.6000 419.6000 207.7000 ;
	    RECT 430.0000 207.6000 430.8000 207.7000 ;
	    RECT 465.2000 208.3000 466.0000 208.4000 ;
	    RECT 478.0000 208.3000 478.8000 208.4000 ;
	    RECT 465.2000 207.7000 478.8000 208.3000 ;
	    RECT 465.2000 207.6000 466.0000 207.7000 ;
	    RECT 478.0000 207.6000 478.8000 207.7000 ;
	    RECT 311.6000 206.3000 312.4000 206.4000 ;
	    RECT 268.5000 205.7000 312.4000 206.3000 ;
	    RECT 231.6000 205.6000 232.4000 205.7000 ;
	    RECT 266.8000 205.6000 267.6000 205.7000 ;
	    RECT 311.6000 205.6000 312.4000 205.7000 ;
	    RECT 327.6000 206.3000 328.4000 206.4000 ;
	    RECT 353.2000 206.3000 354.0000 206.4000 ;
	    RECT 327.6000 205.7000 354.0000 206.3000 ;
	    RECT 327.6000 205.6000 328.4000 205.7000 ;
	    RECT 353.2000 205.6000 354.0000 205.7000 ;
	    RECT 356.4000 205.6000 357.2000 206.4000 ;
	    RECT 402.8000 206.3000 403.6000 206.4000 ;
	    RECT 415.6000 206.3000 416.4000 206.4000 ;
	    RECT 402.8000 205.7000 416.4000 206.3000 ;
	    RECT 402.8000 205.6000 403.6000 205.7000 ;
	    RECT 415.6000 205.6000 416.4000 205.7000 ;
	    RECT 446.0000 206.3000 446.8000 206.4000 ;
	    RECT 457.2000 206.3000 458.0000 206.4000 ;
	    RECT 446.0000 205.7000 458.0000 206.3000 ;
	    RECT 446.0000 205.6000 446.8000 205.7000 ;
	    RECT 457.2000 205.6000 458.0000 205.7000 ;
	    RECT 471.6000 206.3000 472.4000 206.4000 ;
	    RECT 492.4000 206.3000 493.2000 206.4000 ;
	    RECT 471.6000 205.7000 493.2000 206.3000 ;
	    RECT 471.6000 205.6000 472.4000 205.7000 ;
	    RECT 492.4000 205.6000 493.2000 205.7000 ;
	    RECT 14.0000 204.3000 14.8000 204.4000 ;
	    RECT 17.2000 204.3000 18.0000 204.4000 ;
	    RECT 14.0000 203.7000 18.0000 204.3000 ;
	    RECT 14.0000 203.6000 14.8000 203.7000 ;
	    RECT 17.2000 203.6000 18.0000 203.7000 ;
	    RECT 94.0000 204.3000 94.8000 204.4000 ;
	    RECT 106.8000 204.3000 107.6000 204.4000 ;
	    RECT 153.2000 204.3000 154.0000 204.4000 ;
	    RECT 175.6000 204.3000 176.4000 204.4000 ;
	    RECT 193.2000 204.3000 194.0000 204.4000 ;
	    RECT 298.8000 204.3000 299.6000 204.4000 ;
	    RECT 94.0000 203.7000 299.6000 204.3000 ;
	    RECT 94.0000 203.6000 94.8000 203.7000 ;
	    RECT 106.8000 203.6000 107.6000 203.7000 ;
	    RECT 153.2000 203.6000 154.0000 203.7000 ;
	    RECT 175.6000 203.6000 176.4000 203.7000 ;
	    RECT 193.2000 203.6000 194.0000 203.7000 ;
	    RECT 298.8000 203.6000 299.6000 203.7000 ;
	    RECT 302.0000 204.3000 302.8000 204.4000 ;
	    RECT 343.6000 204.3000 344.4000 204.4000 ;
	    RECT 362.8000 204.3000 363.6000 204.4000 ;
	    RECT 394.8000 204.3000 395.6000 204.4000 ;
	    RECT 302.0000 203.7000 395.6000 204.3000 ;
	    RECT 302.0000 203.6000 302.8000 203.7000 ;
	    RECT 343.6000 203.6000 344.4000 203.7000 ;
	    RECT 362.8000 203.6000 363.6000 203.7000 ;
	    RECT 394.8000 203.6000 395.6000 203.7000 ;
	    RECT 148.4000 202.3000 149.2000 202.4000 ;
	    RECT 156.4000 202.3000 157.2000 202.4000 ;
	    RECT 148.4000 201.7000 157.2000 202.3000 ;
	    RECT 148.4000 201.6000 149.2000 201.7000 ;
	    RECT 156.4000 201.6000 157.2000 201.7000 ;
	    RECT 162.8000 202.3000 163.6000 202.4000 ;
	    RECT 188.4000 202.3000 189.2000 202.4000 ;
	    RECT 162.8000 201.7000 189.2000 202.3000 ;
	    RECT 162.8000 201.6000 163.6000 201.7000 ;
	    RECT 188.4000 201.6000 189.2000 201.7000 ;
	    RECT 193.2000 202.3000 194.0000 202.4000 ;
	    RECT 274.8000 202.3000 275.6000 202.4000 ;
	    RECT 282.8000 202.3000 283.6000 202.4000 ;
	    RECT 193.2000 201.7000 275.6000 202.3000 ;
	    RECT 193.2000 201.6000 194.0000 201.7000 ;
	    RECT 274.8000 201.6000 275.6000 201.7000 ;
	    RECT 278.1000 201.7000 283.6000 202.3000 ;
	    RECT 278.1000 200.4000 278.7000 201.7000 ;
	    RECT 282.8000 201.6000 283.6000 201.7000 ;
	    RECT 287.6000 202.3000 288.4000 202.4000 ;
	    RECT 308.4000 202.3000 309.2000 202.4000 ;
	    RECT 287.6000 201.7000 309.2000 202.3000 ;
	    RECT 287.6000 201.6000 288.4000 201.7000 ;
	    RECT 308.4000 201.6000 309.2000 201.7000 ;
	    RECT 356.4000 202.3000 357.2000 202.4000 ;
	    RECT 362.8000 202.3000 363.6000 202.4000 ;
	    RECT 386.8000 202.3000 387.6000 202.4000 ;
	    RECT 391.6000 202.3000 392.4000 202.4000 ;
	    RECT 402.8000 202.3000 403.6000 202.4000 ;
	    RECT 356.4000 201.7000 403.6000 202.3000 ;
	    RECT 356.4000 201.6000 357.2000 201.7000 ;
	    RECT 362.8000 201.6000 363.6000 201.7000 ;
	    RECT 386.8000 201.6000 387.6000 201.7000 ;
	    RECT 391.6000 201.6000 392.4000 201.7000 ;
	    RECT 402.8000 201.6000 403.6000 201.7000 ;
	    RECT 417.2000 202.3000 418.0000 202.4000 ;
	    RECT 446.0000 202.3000 446.8000 202.4000 ;
	    RECT 417.2000 201.7000 446.8000 202.3000 ;
	    RECT 417.2000 201.6000 418.0000 201.7000 ;
	    RECT 446.0000 201.6000 446.8000 201.7000 ;
	    RECT 58.8000 200.3000 59.6000 200.4000 ;
	    RECT 81.2000 200.3000 82.0000 200.4000 ;
	    RECT 191.6000 200.3000 192.4000 200.4000 ;
	    RECT 58.8000 199.7000 82.0000 200.3000 ;
	    RECT 58.8000 199.6000 59.6000 199.7000 ;
	    RECT 81.2000 199.6000 82.0000 199.7000 ;
	    RECT 111.7000 199.7000 192.4000 200.3000 ;
	    RECT 54.0000 198.3000 54.8000 198.4000 ;
	    RECT 111.7000 198.3000 112.3000 199.7000 ;
	    RECT 191.6000 199.6000 192.4000 199.7000 ;
	    RECT 194.8000 200.3000 195.6000 200.4000 ;
	    RECT 196.4000 200.3000 197.2000 200.4000 ;
	    RECT 194.8000 199.7000 197.2000 200.3000 ;
	    RECT 194.8000 199.6000 195.6000 199.7000 ;
	    RECT 196.4000 199.6000 197.2000 199.7000 ;
	    RECT 199.6000 200.3000 200.4000 200.4000 ;
	    RECT 204.4000 200.3000 205.2000 200.4000 ;
	    RECT 206.0000 200.3000 206.8000 200.4000 ;
	    RECT 199.6000 199.7000 206.8000 200.3000 ;
	    RECT 199.6000 199.6000 200.4000 199.7000 ;
	    RECT 204.4000 199.6000 205.2000 199.7000 ;
	    RECT 206.0000 199.6000 206.8000 199.7000 ;
	    RECT 217.2000 200.3000 218.0000 200.4000 ;
	    RECT 222.0000 200.3000 222.8000 200.4000 ;
	    RECT 217.2000 199.7000 222.8000 200.3000 ;
	    RECT 217.2000 199.6000 218.0000 199.7000 ;
	    RECT 222.0000 199.6000 222.8000 199.7000 ;
	    RECT 230.0000 200.3000 230.8000 200.4000 ;
	    RECT 244.4000 200.3000 245.2000 200.4000 ;
	    RECT 230.0000 199.7000 245.2000 200.3000 ;
	    RECT 230.0000 199.6000 230.8000 199.7000 ;
	    RECT 244.4000 199.6000 245.2000 199.7000 ;
	    RECT 247.6000 200.3000 248.4000 200.4000 ;
	    RECT 255.6000 200.3000 256.4000 200.4000 ;
	    RECT 247.6000 199.7000 256.4000 200.3000 ;
	    RECT 247.6000 199.6000 248.4000 199.7000 ;
	    RECT 255.6000 199.6000 256.4000 199.7000 ;
	    RECT 263.6000 200.3000 264.4000 200.4000 ;
	    RECT 271.6000 200.3000 272.4000 200.4000 ;
	    RECT 263.6000 199.7000 272.4000 200.3000 ;
	    RECT 263.6000 199.6000 264.4000 199.7000 ;
	    RECT 271.6000 199.6000 272.4000 199.7000 ;
	    RECT 273.2000 200.3000 274.0000 200.4000 ;
	    RECT 278.0000 200.3000 278.8000 200.4000 ;
	    RECT 273.2000 199.7000 278.8000 200.3000 ;
	    RECT 273.2000 199.6000 274.0000 199.7000 ;
	    RECT 278.0000 199.6000 278.8000 199.7000 ;
	    RECT 281.2000 200.3000 282.0000 200.4000 ;
	    RECT 282.8000 200.3000 283.6000 200.4000 ;
	    RECT 298.8000 200.3000 299.6000 200.4000 ;
	    RECT 281.2000 199.7000 299.6000 200.3000 ;
	    RECT 281.2000 199.6000 282.0000 199.7000 ;
	    RECT 282.8000 199.6000 283.6000 199.7000 ;
	    RECT 298.8000 199.6000 299.6000 199.7000 ;
	    RECT 345.2000 200.3000 346.0000 200.4000 ;
	    RECT 474.8000 200.3000 475.6000 200.4000 ;
	    RECT 345.2000 199.7000 401.9000 200.3000 ;
	    RECT 345.2000 199.6000 346.0000 199.7000 ;
	    RECT 54.0000 197.7000 112.3000 198.3000 ;
	    RECT 113.2000 198.3000 114.0000 198.4000 ;
	    RECT 212.4000 198.3000 213.2000 198.4000 ;
	    RECT 113.2000 197.7000 213.2000 198.3000 ;
	    RECT 54.0000 197.6000 54.8000 197.7000 ;
	    RECT 113.2000 197.6000 114.0000 197.7000 ;
	    RECT 212.4000 197.6000 213.2000 197.7000 ;
	    RECT 214.0000 198.3000 214.8000 198.4000 ;
	    RECT 217.2000 198.3000 218.0000 198.4000 ;
	    RECT 225.2000 198.3000 226.0000 198.4000 ;
	    RECT 241.2000 198.3000 242.0000 198.4000 ;
	    RECT 214.0000 197.7000 221.1000 198.3000 ;
	    RECT 214.0000 197.6000 214.8000 197.7000 ;
	    RECT 217.2000 197.6000 218.0000 197.7000 ;
	    RECT 46.0000 196.3000 46.8000 196.4000 ;
	    RECT 52.4000 196.3000 53.2000 196.4000 ;
	    RECT 55.6000 196.3000 56.4000 196.4000 ;
	    RECT 58.8000 196.3000 59.6000 196.4000 ;
	    RECT 46.0000 195.7000 59.6000 196.3000 ;
	    RECT 46.0000 195.6000 46.8000 195.7000 ;
	    RECT 52.4000 195.6000 53.2000 195.7000 ;
	    RECT 55.6000 195.6000 56.4000 195.7000 ;
	    RECT 58.8000 195.6000 59.6000 195.7000 ;
	    RECT 68.4000 196.3000 69.2000 196.4000 ;
	    RECT 150.0000 196.3000 150.8000 196.4000 ;
	    RECT 68.4000 195.7000 150.8000 196.3000 ;
	    RECT 68.4000 195.6000 69.2000 195.7000 ;
	    RECT 150.0000 195.6000 150.8000 195.7000 ;
	    RECT 170.8000 196.3000 171.6000 196.4000 ;
	    RECT 180.4000 196.3000 181.2000 196.4000 ;
	    RECT 170.8000 195.7000 181.2000 196.3000 ;
	    RECT 170.8000 195.6000 171.6000 195.7000 ;
	    RECT 180.4000 195.6000 181.2000 195.7000 ;
	    RECT 191.6000 196.3000 192.4000 196.4000 ;
	    RECT 198.0000 196.3000 198.8000 196.4000 ;
	    RECT 191.6000 195.7000 198.8000 196.3000 ;
	    RECT 191.6000 195.6000 192.4000 195.7000 ;
	    RECT 198.0000 195.6000 198.8000 195.7000 ;
	    RECT 199.6000 195.6000 200.4000 196.4000 ;
	    RECT 202.8000 196.3000 203.6000 196.4000 ;
	    RECT 206.0000 196.3000 206.8000 196.4000 ;
	    RECT 202.8000 195.7000 206.8000 196.3000 ;
	    RECT 202.8000 195.6000 203.6000 195.7000 ;
	    RECT 206.0000 195.6000 206.8000 195.7000 ;
	    RECT 210.8000 196.3000 211.6000 196.4000 ;
	    RECT 218.8000 196.3000 219.6000 196.4000 ;
	    RECT 210.8000 195.7000 219.6000 196.3000 ;
	    RECT 220.5000 196.3000 221.1000 197.7000 ;
	    RECT 225.2000 197.7000 242.0000 198.3000 ;
	    RECT 225.2000 197.6000 226.0000 197.7000 ;
	    RECT 241.2000 197.6000 242.0000 197.7000 ;
	    RECT 242.8000 198.3000 243.6000 198.4000 ;
	    RECT 250.8000 198.3000 251.6000 198.4000 ;
	    RECT 268.4000 198.3000 269.2000 198.4000 ;
	    RECT 242.8000 197.7000 269.2000 198.3000 ;
	    RECT 242.8000 197.6000 243.6000 197.7000 ;
	    RECT 250.8000 197.6000 251.6000 197.7000 ;
	    RECT 268.4000 197.6000 269.2000 197.7000 ;
	    RECT 270.0000 198.3000 270.8000 198.4000 ;
	    RECT 287.6000 198.3000 288.4000 198.4000 ;
	    RECT 270.0000 197.7000 288.4000 198.3000 ;
	    RECT 270.0000 197.6000 270.8000 197.7000 ;
	    RECT 287.6000 197.6000 288.4000 197.7000 ;
	    RECT 289.2000 198.3000 290.0000 198.4000 ;
	    RECT 303.6000 198.3000 304.4000 198.4000 ;
	    RECT 289.2000 197.7000 304.4000 198.3000 ;
	    RECT 289.2000 197.6000 290.0000 197.7000 ;
	    RECT 303.6000 197.6000 304.4000 197.7000 ;
	    RECT 308.4000 198.3000 309.2000 198.4000 ;
	    RECT 319.6000 198.3000 320.4000 198.4000 ;
	    RECT 308.4000 197.7000 320.4000 198.3000 ;
	    RECT 308.4000 197.6000 309.2000 197.7000 ;
	    RECT 319.6000 197.6000 320.4000 197.7000 ;
	    RECT 326.0000 198.3000 326.8000 198.4000 ;
	    RECT 338.8000 198.3000 339.6000 198.4000 ;
	    RECT 326.0000 197.7000 339.6000 198.3000 ;
	    RECT 326.0000 197.6000 326.8000 197.7000 ;
	    RECT 338.8000 197.6000 339.6000 197.7000 ;
	    RECT 351.6000 198.3000 352.4000 198.4000 ;
	    RECT 358.0000 198.3000 358.8000 198.4000 ;
	    RECT 351.6000 197.7000 358.8000 198.3000 ;
	    RECT 351.6000 197.6000 352.4000 197.7000 ;
	    RECT 358.0000 197.6000 358.8000 197.7000 ;
	    RECT 367.6000 198.3000 368.4000 198.4000 ;
	    RECT 399.6000 198.3000 400.4000 198.4000 ;
	    RECT 367.6000 197.7000 400.4000 198.3000 ;
	    RECT 401.3000 198.3000 401.9000 199.7000 ;
	    RECT 412.5000 199.7000 475.6000 200.3000 ;
	    RECT 412.5000 198.3000 413.1000 199.7000 ;
	    RECT 474.8000 199.6000 475.6000 199.7000 ;
	    RECT 401.3000 197.7000 413.1000 198.3000 ;
	    RECT 414.0000 198.3000 414.8000 198.4000 ;
	    RECT 431.6000 198.3000 432.4000 198.4000 ;
	    RECT 439.6000 198.3000 440.4000 198.4000 ;
	    RECT 414.0000 197.7000 440.4000 198.3000 ;
	    RECT 367.6000 197.6000 368.4000 197.7000 ;
	    RECT 399.6000 197.6000 400.4000 197.7000 ;
	    RECT 414.0000 197.6000 414.8000 197.7000 ;
	    RECT 431.6000 197.6000 432.4000 197.7000 ;
	    RECT 439.6000 197.6000 440.4000 197.7000 ;
	    RECT 225.2000 196.3000 226.0000 196.4000 ;
	    RECT 231.6000 196.3000 232.4000 196.4000 ;
	    RECT 220.5000 195.7000 232.4000 196.3000 ;
	    RECT 210.8000 195.6000 211.6000 195.7000 ;
	    RECT 218.8000 195.6000 219.6000 195.7000 ;
	    RECT 225.2000 195.6000 226.0000 195.7000 ;
	    RECT 231.6000 195.6000 232.4000 195.7000 ;
	    RECT 238.0000 196.3000 238.8000 196.4000 ;
	    RECT 252.4000 196.3000 253.2000 196.4000 ;
	    RECT 276.4000 196.3000 277.2000 196.4000 ;
	    RECT 238.0000 195.7000 277.2000 196.3000 ;
	    RECT 238.0000 195.6000 238.8000 195.7000 ;
	    RECT 252.4000 195.6000 253.2000 195.7000 ;
	    RECT 276.4000 195.6000 277.2000 195.7000 ;
	    RECT 284.4000 196.3000 285.2000 196.4000 ;
	    RECT 359.6000 196.3000 360.4000 196.4000 ;
	    RECT 284.4000 195.7000 360.4000 196.3000 ;
	    RECT 284.4000 195.6000 285.2000 195.7000 ;
	    RECT 359.6000 195.6000 360.4000 195.7000 ;
	    RECT 394.8000 196.3000 395.6000 196.4000 ;
	    RECT 423.6000 196.3000 424.4000 196.4000 ;
	    RECT 438.0000 196.3000 438.8000 196.4000 ;
	    RECT 394.8000 195.7000 438.8000 196.3000 ;
	    RECT 394.8000 195.6000 395.6000 195.7000 ;
	    RECT 423.6000 195.6000 424.4000 195.7000 ;
	    RECT 438.0000 195.6000 438.8000 195.7000 ;
	    RECT 458.8000 196.3000 459.6000 196.4000 ;
	    RECT 482.8000 196.3000 483.6000 196.4000 ;
	    RECT 458.8000 195.7000 483.6000 196.3000 ;
	    RECT 458.8000 195.6000 459.6000 195.7000 ;
	    RECT 482.8000 195.6000 483.6000 195.7000 ;
	    RECT 510.0000 195.6000 510.8000 196.4000 ;
	    RECT 28.4000 194.3000 29.2000 194.4000 ;
	    RECT 156.4000 194.3000 157.2000 194.4000 ;
	    RECT 177.2000 194.3000 178.0000 194.4000 ;
	    RECT 306.8000 194.3000 307.6000 194.4000 ;
	    RECT 330.8000 194.3000 331.6000 194.4000 ;
	    RECT 343.6000 194.3000 344.4000 194.4000 ;
	    RECT 28.4000 193.7000 344.4000 194.3000 ;
	    RECT 28.4000 193.6000 29.2000 193.7000 ;
	    RECT 156.4000 193.6000 157.2000 193.7000 ;
	    RECT 177.2000 193.6000 178.0000 193.7000 ;
	    RECT 306.8000 193.6000 307.6000 193.7000 ;
	    RECT 330.8000 193.6000 331.6000 193.7000 ;
	    RECT 343.6000 193.6000 344.4000 193.7000 ;
	    RECT 346.8000 194.3000 347.6000 194.4000 ;
	    RECT 356.4000 194.3000 357.2000 194.4000 ;
	    RECT 346.8000 193.7000 357.2000 194.3000 ;
	    RECT 359.7000 194.3000 360.3000 195.6000 ;
	    RECT 385.2000 194.3000 386.0000 194.4000 ;
	    RECT 426.8000 194.3000 427.6000 194.4000 ;
	    RECT 359.7000 193.7000 427.6000 194.3000 ;
	    RECT 346.8000 193.6000 347.6000 193.7000 ;
	    RECT 356.4000 193.6000 357.2000 193.7000 ;
	    RECT 385.2000 193.6000 386.0000 193.7000 ;
	    RECT 426.8000 193.6000 427.6000 193.7000 ;
	    RECT 457.2000 194.3000 458.0000 194.4000 ;
	    RECT 463.6000 194.3000 464.4000 194.4000 ;
	    RECT 470.0000 194.3000 470.8000 194.4000 ;
	    RECT 457.2000 193.7000 470.8000 194.3000 ;
	    RECT 457.2000 193.6000 458.0000 193.7000 ;
	    RECT 463.6000 193.6000 464.4000 193.7000 ;
	    RECT 470.0000 193.6000 470.8000 193.7000 ;
	    RECT 474.8000 194.3000 475.6000 194.4000 ;
	    RECT 484.4000 194.3000 485.2000 194.4000 ;
	    RECT 474.8000 193.7000 485.2000 194.3000 ;
	    RECT 474.8000 193.6000 475.6000 193.7000 ;
	    RECT 484.4000 193.6000 485.2000 193.7000 ;
	    RECT 487.6000 194.3000 488.4000 194.4000 ;
	    RECT 505.2000 194.3000 506.0000 194.4000 ;
	    RECT 506.8000 194.3000 507.6000 194.4000 ;
	    RECT 487.6000 193.7000 507.6000 194.3000 ;
	    RECT 487.6000 193.6000 488.4000 193.7000 ;
	    RECT 505.2000 193.6000 506.0000 193.7000 ;
	    RECT 506.8000 193.6000 507.6000 193.7000 ;
	    RECT 4.4000 192.3000 5.2000 192.4000 ;
	    RECT 20.4000 192.3000 21.2000 192.4000 ;
	    RECT 4.4000 191.7000 21.2000 192.3000 ;
	    RECT 4.4000 191.6000 5.2000 191.7000 ;
	    RECT 20.4000 191.6000 21.2000 191.7000 ;
	    RECT 36.4000 192.3000 37.2000 192.4000 ;
	    RECT 41.2000 192.3000 42.0000 192.4000 ;
	    RECT 36.4000 191.7000 42.0000 192.3000 ;
	    RECT 36.4000 191.6000 37.2000 191.7000 ;
	    RECT 41.2000 191.6000 42.0000 191.7000 ;
	    RECT 87.6000 192.3000 88.4000 192.4000 ;
	    RECT 100.4000 192.3000 101.2000 192.4000 ;
	    RECT 105.2000 192.3000 106.0000 192.4000 ;
	    RECT 129.2000 192.3000 130.0000 192.4000 ;
	    RECT 87.6000 191.7000 130.0000 192.3000 ;
	    RECT 87.6000 191.6000 88.4000 191.7000 ;
	    RECT 100.4000 191.6000 101.2000 191.7000 ;
	    RECT 105.2000 191.6000 106.0000 191.7000 ;
	    RECT 129.2000 191.6000 130.0000 191.7000 ;
	    RECT 130.8000 192.3000 131.6000 192.4000 ;
	    RECT 134.0000 192.3000 134.8000 192.4000 ;
	    RECT 130.8000 191.7000 134.8000 192.3000 ;
	    RECT 130.8000 191.6000 131.6000 191.7000 ;
	    RECT 134.0000 191.6000 134.8000 191.7000 ;
	    RECT 145.2000 192.3000 146.0000 192.4000 ;
	    RECT 146.8000 192.3000 147.6000 192.4000 ;
	    RECT 154.8000 192.3000 155.6000 192.4000 ;
	    RECT 145.2000 191.7000 155.6000 192.3000 ;
	    RECT 145.2000 191.6000 146.0000 191.7000 ;
	    RECT 146.8000 191.6000 147.6000 191.7000 ;
	    RECT 154.8000 191.6000 155.6000 191.7000 ;
	    RECT 164.4000 192.3000 165.2000 192.4000 ;
	    RECT 172.4000 192.3000 173.2000 192.4000 ;
	    RECT 177.2000 192.3000 178.0000 192.4000 ;
	    RECT 164.4000 191.7000 178.0000 192.3000 ;
	    RECT 164.4000 191.6000 165.2000 191.7000 ;
	    RECT 172.4000 191.6000 173.2000 191.7000 ;
	    RECT 177.2000 191.6000 178.0000 191.7000 ;
	    RECT 183.6000 192.3000 184.4000 192.4000 ;
	    RECT 185.2000 192.3000 186.0000 192.4000 ;
	    RECT 196.4000 192.3000 197.2000 192.4000 ;
	    RECT 204.4000 192.3000 205.2000 192.4000 ;
	    RECT 183.6000 191.7000 205.2000 192.3000 ;
	    RECT 183.6000 191.6000 184.4000 191.7000 ;
	    RECT 185.2000 191.6000 186.0000 191.7000 ;
	    RECT 196.4000 191.6000 197.2000 191.7000 ;
	    RECT 204.4000 191.6000 205.2000 191.7000 ;
	    RECT 207.6000 192.3000 208.4000 192.4000 ;
	    RECT 217.2000 192.3000 218.0000 192.4000 ;
	    RECT 207.6000 191.7000 218.0000 192.3000 ;
	    RECT 207.6000 191.6000 208.4000 191.7000 ;
	    RECT 217.2000 191.6000 218.0000 191.7000 ;
	    RECT 220.4000 192.3000 221.2000 192.4000 ;
	    RECT 228.4000 192.3000 229.2000 192.4000 ;
	    RECT 220.4000 191.7000 229.2000 192.3000 ;
	    RECT 220.4000 191.6000 221.2000 191.7000 ;
	    RECT 228.4000 191.6000 229.2000 191.7000 ;
	    RECT 231.6000 192.3000 232.4000 192.4000 ;
	    RECT 239.6000 192.3000 240.4000 192.4000 ;
	    RECT 231.6000 191.7000 240.4000 192.3000 ;
	    RECT 231.6000 191.6000 232.4000 191.7000 ;
	    RECT 239.6000 191.6000 240.4000 191.7000 ;
	    RECT 241.2000 192.3000 242.0000 192.4000 ;
	    RECT 249.2000 192.3000 250.0000 192.4000 ;
	    RECT 241.2000 191.7000 250.0000 192.3000 ;
	    RECT 241.2000 191.6000 242.0000 191.7000 ;
	    RECT 249.2000 191.6000 250.0000 191.7000 ;
	    RECT 263.6000 192.3000 264.4000 192.4000 ;
	    RECT 270.0000 192.3000 270.8000 192.4000 ;
	    RECT 263.6000 191.7000 270.8000 192.3000 ;
	    RECT 263.6000 191.6000 264.4000 191.7000 ;
	    RECT 270.0000 191.6000 270.8000 191.7000 ;
	    RECT 274.8000 192.3000 275.6000 192.4000 ;
	    RECT 441.2000 192.3000 442.0000 192.4000 ;
	    RECT 274.8000 191.7000 442.0000 192.3000 ;
	    RECT 274.8000 191.6000 275.6000 191.7000 ;
	    RECT 441.2000 191.6000 442.0000 191.7000 ;
	    RECT 442.8000 192.3000 443.6000 192.4000 ;
	    RECT 450.8000 192.3000 451.6000 192.4000 ;
	    RECT 458.8000 192.3000 459.6000 192.4000 ;
	    RECT 465.2000 192.3000 466.0000 192.4000 ;
	    RECT 471.6000 192.3000 472.4000 192.4000 ;
	    RECT 442.8000 191.7000 472.4000 192.3000 ;
	    RECT 442.8000 191.6000 443.6000 191.7000 ;
	    RECT 450.8000 191.6000 451.6000 191.7000 ;
	    RECT 458.8000 191.6000 459.6000 191.7000 ;
	    RECT 465.2000 191.6000 466.0000 191.7000 ;
	    RECT 471.6000 191.6000 472.4000 191.7000 ;
	    RECT 9.2000 190.3000 10.0000 190.4000 ;
	    RECT 12.4000 190.3000 13.2000 190.4000 ;
	    RECT 17.2000 190.3000 18.0000 190.4000 ;
	    RECT 9.2000 189.7000 18.0000 190.3000 ;
	    RECT 9.2000 189.6000 10.0000 189.7000 ;
	    RECT 12.4000 189.6000 13.2000 189.7000 ;
	    RECT 17.2000 189.6000 18.0000 189.7000 ;
	    RECT 34.8000 190.3000 35.6000 190.4000 ;
	    RECT 47.6000 190.3000 48.4000 190.4000 ;
	    RECT 34.8000 189.7000 48.4000 190.3000 ;
	    RECT 34.8000 189.6000 35.6000 189.7000 ;
	    RECT 47.6000 189.6000 48.4000 189.7000 ;
	    RECT 50.8000 190.3000 51.6000 190.4000 ;
	    RECT 63.6000 190.3000 64.4000 190.4000 ;
	    RECT 50.8000 189.7000 64.4000 190.3000 ;
	    RECT 50.8000 189.6000 51.6000 189.7000 ;
	    RECT 63.6000 189.6000 64.4000 189.7000 ;
	    RECT 78.0000 190.3000 78.8000 190.4000 ;
	    RECT 97.2000 190.3000 98.0000 190.4000 ;
	    RECT 78.0000 189.7000 98.0000 190.3000 ;
	    RECT 78.0000 189.6000 78.8000 189.7000 ;
	    RECT 97.2000 189.6000 98.0000 189.7000 ;
	    RECT 122.8000 190.3000 123.6000 190.4000 ;
	    RECT 138.8000 190.3000 139.6000 190.4000 ;
	    RECT 122.8000 189.7000 139.6000 190.3000 ;
	    RECT 122.8000 189.6000 123.6000 189.7000 ;
	    RECT 138.8000 189.6000 139.6000 189.7000 ;
	    RECT 161.2000 190.3000 162.0000 190.4000 ;
	    RECT 177.2000 190.3000 178.0000 190.4000 ;
	    RECT 161.2000 189.7000 178.0000 190.3000 ;
	    RECT 161.2000 189.6000 162.0000 189.7000 ;
	    RECT 177.2000 189.6000 178.0000 189.7000 ;
	    RECT 188.4000 190.3000 189.2000 190.4000 ;
	    RECT 196.4000 190.3000 197.2000 190.4000 ;
	    RECT 209.2000 190.3000 210.0000 190.4000 ;
	    RECT 188.4000 189.7000 210.0000 190.3000 ;
	    RECT 188.4000 189.6000 189.2000 189.7000 ;
	    RECT 196.4000 189.6000 197.2000 189.7000 ;
	    RECT 209.2000 189.6000 210.0000 189.7000 ;
	    RECT 215.6000 190.3000 216.4000 190.4000 ;
	    RECT 234.8000 190.3000 235.6000 190.4000 ;
	    RECT 215.6000 189.7000 235.6000 190.3000 ;
	    RECT 215.6000 189.6000 216.4000 189.7000 ;
	    RECT 234.8000 189.6000 235.6000 189.7000 ;
	    RECT 241.2000 190.3000 242.0000 190.4000 ;
	    RECT 244.4000 190.3000 245.2000 190.4000 ;
	    RECT 241.2000 189.7000 245.2000 190.3000 ;
	    RECT 241.2000 189.6000 242.0000 189.7000 ;
	    RECT 244.4000 189.6000 245.2000 189.7000 ;
	    RECT 249.2000 190.3000 250.0000 190.4000 ;
	    RECT 265.2000 190.3000 266.0000 190.4000 ;
	    RECT 249.2000 189.7000 266.0000 190.3000 ;
	    RECT 249.2000 189.6000 250.0000 189.7000 ;
	    RECT 265.2000 189.6000 266.0000 189.7000 ;
	    RECT 274.8000 190.3000 275.6000 190.4000 ;
	    RECT 292.4000 190.3000 293.2000 190.4000 ;
	    RECT 274.8000 189.7000 293.2000 190.3000 ;
	    RECT 274.8000 189.6000 275.6000 189.7000 ;
	    RECT 292.4000 189.6000 293.2000 189.7000 ;
	    RECT 297.2000 190.3000 298.0000 190.4000 ;
	    RECT 311.6000 190.3000 312.4000 190.4000 ;
	    RECT 316.4000 190.3000 317.2000 190.4000 ;
	    RECT 297.2000 189.7000 310.7000 190.3000 ;
	    RECT 297.2000 189.6000 298.0000 189.7000 ;
	    RECT 20.4000 188.3000 21.2000 188.4000 ;
	    RECT 46.0000 188.3000 46.8000 188.4000 ;
	    RECT 20.4000 187.7000 46.8000 188.3000 ;
	    RECT 20.4000 187.6000 21.2000 187.7000 ;
	    RECT 46.0000 187.6000 46.8000 187.7000 ;
	    RECT 57.2000 188.3000 58.0000 188.4000 ;
	    RECT 63.6000 188.3000 64.4000 188.4000 ;
	    RECT 68.4000 188.3000 69.2000 188.4000 ;
	    RECT 57.2000 187.7000 69.2000 188.3000 ;
	    RECT 57.2000 187.6000 58.0000 187.7000 ;
	    RECT 63.6000 187.6000 64.4000 187.7000 ;
	    RECT 68.4000 187.6000 69.2000 187.7000 ;
	    RECT 100.4000 188.3000 101.2000 188.4000 ;
	    RECT 103.6000 188.3000 104.4000 188.4000 ;
	    RECT 100.4000 187.7000 104.4000 188.3000 ;
	    RECT 100.4000 187.6000 101.2000 187.7000 ;
	    RECT 103.6000 187.6000 104.4000 187.7000 ;
	    RECT 105.2000 188.3000 106.0000 188.4000 ;
	    RECT 113.2000 188.3000 114.0000 188.4000 ;
	    RECT 105.2000 187.7000 114.0000 188.3000 ;
	    RECT 105.2000 187.6000 106.0000 187.7000 ;
	    RECT 113.2000 187.6000 114.0000 187.7000 ;
	    RECT 119.6000 188.3000 120.4000 188.4000 ;
	    RECT 124.4000 188.3000 125.2000 188.4000 ;
	    RECT 119.6000 187.7000 125.2000 188.3000 ;
	    RECT 119.6000 187.6000 120.4000 187.7000 ;
	    RECT 124.4000 187.6000 125.2000 187.7000 ;
	    RECT 127.6000 188.3000 128.4000 188.4000 ;
	    RECT 142.0000 188.3000 142.8000 188.4000 ;
	    RECT 183.6000 188.3000 184.4000 188.4000 ;
	    RECT 127.6000 187.7000 142.8000 188.3000 ;
	    RECT 127.6000 187.6000 128.4000 187.7000 ;
	    RECT 142.0000 187.6000 142.8000 187.7000 ;
	    RECT 145.3000 187.7000 184.4000 188.3000 ;
	    RECT 145.3000 186.4000 145.9000 187.7000 ;
	    RECT 183.6000 187.6000 184.4000 187.7000 ;
	    RECT 199.6000 188.3000 200.4000 188.4000 ;
	    RECT 207.6000 188.3000 208.4000 188.4000 ;
	    RECT 199.6000 187.7000 208.4000 188.3000 ;
	    RECT 199.6000 187.6000 200.4000 187.7000 ;
	    RECT 207.6000 187.6000 208.4000 187.7000 ;
	    RECT 214.0000 188.3000 214.8000 188.4000 ;
	    RECT 246.0000 188.3000 246.8000 188.4000 ;
	    RECT 214.0000 187.7000 246.8000 188.3000 ;
	    RECT 214.0000 187.6000 214.8000 187.7000 ;
	    RECT 246.0000 187.6000 246.8000 187.7000 ;
	    RECT 249.2000 188.3000 250.0000 188.4000 ;
	    RECT 284.4000 188.3000 285.2000 188.4000 ;
	    RECT 249.2000 187.7000 285.2000 188.3000 ;
	    RECT 310.1000 188.3000 310.7000 189.7000 ;
	    RECT 311.6000 189.7000 317.2000 190.3000 ;
	    RECT 311.6000 189.6000 312.4000 189.7000 ;
	    RECT 316.4000 189.6000 317.2000 189.7000 ;
	    RECT 318.0000 190.3000 318.8000 190.4000 ;
	    RECT 330.8000 190.3000 331.6000 190.4000 ;
	    RECT 318.0000 189.7000 331.6000 190.3000 ;
	    RECT 318.0000 189.6000 318.8000 189.7000 ;
	    RECT 330.8000 189.6000 331.6000 189.7000 ;
	    RECT 353.2000 190.3000 354.0000 190.4000 ;
	    RECT 364.4000 190.3000 365.2000 190.4000 ;
	    RECT 353.2000 189.7000 365.2000 190.3000 ;
	    RECT 353.2000 189.6000 354.0000 189.7000 ;
	    RECT 364.4000 189.6000 365.2000 189.7000 ;
	    RECT 385.2000 190.3000 386.0000 190.4000 ;
	    RECT 410.8000 190.3000 411.6000 190.4000 ;
	    RECT 385.2000 189.7000 411.6000 190.3000 ;
	    RECT 385.2000 189.6000 386.0000 189.7000 ;
	    RECT 410.8000 189.6000 411.6000 189.7000 ;
	    RECT 414.0000 190.3000 414.8000 190.4000 ;
	    RECT 454.0000 190.3000 454.8000 190.4000 ;
	    RECT 414.0000 189.7000 454.8000 190.3000 ;
	    RECT 414.0000 189.6000 414.8000 189.7000 ;
	    RECT 454.0000 189.6000 454.8000 189.7000 ;
	    RECT 482.8000 190.3000 483.6000 190.4000 ;
	    RECT 492.4000 190.3000 493.2000 190.4000 ;
	    RECT 482.8000 189.7000 493.2000 190.3000 ;
	    RECT 482.8000 189.6000 483.6000 189.7000 ;
	    RECT 492.4000 189.6000 493.2000 189.7000 ;
	    RECT 494.0000 190.3000 494.8000 190.4000 ;
	    RECT 513.2000 190.3000 514.0000 190.4000 ;
	    RECT 494.0000 189.7000 514.0000 190.3000 ;
	    RECT 494.0000 189.6000 494.8000 189.7000 ;
	    RECT 513.2000 189.6000 514.0000 189.7000 ;
	    RECT 314.8000 188.3000 315.6000 188.4000 ;
	    RECT 310.1000 187.7000 315.6000 188.3000 ;
	    RECT 249.2000 187.6000 250.0000 187.7000 ;
	    RECT 284.4000 187.6000 285.2000 187.7000 ;
	    RECT 314.8000 187.6000 315.6000 187.7000 ;
	    RECT 318.0000 188.3000 318.8000 188.4000 ;
	    RECT 329.2000 188.3000 330.0000 188.4000 ;
	    RECT 318.0000 187.7000 330.0000 188.3000 ;
	    RECT 318.0000 187.6000 318.8000 187.7000 ;
	    RECT 329.2000 187.6000 330.0000 187.7000 ;
	    RECT 359.6000 188.3000 360.4000 188.4000 ;
	    RECT 375.6000 188.3000 376.4000 188.4000 ;
	    RECT 359.6000 187.7000 376.4000 188.3000 ;
	    RECT 359.6000 187.6000 360.4000 187.7000 ;
	    RECT 375.6000 187.6000 376.4000 187.7000 ;
	    RECT 383.6000 188.3000 384.4000 188.4000 ;
	    RECT 386.8000 188.3000 387.6000 188.4000 ;
	    RECT 383.6000 187.7000 387.6000 188.3000 ;
	    RECT 383.6000 187.6000 384.4000 187.7000 ;
	    RECT 386.8000 187.6000 387.6000 187.7000 ;
	    RECT 506.8000 187.6000 507.6000 188.4000 ;
	    RECT 6.0000 186.3000 6.8000 186.4000 ;
	    RECT 41.2000 186.3000 42.0000 186.4000 ;
	    RECT 46.0000 186.3000 46.8000 186.4000 ;
	    RECT 6.0000 185.7000 46.8000 186.3000 ;
	    RECT 6.0000 185.6000 6.8000 185.7000 ;
	    RECT 41.2000 185.6000 42.0000 185.7000 ;
	    RECT 46.0000 185.6000 46.8000 185.7000 ;
	    RECT 55.6000 186.3000 56.4000 186.4000 ;
	    RECT 129.2000 186.3000 130.0000 186.4000 ;
	    RECT 145.2000 186.3000 146.0000 186.4000 ;
	    RECT 55.6000 185.7000 121.9000 186.3000 ;
	    RECT 55.6000 185.6000 56.4000 185.7000 ;
	    RECT 55.6000 184.3000 56.4000 184.4000 ;
	    RECT 74.8000 184.3000 75.6000 184.4000 ;
	    RECT 119.6000 184.3000 120.4000 184.4000 ;
	    RECT 55.6000 183.7000 120.4000 184.3000 ;
	    RECT 121.3000 184.3000 121.9000 185.7000 ;
	    RECT 129.2000 185.7000 146.0000 186.3000 ;
	    RECT 129.2000 185.6000 130.0000 185.7000 ;
	    RECT 145.2000 185.6000 146.0000 185.7000 ;
	    RECT 154.8000 186.3000 155.6000 186.4000 ;
	    RECT 180.4000 186.3000 181.2000 186.4000 ;
	    RECT 154.8000 185.7000 181.2000 186.3000 ;
	    RECT 154.8000 185.6000 155.6000 185.7000 ;
	    RECT 180.4000 185.6000 181.2000 185.7000 ;
	    RECT 196.4000 186.3000 197.2000 186.4000 ;
	    RECT 222.0000 186.3000 222.8000 186.4000 ;
	    RECT 196.4000 185.7000 222.8000 186.3000 ;
	    RECT 196.4000 185.6000 197.2000 185.7000 ;
	    RECT 222.0000 185.6000 222.8000 185.7000 ;
	    RECT 223.6000 186.3000 224.4000 186.4000 ;
	    RECT 238.0000 186.3000 238.8000 186.4000 ;
	    RECT 223.6000 185.7000 238.8000 186.3000 ;
	    RECT 223.6000 185.6000 224.4000 185.7000 ;
	    RECT 238.0000 185.6000 238.8000 185.7000 ;
	    RECT 241.2000 186.3000 242.0000 186.4000 ;
	    RECT 279.6000 186.3000 280.4000 186.4000 ;
	    RECT 297.2000 186.3000 298.0000 186.4000 ;
	    RECT 343.6000 186.3000 344.4000 186.4000 ;
	    RECT 350.0000 186.3000 350.8000 186.4000 ;
	    RECT 241.2000 185.7000 350.8000 186.3000 ;
	    RECT 241.2000 185.6000 242.0000 185.7000 ;
	    RECT 279.6000 185.6000 280.4000 185.7000 ;
	    RECT 297.2000 185.6000 298.0000 185.7000 ;
	    RECT 343.6000 185.6000 344.4000 185.7000 ;
	    RECT 350.0000 185.6000 350.8000 185.7000 ;
	    RECT 180.5000 184.4000 181.1000 185.6000 ;
	    RECT 134.0000 184.3000 134.8000 184.4000 ;
	    RECT 121.3000 183.7000 134.8000 184.3000 ;
	    RECT 55.6000 183.6000 56.4000 183.7000 ;
	    RECT 74.8000 183.6000 75.6000 183.7000 ;
	    RECT 119.6000 183.6000 120.4000 183.7000 ;
	    RECT 134.0000 183.6000 134.8000 183.7000 ;
	    RECT 151.6000 184.3000 152.4000 184.4000 ;
	    RECT 162.8000 184.3000 163.6000 184.4000 ;
	    RECT 151.6000 183.7000 163.6000 184.3000 ;
	    RECT 151.6000 183.6000 152.4000 183.7000 ;
	    RECT 162.8000 183.6000 163.6000 183.7000 ;
	    RECT 180.4000 183.6000 181.2000 184.4000 ;
	    RECT 182.0000 184.3000 182.8000 184.4000 ;
	    RECT 188.4000 184.3000 189.2000 184.4000 ;
	    RECT 182.0000 183.7000 189.2000 184.3000 ;
	    RECT 182.0000 183.6000 182.8000 183.7000 ;
	    RECT 188.4000 183.6000 189.2000 183.7000 ;
	    RECT 194.8000 184.3000 195.6000 184.4000 ;
	    RECT 215.6000 184.3000 216.4000 184.4000 ;
	    RECT 226.8000 184.3000 227.6000 184.4000 ;
	    RECT 194.8000 183.7000 216.4000 184.3000 ;
	    RECT 194.8000 183.6000 195.6000 183.7000 ;
	    RECT 215.6000 183.6000 216.4000 183.7000 ;
	    RECT 217.3000 183.7000 227.6000 184.3000 ;
	    RECT 22.0000 182.3000 22.8000 182.4000 ;
	    RECT 113.2000 182.3000 114.0000 182.4000 ;
	    RECT 22.0000 181.7000 114.0000 182.3000 ;
	    RECT 22.0000 181.6000 22.8000 181.7000 ;
	    RECT 113.2000 181.6000 114.0000 181.7000 ;
	    RECT 170.8000 182.3000 171.6000 182.4000 ;
	    RECT 185.2000 182.3000 186.0000 182.4000 ;
	    RECT 194.8000 182.3000 195.6000 182.4000 ;
	    RECT 170.8000 181.7000 195.6000 182.3000 ;
	    RECT 170.8000 181.6000 171.6000 181.7000 ;
	    RECT 185.2000 181.6000 186.0000 181.7000 ;
	    RECT 194.8000 181.6000 195.6000 181.7000 ;
	    RECT 199.6000 182.3000 200.4000 182.4000 ;
	    RECT 217.3000 182.3000 217.9000 183.7000 ;
	    RECT 226.8000 183.6000 227.6000 183.7000 ;
	    RECT 228.4000 184.3000 229.2000 184.4000 ;
	    RECT 233.2000 184.3000 234.0000 184.4000 ;
	    RECT 228.4000 183.7000 234.0000 184.3000 ;
	    RECT 228.4000 183.6000 229.2000 183.7000 ;
	    RECT 233.2000 183.6000 234.0000 183.7000 ;
	    RECT 234.8000 184.3000 235.6000 184.4000 ;
	    RECT 244.4000 184.3000 245.2000 184.4000 ;
	    RECT 258.8000 184.3000 259.6000 184.4000 ;
	    RECT 278.0000 184.3000 278.8000 184.4000 ;
	    RECT 234.8000 183.7000 278.8000 184.3000 ;
	    RECT 234.8000 183.6000 235.6000 183.7000 ;
	    RECT 244.4000 183.6000 245.2000 183.7000 ;
	    RECT 258.8000 183.6000 259.6000 183.7000 ;
	    RECT 278.0000 183.6000 278.8000 183.7000 ;
	    RECT 284.4000 184.3000 285.2000 184.4000 ;
	    RECT 327.6000 184.3000 328.4000 184.4000 ;
	    RECT 284.4000 183.7000 328.4000 184.3000 ;
	    RECT 284.4000 183.6000 285.2000 183.7000 ;
	    RECT 327.6000 183.6000 328.4000 183.7000 ;
	    RECT 329.2000 184.3000 330.0000 184.4000 ;
	    RECT 362.8000 184.3000 363.6000 184.4000 ;
	    RECT 380.4000 184.3000 381.2000 184.4000 ;
	    RECT 329.2000 183.7000 381.2000 184.3000 ;
	    RECT 329.2000 183.6000 330.0000 183.7000 ;
	    RECT 362.8000 183.6000 363.6000 183.7000 ;
	    RECT 380.4000 183.6000 381.2000 183.7000 ;
	    RECT 382.0000 184.3000 382.8000 184.4000 ;
	    RECT 436.4000 184.3000 437.2000 184.4000 ;
	    RECT 382.0000 183.7000 437.2000 184.3000 ;
	    RECT 382.0000 183.6000 382.8000 183.7000 ;
	    RECT 436.4000 183.6000 437.2000 183.7000 ;
	    RECT 452.4000 183.6000 453.2000 184.4000 ;
	    RECT 481.2000 184.3000 482.0000 184.4000 ;
	    RECT 495.6000 184.3000 496.4000 184.4000 ;
	    RECT 481.2000 183.7000 496.4000 184.3000 ;
	    RECT 481.2000 183.6000 482.0000 183.7000 ;
	    RECT 495.6000 183.6000 496.4000 183.7000 ;
	    RECT 199.6000 181.7000 217.9000 182.3000 ;
	    RECT 220.4000 182.3000 221.2000 182.4000 ;
	    RECT 223.6000 182.3000 224.4000 182.4000 ;
	    RECT 220.4000 181.7000 224.4000 182.3000 ;
	    RECT 199.6000 181.6000 200.4000 181.7000 ;
	    RECT 220.4000 181.6000 221.2000 181.7000 ;
	    RECT 223.6000 181.6000 224.4000 181.7000 ;
	    RECT 230.0000 182.3000 230.8000 182.4000 ;
	    RECT 234.8000 182.3000 235.6000 182.4000 ;
	    RECT 230.0000 181.7000 235.6000 182.3000 ;
	    RECT 230.0000 181.6000 230.8000 181.7000 ;
	    RECT 234.8000 181.6000 235.6000 181.7000 ;
	    RECT 236.4000 182.3000 237.2000 182.4000 ;
	    RECT 263.6000 182.3000 264.4000 182.4000 ;
	    RECT 274.8000 182.3000 275.6000 182.4000 ;
	    RECT 236.4000 181.7000 251.5000 182.3000 ;
	    RECT 236.4000 181.6000 237.2000 181.7000 ;
	    RECT 122.8000 180.3000 123.6000 180.4000 ;
	    RECT 127.6000 180.3000 128.4000 180.4000 ;
	    RECT 122.8000 179.7000 128.4000 180.3000 ;
	    RECT 122.8000 179.6000 123.6000 179.7000 ;
	    RECT 127.6000 179.6000 128.4000 179.7000 ;
	    RECT 132.4000 180.3000 133.2000 180.4000 ;
	    RECT 146.8000 180.3000 147.6000 180.4000 ;
	    RECT 132.4000 179.7000 147.6000 180.3000 ;
	    RECT 132.4000 179.6000 133.2000 179.7000 ;
	    RECT 146.8000 179.6000 147.6000 179.7000 ;
	    RECT 174.0000 180.3000 174.8000 180.4000 ;
	    RECT 199.6000 180.3000 200.4000 180.4000 ;
	    RECT 174.0000 179.7000 200.4000 180.3000 ;
	    RECT 174.0000 179.6000 174.8000 179.7000 ;
	    RECT 199.6000 179.6000 200.4000 179.7000 ;
	    RECT 201.2000 180.3000 202.0000 180.4000 ;
	    RECT 217.2000 180.3000 218.0000 180.4000 ;
	    RECT 249.2000 180.3000 250.0000 180.4000 ;
	    RECT 201.2000 179.7000 250.0000 180.3000 ;
	    RECT 250.9000 180.3000 251.5000 181.7000 ;
	    RECT 263.6000 181.7000 275.6000 182.3000 ;
	    RECT 263.6000 181.6000 264.4000 181.7000 ;
	    RECT 274.8000 181.6000 275.6000 181.7000 ;
	    RECT 279.6000 182.3000 280.4000 182.4000 ;
	    RECT 292.4000 182.3000 293.2000 182.4000 ;
	    RECT 279.6000 181.7000 293.2000 182.3000 ;
	    RECT 279.6000 181.6000 280.4000 181.7000 ;
	    RECT 292.4000 181.6000 293.2000 181.7000 ;
	    RECT 295.6000 182.3000 296.4000 182.4000 ;
	    RECT 335.6000 182.3000 336.4000 182.4000 ;
	    RECT 295.6000 181.7000 336.4000 182.3000 ;
	    RECT 295.6000 181.6000 296.4000 181.7000 ;
	    RECT 335.6000 181.6000 336.4000 181.7000 ;
	    RECT 338.8000 182.3000 339.6000 182.4000 ;
	    RECT 350.0000 182.3000 350.8000 182.4000 ;
	    RECT 353.2000 182.3000 354.0000 182.4000 ;
	    RECT 338.8000 181.7000 354.0000 182.3000 ;
	    RECT 338.8000 181.6000 339.6000 181.7000 ;
	    RECT 350.0000 181.6000 350.8000 181.7000 ;
	    RECT 353.2000 181.6000 354.0000 181.7000 ;
	    RECT 399.6000 182.3000 400.4000 182.4000 ;
	    RECT 417.2000 182.3000 418.0000 182.4000 ;
	    RECT 399.6000 181.7000 418.0000 182.3000 ;
	    RECT 399.6000 181.6000 400.4000 181.7000 ;
	    RECT 417.2000 181.6000 418.0000 181.7000 ;
	    RECT 265.2000 180.3000 266.0000 180.4000 ;
	    RECT 284.4000 180.3000 285.2000 180.4000 ;
	    RECT 250.9000 179.7000 253.1000 180.3000 ;
	    RECT 201.2000 179.6000 202.0000 179.7000 ;
	    RECT 217.2000 179.6000 218.0000 179.7000 ;
	    RECT 249.2000 179.6000 250.0000 179.7000 ;
	    RECT 34.8000 178.3000 35.6000 178.4000 ;
	    RECT 103.6000 178.3000 104.4000 178.4000 ;
	    RECT 121.2000 178.3000 122.0000 178.4000 ;
	    RECT 34.8000 177.7000 96.3000 178.3000 ;
	    RECT 34.8000 177.6000 35.6000 177.7000 ;
	    RECT 84.4000 176.3000 85.2000 176.4000 ;
	    RECT 94.0000 176.3000 94.8000 176.4000 ;
	    RECT 84.4000 175.7000 94.8000 176.3000 ;
	    RECT 95.7000 176.3000 96.3000 177.7000 ;
	    RECT 103.6000 177.7000 122.0000 178.3000 ;
	    RECT 103.6000 177.6000 104.4000 177.7000 ;
	    RECT 121.2000 177.6000 122.0000 177.7000 ;
	    RECT 158.0000 178.3000 158.8000 178.4000 ;
	    RECT 164.4000 178.3000 165.2000 178.4000 ;
	    RECT 158.0000 177.7000 165.2000 178.3000 ;
	    RECT 158.0000 177.6000 158.8000 177.7000 ;
	    RECT 164.4000 177.6000 165.2000 177.7000 ;
	    RECT 188.4000 178.3000 189.2000 178.4000 ;
	    RECT 198.0000 178.3000 198.8000 178.4000 ;
	    RECT 214.0000 178.3000 214.8000 178.4000 ;
	    RECT 225.2000 178.3000 226.0000 178.4000 ;
	    RECT 188.4000 177.7000 226.0000 178.3000 ;
	    RECT 188.4000 177.6000 189.2000 177.7000 ;
	    RECT 198.0000 177.6000 198.8000 177.7000 ;
	    RECT 214.0000 177.6000 214.8000 177.7000 ;
	    RECT 225.2000 177.6000 226.0000 177.7000 ;
	    RECT 228.4000 178.3000 229.2000 178.4000 ;
	    RECT 246.0000 178.3000 246.8000 178.4000 ;
	    RECT 228.4000 177.7000 246.8000 178.3000 ;
	    RECT 228.4000 177.6000 229.2000 177.7000 ;
	    RECT 246.0000 177.6000 246.8000 177.7000 ;
	    RECT 247.6000 178.3000 248.4000 178.4000 ;
	    RECT 250.8000 178.3000 251.6000 178.4000 ;
	    RECT 247.6000 177.7000 251.6000 178.3000 ;
	    RECT 252.5000 178.3000 253.1000 179.7000 ;
	    RECT 265.2000 179.7000 285.2000 180.3000 ;
	    RECT 265.2000 179.6000 266.0000 179.7000 ;
	    RECT 284.4000 179.6000 285.2000 179.7000 ;
	    RECT 286.0000 180.3000 286.8000 180.4000 ;
	    RECT 292.4000 180.3000 293.2000 180.4000 ;
	    RECT 286.0000 179.7000 293.2000 180.3000 ;
	    RECT 286.0000 179.6000 286.8000 179.7000 ;
	    RECT 292.4000 179.6000 293.2000 179.7000 ;
	    RECT 294.0000 180.3000 294.8000 180.4000 ;
	    RECT 305.2000 180.3000 306.0000 180.4000 ;
	    RECT 294.0000 179.7000 306.0000 180.3000 ;
	    RECT 294.0000 179.6000 294.8000 179.7000 ;
	    RECT 305.2000 179.6000 306.0000 179.7000 ;
	    RECT 319.6000 180.3000 320.4000 180.4000 ;
	    RECT 346.8000 180.3000 347.6000 180.4000 ;
	    RECT 319.6000 179.7000 347.6000 180.3000 ;
	    RECT 319.6000 179.6000 320.4000 179.7000 ;
	    RECT 346.8000 179.6000 347.6000 179.7000 ;
	    RECT 353.2000 180.3000 354.0000 180.4000 ;
	    RECT 361.2000 180.3000 362.0000 180.4000 ;
	    RECT 353.2000 179.7000 362.0000 180.3000 ;
	    RECT 353.2000 179.6000 354.0000 179.7000 ;
	    RECT 361.2000 179.6000 362.0000 179.7000 ;
	    RECT 414.0000 180.3000 414.8000 180.4000 ;
	    RECT 444.4000 180.3000 445.2000 180.4000 ;
	    RECT 414.0000 179.7000 445.2000 180.3000 ;
	    RECT 414.0000 179.6000 414.8000 179.7000 ;
	    RECT 444.4000 179.6000 445.2000 179.7000 ;
	    RECT 255.6000 178.3000 256.4000 178.4000 ;
	    RECT 252.5000 177.7000 256.4000 178.3000 ;
	    RECT 247.6000 177.6000 248.4000 177.7000 ;
	    RECT 250.8000 177.6000 251.6000 177.7000 ;
	    RECT 255.6000 177.6000 256.4000 177.7000 ;
	    RECT 263.6000 178.3000 264.4000 178.4000 ;
	    RECT 268.4000 178.3000 269.2000 178.4000 ;
	    RECT 263.6000 177.7000 269.2000 178.3000 ;
	    RECT 263.6000 177.6000 264.4000 177.7000 ;
	    RECT 268.4000 177.6000 269.2000 177.7000 ;
	    RECT 274.8000 178.3000 275.6000 178.4000 ;
	    RECT 290.8000 178.3000 291.6000 178.4000 ;
	    RECT 274.8000 177.7000 291.6000 178.3000 ;
	    RECT 274.8000 177.6000 275.6000 177.7000 ;
	    RECT 290.8000 177.6000 291.6000 177.7000 ;
	    RECT 295.6000 178.3000 296.4000 178.4000 ;
	    RECT 316.4000 178.3000 317.2000 178.4000 ;
	    RECT 342.0000 178.3000 342.8000 178.4000 ;
	    RECT 375.6000 178.3000 376.4000 178.4000 ;
	    RECT 295.6000 177.7000 376.4000 178.3000 ;
	    RECT 295.6000 177.6000 296.4000 177.7000 ;
	    RECT 316.4000 177.6000 317.2000 177.7000 ;
	    RECT 342.0000 177.6000 342.8000 177.7000 ;
	    RECT 375.6000 177.6000 376.4000 177.7000 ;
	    RECT 167.6000 176.3000 168.4000 176.4000 ;
	    RECT 95.7000 175.7000 168.4000 176.3000 ;
	    RECT 84.4000 175.6000 85.2000 175.7000 ;
	    RECT 94.0000 175.6000 94.8000 175.7000 ;
	    RECT 167.6000 175.6000 168.4000 175.7000 ;
	    RECT 169.2000 176.3000 170.0000 176.4000 ;
	    RECT 212.4000 176.3000 213.2000 176.4000 ;
	    RECT 169.2000 175.7000 213.2000 176.3000 ;
	    RECT 169.2000 175.6000 170.0000 175.7000 ;
	    RECT 212.4000 175.6000 213.2000 175.7000 ;
	    RECT 215.6000 176.3000 216.4000 176.4000 ;
	    RECT 271.6000 176.3000 272.4000 176.4000 ;
	    RECT 215.6000 175.7000 272.4000 176.3000 ;
	    RECT 290.9000 176.3000 291.5000 177.6000 ;
	    RECT 348.4000 176.3000 349.2000 176.4000 ;
	    RECT 370.8000 176.3000 371.6000 176.4000 ;
	    RECT 434.8000 176.3000 435.6000 176.4000 ;
	    RECT 290.9000 175.7000 435.6000 176.3000 ;
	    RECT 215.6000 175.6000 216.4000 175.7000 ;
	    RECT 271.6000 175.6000 272.4000 175.7000 ;
	    RECT 348.4000 175.6000 349.2000 175.7000 ;
	    RECT 370.8000 175.6000 371.6000 175.7000 ;
	    RECT 434.8000 175.6000 435.6000 175.7000 ;
	    RECT 436.4000 176.3000 437.2000 176.4000 ;
	    RECT 439.6000 176.3000 440.4000 176.4000 ;
	    RECT 436.4000 175.7000 440.4000 176.3000 ;
	    RECT 436.4000 175.6000 437.2000 175.7000 ;
	    RECT 439.6000 175.6000 440.4000 175.7000 ;
	    RECT 450.8000 176.3000 451.6000 176.4000 ;
	    RECT 465.2000 176.3000 466.0000 176.4000 ;
	    RECT 494.0000 176.3000 494.8000 176.4000 ;
	    RECT 450.8000 175.7000 494.8000 176.3000 ;
	    RECT 450.8000 175.6000 451.6000 175.7000 ;
	    RECT 465.2000 175.6000 466.0000 175.7000 ;
	    RECT 494.0000 175.6000 494.8000 175.7000 ;
	    RECT 71.6000 174.3000 72.4000 174.4000 ;
	    RECT 87.6000 174.3000 88.4000 174.4000 ;
	    RECT 111.6000 174.3000 112.4000 174.4000 ;
	    RECT 132.4000 174.3000 133.2000 174.4000 ;
	    RECT 164.4000 174.3000 165.2000 174.4000 ;
	    RECT 71.6000 173.7000 165.2000 174.3000 ;
	    RECT 71.6000 173.6000 72.4000 173.7000 ;
	    RECT 87.6000 173.6000 88.4000 173.7000 ;
	    RECT 111.6000 173.6000 112.4000 173.7000 ;
	    RECT 132.4000 173.6000 133.2000 173.7000 ;
	    RECT 164.4000 173.6000 165.2000 173.7000 ;
	    RECT 183.6000 174.3000 184.4000 174.4000 ;
	    RECT 249.2000 174.3000 250.0000 174.4000 ;
	    RECT 252.4000 174.3000 253.2000 174.4000 ;
	    RECT 183.6000 173.7000 193.9000 174.3000 ;
	    RECT 183.6000 173.6000 184.4000 173.7000 ;
	    RECT 193.3000 172.4000 193.9000 173.7000 ;
	    RECT 249.2000 173.7000 253.2000 174.3000 ;
	    RECT 249.2000 173.6000 250.0000 173.7000 ;
	    RECT 252.4000 173.6000 253.2000 173.7000 ;
	    RECT 254.0000 174.3000 254.8000 174.4000 ;
	    RECT 257.2000 174.3000 258.0000 174.4000 ;
	    RECT 254.0000 173.7000 258.0000 174.3000 ;
	    RECT 254.0000 173.6000 254.8000 173.7000 ;
	    RECT 257.2000 173.6000 258.0000 173.7000 ;
	    RECT 258.8000 174.3000 259.6000 174.4000 ;
	    RECT 287.6000 174.3000 288.4000 174.4000 ;
	    RECT 258.8000 173.7000 288.4000 174.3000 ;
	    RECT 258.8000 173.6000 259.6000 173.7000 ;
	    RECT 287.6000 173.6000 288.4000 173.7000 ;
	    RECT 298.8000 174.3000 299.6000 174.4000 ;
	    RECT 329.2000 174.3000 330.0000 174.4000 ;
	    RECT 298.8000 173.7000 330.0000 174.3000 ;
	    RECT 298.8000 173.6000 299.6000 173.7000 ;
	    RECT 329.2000 173.6000 330.0000 173.7000 ;
	    RECT 334.0000 174.3000 334.8000 174.4000 ;
	    RECT 343.6000 174.3000 344.4000 174.4000 ;
	    RECT 334.0000 173.7000 344.4000 174.3000 ;
	    RECT 334.0000 173.6000 334.8000 173.7000 ;
	    RECT 343.6000 173.6000 344.4000 173.7000 ;
	    RECT 358.0000 174.3000 358.8000 174.4000 ;
	    RECT 367.6000 174.3000 368.4000 174.4000 ;
	    RECT 358.0000 173.7000 368.4000 174.3000 ;
	    RECT 358.0000 173.6000 358.8000 173.7000 ;
	    RECT 367.6000 173.6000 368.4000 173.7000 ;
	    RECT 430.0000 174.3000 430.8000 174.4000 ;
	    RECT 439.6000 174.3000 440.4000 174.4000 ;
	    RECT 430.0000 173.7000 440.4000 174.3000 ;
	    RECT 430.0000 173.6000 430.8000 173.7000 ;
	    RECT 439.6000 173.6000 440.4000 173.7000 ;
	    RECT 447.6000 174.3000 448.4000 174.4000 ;
	    RECT 478.0000 174.3000 478.8000 174.4000 ;
	    RECT 481.2000 174.3000 482.0000 174.4000 ;
	    RECT 447.6000 173.7000 482.0000 174.3000 ;
	    RECT 447.6000 173.6000 448.4000 173.7000 ;
	    RECT 478.0000 173.6000 478.8000 173.7000 ;
	    RECT 481.2000 173.6000 482.0000 173.7000 ;
	    RECT 498.8000 174.3000 499.6000 174.4000 ;
	    RECT 511.6000 174.3000 512.4000 174.4000 ;
	    RECT 498.8000 173.7000 512.4000 174.3000 ;
	    RECT 498.8000 173.6000 499.6000 173.7000 ;
	    RECT 511.6000 173.6000 512.4000 173.7000 ;
	    RECT 12.4000 172.3000 13.2000 172.4000 ;
	    RECT 20.4000 172.3000 21.2000 172.4000 ;
	    RECT 12.4000 171.7000 21.2000 172.3000 ;
	    RECT 12.4000 171.6000 13.2000 171.7000 ;
	    RECT 20.4000 171.6000 21.2000 171.7000 ;
	    RECT 33.2000 172.3000 34.0000 172.4000 ;
	    RECT 58.8000 172.3000 59.6000 172.4000 ;
	    RECT 33.2000 171.7000 59.6000 172.3000 ;
	    RECT 33.2000 171.6000 34.0000 171.7000 ;
	    RECT 58.8000 171.6000 59.6000 171.7000 ;
	    RECT 66.8000 172.3000 67.6000 172.4000 ;
	    RECT 79.6000 172.3000 80.4000 172.4000 ;
	    RECT 66.8000 171.7000 80.4000 172.3000 ;
	    RECT 66.8000 171.6000 67.6000 171.7000 ;
	    RECT 79.6000 171.6000 80.4000 171.7000 ;
	    RECT 94.0000 172.3000 94.8000 172.4000 ;
	    RECT 114.8000 172.3000 115.6000 172.4000 ;
	    RECT 94.0000 171.7000 115.6000 172.3000 ;
	    RECT 94.0000 171.6000 94.8000 171.7000 ;
	    RECT 114.8000 171.6000 115.6000 171.7000 ;
	    RECT 135.6000 172.3000 136.4000 172.4000 ;
	    RECT 146.8000 172.3000 147.6000 172.4000 ;
	    RECT 135.6000 171.7000 147.6000 172.3000 ;
	    RECT 135.6000 171.6000 136.4000 171.7000 ;
	    RECT 146.8000 171.6000 147.6000 171.7000 ;
	    RECT 150.0000 172.3000 150.8000 172.4000 ;
	    RECT 154.8000 172.3000 155.6000 172.4000 ;
	    RECT 150.0000 171.7000 155.6000 172.3000 ;
	    RECT 150.0000 171.6000 150.8000 171.7000 ;
	    RECT 154.8000 171.6000 155.6000 171.7000 ;
	    RECT 159.6000 172.3000 160.4000 172.4000 ;
	    RECT 190.0000 172.3000 190.8000 172.4000 ;
	    RECT 159.6000 171.7000 190.8000 172.3000 ;
	    RECT 159.6000 171.6000 160.4000 171.7000 ;
	    RECT 190.0000 171.6000 190.8000 171.7000 ;
	    RECT 193.2000 171.6000 194.0000 172.4000 ;
	    RECT 202.8000 172.3000 203.6000 172.4000 ;
	    RECT 215.6000 172.3000 216.4000 172.4000 ;
	    RECT 202.8000 171.7000 216.4000 172.3000 ;
	    RECT 202.8000 171.6000 203.6000 171.7000 ;
	    RECT 215.6000 171.6000 216.4000 171.7000 ;
	    RECT 217.2000 172.3000 218.0000 172.4000 ;
	    RECT 222.0000 172.3000 222.8000 172.4000 ;
	    RECT 217.2000 171.7000 222.8000 172.3000 ;
	    RECT 217.2000 171.6000 218.0000 171.7000 ;
	    RECT 222.0000 171.6000 222.8000 171.7000 ;
	    RECT 234.8000 172.3000 235.6000 172.4000 ;
	    RECT 246.0000 172.3000 246.8000 172.4000 ;
	    RECT 234.8000 171.7000 246.8000 172.3000 ;
	    RECT 234.8000 171.6000 235.6000 171.7000 ;
	    RECT 246.0000 171.6000 246.8000 171.7000 ;
	    RECT 340.4000 172.3000 341.2000 172.4000 ;
	    RECT 359.6000 172.3000 360.4000 172.4000 ;
	    RECT 340.4000 171.7000 360.4000 172.3000 ;
	    RECT 340.4000 171.6000 341.2000 171.7000 ;
	    RECT 359.6000 171.6000 360.4000 171.7000 ;
	    RECT 372.4000 172.3000 373.2000 172.4000 ;
	    RECT 388.4000 172.3000 389.2000 172.4000 ;
	    RECT 372.4000 171.7000 389.2000 172.3000 ;
	    RECT 372.4000 171.6000 373.2000 171.7000 ;
	    RECT 388.4000 171.6000 389.2000 171.7000 ;
	    RECT 407.6000 172.3000 408.4000 172.4000 ;
	    RECT 414.0000 172.3000 414.8000 172.4000 ;
	    RECT 407.6000 171.7000 414.8000 172.3000 ;
	    RECT 407.6000 171.6000 408.4000 171.7000 ;
	    RECT 414.0000 171.6000 414.8000 171.7000 ;
	    RECT 455.6000 172.3000 456.4000 172.4000 ;
	    RECT 470.0000 172.3000 470.8000 172.4000 ;
	    RECT 455.6000 171.7000 470.8000 172.3000 ;
	    RECT 455.6000 171.6000 456.4000 171.7000 ;
	    RECT 470.0000 171.6000 470.8000 171.7000 ;
	    RECT 486.0000 172.3000 486.8000 172.4000 ;
	    RECT 505.2000 172.3000 506.0000 172.4000 ;
	    RECT 486.0000 171.7000 506.0000 172.3000 ;
	    RECT 486.0000 171.6000 486.8000 171.7000 ;
	    RECT 505.2000 171.6000 506.0000 171.7000 ;
	    RECT 506.8000 172.3000 507.6000 172.4000 ;
	    RECT 513.2000 172.3000 514.0000 172.4000 ;
	    RECT 506.8000 171.7000 514.0000 172.3000 ;
	    RECT 506.8000 171.6000 507.6000 171.7000 ;
	    RECT 513.2000 171.6000 514.0000 171.7000 ;
	    RECT 17.2000 170.3000 18.0000 170.4000 ;
	    RECT 30.0000 170.3000 30.8000 170.4000 ;
	    RECT 17.2000 169.7000 30.8000 170.3000 ;
	    RECT 17.2000 169.6000 18.0000 169.7000 ;
	    RECT 30.0000 169.6000 30.8000 169.7000 ;
	    RECT 81.2000 170.3000 82.0000 170.4000 ;
	    RECT 129.2000 170.3000 130.0000 170.4000 ;
	    RECT 81.2000 169.7000 130.0000 170.3000 ;
	    RECT 81.2000 169.6000 82.0000 169.7000 ;
	    RECT 129.2000 169.6000 130.0000 169.7000 ;
	    RECT 180.4000 170.3000 181.2000 170.4000 ;
	    RECT 191.6000 170.3000 192.4000 170.4000 ;
	    RECT 180.4000 169.7000 192.4000 170.3000 ;
	    RECT 180.4000 169.6000 181.2000 169.7000 ;
	    RECT 191.6000 169.6000 192.4000 169.7000 ;
	    RECT 202.8000 170.3000 203.6000 170.4000 ;
	    RECT 228.4000 170.3000 229.2000 170.4000 ;
	    RECT 202.8000 169.7000 229.2000 170.3000 ;
	    RECT 202.8000 169.6000 203.6000 169.7000 ;
	    RECT 228.4000 169.6000 229.2000 169.7000 ;
	    RECT 284.4000 170.3000 285.2000 170.4000 ;
	    RECT 310.0000 170.3000 310.8000 170.4000 ;
	    RECT 284.4000 169.7000 310.8000 170.3000 ;
	    RECT 284.4000 169.6000 285.2000 169.7000 ;
	    RECT 310.0000 169.6000 310.8000 169.7000 ;
	    RECT 311.6000 170.3000 312.4000 170.4000 ;
	    RECT 332.4000 170.3000 333.2000 170.4000 ;
	    RECT 311.6000 169.7000 333.2000 170.3000 ;
	    RECT 311.6000 169.6000 312.4000 169.7000 ;
	    RECT 332.4000 169.6000 333.2000 169.7000 ;
	    RECT 351.6000 170.3000 352.4000 170.4000 ;
	    RECT 369.2000 170.3000 370.0000 170.4000 ;
	    RECT 351.6000 169.7000 370.0000 170.3000 ;
	    RECT 351.6000 169.6000 352.4000 169.7000 ;
	    RECT 369.2000 169.6000 370.0000 169.7000 ;
	    RECT 375.6000 170.3000 376.4000 170.4000 ;
	    RECT 390.0000 170.3000 390.8000 170.4000 ;
	    RECT 375.6000 169.7000 390.8000 170.3000 ;
	    RECT 375.6000 169.6000 376.4000 169.7000 ;
	    RECT 390.0000 169.6000 390.8000 169.7000 ;
	    RECT 391.6000 170.3000 392.4000 170.4000 ;
	    RECT 420.4000 170.3000 421.2000 170.4000 ;
	    RECT 391.6000 169.7000 421.2000 170.3000 ;
	    RECT 391.6000 169.6000 392.4000 169.7000 ;
	    RECT 420.4000 169.6000 421.2000 169.7000 ;
	    RECT 426.8000 170.3000 427.6000 170.4000 ;
	    RECT 430.0000 170.3000 430.8000 170.4000 ;
	    RECT 438.0000 170.3000 438.8000 170.4000 ;
	    RECT 447.6000 170.3000 448.4000 170.4000 ;
	    RECT 426.8000 169.7000 448.4000 170.3000 ;
	    RECT 426.8000 169.6000 427.6000 169.7000 ;
	    RECT 430.0000 169.6000 430.8000 169.7000 ;
	    RECT 438.0000 169.6000 438.8000 169.7000 ;
	    RECT 447.6000 169.6000 448.4000 169.7000 ;
	    RECT 460.4000 170.3000 461.2000 170.4000 ;
	    RECT 468.4000 170.3000 469.2000 170.4000 ;
	    RECT 478.0000 170.3000 478.8000 170.4000 ;
	    RECT 489.2000 170.3000 490.0000 170.4000 ;
	    RECT 506.8000 170.3000 507.6000 170.4000 ;
	    RECT 460.4000 169.7000 507.6000 170.3000 ;
	    RECT 460.4000 169.6000 461.2000 169.7000 ;
	    RECT 468.4000 169.6000 469.2000 169.7000 ;
	    RECT 478.0000 169.6000 478.8000 169.7000 ;
	    RECT 489.2000 169.6000 490.0000 169.7000 ;
	    RECT 506.8000 169.6000 507.6000 169.7000 ;
	    RECT 18.8000 168.3000 19.6000 168.4000 ;
	    RECT 28.4000 168.3000 29.2000 168.4000 ;
	    RECT 18.8000 167.7000 29.2000 168.3000 ;
	    RECT 18.8000 167.6000 19.6000 167.7000 ;
	    RECT 28.4000 167.6000 29.2000 167.7000 ;
	    RECT 78.0000 168.3000 78.8000 168.4000 ;
	    RECT 82.8000 168.3000 83.6000 168.4000 ;
	    RECT 86.0000 168.3000 86.8000 168.4000 ;
	    RECT 113.2000 168.3000 114.0000 168.4000 ;
	    RECT 118.0000 168.3000 118.8000 168.4000 ;
	    RECT 78.0000 167.7000 118.8000 168.3000 ;
	    RECT 78.0000 167.6000 78.8000 167.7000 ;
	    RECT 82.8000 167.6000 83.6000 167.7000 ;
	    RECT 86.0000 167.6000 86.8000 167.7000 ;
	    RECT 113.2000 167.6000 114.0000 167.7000 ;
	    RECT 118.0000 167.6000 118.8000 167.7000 ;
	    RECT 140.4000 168.3000 141.2000 168.4000 ;
	    RECT 158.0000 168.3000 158.8000 168.4000 ;
	    RECT 206.0000 168.3000 206.8000 168.4000 ;
	    RECT 262.0000 168.3000 262.8000 168.4000 ;
	    RECT 140.4000 167.7000 262.8000 168.3000 ;
	    RECT 140.4000 167.6000 141.2000 167.7000 ;
	    RECT 158.0000 167.6000 158.8000 167.7000 ;
	    RECT 206.0000 167.6000 206.8000 167.7000 ;
	    RECT 262.0000 167.6000 262.8000 167.7000 ;
	    RECT 266.8000 168.3000 267.6000 168.4000 ;
	    RECT 284.4000 168.3000 285.2000 168.4000 ;
	    RECT 266.8000 167.7000 285.2000 168.3000 ;
	    RECT 266.8000 167.6000 267.6000 167.7000 ;
	    RECT 284.4000 167.6000 285.2000 167.7000 ;
	    RECT 286.0000 168.3000 286.8000 168.4000 ;
	    RECT 289.2000 168.3000 290.0000 168.4000 ;
	    RECT 354.8000 168.3000 355.6000 168.4000 ;
	    RECT 356.4000 168.3000 357.2000 168.4000 ;
	    RECT 361.2000 168.3000 362.0000 168.4000 ;
	    RECT 286.0000 167.7000 362.0000 168.3000 ;
	    RECT 286.0000 167.6000 286.8000 167.7000 ;
	    RECT 289.2000 167.6000 290.0000 167.7000 ;
	    RECT 354.8000 167.6000 355.6000 167.7000 ;
	    RECT 356.4000 167.6000 357.2000 167.7000 ;
	    RECT 361.2000 167.6000 362.0000 167.7000 ;
	    RECT 362.8000 168.3000 363.6000 168.4000 ;
	    RECT 396.4000 168.3000 397.2000 168.4000 ;
	    RECT 362.8000 167.7000 397.2000 168.3000 ;
	    RECT 362.8000 167.6000 363.6000 167.7000 ;
	    RECT 396.4000 167.6000 397.2000 167.7000 ;
	    RECT 401.2000 168.3000 402.0000 168.4000 ;
	    RECT 425.2000 168.3000 426.0000 168.4000 ;
	    RECT 457.2000 168.3000 458.0000 168.4000 ;
	    RECT 401.2000 167.7000 458.0000 168.3000 ;
	    RECT 401.2000 167.6000 402.0000 167.7000 ;
	    RECT 425.2000 167.6000 426.0000 167.7000 ;
	    RECT 457.2000 167.6000 458.0000 167.7000 ;
	    RECT 473.2000 168.3000 474.0000 168.4000 ;
	    RECT 476.4000 168.3000 477.2000 168.4000 ;
	    RECT 487.6000 168.3000 488.4000 168.4000 ;
	    RECT 473.2000 167.7000 488.4000 168.3000 ;
	    RECT 473.2000 167.6000 474.0000 167.7000 ;
	    RECT 476.4000 167.6000 477.2000 167.7000 ;
	    RECT 487.6000 167.6000 488.4000 167.7000 ;
	    RECT 81.2000 166.3000 82.0000 166.4000 ;
	    RECT 164.4000 166.3000 165.2000 166.4000 ;
	    RECT 81.2000 165.7000 165.2000 166.3000 ;
	    RECT 81.2000 165.6000 82.0000 165.7000 ;
	    RECT 164.4000 165.6000 165.2000 165.7000 ;
	    RECT 194.8000 166.3000 195.6000 166.4000 ;
	    RECT 198.0000 166.3000 198.8000 166.4000 ;
	    RECT 206.0000 166.3000 206.8000 166.4000 ;
	    RECT 225.2000 166.3000 226.0000 166.4000 ;
	    RECT 194.8000 165.7000 226.0000 166.3000 ;
	    RECT 194.8000 165.6000 195.6000 165.7000 ;
	    RECT 198.0000 165.6000 198.8000 165.7000 ;
	    RECT 206.0000 165.6000 206.8000 165.7000 ;
	    RECT 225.2000 165.6000 226.0000 165.7000 ;
	    RECT 238.0000 166.3000 238.8000 166.4000 ;
	    RECT 258.8000 166.3000 259.6000 166.4000 ;
	    RECT 238.0000 165.7000 259.6000 166.3000 ;
	    RECT 238.0000 165.6000 238.8000 165.7000 ;
	    RECT 258.8000 165.6000 259.6000 165.7000 ;
	    RECT 260.4000 166.3000 261.2000 166.4000 ;
	    RECT 286.0000 166.3000 286.8000 166.4000 ;
	    RECT 348.4000 166.3000 349.2000 166.4000 ;
	    RECT 353.2000 166.3000 354.0000 166.4000 ;
	    RECT 260.4000 165.7000 286.8000 166.3000 ;
	    RECT 260.4000 165.6000 261.2000 165.7000 ;
	    RECT 286.0000 165.6000 286.8000 165.7000 ;
	    RECT 287.7000 165.7000 344.3000 166.3000 ;
	    RECT 65.2000 164.3000 66.0000 164.4000 ;
	    RECT 124.4000 164.3000 125.2000 164.4000 ;
	    RECT 132.4000 164.3000 133.2000 164.4000 ;
	    RECT 151.6000 164.3000 152.4000 164.4000 ;
	    RECT 159.6000 164.3000 160.4000 164.4000 ;
	    RECT 166.0000 164.3000 166.8000 164.4000 ;
	    RECT 218.8000 164.3000 219.6000 164.4000 ;
	    RECT 65.2000 163.7000 219.6000 164.3000 ;
	    RECT 65.2000 163.6000 66.0000 163.7000 ;
	    RECT 124.4000 163.6000 125.2000 163.7000 ;
	    RECT 132.4000 163.6000 133.2000 163.7000 ;
	    RECT 151.6000 163.6000 152.4000 163.7000 ;
	    RECT 159.6000 163.6000 160.4000 163.7000 ;
	    RECT 166.0000 163.6000 166.8000 163.7000 ;
	    RECT 218.8000 163.6000 219.6000 163.7000 ;
	    RECT 222.0000 164.3000 222.8000 164.4000 ;
	    RECT 234.8000 164.3000 235.6000 164.4000 ;
	    RECT 222.0000 163.7000 235.6000 164.3000 ;
	    RECT 222.0000 163.6000 222.8000 163.7000 ;
	    RECT 234.8000 163.6000 235.6000 163.7000 ;
	    RECT 239.6000 164.3000 240.4000 164.4000 ;
	    RECT 242.8000 164.3000 243.6000 164.4000 ;
	    RECT 239.6000 163.7000 243.6000 164.3000 ;
	    RECT 239.6000 163.6000 240.4000 163.7000 ;
	    RECT 242.8000 163.6000 243.6000 163.7000 ;
	    RECT 244.4000 164.3000 245.2000 164.4000 ;
	    RECT 257.2000 164.3000 258.0000 164.4000 ;
	    RECT 287.7000 164.3000 288.3000 165.7000 ;
	    RECT 244.4000 163.7000 288.3000 164.3000 ;
	    RECT 292.4000 164.3000 293.2000 164.4000 ;
	    RECT 302.0000 164.3000 302.8000 164.4000 ;
	    RECT 322.8000 164.3000 323.6000 164.4000 ;
	    RECT 342.0000 164.3000 342.8000 164.4000 ;
	    RECT 292.4000 163.7000 301.1000 164.3000 ;
	    RECT 244.4000 163.6000 245.2000 163.7000 ;
	    RECT 257.2000 163.6000 258.0000 163.7000 ;
	    RECT 292.4000 163.6000 293.2000 163.7000 ;
	    RECT 54.0000 162.3000 54.8000 162.4000 ;
	    RECT 102.0000 162.3000 102.8000 162.4000 ;
	    RECT 54.0000 161.7000 102.8000 162.3000 ;
	    RECT 54.0000 161.6000 54.8000 161.7000 ;
	    RECT 102.0000 161.6000 102.8000 161.7000 ;
	    RECT 167.6000 162.3000 168.4000 162.4000 ;
	    RECT 263.6000 162.3000 264.4000 162.4000 ;
	    RECT 265.2000 162.3000 266.0000 162.4000 ;
	    RECT 167.6000 161.7000 251.5000 162.3000 ;
	    RECT 167.6000 161.6000 168.4000 161.7000 ;
	    RECT 127.6000 160.3000 128.4000 160.4000 ;
	    RECT 153.2000 160.3000 154.0000 160.4000 ;
	    RECT 127.6000 159.7000 154.0000 160.3000 ;
	    RECT 127.6000 159.6000 128.4000 159.7000 ;
	    RECT 153.2000 159.6000 154.0000 159.7000 ;
	    RECT 164.4000 160.3000 165.2000 160.4000 ;
	    RECT 174.0000 160.3000 174.8000 160.4000 ;
	    RECT 164.4000 159.7000 174.8000 160.3000 ;
	    RECT 164.4000 159.6000 165.2000 159.7000 ;
	    RECT 174.0000 159.6000 174.8000 159.7000 ;
	    RECT 180.4000 160.3000 181.2000 160.4000 ;
	    RECT 190.0000 160.3000 190.8000 160.4000 ;
	    RECT 199.6000 160.3000 200.4000 160.4000 ;
	    RECT 180.4000 159.7000 187.5000 160.3000 ;
	    RECT 180.4000 159.6000 181.2000 159.7000 ;
	    RECT 58.8000 158.3000 59.6000 158.4000 ;
	    RECT 156.4000 158.3000 157.2000 158.4000 ;
	    RECT 185.2000 158.3000 186.0000 158.4000 ;
	    RECT 58.8000 157.7000 144.3000 158.3000 ;
	    RECT 58.8000 157.6000 59.6000 157.7000 ;
	    RECT 143.7000 156.4000 144.3000 157.7000 ;
	    RECT 156.4000 157.7000 186.0000 158.3000 ;
	    RECT 186.9000 158.3000 187.5000 159.7000 ;
	    RECT 190.0000 159.7000 200.4000 160.3000 ;
	    RECT 190.0000 159.6000 190.8000 159.7000 ;
	    RECT 199.6000 159.6000 200.4000 159.7000 ;
	    RECT 201.2000 160.3000 202.0000 160.4000 ;
	    RECT 202.8000 160.3000 203.6000 160.4000 ;
	    RECT 201.2000 159.7000 203.6000 160.3000 ;
	    RECT 201.2000 159.6000 202.0000 159.7000 ;
	    RECT 202.8000 159.6000 203.6000 159.7000 ;
	    RECT 217.2000 160.3000 218.0000 160.4000 ;
	    RECT 222.0000 160.3000 222.8000 160.4000 ;
	    RECT 217.2000 159.7000 222.8000 160.3000 ;
	    RECT 217.2000 159.6000 218.0000 159.7000 ;
	    RECT 222.0000 159.6000 222.8000 159.7000 ;
	    RECT 223.6000 160.3000 224.4000 160.4000 ;
	    RECT 239.6000 160.3000 240.4000 160.4000 ;
	    RECT 223.6000 159.7000 240.4000 160.3000 ;
	    RECT 223.6000 159.6000 224.4000 159.7000 ;
	    RECT 239.6000 159.6000 240.4000 159.7000 ;
	    RECT 242.8000 160.3000 243.6000 160.4000 ;
	    RECT 244.4000 160.3000 245.2000 160.4000 ;
	    RECT 242.8000 159.7000 245.2000 160.3000 ;
	    RECT 242.8000 159.6000 243.6000 159.7000 ;
	    RECT 244.4000 159.6000 245.2000 159.7000 ;
	    RECT 246.0000 160.3000 246.8000 160.4000 ;
	    RECT 249.2000 160.3000 250.0000 160.4000 ;
	    RECT 246.0000 159.7000 250.0000 160.3000 ;
	    RECT 250.9000 160.3000 251.5000 161.7000 ;
	    RECT 263.6000 161.7000 266.0000 162.3000 ;
	    RECT 300.5000 162.3000 301.1000 163.7000 ;
	    RECT 302.0000 163.7000 342.8000 164.3000 ;
	    RECT 343.7000 164.3000 344.3000 165.7000 ;
	    RECT 348.4000 165.7000 354.0000 166.3000 ;
	    RECT 348.4000 165.6000 349.2000 165.7000 ;
	    RECT 353.2000 165.6000 354.0000 165.7000 ;
	    RECT 359.6000 166.3000 360.4000 166.4000 ;
	    RECT 374.0000 166.3000 374.8000 166.4000 ;
	    RECT 359.6000 165.7000 374.8000 166.3000 ;
	    RECT 359.6000 165.6000 360.4000 165.7000 ;
	    RECT 374.0000 165.6000 374.8000 165.7000 ;
	    RECT 380.4000 166.3000 381.2000 166.4000 ;
	    RECT 452.4000 166.3000 453.2000 166.4000 ;
	    RECT 380.4000 165.7000 453.2000 166.3000 ;
	    RECT 380.4000 165.6000 381.2000 165.7000 ;
	    RECT 452.4000 165.6000 453.2000 165.7000 ;
	    RECT 394.8000 164.3000 395.6000 164.4000 ;
	    RECT 343.7000 163.7000 395.6000 164.3000 ;
	    RECT 302.0000 163.6000 302.8000 163.7000 ;
	    RECT 322.8000 163.6000 323.6000 163.7000 ;
	    RECT 342.0000 163.6000 342.8000 163.7000 ;
	    RECT 394.8000 163.6000 395.6000 163.7000 ;
	    RECT 316.4000 162.3000 317.2000 162.4000 ;
	    RECT 300.5000 161.7000 317.2000 162.3000 ;
	    RECT 263.6000 161.6000 264.4000 161.7000 ;
	    RECT 265.2000 161.6000 266.0000 161.7000 ;
	    RECT 316.4000 161.6000 317.2000 161.7000 ;
	    RECT 318.0000 162.3000 318.8000 162.4000 ;
	    RECT 383.6000 162.3000 384.4000 162.4000 ;
	    RECT 318.0000 161.7000 384.4000 162.3000 ;
	    RECT 318.0000 161.6000 318.8000 161.7000 ;
	    RECT 383.6000 161.6000 384.4000 161.7000 ;
	    RECT 250.9000 159.7000 385.9000 160.3000 ;
	    RECT 246.0000 159.6000 246.8000 159.7000 ;
	    RECT 249.2000 159.6000 250.0000 159.7000 ;
	    RECT 194.8000 158.3000 195.6000 158.4000 ;
	    RECT 186.9000 157.7000 195.6000 158.3000 ;
	    RECT 156.4000 157.6000 157.2000 157.7000 ;
	    RECT 185.2000 157.6000 186.0000 157.7000 ;
	    RECT 194.8000 157.6000 195.6000 157.7000 ;
	    RECT 198.0000 158.3000 198.8000 158.4000 ;
	    RECT 212.4000 158.3000 213.2000 158.4000 ;
	    RECT 198.0000 157.7000 213.2000 158.3000 ;
	    RECT 198.0000 157.6000 198.8000 157.7000 ;
	    RECT 212.4000 157.6000 213.2000 157.7000 ;
	    RECT 217.2000 158.3000 218.0000 158.4000 ;
	    RECT 231.6000 158.3000 232.4000 158.4000 ;
	    RECT 241.2000 158.3000 242.0000 158.4000 ;
	    RECT 246.0000 158.3000 246.8000 158.4000 ;
	    RECT 262.0000 158.3000 262.8000 158.4000 ;
	    RECT 281.2000 158.3000 282.0000 158.4000 ;
	    RECT 311.6000 158.3000 312.4000 158.4000 ;
	    RECT 217.2000 157.7000 312.4000 158.3000 ;
	    RECT 217.2000 157.6000 218.0000 157.7000 ;
	    RECT 231.6000 157.6000 232.4000 157.7000 ;
	    RECT 241.2000 157.6000 242.0000 157.7000 ;
	    RECT 246.0000 157.6000 246.8000 157.7000 ;
	    RECT 262.0000 157.6000 262.8000 157.7000 ;
	    RECT 281.2000 157.6000 282.0000 157.7000 ;
	    RECT 311.6000 157.6000 312.4000 157.7000 ;
	    RECT 314.8000 158.3000 315.6000 158.4000 ;
	    RECT 321.2000 158.3000 322.0000 158.4000 ;
	    RECT 314.8000 157.7000 322.0000 158.3000 ;
	    RECT 314.8000 157.6000 315.6000 157.7000 ;
	    RECT 321.2000 157.6000 322.0000 157.7000 ;
	    RECT 326.0000 158.3000 326.8000 158.4000 ;
	    RECT 332.4000 158.3000 333.2000 158.4000 ;
	    RECT 346.8000 158.3000 347.6000 158.4000 ;
	    RECT 377.2000 158.3000 378.0000 158.4000 ;
	    RECT 383.6000 158.3000 384.4000 158.4000 ;
	    RECT 326.0000 157.7000 329.9000 158.3000 ;
	    RECT 326.0000 157.6000 326.8000 157.7000 ;
	    RECT 47.6000 156.3000 48.4000 156.4000 ;
	    RECT 135.6000 156.3000 136.4000 156.4000 ;
	    RECT 47.6000 155.7000 136.4000 156.3000 ;
	    RECT 47.6000 155.6000 48.4000 155.7000 ;
	    RECT 135.6000 155.6000 136.4000 155.7000 ;
	    RECT 143.6000 156.3000 144.4000 156.4000 ;
	    RECT 169.2000 156.3000 170.0000 156.4000 ;
	    RECT 143.6000 155.7000 170.0000 156.3000 ;
	    RECT 143.6000 155.6000 144.4000 155.7000 ;
	    RECT 169.2000 155.6000 170.0000 155.7000 ;
	    RECT 170.8000 156.3000 171.6000 156.4000 ;
	    RECT 174.0000 156.3000 174.8000 156.4000 ;
	    RECT 170.8000 155.7000 174.8000 156.3000 ;
	    RECT 170.8000 155.6000 171.6000 155.7000 ;
	    RECT 174.0000 155.6000 174.8000 155.7000 ;
	    RECT 175.6000 156.3000 176.4000 156.4000 ;
	    RECT 185.2000 156.3000 186.0000 156.4000 ;
	    RECT 175.6000 155.7000 186.0000 156.3000 ;
	    RECT 175.6000 155.6000 176.4000 155.7000 ;
	    RECT 185.2000 155.6000 186.0000 155.7000 ;
	    RECT 191.6000 156.3000 192.4000 156.4000 ;
	    RECT 204.4000 156.3000 205.2000 156.4000 ;
	    RECT 191.6000 155.7000 205.2000 156.3000 ;
	    RECT 191.6000 155.6000 192.4000 155.7000 ;
	    RECT 204.4000 155.6000 205.2000 155.7000 ;
	    RECT 206.0000 156.3000 206.8000 156.4000 ;
	    RECT 228.4000 156.3000 229.2000 156.4000 ;
	    RECT 206.0000 155.7000 229.2000 156.3000 ;
	    RECT 206.0000 155.6000 206.8000 155.7000 ;
	    RECT 228.4000 155.6000 229.2000 155.7000 ;
	    RECT 238.0000 156.3000 238.8000 156.4000 ;
	    RECT 294.0000 156.3000 294.8000 156.4000 ;
	    RECT 238.0000 155.7000 294.8000 156.3000 ;
	    RECT 238.0000 155.6000 238.8000 155.7000 ;
	    RECT 294.0000 155.6000 294.8000 155.7000 ;
	    RECT 295.6000 156.3000 296.4000 156.4000 ;
	    RECT 302.0000 156.3000 302.8000 156.4000 ;
	    RECT 295.6000 155.7000 302.8000 156.3000 ;
	    RECT 295.6000 155.6000 296.4000 155.7000 ;
	    RECT 302.0000 155.6000 302.8000 155.7000 ;
	    RECT 303.6000 156.3000 304.4000 156.4000 ;
	    RECT 327.6000 156.3000 328.4000 156.4000 ;
	    RECT 303.6000 155.7000 328.4000 156.3000 ;
	    RECT 329.3000 156.3000 329.9000 157.7000 ;
	    RECT 332.4000 157.7000 384.4000 158.3000 ;
	    RECT 385.3000 158.3000 385.9000 159.7000 ;
	    RECT 486.0000 158.3000 486.8000 158.4000 ;
	    RECT 385.3000 157.7000 486.8000 158.3000 ;
	    RECT 332.4000 157.6000 333.2000 157.7000 ;
	    RECT 346.8000 157.6000 347.6000 157.7000 ;
	    RECT 377.2000 157.6000 378.0000 157.7000 ;
	    RECT 383.6000 157.6000 384.4000 157.7000 ;
	    RECT 486.0000 157.6000 486.8000 157.7000 ;
	    RECT 334.0000 156.3000 334.8000 156.4000 ;
	    RECT 329.3000 155.7000 334.8000 156.3000 ;
	    RECT 303.6000 155.6000 304.4000 155.7000 ;
	    RECT 327.6000 155.6000 328.4000 155.7000 ;
	    RECT 334.0000 155.6000 334.8000 155.7000 ;
	    RECT 350.0000 156.3000 350.8000 156.4000 ;
	    RECT 364.4000 156.3000 365.2000 156.4000 ;
	    RECT 350.0000 155.7000 365.2000 156.3000 ;
	    RECT 350.0000 155.6000 350.8000 155.7000 ;
	    RECT 364.4000 155.6000 365.2000 155.7000 ;
	    RECT 366.0000 156.3000 366.8000 156.4000 ;
	    RECT 409.2000 156.3000 410.0000 156.4000 ;
	    RECT 366.0000 155.7000 410.0000 156.3000 ;
	    RECT 366.0000 155.6000 366.8000 155.7000 ;
	    RECT 409.2000 155.6000 410.0000 155.7000 ;
	    RECT 70.0000 154.3000 70.8000 154.4000 ;
	    RECT 90.8000 154.3000 91.6000 154.4000 ;
	    RECT 70.0000 153.7000 91.6000 154.3000 ;
	    RECT 70.0000 153.6000 70.8000 153.7000 ;
	    RECT 90.8000 153.6000 91.6000 153.7000 ;
	    RECT 94.0000 154.3000 94.8000 154.4000 ;
	    RECT 111.6000 154.3000 112.4000 154.4000 ;
	    RECT 135.6000 154.3000 136.4000 154.4000 ;
	    RECT 199.6000 154.3000 200.4000 154.4000 ;
	    RECT 222.0000 154.3000 222.8000 154.4000 ;
	    RECT 329.2000 154.3000 330.0000 154.4000 ;
	    RECT 94.0000 153.7000 330.0000 154.3000 ;
	    RECT 94.0000 153.6000 94.8000 153.7000 ;
	    RECT 111.6000 153.6000 112.4000 153.7000 ;
	    RECT 135.6000 153.6000 136.4000 153.7000 ;
	    RECT 199.6000 153.6000 200.4000 153.7000 ;
	    RECT 222.0000 153.6000 222.8000 153.7000 ;
	    RECT 329.2000 153.6000 330.0000 153.7000 ;
	    RECT 330.8000 154.3000 331.6000 154.4000 ;
	    RECT 393.2000 154.3000 394.0000 154.4000 ;
	    RECT 330.8000 153.7000 394.0000 154.3000 ;
	    RECT 330.8000 153.6000 331.6000 153.7000 ;
	    RECT 393.2000 153.6000 394.0000 153.7000 ;
	    RECT 4.4000 152.3000 5.2000 152.4000 ;
	    RECT 20.4000 152.3000 21.2000 152.4000 ;
	    RECT 4.4000 151.7000 21.2000 152.3000 ;
	    RECT 4.4000 151.6000 5.2000 151.7000 ;
	    RECT 20.4000 151.6000 21.2000 151.7000 ;
	    RECT 42.8000 152.3000 43.6000 152.4000 ;
	    RECT 98.8000 152.3000 99.6000 152.4000 ;
	    RECT 42.8000 151.7000 99.6000 152.3000 ;
	    RECT 42.8000 151.6000 43.6000 151.7000 ;
	    RECT 98.8000 151.6000 99.6000 151.7000 ;
	    RECT 108.4000 152.3000 109.2000 152.4000 ;
	    RECT 130.8000 152.3000 131.6000 152.4000 ;
	    RECT 108.4000 151.7000 131.6000 152.3000 ;
	    RECT 108.4000 151.6000 109.2000 151.7000 ;
	    RECT 130.8000 151.6000 131.6000 151.7000 ;
	    RECT 134.0000 152.3000 134.8000 152.4000 ;
	    RECT 140.4000 152.3000 141.2000 152.4000 ;
	    RECT 134.0000 151.7000 141.2000 152.3000 ;
	    RECT 134.0000 151.6000 134.8000 151.7000 ;
	    RECT 140.4000 151.6000 141.2000 151.7000 ;
	    RECT 142.0000 152.3000 142.8000 152.4000 ;
	    RECT 170.8000 152.3000 171.6000 152.4000 ;
	    RECT 142.0000 151.7000 171.6000 152.3000 ;
	    RECT 142.0000 151.6000 142.8000 151.7000 ;
	    RECT 170.8000 151.6000 171.6000 151.7000 ;
	    RECT 174.0000 152.3000 174.8000 152.4000 ;
	    RECT 182.0000 152.3000 182.8000 152.4000 ;
	    RECT 174.0000 151.7000 182.8000 152.3000 ;
	    RECT 174.0000 151.6000 174.8000 151.7000 ;
	    RECT 182.0000 151.6000 182.8000 151.7000 ;
	    RECT 183.6000 152.3000 184.4000 152.4000 ;
	    RECT 188.4000 152.3000 189.2000 152.4000 ;
	    RECT 201.2000 152.3000 202.0000 152.4000 ;
	    RECT 183.6000 151.7000 202.0000 152.3000 ;
	    RECT 183.6000 151.6000 184.4000 151.7000 ;
	    RECT 188.4000 151.6000 189.2000 151.7000 ;
	    RECT 201.2000 151.6000 202.0000 151.7000 ;
	    RECT 209.2000 152.3000 210.0000 152.4000 ;
	    RECT 223.6000 152.3000 224.4000 152.4000 ;
	    RECT 209.2000 151.7000 224.4000 152.3000 ;
	    RECT 209.2000 151.6000 210.0000 151.7000 ;
	    RECT 223.6000 151.6000 224.4000 151.7000 ;
	    RECT 225.2000 152.3000 226.0000 152.4000 ;
	    RECT 233.2000 152.3000 234.0000 152.4000 ;
	    RECT 255.6000 152.3000 256.4000 152.4000 ;
	    RECT 225.2000 151.7000 256.4000 152.3000 ;
	    RECT 225.2000 151.6000 226.0000 151.7000 ;
	    RECT 233.2000 151.6000 234.0000 151.7000 ;
	    RECT 255.6000 151.6000 256.4000 151.7000 ;
	    RECT 258.8000 152.3000 259.6000 152.4000 ;
	    RECT 266.8000 152.3000 267.6000 152.4000 ;
	    RECT 290.8000 152.3000 291.6000 152.4000 ;
	    RECT 258.8000 151.7000 267.6000 152.3000 ;
	    RECT 258.8000 151.6000 259.6000 151.7000 ;
	    RECT 266.8000 151.6000 267.6000 151.7000 ;
	    RECT 268.5000 151.7000 291.6000 152.3000 ;
	    RECT 9.2000 150.3000 10.0000 150.4000 ;
	    RECT 17.2000 150.3000 18.0000 150.4000 ;
	    RECT 33.2000 150.3000 34.0000 150.4000 ;
	    RECT 9.2000 149.7000 34.0000 150.3000 ;
	    RECT 9.2000 149.6000 10.0000 149.7000 ;
	    RECT 17.2000 149.6000 18.0000 149.7000 ;
	    RECT 33.2000 149.6000 34.0000 149.7000 ;
	    RECT 87.6000 150.3000 88.4000 150.4000 ;
	    RECT 92.4000 150.3000 93.2000 150.4000 ;
	    RECT 87.6000 149.7000 93.2000 150.3000 ;
	    RECT 87.6000 149.6000 88.4000 149.7000 ;
	    RECT 92.4000 149.6000 93.2000 149.7000 ;
	    RECT 111.6000 150.3000 112.4000 150.4000 ;
	    RECT 121.2000 150.3000 122.0000 150.4000 ;
	    RECT 111.6000 149.7000 122.0000 150.3000 ;
	    RECT 111.6000 149.6000 112.4000 149.7000 ;
	    RECT 121.2000 149.6000 122.0000 149.7000 ;
	    RECT 122.8000 150.3000 123.6000 150.4000 ;
	    RECT 145.2000 150.3000 146.0000 150.4000 ;
	    RECT 122.8000 149.7000 146.0000 150.3000 ;
	    RECT 122.8000 149.6000 123.6000 149.7000 ;
	    RECT 145.2000 149.6000 146.0000 149.7000 ;
	    RECT 150.0000 150.3000 150.8000 150.4000 ;
	    RECT 158.0000 150.3000 158.8000 150.4000 ;
	    RECT 150.0000 149.7000 158.8000 150.3000 ;
	    RECT 150.0000 149.6000 150.8000 149.7000 ;
	    RECT 158.0000 149.6000 158.8000 149.7000 ;
	    RECT 164.4000 149.6000 165.2000 150.4000 ;
	    RECT 170.8000 149.6000 171.6000 150.4000 ;
	    RECT 172.4000 150.3000 173.2000 150.4000 ;
	    RECT 183.6000 150.3000 184.4000 150.4000 ;
	    RECT 172.4000 149.7000 184.4000 150.3000 ;
	    RECT 172.4000 149.6000 173.2000 149.7000 ;
	    RECT 183.6000 149.6000 184.4000 149.7000 ;
	    RECT 190.0000 150.3000 190.8000 150.4000 ;
	    RECT 194.8000 150.3000 195.6000 150.4000 ;
	    RECT 190.0000 149.7000 195.6000 150.3000 ;
	    RECT 190.0000 149.6000 190.8000 149.7000 ;
	    RECT 194.8000 149.6000 195.6000 149.7000 ;
	    RECT 198.0000 150.3000 198.8000 150.4000 ;
	    RECT 199.6000 150.3000 200.4000 150.4000 ;
	    RECT 215.6000 150.3000 216.4000 150.4000 ;
	    RECT 198.0000 149.7000 216.4000 150.3000 ;
	    RECT 198.0000 149.6000 198.8000 149.7000 ;
	    RECT 199.6000 149.6000 200.4000 149.7000 ;
	    RECT 215.6000 149.6000 216.4000 149.7000 ;
	    RECT 249.2000 150.3000 250.0000 150.4000 ;
	    RECT 268.5000 150.3000 269.1000 151.7000 ;
	    RECT 290.8000 151.6000 291.6000 151.7000 ;
	    RECT 295.6000 152.3000 296.4000 152.4000 ;
	    RECT 300.4000 152.3000 301.2000 152.4000 ;
	    RECT 295.6000 151.7000 301.2000 152.3000 ;
	    RECT 295.6000 151.6000 296.4000 151.7000 ;
	    RECT 300.4000 151.6000 301.2000 151.7000 ;
	    RECT 311.6000 152.3000 312.4000 152.4000 ;
	    RECT 329.2000 152.3000 330.0000 152.4000 ;
	    RECT 311.6000 151.7000 330.0000 152.3000 ;
	    RECT 311.6000 151.6000 312.4000 151.7000 ;
	    RECT 329.2000 151.6000 330.0000 151.7000 ;
	    RECT 337.2000 152.3000 338.0000 152.4000 ;
	    RECT 369.2000 152.3000 370.0000 152.4000 ;
	    RECT 375.6000 152.3000 376.4000 152.4000 ;
	    RECT 337.2000 151.7000 358.7000 152.3000 ;
	    RECT 337.2000 151.6000 338.0000 151.7000 ;
	    RECT 358.1000 150.4000 358.7000 151.7000 ;
	    RECT 369.2000 151.7000 376.4000 152.3000 ;
	    RECT 369.2000 151.6000 370.0000 151.7000 ;
	    RECT 375.6000 151.6000 376.4000 151.7000 ;
	    RECT 431.6000 152.3000 432.4000 152.4000 ;
	    RECT 450.8000 152.3000 451.6000 152.4000 ;
	    RECT 455.6000 152.3000 456.4000 152.4000 ;
	    RECT 431.6000 151.7000 456.4000 152.3000 ;
	    RECT 431.6000 151.6000 432.4000 151.7000 ;
	    RECT 450.8000 151.6000 451.6000 151.7000 ;
	    RECT 455.6000 151.6000 456.4000 151.7000 ;
	    RECT 249.2000 149.7000 269.1000 150.3000 ;
	    RECT 270.0000 150.3000 270.8000 150.4000 ;
	    RECT 276.4000 150.3000 277.2000 150.4000 ;
	    RECT 270.0000 149.7000 277.2000 150.3000 ;
	    RECT 249.2000 149.6000 250.0000 149.7000 ;
	    RECT 270.0000 149.6000 270.8000 149.7000 ;
	    RECT 276.4000 149.6000 277.2000 149.7000 ;
	    RECT 279.6000 149.6000 280.4000 150.4000 ;
	    RECT 284.4000 150.3000 285.2000 150.4000 ;
	    RECT 287.6000 150.3000 288.4000 150.4000 ;
	    RECT 284.4000 149.7000 288.4000 150.3000 ;
	    RECT 284.4000 149.6000 285.2000 149.7000 ;
	    RECT 287.6000 149.6000 288.4000 149.7000 ;
	    RECT 289.2000 150.3000 290.0000 150.4000 ;
	    RECT 294.0000 150.3000 294.8000 150.4000 ;
	    RECT 289.2000 149.7000 294.8000 150.3000 ;
	    RECT 289.2000 149.6000 290.0000 149.7000 ;
	    RECT 294.0000 149.6000 294.8000 149.7000 ;
	    RECT 295.6000 150.3000 296.4000 150.4000 ;
	    RECT 297.2000 150.3000 298.0000 150.4000 ;
	    RECT 295.6000 149.7000 298.0000 150.3000 ;
	    RECT 295.6000 149.6000 296.4000 149.7000 ;
	    RECT 297.2000 149.6000 298.0000 149.7000 ;
	    RECT 305.2000 150.3000 306.0000 150.4000 ;
	    RECT 308.4000 150.3000 309.2000 150.4000 ;
	    RECT 305.2000 149.7000 309.2000 150.3000 ;
	    RECT 305.2000 149.6000 306.0000 149.7000 ;
	    RECT 308.4000 149.6000 309.2000 149.7000 ;
	    RECT 310.0000 150.3000 310.8000 150.4000 ;
	    RECT 324.4000 150.3000 325.2000 150.4000 ;
	    RECT 351.6000 150.3000 352.4000 150.4000 ;
	    RECT 356.4000 150.3000 357.2000 150.4000 ;
	    RECT 310.0000 149.7000 357.2000 150.3000 ;
	    RECT 310.0000 149.6000 310.8000 149.7000 ;
	    RECT 324.4000 149.6000 325.2000 149.7000 ;
	    RECT 351.6000 149.6000 352.4000 149.7000 ;
	    RECT 356.4000 149.6000 357.2000 149.7000 ;
	    RECT 358.0000 150.3000 358.8000 150.4000 ;
	    RECT 366.0000 150.3000 366.8000 150.4000 ;
	    RECT 377.2000 150.3000 378.0000 150.4000 ;
	    RECT 358.0000 149.7000 378.0000 150.3000 ;
	    RECT 358.0000 149.6000 358.8000 149.7000 ;
	    RECT 366.0000 149.6000 366.8000 149.7000 ;
	    RECT 377.2000 149.6000 378.0000 149.7000 ;
	    RECT 398.0000 150.3000 398.8000 150.4000 ;
	    RECT 420.4000 150.3000 421.2000 150.4000 ;
	    RECT 398.0000 149.7000 421.2000 150.3000 ;
	    RECT 398.0000 149.6000 398.8000 149.7000 ;
	    RECT 420.4000 149.6000 421.2000 149.7000 ;
	    RECT 441.2000 150.3000 442.0000 150.4000 ;
	    RECT 450.8000 150.3000 451.6000 150.4000 ;
	    RECT 441.2000 149.7000 451.6000 150.3000 ;
	    RECT 441.2000 149.6000 442.0000 149.7000 ;
	    RECT 450.8000 149.6000 451.6000 149.7000 ;
	    RECT 471.6000 150.3000 472.4000 150.4000 ;
	    RECT 478.0000 150.3000 478.8000 150.4000 ;
	    RECT 471.6000 149.7000 478.8000 150.3000 ;
	    RECT 471.6000 149.6000 472.4000 149.7000 ;
	    RECT 478.0000 149.6000 478.8000 149.7000 ;
	    RECT 481.2000 150.3000 482.0000 150.4000 ;
	    RECT 492.4000 150.3000 493.2000 150.4000 ;
	    RECT 497.2000 150.3000 498.0000 150.4000 ;
	    RECT 503.6000 150.3000 504.4000 150.4000 ;
	    RECT 510.0000 150.3000 510.8000 150.4000 ;
	    RECT 481.2000 149.7000 510.8000 150.3000 ;
	    RECT 481.2000 149.6000 482.0000 149.7000 ;
	    RECT 492.4000 149.6000 493.2000 149.7000 ;
	    RECT 497.2000 149.6000 498.0000 149.7000 ;
	    RECT 503.6000 149.6000 504.4000 149.7000 ;
	    RECT 510.0000 149.6000 510.8000 149.7000 ;
	    RECT 52.4000 148.3000 53.2000 148.4000 ;
	    RECT 62.0000 148.3000 62.8000 148.4000 ;
	    RECT 52.4000 147.7000 62.8000 148.3000 ;
	    RECT 52.4000 147.6000 53.2000 147.7000 ;
	    RECT 62.0000 147.6000 62.8000 147.7000 ;
	    RECT 65.2000 148.3000 66.0000 148.4000 ;
	    RECT 70.0000 148.3000 70.8000 148.4000 ;
	    RECT 65.2000 147.7000 70.8000 148.3000 ;
	    RECT 65.2000 147.6000 66.0000 147.7000 ;
	    RECT 70.0000 147.6000 70.8000 147.7000 ;
	    RECT 97.2000 148.3000 98.0000 148.4000 ;
	    RECT 103.6000 148.3000 104.4000 148.4000 ;
	    RECT 161.2000 148.3000 162.0000 148.4000 ;
	    RECT 209.2000 148.3000 210.0000 148.4000 ;
	    RECT 265.2000 148.3000 266.0000 148.4000 ;
	    RECT 271.6000 148.3000 272.4000 148.4000 ;
	    RECT 97.2000 147.7000 264.3000 148.3000 ;
	    RECT 97.2000 147.6000 98.0000 147.7000 ;
	    RECT 103.6000 147.6000 104.4000 147.7000 ;
	    RECT 161.2000 147.6000 162.0000 147.7000 ;
	    RECT 209.2000 147.6000 210.0000 147.7000 ;
	    RECT 263.7000 146.4000 264.3000 147.7000 ;
	    RECT 265.2000 147.7000 272.4000 148.3000 ;
	    RECT 265.2000 147.6000 266.0000 147.7000 ;
	    RECT 271.6000 147.6000 272.4000 147.7000 ;
	    RECT 287.6000 148.3000 288.4000 148.4000 ;
	    RECT 294.0000 148.3000 294.8000 148.4000 ;
	    RECT 306.8000 148.3000 307.6000 148.4000 ;
	    RECT 319.6000 148.3000 320.4000 148.4000 ;
	    RECT 337.2000 148.3000 338.0000 148.4000 ;
	    RECT 351.6000 148.3000 352.4000 148.4000 ;
	    RECT 287.6000 147.7000 352.4000 148.3000 ;
	    RECT 287.6000 147.6000 288.4000 147.7000 ;
	    RECT 294.0000 147.6000 294.8000 147.7000 ;
	    RECT 306.8000 147.6000 307.6000 147.7000 ;
	    RECT 319.6000 147.6000 320.4000 147.7000 ;
	    RECT 337.2000 147.6000 338.0000 147.7000 ;
	    RECT 351.6000 147.6000 352.4000 147.7000 ;
	    RECT 362.8000 148.3000 363.6000 148.4000 ;
	    RECT 383.6000 148.3000 384.4000 148.4000 ;
	    RECT 362.8000 147.7000 384.4000 148.3000 ;
	    RECT 362.8000 147.6000 363.6000 147.7000 ;
	    RECT 383.6000 147.6000 384.4000 147.7000 ;
	    RECT 425.2000 148.3000 426.0000 148.4000 ;
	    RECT 444.4000 148.3000 445.2000 148.4000 ;
	    RECT 470.0000 148.3000 470.8000 148.4000 ;
	    RECT 425.2000 147.7000 470.8000 148.3000 ;
	    RECT 425.2000 147.6000 426.0000 147.7000 ;
	    RECT 444.4000 147.6000 445.2000 147.7000 ;
	    RECT 470.0000 147.6000 470.8000 147.7000 ;
	    RECT 100.4000 146.3000 101.2000 146.4000 ;
	    RECT 105.2000 146.3000 106.0000 146.4000 ;
	    RECT 116.4000 146.3000 117.2000 146.4000 ;
	    RECT 180.4000 146.3000 181.2000 146.4000 ;
	    RECT 191.6000 146.3000 192.4000 146.4000 ;
	    RECT 201.2000 146.3000 202.0000 146.4000 ;
	    RECT 207.6000 146.3000 208.4000 146.4000 ;
	    RECT 100.4000 145.7000 208.4000 146.3000 ;
	    RECT 100.4000 145.6000 101.2000 145.7000 ;
	    RECT 105.2000 145.6000 106.0000 145.7000 ;
	    RECT 116.4000 145.6000 117.2000 145.7000 ;
	    RECT 180.4000 145.6000 181.2000 145.7000 ;
	    RECT 191.6000 145.6000 192.4000 145.7000 ;
	    RECT 201.2000 145.6000 202.0000 145.7000 ;
	    RECT 207.6000 145.6000 208.4000 145.7000 ;
	    RECT 215.6000 146.3000 216.4000 146.4000 ;
	    RECT 228.4000 146.3000 229.2000 146.4000 ;
	    RECT 215.6000 145.7000 229.2000 146.3000 ;
	    RECT 215.6000 145.6000 216.4000 145.7000 ;
	    RECT 228.4000 145.6000 229.2000 145.7000 ;
	    RECT 234.8000 146.3000 235.6000 146.4000 ;
	    RECT 260.4000 146.3000 261.2000 146.4000 ;
	    RECT 234.8000 145.7000 261.2000 146.3000 ;
	    RECT 234.8000 145.6000 235.6000 145.7000 ;
	    RECT 260.4000 145.6000 261.2000 145.7000 ;
	    RECT 263.6000 146.3000 264.4000 146.4000 ;
	    RECT 362.9000 146.3000 363.5000 147.6000 ;
	    RECT 263.6000 145.7000 363.5000 146.3000 ;
	    RECT 374.0000 146.3000 374.8000 146.4000 ;
	    RECT 374.0000 145.7000 429.1000 146.3000 ;
	    RECT 263.6000 145.6000 264.4000 145.7000 ;
	    RECT 374.0000 145.6000 374.8000 145.7000 ;
	    RECT 428.5000 144.4000 429.1000 145.7000 ;
	    RECT 66.8000 144.3000 67.6000 144.4000 ;
	    RECT 87.6000 144.3000 88.4000 144.4000 ;
	    RECT 66.8000 143.7000 88.4000 144.3000 ;
	    RECT 66.8000 143.6000 67.6000 143.7000 ;
	    RECT 87.6000 143.6000 88.4000 143.7000 ;
	    RECT 102.0000 144.3000 102.8000 144.4000 ;
	    RECT 116.4000 144.3000 117.2000 144.4000 ;
	    RECT 102.0000 143.7000 117.2000 144.3000 ;
	    RECT 102.0000 143.6000 102.8000 143.7000 ;
	    RECT 116.4000 143.6000 117.2000 143.7000 ;
	    RECT 118.0000 144.3000 118.8000 144.4000 ;
	    RECT 202.8000 144.3000 203.6000 144.4000 ;
	    RECT 244.4000 144.3000 245.2000 144.4000 ;
	    RECT 118.0000 143.7000 245.2000 144.3000 ;
	    RECT 118.0000 143.6000 118.8000 143.7000 ;
	    RECT 202.8000 143.6000 203.6000 143.7000 ;
	    RECT 244.4000 143.6000 245.2000 143.7000 ;
	    RECT 250.8000 144.3000 251.6000 144.4000 ;
	    RECT 266.8000 144.3000 267.6000 144.4000 ;
	    RECT 286.0000 144.3000 286.8000 144.4000 ;
	    RECT 250.8000 143.7000 286.8000 144.3000 ;
	    RECT 250.8000 143.6000 251.6000 143.7000 ;
	    RECT 266.8000 143.6000 267.6000 143.7000 ;
	    RECT 286.0000 143.6000 286.8000 143.7000 ;
	    RECT 287.6000 144.3000 288.4000 144.4000 ;
	    RECT 318.0000 144.3000 318.8000 144.4000 ;
	    RECT 287.6000 143.7000 318.8000 144.3000 ;
	    RECT 287.6000 143.6000 288.4000 143.7000 ;
	    RECT 318.0000 143.6000 318.8000 143.7000 ;
	    RECT 324.4000 144.3000 325.2000 144.4000 ;
	    RECT 340.4000 144.3000 341.2000 144.4000 ;
	    RECT 324.4000 143.7000 341.2000 144.3000 ;
	    RECT 324.4000 143.6000 325.2000 143.7000 ;
	    RECT 340.4000 143.6000 341.2000 143.7000 ;
	    RECT 345.2000 144.3000 346.0000 144.4000 ;
	    RECT 353.2000 144.3000 354.0000 144.4000 ;
	    RECT 345.2000 143.7000 354.0000 144.3000 ;
	    RECT 345.2000 143.6000 346.0000 143.7000 ;
	    RECT 353.2000 143.6000 354.0000 143.7000 ;
	    RECT 385.2000 143.6000 386.0000 144.4000 ;
	    RECT 428.4000 144.3000 429.2000 144.4000 ;
	    RECT 447.6000 144.3000 448.4000 144.4000 ;
	    RECT 428.4000 143.7000 448.4000 144.3000 ;
	    RECT 428.4000 143.6000 429.2000 143.7000 ;
	    RECT 447.6000 143.6000 448.4000 143.7000 ;
	    RECT 450.8000 144.3000 451.6000 144.4000 ;
	    RECT 458.8000 144.3000 459.6000 144.4000 ;
	    RECT 486.0000 144.3000 486.8000 144.4000 ;
	    RECT 450.8000 143.7000 486.8000 144.3000 ;
	    RECT 450.8000 143.6000 451.6000 143.7000 ;
	    RECT 458.8000 143.6000 459.6000 143.7000 ;
	    RECT 486.0000 143.6000 486.8000 143.7000 ;
	    RECT 68.4000 142.3000 69.2000 142.4000 ;
	    RECT 79.6000 142.3000 80.4000 142.4000 ;
	    RECT 68.4000 141.7000 80.4000 142.3000 ;
	    RECT 68.4000 141.6000 69.2000 141.7000 ;
	    RECT 79.6000 141.6000 80.4000 141.7000 ;
	    RECT 95.6000 142.3000 96.4000 142.4000 ;
	    RECT 108.4000 142.3000 109.2000 142.4000 ;
	    RECT 95.6000 141.7000 109.2000 142.3000 ;
	    RECT 95.6000 141.6000 96.4000 141.7000 ;
	    RECT 108.4000 141.6000 109.2000 141.7000 ;
	    RECT 110.0000 142.3000 110.8000 142.4000 ;
	    RECT 132.4000 142.3000 133.2000 142.4000 ;
	    RECT 110.0000 141.7000 133.2000 142.3000 ;
	    RECT 110.0000 141.6000 110.8000 141.7000 ;
	    RECT 132.4000 141.6000 133.2000 141.7000 ;
	    RECT 134.0000 142.3000 134.8000 142.4000 ;
	    RECT 142.0000 142.3000 142.8000 142.4000 ;
	    RECT 134.0000 141.7000 142.8000 142.3000 ;
	    RECT 134.0000 141.6000 134.8000 141.7000 ;
	    RECT 142.0000 141.6000 142.8000 141.7000 ;
	    RECT 167.6000 142.3000 168.4000 142.4000 ;
	    RECT 172.4000 142.3000 173.2000 142.4000 ;
	    RECT 167.6000 141.7000 173.2000 142.3000 ;
	    RECT 167.6000 141.6000 168.4000 141.7000 ;
	    RECT 172.4000 141.6000 173.2000 141.7000 ;
	    RECT 174.0000 142.3000 174.8000 142.4000 ;
	    RECT 180.4000 142.3000 181.2000 142.4000 ;
	    RECT 174.0000 141.7000 181.2000 142.3000 ;
	    RECT 174.0000 141.6000 174.8000 141.7000 ;
	    RECT 180.4000 141.6000 181.2000 141.7000 ;
	    RECT 188.4000 142.3000 189.2000 142.4000 ;
	    RECT 194.8000 142.3000 195.6000 142.4000 ;
	    RECT 188.4000 141.7000 195.6000 142.3000 ;
	    RECT 188.4000 141.6000 189.2000 141.7000 ;
	    RECT 194.8000 141.6000 195.6000 141.7000 ;
	    RECT 198.0000 142.3000 198.8000 142.4000 ;
	    RECT 249.2000 142.3000 250.0000 142.4000 ;
	    RECT 198.0000 141.7000 250.0000 142.3000 ;
	    RECT 198.0000 141.6000 198.8000 141.7000 ;
	    RECT 249.2000 141.6000 250.0000 141.7000 ;
	    RECT 266.8000 142.3000 267.6000 142.4000 ;
	    RECT 289.2000 142.3000 290.0000 142.4000 ;
	    RECT 266.8000 141.7000 290.0000 142.3000 ;
	    RECT 266.8000 141.6000 267.6000 141.7000 ;
	    RECT 289.2000 141.6000 290.0000 141.7000 ;
	    RECT 292.4000 142.3000 293.2000 142.4000 ;
	    RECT 295.6000 142.3000 296.4000 142.4000 ;
	    RECT 292.4000 141.7000 296.4000 142.3000 ;
	    RECT 292.4000 141.6000 293.2000 141.7000 ;
	    RECT 295.6000 141.6000 296.4000 141.7000 ;
	    RECT 297.2000 142.3000 298.0000 142.4000 ;
	    RECT 318.0000 142.3000 318.8000 142.4000 ;
	    RECT 297.2000 141.7000 318.8000 142.3000 ;
	    RECT 297.2000 141.6000 298.0000 141.7000 ;
	    RECT 318.0000 141.6000 318.8000 141.7000 ;
	    RECT 330.8000 142.3000 331.6000 142.4000 ;
	    RECT 348.4000 142.3000 349.2000 142.4000 ;
	    RECT 330.8000 141.7000 349.2000 142.3000 ;
	    RECT 330.8000 141.6000 331.6000 141.7000 ;
	    RECT 348.4000 141.6000 349.2000 141.7000 ;
	    RECT 356.4000 142.3000 357.2000 142.4000 ;
	    RECT 369.2000 142.3000 370.0000 142.4000 ;
	    RECT 372.4000 142.3000 373.2000 142.4000 ;
	    RECT 356.4000 141.7000 373.2000 142.3000 ;
	    RECT 356.4000 141.6000 357.2000 141.7000 ;
	    RECT 369.2000 141.6000 370.0000 141.7000 ;
	    RECT 372.4000 141.6000 373.2000 141.7000 ;
	    RECT 375.6000 142.3000 376.4000 142.4000 ;
	    RECT 414.0000 142.3000 414.8000 142.4000 ;
	    RECT 375.6000 141.7000 414.8000 142.3000 ;
	    RECT 375.6000 141.6000 376.4000 141.7000 ;
	    RECT 414.0000 141.6000 414.8000 141.7000 ;
	    RECT 65.2000 140.3000 66.0000 140.4000 ;
	    RECT 82.8000 140.3000 83.6000 140.4000 ;
	    RECT 65.2000 139.7000 83.6000 140.3000 ;
	    RECT 65.2000 139.6000 66.0000 139.7000 ;
	    RECT 82.8000 139.6000 83.6000 139.7000 ;
	    RECT 87.6000 140.3000 88.4000 140.4000 ;
	    RECT 226.8000 140.3000 227.6000 140.4000 ;
	    RECT 87.6000 139.7000 227.6000 140.3000 ;
	    RECT 87.6000 139.6000 88.4000 139.7000 ;
	    RECT 226.8000 139.6000 227.6000 139.7000 ;
	    RECT 228.4000 140.3000 229.2000 140.4000 ;
	    RECT 250.8000 140.3000 251.6000 140.4000 ;
	    RECT 228.4000 139.7000 251.6000 140.3000 ;
	    RECT 228.4000 139.6000 229.2000 139.7000 ;
	    RECT 250.8000 139.6000 251.6000 139.7000 ;
	    RECT 266.8000 140.3000 267.6000 140.4000 ;
	    RECT 281.2000 140.3000 282.0000 140.4000 ;
	    RECT 266.8000 139.7000 282.0000 140.3000 ;
	    RECT 266.8000 139.6000 267.6000 139.7000 ;
	    RECT 281.2000 139.6000 282.0000 139.7000 ;
	    RECT 287.6000 140.3000 288.4000 140.4000 ;
	    RECT 292.4000 140.3000 293.2000 140.4000 ;
	    RECT 287.6000 139.7000 293.2000 140.3000 ;
	    RECT 287.6000 139.6000 288.4000 139.7000 ;
	    RECT 292.4000 139.6000 293.2000 139.7000 ;
	    RECT 295.6000 140.3000 296.4000 140.4000 ;
	    RECT 302.0000 140.3000 302.8000 140.4000 ;
	    RECT 295.6000 139.7000 302.8000 140.3000 ;
	    RECT 295.6000 139.6000 296.4000 139.7000 ;
	    RECT 302.0000 139.6000 302.8000 139.7000 ;
	    RECT 311.6000 139.6000 312.4000 140.4000 ;
	    RECT 313.2000 140.3000 314.0000 140.4000 ;
	    RECT 364.4000 140.3000 365.2000 140.4000 ;
	    RECT 377.2000 140.3000 378.0000 140.4000 ;
	    RECT 313.2000 139.7000 365.2000 140.3000 ;
	    RECT 313.2000 139.6000 314.0000 139.7000 ;
	    RECT 364.4000 139.6000 365.2000 139.7000 ;
	    RECT 366.1000 139.7000 378.0000 140.3000 ;
	    RECT 4.4000 138.3000 5.2000 138.4000 ;
	    RECT 10.8000 138.3000 11.6000 138.4000 ;
	    RECT 30.0000 138.3000 30.8000 138.4000 ;
	    RECT 4.4000 137.7000 30.8000 138.3000 ;
	    RECT 4.4000 137.6000 5.2000 137.7000 ;
	    RECT 10.8000 137.6000 11.6000 137.7000 ;
	    RECT 30.0000 137.6000 30.8000 137.7000 ;
	    RECT 78.0000 138.3000 78.8000 138.4000 ;
	    RECT 84.4000 138.3000 85.2000 138.4000 ;
	    RECT 132.4000 138.3000 133.2000 138.4000 ;
	    RECT 151.6000 138.3000 152.4000 138.4000 ;
	    RECT 78.0000 137.7000 152.4000 138.3000 ;
	    RECT 78.0000 137.6000 78.8000 137.7000 ;
	    RECT 84.4000 137.6000 85.2000 137.7000 ;
	    RECT 132.4000 137.6000 133.2000 137.7000 ;
	    RECT 151.6000 137.6000 152.4000 137.7000 ;
	    RECT 154.8000 138.3000 155.6000 138.4000 ;
	    RECT 172.4000 138.3000 173.2000 138.4000 ;
	    RECT 154.8000 137.7000 173.2000 138.3000 ;
	    RECT 154.8000 137.6000 155.6000 137.7000 ;
	    RECT 172.4000 137.6000 173.2000 137.7000 ;
	    RECT 174.0000 138.3000 174.8000 138.4000 ;
	    RECT 177.2000 138.3000 178.0000 138.4000 ;
	    RECT 178.8000 138.3000 179.6000 138.4000 ;
	    RECT 174.0000 137.7000 179.6000 138.3000 ;
	    RECT 174.0000 137.6000 174.8000 137.7000 ;
	    RECT 177.2000 137.6000 178.0000 137.7000 ;
	    RECT 178.8000 137.6000 179.6000 137.7000 ;
	    RECT 193.2000 138.3000 194.0000 138.4000 ;
	    RECT 199.6000 138.3000 200.4000 138.4000 ;
	    RECT 206.0000 138.3000 206.8000 138.4000 ;
	    RECT 228.4000 138.3000 229.2000 138.4000 ;
	    RECT 241.2000 138.3000 242.0000 138.4000 ;
	    RECT 193.2000 137.7000 227.5000 138.3000 ;
	    RECT 193.2000 137.6000 194.0000 137.7000 ;
	    RECT 199.6000 137.6000 200.4000 137.7000 ;
	    RECT 206.0000 137.6000 206.8000 137.7000 ;
	    RECT 23.6000 136.3000 24.4000 136.4000 ;
	    RECT 62.0000 136.3000 62.8000 136.4000 ;
	    RECT 23.6000 135.7000 62.8000 136.3000 ;
	    RECT 23.6000 135.6000 24.4000 135.7000 ;
	    RECT 62.0000 135.6000 62.8000 135.7000 ;
	    RECT 74.8000 136.3000 75.6000 136.4000 ;
	    RECT 79.6000 136.3000 80.4000 136.4000 ;
	    RECT 74.8000 135.7000 80.4000 136.3000 ;
	    RECT 74.8000 135.6000 75.6000 135.7000 ;
	    RECT 79.6000 135.6000 80.4000 135.7000 ;
	    RECT 81.2000 136.3000 82.0000 136.4000 ;
	    RECT 110.0000 136.3000 110.8000 136.4000 ;
	    RECT 81.2000 135.7000 110.8000 136.3000 ;
	    RECT 81.2000 135.6000 82.0000 135.7000 ;
	    RECT 110.0000 135.6000 110.8000 135.7000 ;
	    RECT 113.2000 136.3000 114.0000 136.4000 ;
	    RECT 145.2000 136.3000 146.0000 136.4000 ;
	    RECT 150.0000 136.3000 150.8000 136.4000 ;
	    RECT 180.4000 136.3000 181.2000 136.4000 ;
	    RECT 113.2000 135.7000 144.3000 136.3000 ;
	    RECT 113.2000 135.6000 114.0000 135.7000 ;
	    RECT 14.0000 134.3000 14.8000 134.4000 ;
	    RECT 34.8000 134.3000 35.6000 134.4000 ;
	    RECT 14.0000 133.7000 35.6000 134.3000 ;
	    RECT 14.0000 133.6000 14.8000 133.7000 ;
	    RECT 34.8000 133.6000 35.6000 133.7000 ;
	    RECT 68.4000 134.3000 69.2000 134.4000 ;
	    RECT 78.0000 134.3000 78.8000 134.4000 ;
	    RECT 68.4000 133.7000 78.8000 134.3000 ;
	    RECT 68.4000 133.6000 69.2000 133.7000 ;
	    RECT 78.0000 133.6000 78.8000 133.7000 ;
	    RECT 89.2000 134.3000 90.0000 134.4000 ;
	    RECT 97.2000 134.3000 98.0000 134.4000 ;
	    RECT 89.2000 133.7000 98.0000 134.3000 ;
	    RECT 89.2000 133.6000 90.0000 133.7000 ;
	    RECT 97.2000 133.6000 98.0000 133.7000 ;
	    RECT 114.8000 134.3000 115.6000 134.4000 ;
	    RECT 121.2000 134.3000 122.0000 134.4000 ;
	    RECT 114.8000 133.7000 122.0000 134.3000 ;
	    RECT 114.8000 133.6000 115.6000 133.7000 ;
	    RECT 121.2000 133.6000 122.0000 133.7000 ;
	    RECT 134.0000 134.3000 134.8000 134.4000 ;
	    RECT 142.0000 134.3000 142.8000 134.4000 ;
	    RECT 134.0000 133.7000 142.8000 134.3000 ;
	    RECT 143.7000 134.3000 144.3000 135.7000 ;
	    RECT 145.2000 135.7000 181.2000 136.3000 ;
	    RECT 145.2000 135.6000 146.0000 135.7000 ;
	    RECT 150.0000 135.6000 150.8000 135.7000 ;
	    RECT 180.4000 135.6000 181.2000 135.7000 ;
	    RECT 186.8000 136.3000 187.6000 136.4000 ;
	    RECT 218.8000 136.3000 219.6000 136.4000 ;
	    RECT 186.8000 135.7000 219.6000 136.3000 ;
	    RECT 226.9000 136.3000 227.5000 137.7000 ;
	    RECT 228.4000 137.7000 242.0000 138.3000 ;
	    RECT 228.4000 137.6000 229.2000 137.7000 ;
	    RECT 241.2000 137.6000 242.0000 137.7000 ;
	    RECT 242.8000 138.3000 243.6000 138.4000 ;
	    RECT 247.6000 138.3000 248.4000 138.4000 ;
	    RECT 242.8000 137.7000 248.4000 138.3000 ;
	    RECT 242.8000 137.6000 243.6000 137.7000 ;
	    RECT 247.6000 137.6000 248.4000 137.7000 ;
	    RECT 249.2000 138.3000 250.0000 138.4000 ;
	    RECT 268.4000 138.3000 269.2000 138.4000 ;
	    RECT 249.2000 137.7000 269.2000 138.3000 ;
	    RECT 249.2000 137.6000 250.0000 137.7000 ;
	    RECT 268.4000 137.6000 269.2000 137.7000 ;
	    RECT 271.6000 138.3000 272.4000 138.4000 ;
	    RECT 278.0000 138.3000 278.8000 138.4000 ;
	    RECT 271.6000 137.7000 278.8000 138.3000 ;
	    RECT 271.6000 137.6000 272.4000 137.7000 ;
	    RECT 278.0000 137.6000 278.8000 137.7000 ;
	    RECT 282.8000 138.3000 283.6000 138.4000 ;
	    RECT 305.2000 138.3000 306.0000 138.4000 ;
	    RECT 308.4000 138.3000 309.2000 138.4000 ;
	    RECT 282.8000 137.7000 309.2000 138.3000 ;
	    RECT 282.8000 137.6000 283.6000 137.7000 ;
	    RECT 305.2000 137.6000 306.0000 137.7000 ;
	    RECT 308.4000 137.6000 309.2000 137.7000 ;
	    RECT 318.0000 138.3000 318.8000 138.4000 ;
	    RECT 326.0000 138.3000 326.8000 138.4000 ;
	    RECT 318.0000 137.7000 326.8000 138.3000 ;
	    RECT 318.0000 137.6000 318.8000 137.7000 ;
	    RECT 326.0000 137.6000 326.8000 137.7000 ;
	    RECT 327.6000 138.3000 328.4000 138.4000 ;
	    RECT 366.1000 138.3000 366.7000 139.7000 ;
	    RECT 377.2000 139.6000 378.0000 139.7000 ;
	    RECT 422.0000 140.3000 422.8000 140.4000 ;
	    RECT 433.2000 140.3000 434.0000 140.4000 ;
	    RECT 444.4000 140.3000 445.2000 140.4000 ;
	    RECT 422.0000 139.7000 445.2000 140.3000 ;
	    RECT 422.0000 139.6000 422.8000 139.7000 ;
	    RECT 433.2000 139.6000 434.0000 139.7000 ;
	    RECT 444.4000 139.6000 445.2000 139.7000 ;
	    RECT 487.6000 140.3000 488.4000 140.4000 ;
	    RECT 511.6000 140.3000 512.4000 140.4000 ;
	    RECT 487.6000 139.7000 512.4000 140.3000 ;
	    RECT 487.6000 139.6000 488.4000 139.7000 ;
	    RECT 511.6000 139.6000 512.4000 139.7000 ;
	    RECT 327.6000 137.7000 366.7000 138.3000 ;
	    RECT 370.8000 138.3000 371.6000 138.4000 ;
	    RECT 378.8000 138.3000 379.6000 138.4000 ;
	    RECT 473.2000 138.3000 474.0000 138.4000 ;
	    RECT 492.4000 138.3000 493.2000 138.4000 ;
	    RECT 370.8000 137.7000 493.2000 138.3000 ;
	    RECT 327.6000 137.6000 328.4000 137.7000 ;
	    RECT 370.8000 137.6000 371.6000 137.7000 ;
	    RECT 378.8000 137.6000 379.6000 137.7000 ;
	    RECT 473.2000 137.6000 474.0000 137.7000 ;
	    RECT 492.4000 137.6000 493.2000 137.7000 ;
	    RECT 265.2000 136.3000 266.0000 136.4000 ;
	    RECT 226.9000 135.7000 266.0000 136.3000 ;
	    RECT 186.8000 135.6000 187.6000 135.7000 ;
	    RECT 218.8000 135.6000 219.6000 135.7000 ;
	    RECT 265.2000 135.6000 266.0000 135.7000 ;
	    RECT 270.0000 136.3000 270.8000 136.4000 ;
	    RECT 292.4000 136.3000 293.2000 136.4000 ;
	    RECT 270.0000 135.7000 293.2000 136.3000 ;
	    RECT 270.0000 135.6000 270.8000 135.7000 ;
	    RECT 292.4000 135.6000 293.2000 135.7000 ;
	    RECT 295.6000 136.3000 296.4000 136.4000 ;
	    RECT 303.6000 136.3000 304.4000 136.4000 ;
	    RECT 295.6000 135.7000 304.4000 136.3000 ;
	    RECT 295.6000 135.6000 296.4000 135.7000 ;
	    RECT 303.6000 135.6000 304.4000 135.7000 ;
	    RECT 305.2000 136.3000 306.0000 136.4000 ;
	    RECT 313.2000 136.3000 314.0000 136.4000 ;
	    RECT 305.2000 135.7000 314.0000 136.3000 ;
	    RECT 305.2000 135.6000 306.0000 135.7000 ;
	    RECT 313.2000 135.6000 314.0000 135.7000 ;
	    RECT 316.4000 136.3000 317.2000 136.4000 ;
	    RECT 321.2000 136.3000 322.0000 136.4000 ;
	    RECT 316.4000 135.7000 322.0000 136.3000 ;
	    RECT 316.4000 135.6000 317.2000 135.7000 ;
	    RECT 321.2000 135.6000 322.0000 135.7000 ;
	    RECT 343.6000 136.3000 344.4000 136.4000 ;
	    RECT 350.0000 136.3000 350.8000 136.4000 ;
	    RECT 343.6000 135.7000 350.8000 136.3000 ;
	    RECT 343.6000 135.6000 344.4000 135.7000 ;
	    RECT 350.0000 135.6000 350.8000 135.7000 ;
	    RECT 354.8000 136.3000 355.6000 136.4000 ;
	    RECT 359.6000 136.3000 360.4000 136.4000 ;
	    RECT 354.8000 135.7000 360.4000 136.3000 ;
	    RECT 354.8000 135.6000 355.6000 135.7000 ;
	    RECT 359.6000 135.6000 360.4000 135.7000 ;
	    RECT 361.2000 136.3000 362.0000 136.4000 ;
	    RECT 391.6000 136.3000 392.4000 136.4000 ;
	    RECT 361.2000 135.7000 392.4000 136.3000 ;
	    RECT 361.2000 135.6000 362.0000 135.7000 ;
	    RECT 391.6000 135.6000 392.4000 135.7000 ;
	    RECT 412.4000 136.3000 413.2000 136.4000 ;
	    RECT 434.8000 136.3000 435.6000 136.4000 ;
	    RECT 412.4000 135.7000 435.6000 136.3000 ;
	    RECT 412.4000 135.6000 413.2000 135.7000 ;
	    RECT 434.8000 135.6000 435.6000 135.7000 ;
	    RECT 502.0000 136.3000 502.8000 136.4000 ;
	    RECT 506.8000 136.3000 507.6000 136.4000 ;
	    RECT 502.0000 135.7000 507.6000 136.3000 ;
	    RECT 502.0000 135.6000 502.8000 135.7000 ;
	    RECT 506.8000 135.6000 507.6000 135.7000 ;
	    RECT 174.0000 134.3000 174.8000 134.4000 ;
	    RECT 143.7000 133.7000 174.8000 134.3000 ;
	    RECT 134.0000 133.6000 134.8000 133.7000 ;
	    RECT 142.0000 133.6000 142.8000 133.7000 ;
	    RECT 174.0000 133.6000 174.8000 133.7000 ;
	    RECT 204.4000 134.3000 205.2000 134.4000 ;
	    RECT 225.2000 134.3000 226.0000 134.4000 ;
	    RECT 260.4000 134.3000 261.2000 134.4000 ;
	    RECT 204.4000 133.7000 261.2000 134.3000 ;
	    RECT 204.4000 133.6000 205.2000 133.7000 ;
	    RECT 225.2000 133.6000 226.0000 133.7000 ;
	    RECT 260.4000 133.6000 261.2000 133.7000 ;
	    RECT 263.6000 134.3000 264.4000 134.4000 ;
	    RECT 270.0000 134.3000 270.8000 134.4000 ;
	    RECT 297.2000 134.3000 298.0000 134.4000 ;
	    RECT 263.6000 133.7000 267.5000 134.3000 ;
	    RECT 263.6000 133.6000 264.4000 133.7000 ;
	    RECT 266.9000 132.4000 267.5000 133.7000 ;
	    RECT 270.0000 133.7000 298.0000 134.3000 ;
	    RECT 270.0000 133.6000 270.8000 133.7000 ;
	    RECT 297.2000 133.6000 298.0000 133.7000 ;
	    RECT 300.4000 134.3000 301.2000 134.4000 ;
	    RECT 305.2000 134.3000 306.0000 134.4000 ;
	    RECT 300.4000 133.7000 306.0000 134.3000 ;
	    RECT 300.4000 133.6000 301.2000 133.7000 ;
	    RECT 305.2000 133.6000 306.0000 133.7000 ;
	    RECT 308.4000 134.3000 309.2000 134.4000 ;
	    RECT 330.8000 134.3000 331.6000 134.4000 ;
	    RECT 338.8000 134.3000 339.6000 134.4000 ;
	    RECT 362.8000 134.3000 363.6000 134.4000 ;
	    RECT 308.4000 133.7000 363.6000 134.3000 ;
	    RECT 308.4000 133.6000 309.2000 133.7000 ;
	    RECT 330.8000 133.6000 331.6000 133.7000 ;
	    RECT 338.8000 133.6000 339.6000 133.7000 ;
	    RECT 362.8000 133.6000 363.6000 133.7000 ;
	    RECT 398.0000 134.3000 398.8000 134.4000 ;
	    RECT 401.2000 134.3000 402.0000 134.4000 ;
	    RECT 398.0000 133.7000 402.0000 134.3000 ;
	    RECT 398.0000 133.6000 398.8000 133.7000 ;
	    RECT 401.2000 133.6000 402.0000 133.7000 ;
	    RECT 404.4000 134.3000 405.2000 134.4000 ;
	    RECT 442.8000 134.3000 443.6000 134.4000 ;
	    RECT 404.4000 133.7000 443.6000 134.3000 ;
	    RECT 404.4000 133.6000 405.2000 133.7000 ;
	    RECT 442.8000 133.6000 443.6000 133.7000 ;
	    RECT 486.0000 134.3000 486.8000 134.4000 ;
	    RECT 498.8000 134.3000 499.6000 134.4000 ;
	    RECT 486.0000 133.7000 499.6000 134.3000 ;
	    RECT 486.0000 133.6000 486.8000 133.7000 ;
	    RECT 498.8000 133.6000 499.6000 133.7000 ;
	    RECT 502.0000 134.3000 502.8000 134.4000 ;
	    RECT 503.6000 134.3000 504.4000 134.4000 ;
	    RECT 502.0000 133.7000 504.4000 134.3000 ;
	    RECT 502.0000 133.6000 502.8000 133.7000 ;
	    RECT 503.6000 133.6000 504.4000 133.7000 ;
	    RECT 41.2000 132.3000 42.0000 132.4000 ;
	    RECT 90.8000 132.3000 91.6000 132.4000 ;
	    RECT 41.2000 131.7000 91.6000 132.3000 ;
	    RECT 41.2000 131.6000 42.0000 131.7000 ;
	    RECT 90.8000 131.6000 91.6000 131.7000 ;
	    RECT 94.0000 132.3000 94.8000 132.4000 ;
	    RECT 100.4000 132.3000 101.2000 132.4000 ;
	    RECT 94.0000 131.7000 101.2000 132.3000 ;
	    RECT 94.0000 131.6000 94.8000 131.7000 ;
	    RECT 100.4000 131.6000 101.2000 131.7000 ;
	    RECT 110.0000 132.3000 110.8000 132.4000 ;
	    RECT 130.8000 132.3000 131.6000 132.4000 ;
	    RECT 110.0000 131.7000 131.6000 132.3000 ;
	    RECT 110.0000 131.6000 110.8000 131.7000 ;
	    RECT 130.8000 131.6000 131.6000 131.7000 ;
	    RECT 138.8000 132.3000 139.6000 132.4000 ;
	    RECT 154.8000 132.3000 155.6000 132.4000 ;
	    RECT 138.8000 131.7000 155.6000 132.3000 ;
	    RECT 138.8000 131.6000 139.6000 131.7000 ;
	    RECT 154.8000 131.6000 155.6000 131.7000 ;
	    RECT 161.2000 132.3000 162.0000 132.4000 ;
	    RECT 164.4000 132.3000 165.2000 132.4000 ;
	    RECT 170.8000 132.3000 171.6000 132.4000 ;
	    RECT 174.0000 132.3000 174.8000 132.4000 ;
	    RECT 177.2000 132.3000 178.0000 132.4000 ;
	    RECT 161.2000 131.7000 178.0000 132.3000 ;
	    RECT 161.2000 131.6000 162.0000 131.7000 ;
	    RECT 164.4000 131.6000 165.2000 131.7000 ;
	    RECT 170.8000 131.6000 171.6000 131.7000 ;
	    RECT 174.0000 131.6000 174.8000 131.7000 ;
	    RECT 177.2000 131.6000 178.0000 131.7000 ;
	    RECT 178.8000 132.3000 179.6000 132.4000 ;
	    RECT 196.4000 132.3000 197.2000 132.4000 ;
	    RECT 178.8000 131.7000 197.2000 132.3000 ;
	    RECT 178.8000 131.6000 179.6000 131.7000 ;
	    RECT 196.4000 131.6000 197.2000 131.7000 ;
	    RECT 215.6000 131.6000 216.4000 132.4000 ;
	    RECT 218.8000 132.3000 219.6000 132.4000 ;
	    RECT 265.2000 132.3000 266.0000 132.4000 ;
	    RECT 218.8000 131.7000 266.0000 132.3000 ;
	    RECT 218.8000 131.6000 219.6000 131.7000 ;
	    RECT 265.2000 131.6000 266.0000 131.7000 ;
	    RECT 266.8000 131.6000 267.6000 132.4000 ;
	    RECT 268.4000 132.3000 269.2000 132.4000 ;
	    RECT 297.2000 132.3000 298.0000 132.4000 ;
	    RECT 268.4000 131.7000 298.0000 132.3000 ;
	    RECT 268.4000 131.6000 269.2000 131.7000 ;
	    RECT 297.2000 131.6000 298.0000 131.7000 ;
	    RECT 298.8000 132.3000 299.6000 132.4000 ;
	    RECT 324.4000 132.3000 325.2000 132.4000 ;
	    RECT 298.8000 131.7000 325.2000 132.3000 ;
	    RECT 298.8000 131.6000 299.6000 131.7000 ;
	    RECT 324.4000 131.6000 325.2000 131.7000 ;
	    RECT 330.8000 132.3000 331.6000 132.4000 ;
	    RECT 332.4000 132.3000 333.2000 132.4000 ;
	    RECT 330.8000 131.7000 333.2000 132.3000 ;
	    RECT 330.8000 131.6000 331.6000 131.7000 ;
	    RECT 332.4000 131.6000 333.2000 131.7000 ;
	    RECT 335.6000 132.3000 336.4000 132.4000 ;
	    RECT 364.4000 132.3000 365.2000 132.4000 ;
	    RECT 374.0000 132.3000 374.8000 132.4000 ;
	    RECT 335.6000 131.7000 363.5000 132.3000 ;
	    RECT 335.6000 131.6000 336.4000 131.7000 ;
	    RECT 9.2000 130.3000 10.0000 130.4000 ;
	    RECT 41.2000 130.3000 42.0000 130.4000 ;
	    RECT 62.0000 130.3000 62.8000 130.4000 ;
	    RECT 9.2000 129.7000 42.0000 130.3000 ;
	    RECT 9.2000 129.6000 10.0000 129.7000 ;
	    RECT 41.2000 129.6000 42.0000 129.7000 ;
	    RECT 54.1000 129.7000 62.8000 130.3000 ;
	    RECT 33.2000 128.3000 34.0000 128.4000 ;
	    RECT 54.1000 128.3000 54.7000 129.7000 ;
	    RECT 62.0000 129.6000 62.8000 129.7000 ;
	    RECT 73.2000 130.3000 74.0000 130.4000 ;
	    RECT 84.4000 130.3000 85.2000 130.4000 ;
	    RECT 102.0000 130.3000 102.8000 130.4000 ;
	    RECT 73.2000 129.7000 102.8000 130.3000 ;
	    RECT 73.2000 129.6000 74.0000 129.7000 ;
	    RECT 84.4000 129.6000 85.2000 129.7000 ;
	    RECT 102.0000 129.6000 102.8000 129.7000 ;
	    RECT 118.0000 130.3000 118.8000 130.4000 ;
	    RECT 127.6000 130.3000 128.4000 130.4000 ;
	    RECT 118.0000 129.7000 128.4000 130.3000 ;
	    RECT 118.0000 129.6000 118.8000 129.7000 ;
	    RECT 127.6000 129.6000 128.4000 129.7000 ;
	    RECT 129.2000 130.3000 130.0000 130.4000 ;
	    RECT 167.6000 130.3000 168.4000 130.4000 ;
	    RECT 129.2000 129.7000 168.4000 130.3000 ;
	    RECT 129.2000 129.6000 130.0000 129.7000 ;
	    RECT 167.6000 129.6000 168.4000 129.7000 ;
	    RECT 244.4000 129.6000 245.2000 130.4000 ;
	    RECT 282.8000 130.3000 283.6000 130.4000 ;
	    RECT 287.6000 130.3000 288.4000 130.4000 ;
	    RECT 282.8000 129.7000 288.4000 130.3000 ;
	    RECT 282.8000 129.6000 283.6000 129.7000 ;
	    RECT 287.6000 129.6000 288.4000 129.7000 ;
	    RECT 290.8000 130.3000 291.6000 130.4000 ;
	    RECT 298.8000 130.3000 299.6000 130.4000 ;
	    RECT 290.8000 129.7000 299.6000 130.3000 ;
	    RECT 290.8000 129.6000 291.6000 129.7000 ;
	    RECT 298.8000 129.6000 299.6000 129.7000 ;
	    RECT 302.0000 130.3000 302.8000 130.4000 ;
	    RECT 326.0000 130.3000 326.8000 130.4000 ;
	    RECT 332.4000 130.3000 333.2000 130.4000 ;
	    RECT 359.6000 130.3000 360.4000 130.4000 ;
	    RECT 302.0000 129.7000 321.9000 130.3000 ;
	    RECT 302.0000 129.6000 302.8000 129.7000 ;
	    RECT 33.2000 127.7000 54.7000 128.3000 ;
	    RECT 55.6000 128.3000 56.4000 128.4000 ;
	    RECT 94.0000 128.3000 94.8000 128.4000 ;
	    RECT 55.6000 127.7000 94.8000 128.3000 ;
	    RECT 33.2000 127.6000 34.0000 127.7000 ;
	    RECT 55.6000 127.6000 56.4000 127.7000 ;
	    RECT 94.0000 127.6000 94.8000 127.7000 ;
	    RECT 98.8000 128.3000 99.6000 128.4000 ;
	    RECT 121.2000 128.3000 122.0000 128.4000 ;
	    RECT 98.8000 127.7000 122.0000 128.3000 ;
	    RECT 98.8000 127.6000 99.6000 127.7000 ;
	    RECT 121.2000 127.6000 122.0000 127.7000 ;
	    RECT 127.6000 128.3000 128.4000 128.4000 ;
	    RECT 135.6000 128.3000 136.4000 128.4000 ;
	    RECT 127.6000 127.7000 136.4000 128.3000 ;
	    RECT 127.6000 127.6000 128.4000 127.7000 ;
	    RECT 135.6000 127.6000 136.4000 127.7000 ;
	    RECT 142.0000 128.3000 142.8000 128.4000 ;
	    RECT 143.6000 128.3000 144.4000 128.4000 ;
	    RECT 142.0000 127.7000 144.4000 128.3000 ;
	    RECT 142.0000 127.6000 142.8000 127.7000 ;
	    RECT 143.6000 127.6000 144.4000 127.7000 ;
	    RECT 148.4000 128.3000 149.2000 128.4000 ;
	    RECT 151.6000 128.3000 152.4000 128.4000 ;
	    RECT 148.4000 127.7000 152.4000 128.3000 ;
	    RECT 148.4000 127.6000 149.2000 127.7000 ;
	    RECT 151.6000 127.6000 152.4000 127.7000 ;
	    RECT 231.6000 128.3000 232.4000 128.4000 ;
	    RECT 238.0000 128.3000 238.8000 128.4000 ;
	    RECT 231.6000 127.7000 238.8000 128.3000 ;
	    RECT 244.5000 128.3000 245.1000 129.6000 ;
	    RECT 258.8000 128.3000 259.6000 128.4000 ;
	    RECT 244.5000 127.7000 259.6000 128.3000 ;
	    RECT 231.6000 127.6000 232.4000 127.7000 ;
	    RECT 238.0000 127.6000 238.8000 127.7000 ;
	    RECT 258.8000 127.6000 259.6000 127.7000 ;
	    RECT 260.4000 128.3000 261.2000 128.4000 ;
	    RECT 273.2000 128.3000 274.0000 128.4000 ;
	    RECT 260.4000 127.7000 274.0000 128.3000 ;
	    RECT 260.4000 127.6000 261.2000 127.7000 ;
	    RECT 273.2000 127.6000 274.0000 127.7000 ;
	    RECT 278.0000 128.3000 278.8000 128.4000 ;
	    RECT 284.4000 128.3000 285.2000 128.4000 ;
	    RECT 313.2000 128.3000 314.0000 128.4000 ;
	    RECT 278.0000 127.7000 314.0000 128.3000 ;
	    RECT 278.0000 127.6000 278.8000 127.7000 ;
	    RECT 284.4000 127.6000 285.2000 127.7000 ;
	    RECT 313.2000 127.6000 314.0000 127.7000 ;
	    RECT 316.4000 128.3000 317.2000 128.4000 ;
	    RECT 319.6000 128.3000 320.4000 128.4000 ;
	    RECT 316.4000 127.7000 320.4000 128.3000 ;
	    RECT 321.3000 128.3000 321.9000 129.7000 ;
	    RECT 326.0000 129.7000 360.4000 130.3000 ;
	    RECT 362.9000 130.3000 363.5000 131.7000 ;
	    RECT 364.4000 131.7000 374.8000 132.3000 ;
	    RECT 364.4000 131.6000 365.2000 131.7000 ;
	    RECT 374.0000 131.6000 374.8000 131.7000 ;
	    RECT 425.2000 132.3000 426.0000 132.4000 ;
	    RECT 434.8000 132.3000 435.6000 132.4000 ;
	    RECT 425.2000 131.7000 435.6000 132.3000 ;
	    RECT 425.2000 131.6000 426.0000 131.7000 ;
	    RECT 434.8000 131.6000 435.6000 131.7000 ;
	    RECT 449.2000 132.3000 450.0000 132.4000 ;
	    RECT 463.6000 132.3000 464.4000 132.4000 ;
	    RECT 449.2000 131.7000 464.4000 132.3000 ;
	    RECT 449.2000 131.6000 450.0000 131.7000 ;
	    RECT 463.6000 131.6000 464.4000 131.7000 ;
	    RECT 470.0000 132.3000 470.8000 132.4000 ;
	    RECT 489.2000 132.3000 490.0000 132.4000 ;
	    RECT 505.2000 132.3000 506.0000 132.4000 ;
	    RECT 470.0000 131.7000 506.0000 132.3000 ;
	    RECT 470.0000 131.6000 470.8000 131.7000 ;
	    RECT 489.2000 131.6000 490.0000 131.7000 ;
	    RECT 505.2000 131.6000 506.0000 131.7000 ;
	    RECT 510.0000 131.6000 510.8000 132.4000 ;
	    RECT 377.2000 130.3000 378.0000 130.4000 ;
	    RECT 391.6000 130.3000 392.4000 130.4000 ;
	    RECT 362.9000 129.7000 392.4000 130.3000 ;
	    RECT 326.0000 129.6000 326.8000 129.7000 ;
	    RECT 332.4000 129.6000 333.2000 129.7000 ;
	    RECT 359.6000 129.6000 360.4000 129.7000 ;
	    RECT 377.2000 129.6000 378.0000 129.7000 ;
	    RECT 391.6000 129.6000 392.4000 129.7000 ;
	    RECT 430.0000 130.3000 430.8000 130.4000 ;
	    RECT 431.6000 130.3000 432.4000 130.4000 ;
	    RECT 439.6000 130.3000 440.4000 130.4000 ;
	    RECT 430.0000 129.7000 440.4000 130.3000 ;
	    RECT 430.0000 129.6000 430.8000 129.7000 ;
	    RECT 431.6000 129.6000 432.4000 129.7000 ;
	    RECT 439.6000 129.6000 440.4000 129.7000 ;
	    RECT 444.4000 130.3000 445.2000 130.4000 ;
	    RECT 449.2000 130.3000 450.0000 130.4000 ;
	    RECT 457.2000 130.3000 458.0000 130.4000 ;
	    RECT 444.4000 129.7000 458.0000 130.3000 ;
	    RECT 444.4000 129.6000 445.2000 129.7000 ;
	    RECT 449.2000 129.6000 450.0000 129.7000 ;
	    RECT 457.2000 129.6000 458.0000 129.7000 ;
	    RECT 327.6000 128.3000 328.4000 128.4000 ;
	    RECT 321.3000 127.7000 328.4000 128.3000 ;
	    RECT 316.4000 127.6000 317.2000 127.7000 ;
	    RECT 319.6000 127.6000 320.4000 127.7000 ;
	    RECT 327.6000 127.6000 328.4000 127.7000 ;
	    RECT 334.0000 128.3000 334.8000 128.4000 ;
	    RECT 340.4000 128.3000 341.2000 128.4000 ;
	    RECT 356.4000 128.3000 357.2000 128.4000 ;
	    RECT 334.0000 127.7000 357.2000 128.3000 ;
	    RECT 334.0000 127.6000 334.8000 127.7000 ;
	    RECT 340.4000 127.6000 341.2000 127.7000 ;
	    RECT 356.4000 127.6000 357.2000 127.7000 ;
	    RECT 506.8000 128.3000 507.6000 128.4000 ;
	    RECT 510.0000 128.3000 510.8000 128.4000 ;
	    RECT 506.8000 127.7000 510.8000 128.3000 ;
	    RECT 506.8000 127.6000 507.6000 127.7000 ;
	    RECT 510.0000 127.6000 510.8000 127.7000 ;
	    RECT 33.2000 126.3000 34.0000 126.4000 ;
	    RECT 36.4000 126.3000 37.2000 126.4000 ;
	    RECT 33.2000 125.7000 37.2000 126.3000 ;
	    RECT 33.2000 125.6000 34.0000 125.7000 ;
	    RECT 36.4000 125.6000 37.2000 125.7000 ;
	    RECT 82.8000 126.3000 83.6000 126.4000 ;
	    RECT 198.0000 126.3000 198.8000 126.4000 ;
	    RECT 82.8000 125.7000 198.8000 126.3000 ;
	    RECT 82.8000 125.6000 83.6000 125.7000 ;
	    RECT 198.0000 125.6000 198.8000 125.7000 ;
	    RECT 199.6000 126.3000 200.4000 126.4000 ;
	    RECT 209.2000 126.3000 210.0000 126.4000 ;
	    RECT 199.6000 125.7000 210.0000 126.3000 ;
	    RECT 199.6000 125.6000 200.4000 125.7000 ;
	    RECT 209.2000 125.6000 210.0000 125.7000 ;
	    RECT 215.6000 126.3000 216.4000 126.4000 ;
	    RECT 228.4000 126.3000 229.2000 126.4000 ;
	    RECT 215.6000 125.7000 229.2000 126.3000 ;
	    RECT 215.6000 125.6000 216.4000 125.7000 ;
	    RECT 228.4000 125.6000 229.2000 125.7000 ;
	    RECT 230.0000 126.3000 230.8000 126.4000 ;
	    RECT 252.4000 126.3000 253.2000 126.4000 ;
	    RECT 281.2000 126.3000 282.0000 126.4000 ;
	    RECT 230.0000 125.7000 246.7000 126.3000 ;
	    RECT 230.0000 125.6000 230.8000 125.7000 ;
	    RECT 106.8000 124.3000 107.6000 124.4000 ;
	    RECT 119.6000 124.3000 120.4000 124.4000 ;
	    RECT 178.8000 124.3000 179.6000 124.4000 ;
	    RECT 106.8000 123.7000 179.6000 124.3000 ;
	    RECT 106.8000 123.6000 107.6000 123.7000 ;
	    RECT 119.6000 123.6000 120.4000 123.7000 ;
	    RECT 178.8000 123.6000 179.6000 123.7000 ;
	    RECT 180.4000 124.3000 181.2000 124.4000 ;
	    RECT 202.8000 124.3000 203.6000 124.4000 ;
	    RECT 180.4000 123.7000 203.6000 124.3000 ;
	    RECT 180.4000 123.6000 181.2000 123.7000 ;
	    RECT 202.8000 123.6000 203.6000 123.7000 ;
	    RECT 204.4000 124.3000 205.2000 124.4000 ;
	    RECT 241.2000 124.3000 242.0000 124.4000 ;
	    RECT 204.4000 123.7000 242.0000 124.3000 ;
	    RECT 204.4000 123.6000 205.2000 123.7000 ;
	    RECT 241.2000 123.6000 242.0000 123.7000 ;
	    RECT 242.8000 124.3000 243.6000 124.4000 ;
	    RECT 244.4000 124.3000 245.2000 124.4000 ;
	    RECT 242.8000 123.7000 245.2000 124.3000 ;
	    RECT 246.1000 124.3000 246.7000 125.7000 ;
	    RECT 252.4000 125.7000 282.0000 126.3000 ;
	    RECT 252.4000 125.6000 253.2000 125.7000 ;
	    RECT 281.2000 125.6000 282.0000 125.7000 ;
	    RECT 286.0000 126.3000 286.8000 126.4000 ;
	    RECT 318.0000 126.3000 318.8000 126.4000 ;
	    RECT 286.0000 125.7000 318.8000 126.3000 ;
	    RECT 286.0000 125.6000 286.8000 125.7000 ;
	    RECT 318.0000 125.6000 318.8000 125.7000 ;
	    RECT 322.8000 126.3000 323.6000 126.4000 ;
	    RECT 350.0000 126.3000 350.8000 126.4000 ;
	    RECT 322.8000 125.7000 350.8000 126.3000 ;
	    RECT 322.8000 125.6000 323.6000 125.7000 ;
	    RECT 350.0000 125.6000 350.8000 125.7000 ;
	    RECT 354.8000 126.3000 355.6000 126.4000 ;
	    RECT 367.6000 126.3000 368.4000 126.4000 ;
	    RECT 452.4000 126.3000 453.2000 126.4000 ;
	    RECT 354.8000 125.7000 453.2000 126.3000 ;
	    RECT 354.8000 125.6000 355.6000 125.7000 ;
	    RECT 367.6000 125.6000 368.4000 125.7000 ;
	    RECT 452.4000 125.6000 453.2000 125.7000 ;
	    RECT 319.6000 124.3000 320.4000 124.4000 ;
	    RECT 246.1000 123.7000 320.4000 124.3000 ;
	    RECT 242.8000 123.6000 243.6000 123.7000 ;
	    RECT 244.4000 123.6000 245.2000 123.7000 ;
	    RECT 319.6000 123.6000 320.4000 123.7000 ;
	    RECT 348.4000 124.3000 349.2000 124.4000 ;
	    RECT 356.4000 124.3000 357.2000 124.4000 ;
	    RECT 398.0000 124.3000 398.8000 124.4000 ;
	    RECT 348.4000 123.7000 398.8000 124.3000 ;
	    RECT 348.4000 123.6000 349.2000 123.7000 ;
	    RECT 356.4000 123.6000 357.2000 123.7000 ;
	    RECT 398.0000 123.6000 398.8000 123.7000 ;
	    RECT 487.6000 124.3000 488.4000 124.4000 ;
	    RECT 510.0000 124.3000 510.8000 124.4000 ;
	    RECT 487.6000 123.7000 510.8000 124.3000 ;
	    RECT 487.6000 123.6000 488.4000 123.7000 ;
	    RECT 510.0000 123.6000 510.8000 123.7000 ;
	    RECT 134.0000 122.3000 134.8000 122.4000 ;
	    RECT 140.4000 122.3000 141.2000 122.4000 ;
	    RECT 134.0000 121.7000 141.2000 122.3000 ;
	    RECT 134.0000 121.6000 134.8000 121.7000 ;
	    RECT 140.4000 121.6000 141.2000 121.7000 ;
	    RECT 146.8000 122.3000 147.6000 122.4000 ;
	    RECT 222.0000 122.3000 222.8000 122.4000 ;
	    RECT 238.0000 122.3000 238.8000 122.4000 ;
	    RECT 282.8000 122.3000 283.6000 122.4000 ;
	    RECT 146.8000 121.7000 283.6000 122.3000 ;
	    RECT 146.8000 121.6000 147.6000 121.7000 ;
	    RECT 222.0000 121.6000 222.8000 121.7000 ;
	    RECT 238.0000 121.6000 238.8000 121.7000 ;
	    RECT 282.8000 121.6000 283.6000 121.7000 ;
	    RECT 286.0000 122.3000 286.8000 122.4000 ;
	    RECT 346.8000 122.3000 347.6000 122.4000 ;
	    RECT 286.0000 121.7000 347.6000 122.3000 ;
	    RECT 286.0000 121.6000 286.8000 121.7000 ;
	    RECT 346.8000 121.6000 347.6000 121.7000 ;
	    RECT 350.0000 122.3000 350.8000 122.4000 ;
	    RECT 366.0000 122.3000 366.8000 122.4000 ;
	    RECT 350.0000 121.7000 366.8000 122.3000 ;
	    RECT 350.0000 121.6000 350.8000 121.7000 ;
	    RECT 366.0000 121.6000 366.8000 121.7000 ;
	    RECT 111.6000 120.3000 112.4000 120.4000 ;
	    RECT 158.0000 120.3000 158.8000 120.4000 ;
	    RECT 111.6000 119.7000 158.8000 120.3000 ;
	    RECT 111.6000 119.6000 112.4000 119.7000 ;
	    RECT 158.0000 119.6000 158.8000 119.7000 ;
	    RECT 177.2000 120.3000 178.0000 120.4000 ;
	    RECT 210.8000 120.3000 211.6000 120.4000 ;
	    RECT 218.8000 120.3000 219.6000 120.4000 ;
	    RECT 177.2000 119.7000 219.6000 120.3000 ;
	    RECT 177.2000 119.6000 178.0000 119.7000 ;
	    RECT 210.8000 119.6000 211.6000 119.7000 ;
	    RECT 218.8000 119.6000 219.6000 119.7000 ;
	    RECT 247.6000 120.3000 248.4000 120.4000 ;
	    RECT 295.6000 120.3000 296.4000 120.4000 ;
	    RECT 247.6000 119.7000 296.4000 120.3000 ;
	    RECT 247.6000 119.6000 248.4000 119.7000 ;
	    RECT 295.6000 119.6000 296.4000 119.7000 ;
	    RECT 298.8000 120.3000 299.6000 120.4000 ;
	    RECT 303.6000 120.3000 304.4000 120.4000 ;
	    RECT 298.8000 119.7000 304.4000 120.3000 ;
	    RECT 298.8000 119.6000 299.6000 119.7000 ;
	    RECT 303.6000 119.6000 304.4000 119.7000 ;
	    RECT 313.2000 120.3000 314.0000 120.4000 ;
	    RECT 318.0000 120.3000 318.8000 120.4000 ;
	    RECT 313.2000 119.7000 318.8000 120.3000 ;
	    RECT 313.2000 119.6000 314.0000 119.7000 ;
	    RECT 318.0000 119.6000 318.8000 119.7000 ;
	    RECT 321.2000 120.3000 322.0000 120.4000 ;
	    RECT 380.4000 120.3000 381.2000 120.4000 ;
	    RECT 321.2000 119.7000 381.2000 120.3000 ;
	    RECT 321.2000 119.6000 322.0000 119.7000 ;
	    RECT 380.4000 119.6000 381.2000 119.7000 ;
	    RECT 92.4000 118.3000 93.2000 118.4000 ;
	    RECT 113.2000 118.3000 114.0000 118.4000 ;
	    RECT 148.4000 118.3000 149.2000 118.4000 ;
	    RECT 244.4000 118.3000 245.2000 118.4000 ;
	    RECT 92.4000 117.7000 245.2000 118.3000 ;
	    RECT 92.4000 117.6000 93.2000 117.7000 ;
	    RECT 113.2000 117.6000 114.0000 117.7000 ;
	    RECT 148.4000 117.6000 149.2000 117.7000 ;
	    RECT 244.4000 117.6000 245.2000 117.7000 ;
	    RECT 246.0000 118.3000 246.8000 118.4000 ;
	    RECT 282.8000 118.3000 283.6000 118.4000 ;
	    RECT 314.8000 118.3000 315.6000 118.4000 ;
	    RECT 246.0000 117.7000 315.6000 118.3000 ;
	    RECT 246.0000 117.6000 246.8000 117.7000 ;
	    RECT 282.8000 117.6000 283.6000 117.7000 ;
	    RECT 314.8000 117.6000 315.6000 117.7000 ;
	    RECT 316.4000 118.3000 317.2000 118.4000 ;
	    RECT 378.8000 118.3000 379.6000 118.4000 ;
	    RECT 386.8000 118.3000 387.6000 118.4000 ;
	    RECT 316.4000 117.7000 387.6000 118.3000 ;
	    RECT 316.4000 117.6000 317.2000 117.7000 ;
	    RECT 378.8000 117.6000 379.6000 117.7000 ;
	    RECT 386.8000 117.6000 387.6000 117.7000 ;
	    RECT 398.0000 118.3000 398.8000 118.4000 ;
	    RECT 404.4000 118.3000 405.2000 118.4000 ;
	    RECT 398.0000 117.7000 405.2000 118.3000 ;
	    RECT 398.0000 117.6000 398.8000 117.7000 ;
	    RECT 404.4000 117.6000 405.2000 117.7000 ;
	    RECT 442.8000 118.3000 443.6000 118.4000 ;
	    RECT 465.2000 118.3000 466.0000 118.4000 ;
	    RECT 442.8000 117.7000 466.0000 118.3000 ;
	    RECT 442.8000 117.6000 443.6000 117.7000 ;
	    RECT 465.2000 117.6000 466.0000 117.7000 ;
	    RECT 498.8000 118.3000 499.6000 118.4000 ;
	    RECT 508.4000 118.3000 509.2000 118.4000 ;
	    RECT 498.8000 117.7000 509.2000 118.3000 ;
	    RECT 498.8000 117.6000 499.6000 117.7000 ;
	    RECT 508.4000 117.6000 509.2000 117.7000 ;
	    RECT 22.0000 116.3000 22.8000 116.4000 ;
	    RECT 81.2000 116.3000 82.0000 116.4000 ;
	    RECT 22.0000 115.7000 82.0000 116.3000 ;
	    RECT 22.0000 115.6000 22.8000 115.7000 ;
	    RECT 81.2000 115.6000 82.0000 115.7000 ;
	    RECT 87.6000 116.3000 88.4000 116.4000 ;
	    RECT 111.6000 116.3000 112.4000 116.4000 ;
	    RECT 87.6000 115.7000 112.4000 116.3000 ;
	    RECT 87.6000 115.6000 88.4000 115.7000 ;
	    RECT 111.6000 115.6000 112.4000 115.7000 ;
	    RECT 119.6000 116.3000 120.4000 116.4000 ;
	    RECT 142.0000 116.3000 142.8000 116.4000 ;
	    RECT 119.6000 115.7000 142.8000 116.3000 ;
	    RECT 119.6000 115.6000 120.4000 115.7000 ;
	    RECT 142.0000 115.6000 142.8000 115.7000 ;
	    RECT 148.4000 116.3000 149.2000 116.4000 ;
	    RECT 156.4000 116.3000 157.2000 116.4000 ;
	    RECT 148.4000 115.7000 157.2000 116.3000 ;
	    RECT 148.4000 115.6000 149.2000 115.7000 ;
	    RECT 156.4000 115.6000 157.2000 115.7000 ;
	    RECT 158.0000 116.3000 158.8000 116.4000 ;
	    RECT 300.4000 116.3000 301.2000 116.4000 ;
	    RECT 158.0000 115.7000 301.2000 116.3000 ;
	    RECT 158.0000 115.6000 158.8000 115.7000 ;
	    RECT 300.4000 115.6000 301.2000 115.7000 ;
	    RECT 361.2000 116.3000 362.0000 116.4000 ;
	    RECT 370.8000 116.3000 371.6000 116.4000 ;
	    RECT 412.4000 116.3000 413.2000 116.4000 ;
	    RECT 471.6000 116.3000 472.4000 116.4000 ;
	    RECT 361.2000 115.7000 413.2000 116.3000 ;
	    RECT 361.2000 115.6000 362.0000 115.7000 ;
	    RECT 370.8000 115.6000 371.6000 115.7000 ;
	    RECT 412.4000 115.6000 413.2000 115.7000 ;
	    RECT 414.1000 115.7000 472.4000 116.3000 ;
	    RECT 26.8000 114.3000 27.6000 114.4000 ;
	    RECT 55.6000 114.3000 56.4000 114.4000 ;
	    RECT 26.8000 113.7000 56.4000 114.3000 ;
	    RECT 26.8000 113.6000 27.6000 113.7000 ;
	    RECT 55.6000 113.6000 56.4000 113.7000 ;
	    RECT 58.8000 114.3000 59.6000 114.4000 ;
	    RECT 71.6000 114.3000 72.4000 114.4000 ;
	    RECT 58.8000 113.7000 72.4000 114.3000 ;
	    RECT 58.8000 113.6000 59.6000 113.7000 ;
	    RECT 71.6000 113.6000 72.4000 113.7000 ;
	    RECT 79.6000 114.3000 80.4000 114.4000 ;
	    RECT 98.8000 114.3000 99.6000 114.4000 ;
	    RECT 124.4000 114.3000 125.2000 114.4000 ;
	    RECT 79.6000 113.7000 125.2000 114.3000 ;
	    RECT 79.6000 113.6000 80.4000 113.7000 ;
	    RECT 98.8000 113.6000 99.6000 113.7000 ;
	    RECT 124.4000 113.6000 125.2000 113.7000 ;
	    RECT 137.2000 114.3000 138.0000 114.4000 ;
	    RECT 142.0000 114.3000 142.8000 114.4000 ;
	    RECT 154.8000 114.3000 155.6000 114.4000 ;
	    RECT 159.6000 114.3000 160.4000 114.4000 ;
	    RECT 182.0000 114.3000 182.8000 114.4000 ;
	    RECT 185.2000 114.3000 186.0000 114.4000 ;
	    RECT 137.2000 113.7000 186.0000 114.3000 ;
	    RECT 137.2000 113.6000 138.0000 113.7000 ;
	    RECT 142.0000 113.6000 142.8000 113.7000 ;
	    RECT 154.8000 113.6000 155.6000 113.7000 ;
	    RECT 159.6000 113.6000 160.4000 113.7000 ;
	    RECT 182.0000 113.6000 182.8000 113.7000 ;
	    RECT 185.2000 113.6000 186.0000 113.7000 ;
	    RECT 188.4000 114.3000 189.2000 114.4000 ;
	    RECT 193.2000 114.3000 194.0000 114.4000 ;
	    RECT 206.0000 114.3000 206.8000 114.4000 ;
	    RECT 188.4000 113.7000 206.8000 114.3000 ;
	    RECT 188.4000 113.6000 189.2000 113.7000 ;
	    RECT 193.2000 113.6000 194.0000 113.7000 ;
	    RECT 206.0000 113.6000 206.8000 113.7000 ;
	    RECT 214.0000 114.3000 214.8000 114.4000 ;
	    RECT 215.6000 114.3000 216.4000 114.4000 ;
	    RECT 276.4000 114.3000 277.2000 114.4000 ;
	    RECT 214.0000 113.7000 216.4000 114.3000 ;
	    RECT 214.0000 113.6000 214.8000 113.7000 ;
	    RECT 215.6000 113.6000 216.4000 113.7000 ;
	    RECT 226.9000 113.7000 277.2000 114.3000 ;
	    RECT 4.4000 112.3000 5.2000 112.4000 ;
	    RECT 30.0000 112.3000 30.8000 112.4000 ;
	    RECT 36.4000 112.3000 37.2000 112.4000 ;
	    RECT 4.4000 111.7000 37.2000 112.3000 ;
	    RECT 4.4000 111.6000 5.2000 111.7000 ;
	    RECT 30.0000 111.6000 30.8000 111.7000 ;
	    RECT 36.4000 111.6000 37.2000 111.7000 ;
	    RECT 71.6000 112.3000 72.4000 112.4000 ;
	    RECT 86.0000 112.3000 86.8000 112.4000 ;
	    RECT 71.6000 111.7000 86.8000 112.3000 ;
	    RECT 71.6000 111.6000 72.4000 111.7000 ;
	    RECT 86.0000 111.6000 86.8000 111.7000 ;
	    RECT 121.2000 112.3000 122.0000 112.4000 ;
	    RECT 134.0000 112.3000 134.8000 112.4000 ;
	    RECT 121.2000 111.7000 134.8000 112.3000 ;
	    RECT 121.2000 111.6000 122.0000 111.7000 ;
	    RECT 134.0000 111.6000 134.8000 111.7000 ;
	    RECT 135.6000 112.3000 136.4000 112.4000 ;
	    RECT 154.8000 112.3000 155.6000 112.4000 ;
	    RECT 135.6000 111.7000 155.6000 112.3000 ;
	    RECT 135.6000 111.6000 136.4000 111.7000 ;
	    RECT 154.8000 111.6000 155.6000 111.7000 ;
	    RECT 158.0000 112.3000 158.8000 112.4000 ;
	    RECT 161.2000 112.3000 162.0000 112.4000 ;
	    RECT 166.0000 112.3000 166.8000 112.4000 ;
	    RECT 158.0000 111.7000 166.8000 112.3000 ;
	    RECT 158.0000 111.6000 158.8000 111.7000 ;
	    RECT 161.2000 111.6000 162.0000 111.7000 ;
	    RECT 166.0000 111.6000 166.8000 111.7000 ;
	    RECT 169.2000 112.3000 170.0000 112.4000 ;
	    RECT 175.6000 112.3000 176.4000 112.4000 ;
	    RECT 183.6000 112.3000 184.4000 112.4000 ;
	    RECT 188.4000 112.3000 189.2000 112.4000 ;
	    RECT 169.2000 111.7000 181.1000 112.3000 ;
	    RECT 169.2000 111.6000 170.0000 111.7000 ;
	    RECT 175.6000 111.6000 176.4000 111.7000 ;
	    RECT 26.8000 110.3000 27.6000 110.4000 ;
	    RECT 31.6000 110.3000 32.4000 110.4000 ;
	    RECT 26.8000 109.7000 32.4000 110.3000 ;
	    RECT 26.8000 109.6000 27.6000 109.7000 ;
	    RECT 31.6000 109.6000 32.4000 109.7000 ;
	    RECT 49.2000 110.3000 50.0000 110.4000 ;
	    RECT 55.6000 110.3000 56.4000 110.4000 ;
	    RECT 49.2000 109.7000 56.4000 110.3000 ;
	    RECT 49.2000 109.6000 50.0000 109.7000 ;
	    RECT 55.6000 109.6000 56.4000 109.7000 ;
	    RECT 84.4000 110.3000 85.2000 110.4000 ;
	    RECT 89.2000 110.3000 90.0000 110.4000 ;
	    RECT 84.4000 109.7000 90.0000 110.3000 ;
	    RECT 84.4000 109.6000 85.2000 109.7000 ;
	    RECT 89.2000 109.6000 90.0000 109.7000 ;
	    RECT 95.6000 110.3000 96.4000 110.4000 ;
	    RECT 110.0000 110.3000 110.8000 110.4000 ;
	    RECT 95.6000 109.7000 110.8000 110.3000 ;
	    RECT 95.6000 109.6000 96.4000 109.7000 ;
	    RECT 110.0000 109.6000 110.8000 109.7000 ;
	    RECT 122.8000 110.3000 123.6000 110.4000 ;
	    RECT 132.4000 110.3000 133.2000 110.4000 ;
	    RECT 145.2000 110.3000 146.0000 110.4000 ;
	    RECT 122.8000 109.7000 146.0000 110.3000 ;
	    RECT 122.8000 109.6000 123.6000 109.7000 ;
	    RECT 132.4000 109.6000 133.2000 109.7000 ;
	    RECT 145.2000 109.6000 146.0000 109.7000 ;
	    RECT 151.6000 110.3000 152.4000 110.4000 ;
	    RECT 161.2000 110.3000 162.0000 110.4000 ;
	    RECT 151.6000 109.7000 162.0000 110.3000 ;
	    RECT 151.6000 109.6000 152.4000 109.7000 ;
	    RECT 161.2000 109.6000 162.0000 109.7000 ;
	    RECT 174.0000 110.3000 174.8000 110.4000 ;
	    RECT 178.8000 110.3000 179.6000 110.4000 ;
	    RECT 174.0000 109.7000 179.6000 110.3000 ;
	    RECT 180.5000 110.3000 181.1000 111.7000 ;
	    RECT 183.6000 111.7000 189.2000 112.3000 ;
	    RECT 183.6000 111.6000 184.4000 111.7000 ;
	    RECT 188.4000 111.6000 189.2000 111.7000 ;
	    RECT 201.2000 112.3000 202.0000 112.4000 ;
	    RECT 212.4000 112.3000 213.2000 112.4000 ;
	    RECT 201.2000 111.7000 213.2000 112.3000 ;
	    RECT 201.2000 111.6000 202.0000 111.7000 ;
	    RECT 212.4000 111.6000 213.2000 111.7000 ;
	    RECT 215.6000 112.3000 216.4000 112.4000 ;
	    RECT 226.9000 112.3000 227.5000 113.7000 ;
	    RECT 276.4000 113.6000 277.2000 113.7000 ;
	    RECT 294.0000 114.3000 294.8000 114.4000 ;
	    RECT 300.4000 114.3000 301.2000 114.4000 ;
	    RECT 294.0000 113.7000 301.2000 114.3000 ;
	    RECT 294.0000 113.6000 294.8000 113.7000 ;
	    RECT 300.4000 113.6000 301.2000 113.7000 ;
	    RECT 366.0000 114.3000 366.8000 114.4000 ;
	    RECT 375.6000 114.3000 376.4000 114.4000 ;
	    RECT 414.1000 114.3000 414.7000 115.7000 ;
	    RECT 471.6000 115.6000 472.4000 115.7000 ;
	    RECT 366.0000 113.7000 414.7000 114.3000 ;
	    RECT 462.0000 114.3000 462.8000 114.4000 ;
	    RECT 465.2000 114.3000 466.0000 114.4000 ;
	    RECT 462.0000 113.7000 466.0000 114.3000 ;
	    RECT 366.0000 113.6000 366.8000 113.7000 ;
	    RECT 375.6000 113.6000 376.4000 113.7000 ;
	    RECT 462.0000 113.6000 462.8000 113.7000 ;
	    RECT 465.2000 113.6000 466.0000 113.7000 ;
	    RECT 484.4000 114.3000 485.2000 114.4000 ;
	    RECT 502.0000 114.3000 502.8000 114.4000 ;
	    RECT 484.4000 113.7000 502.8000 114.3000 ;
	    RECT 484.4000 113.6000 485.2000 113.7000 ;
	    RECT 502.0000 113.6000 502.8000 113.7000 ;
	    RECT 503.6000 114.3000 504.4000 114.4000 ;
	    RECT 510.0000 114.3000 510.8000 114.4000 ;
	    RECT 503.6000 113.7000 510.8000 114.3000 ;
	    RECT 503.6000 113.6000 504.4000 113.7000 ;
	    RECT 510.0000 113.6000 510.8000 113.7000 ;
	    RECT 215.6000 111.7000 227.5000 112.3000 ;
	    RECT 233.2000 112.3000 234.0000 112.4000 ;
	    RECT 234.8000 112.3000 235.6000 112.4000 ;
	    RECT 233.2000 111.7000 235.6000 112.3000 ;
	    RECT 215.6000 111.6000 216.4000 111.7000 ;
	    RECT 233.2000 111.6000 234.0000 111.7000 ;
	    RECT 234.8000 111.6000 235.6000 111.7000 ;
	    RECT 239.6000 112.3000 240.4000 112.4000 ;
	    RECT 246.0000 112.3000 246.8000 112.4000 ;
	    RECT 239.6000 111.7000 246.8000 112.3000 ;
	    RECT 239.6000 111.6000 240.4000 111.7000 ;
	    RECT 246.0000 111.6000 246.8000 111.7000 ;
	    RECT 247.6000 112.3000 248.4000 112.4000 ;
	    RECT 263.6000 112.3000 264.4000 112.4000 ;
	    RECT 247.6000 111.7000 264.4000 112.3000 ;
	    RECT 247.6000 111.6000 248.4000 111.7000 ;
	    RECT 263.6000 111.6000 264.4000 111.7000 ;
	    RECT 265.2000 112.3000 266.0000 112.4000 ;
	    RECT 270.0000 112.3000 270.8000 112.4000 ;
	    RECT 265.2000 111.7000 270.8000 112.3000 ;
	    RECT 265.2000 111.6000 266.0000 111.7000 ;
	    RECT 270.0000 111.6000 270.8000 111.7000 ;
	    RECT 271.6000 112.3000 272.4000 112.4000 ;
	    RECT 286.0000 112.3000 286.8000 112.4000 ;
	    RECT 271.6000 111.7000 286.8000 112.3000 ;
	    RECT 271.6000 111.6000 272.4000 111.7000 ;
	    RECT 286.0000 111.6000 286.8000 111.7000 ;
	    RECT 289.2000 112.3000 290.0000 112.4000 ;
	    RECT 306.8000 112.3000 307.6000 112.4000 ;
	    RECT 319.6000 112.3000 320.4000 112.4000 ;
	    RECT 324.4000 112.3000 325.2000 112.4000 ;
	    RECT 289.2000 111.7000 325.2000 112.3000 ;
	    RECT 289.2000 111.6000 290.0000 111.7000 ;
	    RECT 306.8000 111.6000 307.6000 111.7000 ;
	    RECT 319.6000 111.6000 320.4000 111.7000 ;
	    RECT 324.4000 111.6000 325.2000 111.7000 ;
	    RECT 346.8000 112.3000 347.6000 112.4000 ;
	    RECT 354.8000 112.3000 355.6000 112.4000 ;
	    RECT 346.8000 111.7000 355.6000 112.3000 ;
	    RECT 346.8000 111.6000 347.6000 111.7000 ;
	    RECT 354.8000 111.6000 355.6000 111.7000 ;
	    RECT 359.6000 112.3000 360.4000 112.4000 ;
	    RECT 362.8000 112.3000 363.6000 112.4000 ;
	    RECT 359.6000 111.7000 363.6000 112.3000 ;
	    RECT 359.6000 111.6000 360.4000 111.7000 ;
	    RECT 362.8000 111.6000 363.6000 111.7000 ;
	    RECT 390.0000 112.3000 390.8000 112.4000 ;
	    RECT 398.0000 112.3000 398.8000 112.4000 ;
	    RECT 390.0000 111.7000 398.8000 112.3000 ;
	    RECT 390.0000 111.6000 390.8000 111.7000 ;
	    RECT 398.0000 111.6000 398.8000 111.7000 ;
	    RECT 401.2000 112.3000 402.0000 112.4000 ;
	    RECT 422.0000 112.3000 422.8000 112.4000 ;
	    RECT 401.2000 111.7000 422.8000 112.3000 ;
	    RECT 401.2000 111.6000 402.0000 111.7000 ;
	    RECT 422.0000 111.6000 422.8000 111.7000 ;
	    RECT 457.2000 112.3000 458.0000 112.4000 ;
	    RECT 462.0000 112.3000 462.8000 112.4000 ;
	    RECT 457.2000 111.7000 462.8000 112.3000 ;
	    RECT 457.2000 111.6000 458.0000 111.7000 ;
	    RECT 462.0000 111.6000 462.8000 111.7000 ;
	    RECT 471.6000 112.3000 472.4000 112.4000 ;
	    RECT 490.8000 112.3000 491.6000 112.4000 ;
	    RECT 471.6000 111.7000 491.6000 112.3000 ;
	    RECT 471.6000 111.6000 472.4000 111.7000 ;
	    RECT 490.8000 111.6000 491.6000 111.7000 ;
	    RECT 191.6000 110.3000 192.4000 110.4000 ;
	    RECT 194.8000 110.3000 195.6000 110.4000 ;
	    RECT 180.5000 109.7000 195.6000 110.3000 ;
	    RECT 174.0000 109.6000 174.8000 109.7000 ;
	    RECT 178.8000 109.6000 179.6000 109.7000 ;
	    RECT 191.6000 109.6000 192.4000 109.7000 ;
	    RECT 194.8000 109.6000 195.6000 109.7000 ;
	    RECT 196.4000 110.3000 197.2000 110.4000 ;
	    RECT 204.4000 110.3000 205.2000 110.4000 ;
	    RECT 196.4000 109.7000 205.2000 110.3000 ;
	    RECT 196.4000 109.6000 197.2000 109.7000 ;
	    RECT 204.4000 109.6000 205.2000 109.7000 ;
	    RECT 206.0000 110.3000 206.8000 110.4000 ;
	    RECT 212.4000 110.3000 213.2000 110.4000 ;
	    RECT 236.4000 110.3000 237.2000 110.4000 ;
	    RECT 206.0000 109.7000 213.2000 110.3000 ;
	    RECT 206.0000 109.6000 206.8000 109.7000 ;
	    RECT 212.4000 109.6000 213.2000 109.7000 ;
	    RECT 214.1000 109.7000 237.2000 110.3000 ;
	    RECT 25.2000 108.3000 26.0000 108.4000 ;
	    RECT 34.8000 108.3000 35.6000 108.4000 ;
	    RECT 25.2000 107.7000 35.6000 108.3000 ;
	    RECT 25.2000 107.6000 26.0000 107.7000 ;
	    RECT 34.8000 107.6000 35.6000 107.7000 ;
	    RECT 60.4000 108.3000 61.2000 108.4000 ;
	    RECT 63.6000 108.3000 64.4000 108.4000 ;
	    RECT 60.4000 107.7000 64.4000 108.3000 ;
	    RECT 60.4000 107.6000 61.2000 107.7000 ;
	    RECT 63.6000 107.6000 64.4000 107.7000 ;
	    RECT 78.0000 108.3000 78.8000 108.4000 ;
	    RECT 108.4000 108.3000 109.2000 108.4000 ;
	    RECT 116.4000 108.3000 117.2000 108.4000 ;
	    RECT 118.0000 108.3000 118.8000 108.4000 ;
	    RECT 137.2000 108.3000 138.0000 108.4000 ;
	    RECT 186.8000 108.3000 187.6000 108.4000 ;
	    RECT 190.0000 108.3000 190.8000 108.4000 ;
	    RECT 78.0000 107.7000 99.5000 108.3000 ;
	    RECT 78.0000 107.6000 78.8000 107.7000 ;
	    RECT 79.6000 106.3000 80.4000 106.4000 ;
	    RECT 97.2000 106.3000 98.0000 106.4000 ;
	    RECT 79.6000 105.7000 98.0000 106.3000 ;
	    RECT 98.9000 106.3000 99.5000 107.7000 ;
	    RECT 108.4000 107.7000 190.8000 108.3000 ;
	    RECT 108.4000 107.6000 109.2000 107.7000 ;
	    RECT 116.4000 107.6000 117.2000 107.7000 ;
	    RECT 118.0000 107.6000 118.8000 107.7000 ;
	    RECT 137.2000 107.6000 138.0000 107.7000 ;
	    RECT 186.8000 107.6000 187.6000 107.7000 ;
	    RECT 190.0000 107.6000 190.8000 107.7000 ;
	    RECT 196.4000 108.3000 197.2000 108.4000 ;
	    RECT 214.1000 108.3000 214.7000 109.7000 ;
	    RECT 236.4000 109.6000 237.2000 109.7000 ;
	    RECT 246.0000 110.3000 246.8000 110.4000 ;
	    RECT 260.4000 110.3000 261.2000 110.4000 ;
	    RECT 246.0000 109.7000 261.2000 110.3000 ;
	    RECT 246.0000 109.6000 246.8000 109.7000 ;
	    RECT 260.4000 109.6000 261.2000 109.7000 ;
	    RECT 286.0000 110.3000 286.8000 110.4000 ;
	    RECT 290.8000 110.3000 291.6000 110.4000 ;
	    RECT 286.0000 109.7000 291.6000 110.3000 ;
	    RECT 286.0000 109.6000 286.8000 109.7000 ;
	    RECT 290.8000 109.6000 291.6000 109.7000 ;
	    RECT 297.2000 110.3000 298.0000 110.4000 ;
	    RECT 311.6000 110.3000 312.4000 110.4000 ;
	    RECT 322.8000 110.3000 323.6000 110.4000 ;
	    RECT 326.0000 110.3000 326.8000 110.4000 ;
	    RECT 297.2000 109.7000 326.8000 110.3000 ;
	    RECT 297.2000 109.6000 298.0000 109.7000 ;
	    RECT 311.6000 109.6000 312.4000 109.7000 ;
	    RECT 322.8000 109.6000 323.6000 109.7000 ;
	    RECT 326.0000 109.6000 326.8000 109.7000 ;
	    RECT 343.6000 110.3000 344.4000 110.4000 ;
	    RECT 354.8000 110.3000 355.6000 110.4000 ;
	    RECT 401.2000 110.3000 402.0000 110.4000 ;
	    RECT 343.6000 109.7000 402.0000 110.3000 ;
	    RECT 343.6000 109.6000 344.4000 109.7000 ;
	    RECT 354.8000 109.6000 355.6000 109.7000 ;
	    RECT 401.2000 109.6000 402.0000 109.7000 ;
	    RECT 447.6000 110.3000 448.4000 110.4000 ;
	    RECT 457.2000 110.3000 458.0000 110.4000 ;
	    RECT 447.6000 109.7000 458.0000 110.3000 ;
	    RECT 447.6000 109.6000 448.4000 109.7000 ;
	    RECT 457.2000 109.6000 458.0000 109.7000 ;
	    RECT 484.4000 110.3000 485.2000 110.4000 ;
	    RECT 495.6000 110.3000 496.4000 110.4000 ;
	    RECT 484.4000 109.7000 496.4000 110.3000 ;
	    RECT 484.4000 109.6000 485.2000 109.7000 ;
	    RECT 495.6000 109.6000 496.4000 109.7000 ;
	    RECT 498.8000 110.3000 499.6000 110.4000 ;
	    RECT 502.0000 110.3000 502.8000 110.4000 ;
	    RECT 506.8000 110.3000 507.6000 110.4000 ;
	    RECT 508.4000 110.3000 509.2000 110.4000 ;
	    RECT 498.8000 109.7000 509.2000 110.3000 ;
	    RECT 498.8000 109.6000 499.6000 109.7000 ;
	    RECT 502.0000 109.6000 502.8000 109.7000 ;
	    RECT 506.8000 109.6000 507.6000 109.7000 ;
	    RECT 508.4000 109.6000 509.2000 109.7000 ;
	    RECT 196.4000 107.7000 214.7000 108.3000 ;
	    RECT 218.8000 108.3000 219.6000 108.4000 ;
	    RECT 223.6000 108.3000 224.4000 108.4000 ;
	    RECT 228.4000 108.3000 229.2000 108.4000 ;
	    RECT 218.8000 107.7000 229.2000 108.3000 ;
	    RECT 196.4000 107.6000 197.2000 107.7000 ;
	    RECT 218.8000 107.6000 219.6000 107.7000 ;
	    RECT 223.6000 107.6000 224.4000 107.7000 ;
	    RECT 228.4000 107.6000 229.2000 107.7000 ;
	    RECT 241.2000 108.3000 242.0000 108.4000 ;
	    RECT 265.2000 108.3000 266.0000 108.4000 ;
	    RECT 241.2000 107.7000 266.0000 108.3000 ;
	    RECT 241.2000 107.6000 242.0000 107.7000 ;
	    RECT 265.2000 107.6000 266.0000 107.7000 ;
	    RECT 281.2000 108.3000 282.0000 108.4000 ;
	    RECT 295.6000 108.3000 296.4000 108.4000 ;
	    RECT 281.2000 107.7000 296.4000 108.3000 ;
	    RECT 281.2000 107.6000 282.0000 107.7000 ;
	    RECT 295.6000 107.6000 296.4000 107.7000 ;
	    RECT 298.8000 108.3000 299.6000 108.4000 ;
	    RECT 340.4000 108.3000 341.2000 108.4000 ;
	    RECT 298.8000 107.7000 341.2000 108.3000 ;
	    RECT 298.8000 107.6000 299.6000 107.7000 ;
	    RECT 340.4000 107.6000 341.2000 107.7000 ;
	    RECT 346.8000 107.6000 347.6000 108.4000 ;
	    RECT 375.6000 108.3000 376.4000 108.4000 ;
	    RECT 382.0000 108.3000 382.8000 108.4000 ;
	    RECT 375.6000 107.7000 382.8000 108.3000 ;
	    RECT 375.6000 107.6000 376.4000 107.7000 ;
	    RECT 382.0000 107.6000 382.8000 107.7000 ;
	    RECT 390.0000 108.3000 390.8000 108.4000 ;
	    RECT 398.0000 108.3000 398.8000 108.4000 ;
	    RECT 390.0000 107.7000 398.8000 108.3000 ;
	    RECT 390.0000 107.6000 390.8000 107.7000 ;
	    RECT 398.0000 107.6000 398.8000 107.7000 ;
	    RECT 110.0000 106.3000 110.8000 106.4000 ;
	    RECT 98.9000 105.7000 110.8000 106.3000 ;
	    RECT 79.6000 105.6000 80.4000 105.7000 ;
	    RECT 97.2000 105.6000 98.0000 105.7000 ;
	    RECT 110.0000 105.6000 110.8000 105.7000 ;
	    RECT 111.6000 106.3000 112.4000 106.4000 ;
	    RECT 129.2000 106.3000 130.0000 106.4000 ;
	    RECT 111.6000 105.7000 130.0000 106.3000 ;
	    RECT 111.6000 105.6000 112.4000 105.7000 ;
	    RECT 129.2000 105.6000 130.0000 105.7000 ;
	    RECT 134.0000 106.3000 134.8000 106.4000 ;
	    RECT 151.6000 106.3000 152.4000 106.4000 ;
	    RECT 134.0000 105.7000 152.4000 106.3000 ;
	    RECT 134.0000 105.6000 134.8000 105.7000 ;
	    RECT 151.6000 105.6000 152.4000 105.7000 ;
	    RECT 154.8000 106.3000 155.6000 106.4000 ;
	    RECT 166.0000 106.3000 166.8000 106.4000 ;
	    RECT 154.8000 105.7000 166.8000 106.3000 ;
	    RECT 154.8000 105.6000 155.6000 105.7000 ;
	    RECT 166.0000 105.6000 166.8000 105.7000 ;
	    RECT 172.4000 106.3000 173.2000 106.4000 ;
	    RECT 177.2000 106.3000 178.0000 106.4000 ;
	    RECT 172.4000 105.7000 178.0000 106.3000 ;
	    RECT 172.4000 105.6000 173.2000 105.7000 ;
	    RECT 177.2000 105.6000 178.0000 105.7000 ;
	    RECT 183.6000 106.3000 184.4000 106.4000 ;
	    RECT 226.8000 106.3000 227.6000 106.4000 ;
	    RECT 236.4000 106.3000 237.2000 106.4000 ;
	    RECT 183.6000 105.7000 237.2000 106.3000 ;
	    RECT 183.6000 105.6000 184.4000 105.7000 ;
	    RECT 226.8000 105.6000 227.6000 105.7000 ;
	    RECT 236.4000 105.6000 237.2000 105.7000 ;
	    RECT 247.6000 106.3000 248.4000 106.4000 ;
	    RECT 263.6000 106.3000 264.4000 106.4000 ;
	    RECT 247.6000 105.7000 264.4000 106.3000 ;
	    RECT 247.6000 105.6000 248.4000 105.7000 ;
	    RECT 263.6000 105.6000 264.4000 105.7000 ;
	    RECT 273.2000 106.3000 274.0000 106.4000 ;
	    RECT 286.0000 106.3000 286.8000 106.4000 ;
	    RECT 273.2000 105.7000 286.8000 106.3000 ;
	    RECT 273.2000 105.6000 274.0000 105.7000 ;
	    RECT 286.0000 105.6000 286.8000 105.7000 ;
	    RECT 295.6000 106.3000 296.4000 106.4000 ;
	    RECT 306.8000 106.3000 307.6000 106.4000 ;
	    RECT 295.6000 105.7000 307.6000 106.3000 ;
	    RECT 295.6000 105.6000 296.4000 105.7000 ;
	    RECT 306.8000 105.6000 307.6000 105.7000 ;
	    RECT 308.4000 106.3000 309.2000 106.4000 ;
	    RECT 313.2000 106.3000 314.0000 106.4000 ;
	    RECT 308.4000 105.7000 314.0000 106.3000 ;
	    RECT 308.4000 105.6000 309.2000 105.7000 ;
	    RECT 313.2000 105.6000 314.0000 105.7000 ;
	    RECT 337.2000 106.3000 338.0000 106.4000 ;
	    RECT 372.4000 106.3000 373.2000 106.4000 ;
	    RECT 337.2000 105.7000 373.2000 106.3000 ;
	    RECT 337.2000 105.6000 338.0000 105.7000 ;
	    RECT 372.4000 105.6000 373.2000 105.7000 ;
	    RECT 380.4000 106.3000 381.2000 106.4000 ;
	    RECT 386.8000 106.3000 387.6000 106.4000 ;
	    RECT 380.4000 105.7000 387.6000 106.3000 ;
	    RECT 380.4000 105.6000 381.2000 105.7000 ;
	    RECT 386.8000 105.6000 387.6000 105.7000 ;
	    RECT 455.6000 106.3000 456.4000 106.4000 ;
	    RECT 460.4000 106.3000 461.2000 106.4000 ;
	    RECT 455.6000 105.7000 461.2000 106.3000 ;
	    RECT 455.6000 105.6000 456.4000 105.7000 ;
	    RECT 460.4000 105.6000 461.2000 105.7000 ;
	    RECT 52.4000 104.3000 53.2000 104.4000 ;
	    RECT 135.6000 104.3000 136.4000 104.4000 ;
	    RECT 52.4000 103.7000 136.4000 104.3000 ;
	    RECT 52.4000 103.6000 53.2000 103.7000 ;
	    RECT 135.6000 103.6000 136.4000 103.7000 ;
	    RECT 142.0000 104.3000 142.8000 104.4000 ;
	    RECT 170.8000 104.3000 171.6000 104.4000 ;
	    RECT 142.0000 103.7000 171.6000 104.3000 ;
	    RECT 142.0000 103.6000 142.8000 103.7000 ;
	    RECT 170.8000 103.6000 171.6000 103.7000 ;
	    RECT 172.4000 104.3000 173.2000 104.4000 ;
	    RECT 185.2000 104.3000 186.0000 104.4000 ;
	    RECT 172.4000 103.7000 186.0000 104.3000 ;
	    RECT 172.4000 103.6000 173.2000 103.7000 ;
	    RECT 185.2000 103.6000 186.0000 103.7000 ;
	    RECT 206.0000 104.3000 206.8000 104.4000 ;
	    RECT 209.2000 104.3000 210.0000 104.4000 ;
	    RECT 212.4000 104.3000 213.2000 104.4000 ;
	    RECT 206.0000 103.7000 208.3000 104.3000 ;
	    RECT 206.0000 103.6000 206.8000 103.7000 ;
	    RECT 55.6000 102.3000 56.4000 102.4000 ;
	    RECT 60.4000 102.3000 61.2000 102.4000 ;
	    RECT 70.0000 102.3000 70.8000 102.4000 ;
	    RECT 74.8000 102.3000 75.6000 102.4000 ;
	    RECT 55.6000 101.7000 75.6000 102.3000 ;
	    RECT 55.6000 101.6000 56.4000 101.7000 ;
	    RECT 60.4000 101.6000 61.2000 101.7000 ;
	    RECT 70.0000 101.6000 70.8000 101.7000 ;
	    RECT 74.8000 101.6000 75.6000 101.7000 ;
	    RECT 94.0000 102.3000 94.8000 102.4000 ;
	    RECT 98.8000 102.3000 99.6000 102.4000 ;
	    RECT 94.0000 101.7000 99.6000 102.3000 ;
	    RECT 94.0000 101.6000 94.8000 101.7000 ;
	    RECT 98.8000 101.6000 99.6000 101.7000 ;
	    RECT 100.4000 102.3000 101.2000 102.4000 ;
	    RECT 119.6000 102.3000 120.4000 102.4000 ;
	    RECT 122.8000 102.3000 123.6000 102.4000 ;
	    RECT 130.8000 102.3000 131.6000 102.4000 ;
	    RECT 148.4000 102.3000 149.2000 102.4000 ;
	    RECT 196.4000 102.3000 197.2000 102.4000 ;
	    RECT 206.0000 102.3000 206.8000 102.4000 ;
	    RECT 100.4000 101.7000 206.8000 102.3000 ;
	    RECT 207.7000 102.3000 208.3000 103.7000 ;
	    RECT 209.2000 103.7000 213.2000 104.3000 ;
	    RECT 209.2000 103.6000 210.0000 103.7000 ;
	    RECT 212.4000 103.6000 213.2000 103.7000 ;
	    RECT 214.0000 104.3000 214.8000 104.4000 ;
	    RECT 265.2000 104.3000 266.0000 104.4000 ;
	    RECT 298.8000 104.3000 299.6000 104.4000 ;
	    RECT 214.0000 103.7000 262.7000 104.3000 ;
	    RECT 214.0000 103.6000 214.8000 103.7000 ;
	    RECT 215.6000 102.3000 216.4000 102.4000 ;
	    RECT 207.7000 101.7000 216.4000 102.3000 ;
	    RECT 100.4000 101.6000 101.2000 101.7000 ;
	    RECT 119.6000 101.6000 120.4000 101.7000 ;
	    RECT 122.8000 101.6000 123.6000 101.7000 ;
	    RECT 130.8000 101.6000 131.6000 101.7000 ;
	    RECT 148.4000 101.6000 149.2000 101.7000 ;
	    RECT 196.4000 101.6000 197.2000 101.7000 ;
	    RECT 206.0000 101.6000 206.8000 101.7000 ;
	    RECT 215.6000 101.6000 216.4000 101.7000 ;
	    RECT 228.4000 102.3000 229.2000 102.4000 ;
	    RECT 247.6000 102.3000 248.4000 102.4000 ;
	    RECT 228.4000 101.7000 248.4000 102.3000 ;
	    RECT 262.1000 102.3000 262.7000 103.7000 ;
	    RECT 265.2000 103.7000 299.6000 104.3000 ;
	    RECT 265.2000 103.6000 266.0000 103.7000 ;
	    RECT 298.8000 103.6000 299.6000 103.7000 ;
	    RECT 305.2000 104.3000 306.0000 104.4000 ;
	    RECT 310.0000 104.3000 310.8000 104.4000 ;
	    RECT 305.2000 103.7000 310.8000 104.3000 ;
	    RECT 305.2000 103.6000 306.0000 103.7000 ;
	    RECT 310.0000 103.6000 310.8000 103.7000 ;
	    RECT 311.6000 104.3000 312.4000 104.4000 ;
	    RECT 318.0000 104.3000 318.8000 104.4000 ;
	    RECT 434.8000 104.3000 435.6000 104.4000 ;
	    RECT 454.0000 104.3000 454.8000 104.4000 ;
	    RECT 311.6000 103.7000 454.8000 104.3000 ;
	    RECT 311.6000 103.6000 312.4000 103.7000 ;
	    RECT 318.0000 103.6000 318.8000 103.7000 ;
	    RECT 434.8000 103.6000 435.6000 103.7000 ;
	    RECT 454.0000 103.6000 454.8000 103.7000 ;
	    RECT 460.4000 104.3000 461.2000 104.4000 ;
	    RECT 468.4000 104.3000 469.2000 104.4000 ;
	    RECT 460.4000 103.7000 469.2000 104.3000 ;
	    RECT 460.4000 103.6000 461.2000 103.7000 ;
	    RECT 468.4000 103.6000 469.2000 103.7000 ;
	    RECT 262.1000 101.7000 414.7000 102.3000 ;
	    RECT 228.4000 101.6000 229.2000 101.7000 ;
	    RECT 247.6000 101.6000 248.4000 101.7000 ;
	    RECT 414.1000 100.4000 414.7000 101.7000 ;
	    RECT 68.4000 100.3000 69.2000 100.4000 ;
	    RECT 244.4000 100.3000 245.2000 100.4000 ;
	    RECT 68.4000 99.7000 245.2000 100.3000 ;
	    RECT 68.4000 99.6000 69.2000 99.7000 ;
	    RECT 244.4000 99.6000 245.2000 99.7000 ;
	    RECT 262.0000 100.3000 262.8000 100.4000 ;
	    RECT 282.8000 100.3000 283.6000 100.4000 ;
	    RECT 262.0000 99.7000 283.6000 100.3000 ;
	    RECT 262.0000 99.6000 262.8000 99.7000 ;
	    RECT 282.8000 99.6000 283.6000 99.7000 ;
	    RECT 286.0000 100.3000 286.8000 100.4000 ;
	    RECT 295.6000 100.3000 296.4000 100.4000 ;
	    RECT 286.0000 99.7000 296.4000 100.3000 ;
	    RECT 286.0000 99.6000 286.8000 99.7000 ;
	    RECT 295.6000 99.6000 296.4000 99.7000 ;
	    RECT 302.0000 100.3000 302.8000 100.4000 ;
	    RECT 345.2000 100.3000 346.0000 100.4000 ;
	    RECT 302.0000 99.7000 346.0000 100.3000 ;
	    RECT 302.0000 99.6000 302.8000 99.7000 ;
	    RECT 345.2000 99.6000 346.0000 99.7000 ;
	    RECT 353.2000 100.3000 354.0000 100.4000 ;
	    RECT 374.0000 100.3000 374.8000 100.4000 ;
	    RECT 394.8000 100.3000 395.6000 100.4000 ;
	    RECT 353.2000 99.7000 395.6000 100.3000 ;
	    RECT 353.2000 99.6000 354.0000 99.7000 ;
	    RECT 374.0000 99.6000 374.8000 99.7000 ;
	    RECT 394.8000 99.6000 395.6000 99.7000 ;
	    RECT 414.0000 100.3000 414.8000 100.4000 ;
	    RECT 430.0000 100.3000 430.8000 100.4000 ;
	    RECT 414.0000 99.7000 430.8000 100.3000 ;
	    RECT 414.0000 99.6000 414.8000 99.7000 ;
	    RECT 430.0000 99.6000 430.8000 99.7000 ;
	    RECT 462.0000 100.3000 462.8000 100.4000 ;
	    RECT 463.6000 100.3000 464.4000 100.4000 ;
	    RECT 462.0000 99.7000 464.4000 100.3000 ;
	    RECT 462.0000 99.6000 462.8000 99.7000 ;
	    RECT 463.6000 99.6000 464.4000 99.7000 ;
	    RECT 68.4000 98.3000 69.2000 98.4000 ;
	    RECT 87.6000 98.3000 88.4000 98.4000 ;
	    RECT 68.4000 97.7000 88.4000 98.3000 ;
	    RECT 68.4000 97.6000 69.2000 97.7000 ;
	    RECT 87.6000 97.6000 88.4000 97.7000 ;
	    RECT 97.2000 98.3000 98.0000 98.4000 ;
	    RECT 119.6000 98.3000 120.4000 98.4000 ;
	    RECT 97.2000 97.7000 120.4000 98.3000 ;
	    RECT 97.2000 97.6000 98.0000 97.7000 ;
	    RECT 119.6000 97.6000 120.4000 97.7000 ;
	    RECT 129.2000 98.3000 130.0000 98.4000 ;
	    RECT 135.6000 98.3000 136.4000 98.4000 ;
	    RECT 129.2000 97.7000 136.4000 98.3000 ;
	    RECT 129.2000 97.6000 130.0000 97.7000 ;
	    RECT 135.6000 97.6000 136.4000 97.7000 ;
	    RECT 138.8000 98.3000 139.6000 98.4000 ;
	    RECT 150.0000 98.3000 150.8000 98.4000 ;
	    RECT 158.0000 98.3000 158.8000 98.4000 ;
	    RECT 162.8000 98.3000 163.6000 98.4000 ;
	    RECT 138.8000 97.7000 163.6000 98.3000 ;
	    RECT 138.8000 97.6000 139.6000 97.7000 ;
	    RECT 150.0000 97.6000 150.8000 97.7000 ;
	    RECT 158.0000 97.6000 158.8000 97.7000 ;
	    RECT 162.8000 97.6000 163.6000 97.7000 ;
	    RECT 166.0000 98.3000 166.8000 98.4000 ;
	    RECT 172.4000 98.3000 173.2000 98.4000 ;
	    RECT 166.0000 97.7000 173.2000 98.3000 ;
	    RECT 166.0000 97.6000 166.8000 97.7000 ;
	    RECT 172.4000 97.6000 173.2000 97.7000 ;
	    RECT 174.0000 98.3000 174.8000 98.4000 ;
	    RECT 210.8000 98.3000 211.6000 98.4000 ;
	    RECT 225.2000 98.3000 226.0000 98.4000 ;
	    RECT 239.6000 98.3000 240.4000 98.4000 ;
	    RECT 174.0000 97.7000 198.7000 98.3000 ;
	    RECT 174.0000 97.6000 174.8000 97.7000 ;
	    RECT 198.1000 96.4000 198.7000 97.7000 ;
	    RECT 210.8000 97.7000 226.0000 98.3000 ;
	    RECT 210.8000 97.6000 211.6000 97.7000 ;
	    RECT 225.2000 97.6000 226.0000 97.7000 ;
	    RECT 226.9000 97.7000 240.4000 98.3000 ;
	    RECT 58.8000 96.3000 59.6000 96.4000 ;
	    RECT 132.4000 96.3000 133.2000 96.4000 ;
	    RECT 166.0000 96.3000 166.8000 96.4000 ;
	    RECT 58.8000 95.7000 121.9000 96.3000 ;
	    RECT 58.8000 95.6000 59.6000 95.7000 ;
	    RECT 15.6000 94.3000 16.4000 94.4000 ;
	    RECT 23.6000 94.3000 24.4000 94.4000 ;
	    RECT 15.6000 93.7000 24.4000 94.3000 ;
	    RECT 15.6000 93.6000 16.4000 93.7000 ;
	    RECT 23.6000 93.6000 24.4000 93.7000 ;
	    RECT 42.8000 94.3000 43.6000 94.4000 ;
	    RECT 49.2000 94.3000 50.0000 94.4000 ;
	    RECT 42.8000 93.7000 50.0000 94.3000 ;
	    RECT 42.8000 93.6000 43.6000 93.7000 ;
	    RECT 49.2000 93.6000 50.0000 93.7000 ;
	    RECT 52.4000 94.3000 53.2000 94.4000 ;
	    RECT 73.2000 94.3000 74.0000 94.4000 ;
	    RECT 52.4000 93.7000 74.0000 94.3000 ;
	    RECT 52.4000 93.6000 53.2000 93.7000 ;
	    RECT 73.2000 93.6000 74.0000 93.7000 ;
	    RECT 89.2000 94.3000 90.0000 94.4000 ;
	    RECT 103.6000 94.3000 104.4000 94.4000 ;
	    RECT 89.2000 93.7000 104.4000 94.3000 ;
	    RECT 89.2000 93.6000 90.0000 93.7000 ;
	    RECT 103.6000 93.6000 104.4000 93.7000 ;
	    RECT 118.0000 94.3000 118.8000 94.4000 ;
	    RECT 119.6000 94.3000 120.4000 94.4000 ;
	    RECT 118.0000 93.7000 120.4000 94.3000 ;
	    RECT 121.3000 94.3000 121.9000 95.7000 ;
	    RECT 132.4000 95.7000 166.8000 96.3000 ;
	    RECT 132.4000 95.6000 133.2000 95.7000 ;
	    RECT 166.0000 95.6000 166.8000 95.7000 ;
	    RECT 167.6000 96.3000 168.4000 96.4000 ;
	    RECT 175.6000 96.3000 176.4000 96.4000 ;
	    RECT 194.8000 96.3000 195.6000 96.4000 ;
	    RECT 167.6000 95.7000 176.4000 96.3000 ;
	    RECT 167.6000 95.6000 168.4000 95.7000 ;
	    RECT 175.6000 95.6000 176.4000 95.7000 ;
	    RECT 182.1000 95.7000 195.6000 96.3000 ;
	    RECT 182.1000 94.4000 182.7000 95.7000 ;
	    RECT 194.8000 95.6000 195.6000 95.7000 ;
	    RECT 198.0000 96.3000 198.8000 96.4000 ;
	    RECT 214.0000 96.3000 214.8000 96.4000 ;
	    RECT 198.0000 95.7000 214.8000 96.3000 ;
	    RECT 198.0000 95.6000 198.8000 95.7000 ;
	    RECT 214.0000 95.6000 214.8000 95.7000 ;
	    RECT 222.0000 96.3000 222.8000 96.4000 ;
	    RECT 226.9000 96.3000 227.5000 97.7000 ;
	    RECT 239.6000 97.6000 240.4000 97.7000 ;
	    RECT 241.2000 98.3000 242.0000 98.4000 ;
	    RECT 450.8000 98.3000 451.6000 98.4000 ;
	    RECT 241.2000 97.7000 451.6000 98.3000 ;
	    RECT 241.2000 97.6000 242.0000 97.7000 ;
	    RECT 450.8000 97.6000 451.6000 97.7000 ;
	    RECT 222.0000 95.7000 227.5000 96.3000 ;
	    RECT 230.0000 96.3000 230.8000 96.4000 ;
	    RECT 241.2000 96.3000 242.0000 96.4000 ;
	    RECT 310.0000 96.3000 310.8000 96.4000 ;
	    RECT 230.0000 95.7000 242.0000 96.3000 ;
	    RECT 222.0000 95.6000 222.8000 95.7000 ;
	    RECT 230.0000 95.6000 230.8000 95.7000 ;
	    RECT 241.2000 95.6000 242.0000 95.7000 ;
	    RECT 242.9000 95.7000 310.8000 96.3000 ;
	    RECT 138.8000 94.3000 139.6000 94.4000 ;
	    RECT 121.3000 93.7000 139.6000 94.3000 ;
	    RECT 118.0000 93.6000 118.8000 93.7000 ;
	    RECT 119.6000 93.6000 120.4000 93.7000 ;
	    RECT 138.8000 93.6000 139.6000 93.7000 ;
	    RECT 145.2000 94.3000 146.0000 94.4000 ;
	    RECT 164.4000 94.3000 165.2000 94.4000 ;
	    RECT 175.6000 94.3000 176.4000 94.4000 ;
	    RECT 145.2000 93.7000 176.4000 94.3000 ;
	    RECT 145.2000 93.6000 146.0000 93.7000 ;
	    RECT 164.4000 93.6000 165.2000 93.7000 ;
	    RECT 175.6000 93.6000 176.4000 93.7000 ;
	    RECT 182.0000 93.6000 182.8000 94.4000 ;
	    RECT 186.8000 94.3000 187.6000 94.4000 ;
	    RECT 209.2000 94.3000 210.0000 94.4000 ;
	    RECT 186.8000 93.7000 210.0000 94.3000 ;
	    RECT 186.8000 93.6000 187.6000 93.7000 ;
	    RECT 209.2000 93.6000 210.0000 93.7000 ;
	    RECT 215.6000 94.3000 216.4000 94.4000 ;
	    RECT 242.9000 94.3000 243.5000 95.7000 ;
	    RECT 310.0000 95.6000 310.8000 95.7000 ;
	    RECT 318.0000 96.3000 318.8000 96.4000 ;
	    RECT 351.6000 96.3000 352.4000 96.4000 ;
	    RECT 439.6000 96.3000 440.4000 96.4000 ;
	    RECT 458.8000 96.3000 459.6000 96.4000 ;
	    RECT 318.0000 95.7000 352.4000 96.3000 ;
	    RECT 318.0000 95.6000 318.8000 95.7000 ;
	    RECT 351.6000 95.6000 352.4000 95.7000 ;
	    RECT 353.3000 95.7000 459.6000 96.3000 ;
	    RECT 215.6000 93.7000 243.5000 94.3000 ;
	    RECT 244.4000 94.3000 245.2000 94.4000 ;
	    RECT 262.0000 94.3000 262.8000 94.4000 ;
	    RECT 244.4000 93.7000 262.8000 94.3000 ;
	    RECT 215.6000 93.6000 216.4000 93.7000 ;
	    RECT 244.4000 93.6000 245.2000 93.7000 ;
	    RECT 262.0000 93.6000 262.8000 93.7000 ;
	    RECT 276.4000 94.3000 277.2000 94.4000 ;
	    RECT 284.4000 94.3000 285.2000 94.4000 ;
	    RECT 276.4000 93.7000 285.2000 94.3000 ;
	    RECT 276.4000 93.6000 277.2000 93.7000 ;
	    RECT 284.4000 93.6000 285.2000 93.7000 ;
	    RECT 287.6000 94.3000 288.4000 94.4000 ;
	    RECT 290.8000 94.3000 291.6000 94.4000 ;
	    RECT 287.6000 93.7000 291.6000 94.3000 ;
	    RECT 287.6000 93.6000 288.4000 93.7000 ;
	    RECT 290.8000 93.6000 291.6000 93.7000 ;
	    RECT 292.4000 94.3000 293.2000 94.4000 ;
	    RECT 295.6000 94.3000 296.4000 94.4000 ;
	    RECT 314.8000 94.3000 315.6000 94.4000 ;
	    RECT 292.4000 93.7000 315.6000 94.3000 ;
	    RECT 292.4000 93.6000 293.2000 93.7000 ;
	    RECT 295.6000 93.6000 296.4000 93.7000 ;
	    RECT 314.8000 93.6000 315.6000 93.7000 ;
	    RECT 324.4000 94.3000 325.2000 94.4000 ;
	    RECT 335.6000 94.3000 336.4000 94.4000 ;
	    RECT 324.4000 93.7000 336.4000 94.3000 ;
	    RECT 324.4000 93.6000 325.2000 93.7000 ;
	    RECT 335.6000 93.6000 336.4000 93.7000 ;
	    RECT 343.6000 94.3000 344.4000 94.4000 ;
	    RECT 353.3000 94.3000 353.9000 95.7000 ;
	    RECT 439.6000 95.6000 440.4000 95.7000 ;
	    RECT 458.8000 95.6000 459.6000 95.7000 ;
	    RECT 481.2000 96.3000 482.0000 96.4000 ;
	    RECT 487.6000 96.3000 488.4000 96.4000 ;
	    RECT 481.2000 95.7000 488.4000 96.3000 ;
	    RECT 481.2000 95.6000 482.0000 95.7000 ;
	    RECT 487.6000 95.6000 488.4000 95.7000 ;
	    RECT 343.6000 93.7000 353.9000 94.3000 ;
	    RECT 359.6000 94.3000 360.4000 94.4000 ;
	    RECT 362.8000 94.3000 363.6000 94.4000 ;
	    RECT 359.6000 93.7000 363.6000 94.3000 ;
	    RECT 343.6000 93.6000 344.4000 93.7000 ;
	    RECT 359.6000 93.6000 360.4000 93.7000 ;
	    RECT 362.8000 93.6000 363.6000 93.7000 ;
	    RECT 404.4000 94.3000 405.2000 94.4000 ;
	    RECT 430.0000 94.3000 430.8000 94.4000 ;
	    RECT 447.6000 94.3000 448.4000 94.4000 ;
	    RECT 404.4000 93.7000 448.4000 94.3000 ;
	    RECT 404.4000 93.6000 405.2000 93.7000 ;
	    RECT 430.0000 93.6000 430.8000 93.7000 ;
	    RECT 447.6000 93.6000 448.4000 93.7000 ;
	    RECT 452.4000 94.3000 453.2000 94.4000 ;
	    RECT 465.2000 94.3000 466.0000 94.4000 ;
	    RECT 452.4000 93.7000 466.0000 94.3000 ;
	    RECT 452.4000 93.6000 453.2000 93.7000 ;
	    RECT 465.2000 93.6000 466.0000 93.7000 ;
	    RECT 468.4000 94.3000 469.2000 94.4000 ;
	    RECT 494.0000 94.3000 494.8000 94.4000 ;
	    RECT 468.4000 93.7000 494.8000 94.3000 ;
	    RECT 468.4000 93.6000 469.2000 93.7000 ;
	    RECT 494.0000 93.6000 494.8000 93.7000 ;
	    RECT 502.0000 94.3000 502.8000 94.4000 ;
	    RECT 505.2000 94.3000 506.0000 94.4000 ;
	    RECT 502.0000 93.7000 506.0000 94.3000 ;
	    RECT 502.0000 93.6000 502.8000 93.7000 ;
	    RECT 505.2000 93.6000 506.0000 93.7000 ;
	    RECT 4.4000 92.3000 5.2000 92.4000 ;
	    RECT 10.8000 92.3000 11.6000 92.4000 ;
	    RECT 4.4000 91.7000 11.6000 92.3000 ;
	    RECT 4.4000 91.6000 5.2000 91.7000 ;
	    RECT 10.8000 91.6000 11.6000 91.7000 ;
	    RECT 14.0000 92.3000 14.8000 92.4000 ;
	    RECT 25.2000 92.3000 26.0000 92.4000 ;
	    RECT 14.0000 91.7000 26.0000 92.3000 ;
	    RECT 14.0000 91.6000 14.8000 91.7000 ;
	    RECT 25.2000 91.6000 26.0000 91.7000 ;
	    RECT 28.4000 92.3000 29.2000 92.4000 ;
	    RECT 49.2000 92.3000 50.0000 92.4000 ;
	    RECT 28.4000 91.7000 50.0000 92.3000 ;
	    RECT 28.4000 91.6000 29.2000 91.7000 ;
	    RECT 49.2000 91.6000 50.0000 91.7000 ;
	    RECT 63.6000 92.3000 64.4000 92.4000 ;
	    RECT 68.4000 92.3000 69.2000 92.4000 ;
	    RECT 63.6000 91.7000 69.2000 92.3000 ;
	    RECT 63.6000 91.6000 64.4000 91.7000 ;
	    RECT 68.4000 91.6000 69.2000 91.7000 ;
	    RECT 73.2000 92.3000 74.0000 92.4000 ;
	    RECT 82.8000 92.3000 83.6000 92.4000 ;
	    RECT 73.2000 91.7000 83.6000 92.3000 ;
	    RECT 73.2000 91.6000 74.0000 91.7000 ;
	    RECT 82.8000 91.6000 83.6000 91.7000 ;
	    RECT 98.8000 92.3000 99.6000 92.4000 ;
	    RECT 111.6000 92.3000 112.4000 92.4000 ;
	    RECT 98.8000 91.7000 112.4000 92.3000 ;
	    RECT 98.8000 91.6000 99.6000 91.7000 ;
	    RECT 111.6000 91.6000 112.4000 91.7000 ;
	    RECT 116.4000 91.6000 117.2000 92.4000 ;
	    RECT 118.0000 92.3000 118.8000 92.4000 ;
	    RECT 121.2000 92.3000 122.0000 92.4000 ;
	    RECT 118.0000 91.7000 122.0000 92.3000 ;
	    RECT 118.0000 91.6000 118.8000 91.7000 ;
	    RECT 121.2000 91.6000 122.0000 91.7000 ;
	    RECT 122.8000 92.3000 123.6000 92.4000 ;
	    RECT 134.0000 92.3000 134.8000 92.4000 ;
	    RECT 122.8000 91.7000 134.8000 92.3000 ;
	    RECT 122.8000 91.6000 123.6000 91.7000 ;
	    RECT 134.0000 91.6000 134.8000 91.7000 ;
	    RECT 137.2000 92.3000 138.0000 92.4000 ;
	    RECT 145.2000 92.3000 146.0000 92.4000 ;
	    RECT 137.2000 91.7000 146.0000 92.3000 ;
	    RECT 137.2000 91.6000 138.0000 91.7000 ;
	    RECT 145.2000 91.6000 146.0000 91.7000 ;
	    RECT 151.6000 92.3000 152.4000 92.4000 ;
	    RECT 159.6000 92.3000 160.4000 92.4000 ;
	    RECT 151.6000 91.7000 160.4000 92.3000 ;
	    RECT 151.6000 91.6000 152.4000 91.7000 ;
	    RECT 159.6000 91.6000 160.4000 91.7000 ;
	    RECT 161.2000 92.3000 162.0000 92.4000 ;
	    RECT 174.0000 92.3000 174.8000 92.4000 ;
	    RECT 177.2000 92.3000 178.0000 92.4000 ;
	    RECT 161.2000 91.7000 173.1000 92.3000 ;
	    RECT 161.2000 91.6000 162.0000 91.7000 ;
	    RECT 9.2000 90.3000 10.0000 90.4000 ;
	    RECT 28.4000 90.3000 29.2000 90.4000 ;
	    RECT 9.2000 89.7000 29.2000 90.3000 ;
	    RECT 9.2000 89.6000 10.0000 89.7000 ;
	    RECT 28.4000 89.6000 29.2000 89.7000 ;
	    RECT 74.8000 90.3000 75.6000 90.4000 ;
	    RECT 126.0000 90.3000 126.8000 90.4000 ;
	    RECT 74.8000 89.7000 126.8000 90.3000 ;
	    RECT 74.8000 89.6000 75.6000 89.7000 ;
	    RECT 126.0000 89.6000 126.8000 89.7000 ;
	    RECT 129.2000 90.3000 130.0000 90.4000 ;
	    RECT 138.8000 90.3000 139.6000 90.4000 ;
	    RECT 129.2000 89.7000 139.6000 90.3000 ;
	    RECT 129.2000 89.6000 130.0000 89.7000 ;
	    RECT 138.8000 89.6000 139.6000 89.7000 ;
	    RECT 140.4000 90.3000 141.2000 90.4000 ;
	    RECT 153.2000 90.3000 154.0000 90.4000 ;
	    RECT 140.4000 89.7000 154.0000 90.3000 ;
	    RECT 140.4000 89.6000 141.2000 89.7000 ;
	    RECT 153.2000 89.6000 154.0000 89.7000 ;
	    RECT 159.6000 90.3000 160.4000 90.4000 ;
	    RECT 170.8000 90.3000 171.6000 90.4000 ;
	    RECT 159.6000 89.7000 171.6000 90.3000 ;
	    RECT 172.5000 90.3000 173.1000 91.7000 ;
	    RECT 174.0000 91.7000 178.0000 92.3000 ;
	    RECT 174.0000 91.6000 174.8000 91.7000 ;
	    RECT 177.2000 91.6000 178.0000 91.7000 ;
	    RECT 185.2000 92.3000 186.0000 92.4000 ;
	    RECT 193.2000 92.3000 194.0000 92.4000 ;
	    RECT 185.2000 91.7000 194.0000 92.3000 ;
	    RECT 185.2000 91.6000 186.0000 91.7000 ;
	    RECT 193.2000 91.6000 194.0000 91.7000 ;
	    RECT 194.8000 92.3000 195.6000 92.4000 ;
	    RECT 194.8000 91.7000 201.9000 92.3000 ;
	    RECT 194.8000 91.6000 195.6000 91.7000 ;
	    RECT 186.8000 90.3000 187.6000 90.4000 ;
	    RECT 172.5000 89.7000 187.6000 90.3000 ;
	    RECT 159.6000 89.6000 160.4000 89.7000 ;
	    RECT 170.8000 89.6000 171.6000 89.7000 ;
	    RECT 186.8000 89.6000 187.6000 89.7000 ;
	    RECT 193.2000 90.3000 194.0000 90.4000 ;
	    RECT 199.6000 90.3000 200.4000 90.4000 ;
	    RECT 193.2000 89.7000 200.4000 90.3000 ;
	    RECT 201.3000 90.3000 201.9000 91.7000 ;
	    RECT 202.8000 91.6000 203.6000 92.4000 ;
	    RECT 207.6000 92.3000 208.4000 92.4000 ;
	    RECT 222.0000 92.3000 222.8000 92.4000 ;
	    RECT 230.0000 92.3000 230.8000 92.4000 ;
	    RECT 207.6000 91.7000 230.8000 92.3000 ;
	    RECT 207.6000 91.6000 208.4000 91.7000 ;
	    RECT 222.0000 91.6000 222.8000 91.7000 ;
	    RECT 230.0000 91.6000 230.8000 91.7000 ;
	    RECT 233.2000 92.3000 234.0000 92.4000 ;
	    RECT 238.0000 92.3000 238.8000 92.4000 ;
	    RECT 233.2000 91.7000 238.8000 92.3000 ;
	    RECT 233.2000 91.6000 234.0000 91.7000 ;
	    RECT 238.0000 91.6000 238.8000 91.7000 ;
	    RECT 247.6000 92.3000 248.4000 92.4000 ;
	    RECT 263.6000 92.3000 264.4000 92.4000 ;
	    RECT 278.0000 92.3000 278.8000 92.4000 ;
	    RECT 247.6000 91.7000 254.7000 92.3000 ;
	    RECT 247.6000 91.6000 248.4000 91.7000 ;
	    RECT 218.8000 90.3000 219.6000 90.4000 ;
	    RECT 201.3000 89.7000 219.6000 90.3000 ;
	    RECT 193.2000 89.6000 194.0000 89.7000 ;
	    RECT 199.6000 89.6000 200.4000 89.7000 ;
	    RECT 218.8000 89.6000 219.6000 89.7000 ;
	    RECT 238.0000 90.3000 238.8000 90.4000 ;
	    RECT 252.4000 90.3000 253.2000 90.4000 ;
	    RECT 238.0000 89.7000 253.2000 90.3000 ;
	    RECT 254.1000 90.3000 254.7000 91.7000 ;
	    RECT 263.6000 91.7000 278.8000 92.3000 ;
	    RECT 263.6000 91.6000 264.4000 91.7000 ;
	    RECT 278.0000 91.6000 278.8000 91.7000 ;
	    RECT 289.2000 92.3000 290.0000 92.4000 ;
	    RECT 322.8000 92.3000 323.6000 92.4000 ;
	    RECT 289.2000 91.7000 323.6000 92.3000 ;
	    RECT 289.2000 91.6000 290.0000 91.7000 ;
	    RECT 322.8000 91.6000 323.6000 91.7000 ;
	    RECT 326.0000 92.3000 326.8000 92.4000 ;
	    RECT 338.8000 92.3000 339.6000 92.4000 ;
	    RECT 326.0000 91.7000 339.6000 92.3000 ;
	    RECT 326.0000 91.6000 326.8000 91.7000 ;
	    RECT 338.8000 91.6000 339.6000 91.7000 ;
	    RECT 356.4000 92.3000 357.2000 92.4000 ;
	    RECT 364.4000 92.3000 365.2000 92.4000 ;
	    RECT 356.4000 91.7000 365.2000 92.3000 ;
	    RECT 356.4000 91.6000 357.2000 91.7000 ;
	    RECT 364.4000 91.6000 365.2000 91.7000 ;
	    RECT 374.0000 92.3000 374.8000 92.4000 ;
	    RECT 382.0000 92.3000 382.8000 92.4000 ;
	    RECT 374.0000 91.7000 382.8000 92.3000 ;
	    RECT 374.0000 91.6000 374.8000 91.7000 ;
	    RECT 382.0000 91.6000 382.8000 91.7000 ;
	    RECT 383.6000 92.3000 384.4000 92.4000 ;
	    RECT 396.4000 92.3000 397.2000 92.4000 ;
	    RECT 383.6000 91.7000 397.2000 92.3000 ;
	    RECT 383.6000 91.6000 384.4000 91.7000 ;
	    RECT 396.4000 91.6000 397.2000 91.7000 ;
	    RECT 426.8000 92.3000 427.6000 92.4000 ;
	    RECT 434.8000 92.3000 435.6000 92.4000 ;
	    RECT 426.8000 91.7000 435.6000 92.3000 ;
	    RECT 426.8000 91.6000 427.6000 91.7000 ;
	    RECT 434.8000 91.6000 435.6000 91.7000 ;
	    RECT 438.0000 92.3000 438.8000 92.4000 ;
	    RECT 462.0000 92.3000 462.8000 92.4000 ;
	    RECT 438.0000 91.7000 462.8000 92.3000 ;
	    RECT 438.0000 91.6000 438.8000 91.7000 ;
	    RECT 462.0000 91.6000 462.8000 91.7000 ;
	    RECT 463.6000 92.3000 464.4000 92.4000 ;
	    RECT 478.0000 92.3000 478.8000 92.4000 ;
	    RECT 492.4000 92.3000 493.2000 92.4000 ;
	    RECT 463.6000 91.7000 493.2000 92.3000 ;
	    RECT 463.6000 91.6000 464.4000 91.7000 ;
	    RECT 478.0000 91.6000 478.8000 91.7000 ;
	    RECT 492.4000 91.6000 493.2000 91.7000 ;
	    RECT 279.6000 90.3000 280.4000 90.4000 ;
	    RECT 254.1000 89.7000 280.4000 90.3000 ;
	    RECT 238.0000 89.6000 238.8000 89.7000 ;
	    RECT 252.4000 89.6000 253.2000 89.7000 ;
	    RECT 279.6000 89.6000 280.4000 89.7000 ;
	    RECT 281.2000 90.3000 282.0000 90.4000 ;
	    RECT 298.8000 90.3000 299.6000 90.4000 ;
	    RECT 308.4000 90.3000 309.2000 90.4000 ;
	    RECT 281.2000 89.7000 309.2000 90.3000 ;
	    RECT 281.2000 89.6000 282.0000 89.7000 ;
	    RECT 298.8000 89.6000 299.6000 89.7000 ;
	    RECT 308.4000 89.6000 309.2000 89.7000 ;
	    RECT 310.0000 90.3000 310.8000 90.4000 ;
	    RECT 468.4000 90.3000 469.2000 90.4000 ;
	    RECT 310.0000 89.7000 469.2000 90.3000 ;
	    RECT 310.0000 89.6000 310.8000 89.7000 ;
	    RECT 468.4000 89.6000 469.2000 89.7000 ;
	    RECT 14.0000 88.3000 14.8000 88.4000 ;
	    RECT 17.2000 88.3000 18.0000 88.4000 ;
	    RECT 14.0000 87.7000 18.0000 88.3000 ;
	    RECT 14.0000 87.6000 14.8000 87.7000 ;
	    RECT 17.2000 87.6000 18.0000 87.7000 ;
	    RECT 55.6000 88.3000 56.4000 88.4000 ;
	    RECT 81.2000 88.3000 82.0000 88.4000 ;
	    RECT 55.6000 87.7000 82.0000 88.3000 ;
	    RECT 55.6000 87.6000 56.4000 87.7000 ;
	    RECT 81.2000 87.6000 82.0000 87.7000 ;
	    RECT 82.8000 88.3000 83.6000 88.4000 ;
	    RECT 161.2000 88.3000 162.0000 88.4000 ;
	    RECT 82.8000 87.7000 162.0000 88.3000 ;
	    RECT 82.8000 87.6000 83.6000 87.7000 ;
	    RECT 161.2000 87.6000 162.0000 87.7000 ;
	    RECT 162.8000 88.3000 163.6000 88.4000 ;
	    RECT 166.0000 88.3000 166.8000 88.4000 ;
	    RECT 169.2000 88.3000 170.0000 88.4000 ;
	    RECT 215.6000 88.3000 216.4000 88.4000 ;
	    RECT 460.4000 88.3000 461.2000 88.4000 ;
	    RECT 162.8000 87.7000 166.8000 88.3000 ;
	    RECT 162.8000 87.6000 163.6000 87.7000 ;
	    RECT 166.0000 87.6000 166.8000 87.7000 ;
	    RECT 167.7000 87.7000 461.2000 88.3000 ;
	    RECT 90.8000 86.3000 91.6000 86.4000 ;
	    RECT 100.4000 86.3000 101.2000 86.4000 ;
	    RECT 153.2000 86.3000 154.0000 86.4000 ;
	    RECT 167.7000 86.3000 168.3000 87.7000 ;
	    RECT 169.2000 87.6000 170.0000 87.7000 ;
	    RECT 215.6000 87.6000 216.4000 87.7000 ;
	    RECT 460.4000 87.6000 461.2000 87.7000 ;
	    RECT 466.8000 88.3000 467.6000 88.4000 ;
	    RECT 498.8000 88.3000 499.6000 88.4000 ;
	    RECT 466.8000 87.7000 499.6000 88.3000 ;
	    RECT 466.8000 87.6000 467.6000 87.7000 ;
	    RECT 498.8000 87.6000 499.6000 87.7000 ;
	    RECT 226.8000 86.3000 227.6000 86.4000 ;
	    RECT 90.8000 85.7000 168.3000 86.3000 ;
	    RECT 169.3000 85.7000 227.6000 86.3000 ;
	    RECT 90.8000 85.6000 91.6000 85.7000 ;
	    RECT 100.4000 85.6000 101.2000 85.7000 ;
	    RECT 153.2000 85.6000 154.0000 85.7000 ;
	    RECT 33.2000 84.3000 34.0000 84.4000 ;
	    RECT 65.2000 84.3000 66.0000 84.4000 ;
	    RECT 33.2000 83.7000 66.0000 84.3000 ;
	    RECT 33.2000 83.6000 34.0000 83.7000 ;
	    RECT 65.2000 83.6000 66.0000 83.7000 ;
	    RECT 74.8000 84.3000 75.6000 84.4000 ;
	    RECT 119.6000 84.3000 120.4000 84.4000 ;
	    RECT 74.8000 83.7000 120.4000 84.3000 ;
	    RECT 74.8000 83.6000 75.6000 83.7000 ;
	    RECT 119.6000 83.6000 120.4000 83.7000 ;
	    RECT 121.2000 84.3000 122.0000 84.4000 ;
	    RECT 169.3000 84.3000 169.9000 85.7000 ;
	    RECT 226.8000 85.6000 227.6000 85.7000 ;
	    RECT 234.8000 86.3000 235.6000 86.4000 ;
	    RECT 249.2000 86.3000 250.0000 86.4000 ;
	    RECT 281.2000 86.3000 282.0000 86.4000 ;
	    RECT 234.8000 85.7000 282.0000 86.3000 ;
	    RECT 234.8000 85.6000 235.6000 85.7000 ;
	    RECT 249.2000 85.6000 250.0000 85.7000 ;
	    RECT 281.2000 85.6000 282.0000 85.7000 ;
	    RECT 282.8000 86.3000 283.6000 86.4000 ;
	    RECT 289.2000 86.3000 290.0000 86.4000 ;
	    RECT 282.8000 85.7000 290.0000 86.3000 ;
	    RECT 282.8000 85.6000 283.6000 85.7000 ;
	    RECT 289.2000 85.6000 290.0000 85.7000 ;
	    RECT 292.4000 86.3000 293.2000 86.4000 ;
	    RECT 313.2000 86.3000 314.0000 86.4000 ;
	    RECT 350.0000 86.3000 350.8000 86.4000 ;
	    RECT 369.2000 86.3000 370.0000 86.4000 ;
	    RECT 292.4000 85.7000 370.0000 86.3000 ;
	    RECT 292.4000 85.6000 293.2000 85.7000 ;
	    RECT 313.2000 85.6000 314.0000 85.7000 ;
	    RECT 350.0000 85.6000 350.8000 85.7000 ;
	    RECT 369.2000 85.6000 370.0000 85.7000 ;
	    RECT 385.2000 86.3000 386.0000 86.4000 ;
	    RECT 388.4000 86.3000 389.2000 86.4000 ;
	    RECT 385.2000 85.7000 389.2000 86.3000 ;
	    RECT 385.2000 85.6000 386.0000 85.7000 ;
	    RECT 388.4000 85.6000 389.2000 85.7000 ;
	    RECT 407.6000 86.3000 408.4000 86.4000 ;
	    RECT 430.0000 86.3000 430.8000 86.4000 ;
	    RECT 407.6000 85.7000 430.8000 86.3000 ;
	    RECT 407.6000 85.6000 408.4000 85.7000 ;
	    RECT 430.0000 85.6000 430.8000 85.7000 ;
	    RECT 462.0000 86.3000 462.8000 86.4000 ;
	    RECT 474.8000 86.3000 475.6000 86.4000 ;
	    RECT 462.0000 85.7000 475.6000 86.3000 ;
	    RECT 462.0000 85.6000 462.8000 85.7000 ;
	    RECT 474.8000 85.6000 475.6000 85.7000 ;
	    RECT 121.2000 83.7000 169.9000 84.3000 ;
	    RECT 121.2000 83.6000 122.0000 83.7000 ;
	    RECT 174.0000 83.6000 174.8000 84.4000 ;
	    RECT 177.2000 84.3000 178.0000 84.4000 ;
	    RECT 220.4000 84.3000 221.2000 84.4000 ;
	    RECT 177.2000 83.7000 221.2000 84.3000 ;
	    RECT 177.2000 83.6000 178.0000 83.7000 ;
	    RECT 220.4000 83.6000 221.2000 83.7000 ;
	    RECT 223.6000 84.3000 224.4000 84.4000 ;
	    RECT 230.0000 84.3000 230.8000 84.4000 ;
	    RECT 255.6000 84.3000 256.4000 84.4000 ;
	    RECT 292.5000 84.3000 293.1000 85.6000 ;
	    RECT 223.6000 83.7000 293.1000 84.3000 ;
	    RECT 294.0000 84.3000 294.8000 84.4000 ;
	    RECT 302.0000 84.3000 302.8000 84.4000 ;
	    RECT 294.0000 83.7000 302.8000 84.3000 ;
	    RECT 223.6000 83.6000 224.4000 83.7000 ;
	    RECT 230.0000 83.6000 230.8000 83.7000 ;
	    RECT 255.6000 83.6000 256.4000 83.7000 ;
	    RECT 294.0000 83.6000 294.8000 83.7000 ;
	    RECT 302.0000 83.6000 302.8000 83.7000 ;
	    RECT 303.6000 84.3000 304.4000 84.4000 ;
	    RECT 358.0000 84.3000 358.8000 84.4000 ;
	    RECT 303.6000 83.7000 358.8000 84.3000 ;
	    RECT 303.6000 83.6000 304.4000 83.7000 ;
	    RECT 358.0000 83.6000 358.8000 83.7000 ;
	    RECT 382.0000 84.3000 382.8000 84.4000 ;
	    RECT 439.6000 84.3000 440.4000 84.4000 ;
	    RECT 382.0000 83.7000 440.4000 84.3000 ;
	    RECT 382.0000 83.6000 382.8000 83.7000 ;
	    RECT 439.6000 83.6000 440.4000 83.7000 ;
	    RECT 78.0000 82.3000 78.8000 82.4000 ;
	    RECT 97.2000 82.3000 98.0000 82.4000 ;
	    RECT 78.0000 81.7000 98.0000 82.3000 ;
	    RECT 78.0000 81.6000 78.8000 81.7000 ;
	    RECT 97.2000 81.6000 98.0000 81.7000 ;
	    RECT 135.6000 82.3000 136.4000 82.4000 ;
	    RECT 246.0000 82.3000 246.8000 82.4000 ;
	    RECT 135.6000 81.7000 246.8000 82.3000 ;
	    RECT 135.6000 81.6000 136.4000 81.7000 ;
	    RECT 246.0000 81.6000 246.8000 81.7000 ;
	    RECT 247.6000 82.3000 248.4000 82.4000 ;
	    RECT 273.2000 82.3000 274.0000 82.4000 ;
	    RECT 297.2000 82.3000 298.0000 82.4000 ;
	    RECT 247.6000 81.7000 298.0000 82.3000 ;
	    RECT 247.6000 81.6000 248.4000 81.7000 ;
	    RECT 273.2000 81.6000 274.0000 81.7000 ;
	    RECT 297.2000 81.6000 298.0000 81.7000 ;
	    RECT 308.4000 82.3000 309.2000 82.4000 ;
	    RECT 361.2000 82.3000 362.0000 82.4000 ;
	    RECT 377.2000 82.3000 378.0000 82.4000 ;
	    RECT 308.4000 81.7000 378.0000 82.3000 ;
	    RECT 308.4000 81.6000 309.2000 81.7000 ;
	    RECT 361.2000 81.6000 362.0000 81.7000 ;
	    RECT 377.2000 81.6000 378.0000 81.7000 ;
	    RECT 68.4000 80.3000 69.2000 80.4000 ;
	    RECT 102.0000 80.3000 102.8000 80.4000 ;
	    RECT 68.4000 79.7000 102.8000 80.3000 ;
	    RECT 68.4000 79.6000 69.2000 79.7000 ;
	    RECT 102.0000 79.6000 102.8000 79.7000 ;
	    RECT 114.8000 80.3000 115.6000 80.4000 ;
	    RECT 167.6000 80.3000 168.4000 80.4000 ;
	    RECT 114.8000 79.7000 168.4000 80.3000 ;
	    RECT 114.8000 79.6000 115.6000 79.7000 ;
	    RECT 167.6000 79.6000 168.4000 79.7000 ;
	    RECT 169.2000 80.3000 170.0000 80.4000 ;
	    RECT 206.0000 80.3000 206.8000 80.4000 ;
	    RECT 169.2000 79.7000 206.8000 80.3000 ;
	    RECT 169.2000 79.6000 170.0000 79.7000 ;
	    RECT 206.0000 79.6000 206.8000 79.7000 ;
	    RECT 209.2000 80.3000 210.0000 80.4000 ;
	    RECT 217.2000 80.3000 218.0000 80.4000 ;
	    RECT 239.6000 80.3000 240.4000 80.4000 ;
	    RECT 209.2000 79.7000 265.9000 80.3000 ;
	    RECT 209.2000 79.6000 210.0000 79.7000 ;
	    RECT 217.2000 79.6000 218.0000 79.7000 ;
	    RECT 239.6000 79.6000 240.4000 79.7000 ;
	    RECT 100.4000 78.3000 101.2000 78.4000 ;
	    RECT 118.0000 78.3000 118.8000 78.4000 ;
	    RECT 100.4000 77.7000 118.8000 78.3000 ;
	    RECT 100.4000 77.6000 101.2000 77.7000 ;
	    RECT 118.0000 77.6000 118.8000 77.7000 ;
	    RECT 119.6000 78.3000 120.4000 78.4000 ;
	    RECT 231.6000 78.3000 232.4000 78.4000 ;
	    RECT 119.6000 77.7000 232.4000 78.3000 ;
	    RECT 119.6000 77.6000 120.4000 77.7000 ;
	    RECT 231.6000 77.6000 232.4000 77.7000 ;
	    RECT 233.2000 78.3000 234.0000 78.4000 ;
	    RECT 234.8000 78.3000 235.6000 78.4000 ;
	    RECT 233.2000 77.7000 235.6000 78.3000 ;
	    RECT 233.2000 77.6000 234.0000 77.7000 ;
	    RECT 234.8000 77.6000 235.6000 77.7000 ;
	    RECT 238.0000 78.3000 238.8000 78.4000 ;
	    RECT 263.6000 78.3000 264.4000 78.4000 ;
	    RECT 238.0000 77.7000 264.4000 78.3000 ;
	    RECT 265.3000 78.3000 265.9000 79.7000 ;
	    RECT 266.8000 79.6000 267.6000 80.4000 ;
	    RECT 268.4000 80.3000 269.2000 80.4000 ;
	    RECT 274.8000 80.3000 275.6000 80.4000 ;
	    RECT 268.4000 79.7000 275.6000 80.3000 ;
	    RECT 268.4000 79.6000 269.2000 79.7000 ;
	    RECT 274.8000 79.6000 275.6000 79.7000 ;
	    RECT 276.4000 79.6000 277.2000 80.4000 ;
	    RECT 278.0000 80.3000 278.8000 80.4000 ;
	    RECT 303.6000 80.3000 304.4000 80.4000 ;
	    RECT 278.0000 79.7000 304.4000 80.3000 ;
	    RECT 278.0000 79.6000 278.8000 79.7000 ;
	    RECT 303.6000 79.6000 304.4000 79.7000 ;
	    RECT 314.8000 80.3000 315.6000 80.4000 ;
	    RECT 380.4000 80.3000 381.2000 80.4000 ;
	    RECT 388.4000 80.3000 389.2000 80.4000 ;
	    RECT 314.8000 79.7000 389.2000 80.3000 ;
	    RECT 314.8000 79.6000 315.6000 79.7000 ;
	    RECT 380.4000 79.6000 381.2000 79.7000 ;
	    RECT 388.4000 79.6000 389.2000 79.7000 ;
	    RECT 455.6000 80.3000 456.4000 80.4000 ;
	    RECT 462.0000 80.3000 462.8000 80.4000 ;
	    RECT 455.6000 79.7000 462.8000 80.3000 ;
	    RECT 455.6000 79.6000 456.4000 79.7000 ;
	    RECT 462.0000 79.6000 462.8000 79.7000 ;
	    RECT 465.2000 80.3000 466.0000 80.4000 ;
	    RECT 486.0000 80.3000 486.8000 80.4000 ;
	    RECT 500.4000 80.3000 501.2000 80.4000 ;
	    RECT 505.2000 80.3000 506.0000 80.4000 ;
	    RECT 465.2000 79.7000 506.0000 80.3000 ;
	    RECT 465.2000 79.6000 466.0000 79.7000 ;
	    RECT 486.0000 79.6000 486.8000 79.7000 ;
	    RECT 500.4000 79.6000 501.2000 79.7000 ;
	    RECT 505.2000 79.6000 506.0000 79.7000 ;
	    RECT 327.6000 78.3000 328.4000 78.4000 ;
	    RECT 436.4000 78.3000 437.2000 78.4000 ;
	    RECT 265.3000 77.7000 437.2000 78.3000 ;
	    RECT 238.0000 77.6000 238.8000 77.7000 ;
	    RECT 263.6000 77.6000 264.4000 77.7000 ;
	    RECT 327.6000 77.6000 328.4000 77.7000 ;
	    RECT 436.4000 77.6000 437.2000 77.7000 ;
	    RECT 22.0000 76.3000 22.8000 76.4000 ;
	    RECT 174.0000 76.3000 174.8000 76.4000 ;
	    RECT 22.0000 75.7000 174.8000 76.3000 ;
	    RECT 22.0000 75.6000 22.8000 75.7000 ;
	    RECT 174.0000 75.6000 174.8000 75.7000 ;
	    RECT 175.6000 76.3000 176.4000 76.4000 ;
	    RECT 236.4000 76.3000 237.2000 76.4000 ;
	    RECT 175.6000 75.7000 237.2000 76.3000 ;
	    RECT 175.6000 75.6000 176.4000 75.7000 ;
	    RECT 236.4000 75.6000 237.2000 75.7000 ;
	    RECT 238.0000 76.3000 238.8000 76.4000 ;
	    RECT 262.0000 76.3000 262.8000 76.4000 ;
	    RECT 238.0000 75.7000 262.8000 76.3000 ;
	    RECT 238.0000 75.6000 238.8000 75.7000 ;
	    RECT 262.0000 75.6000 262.8000 75.7000 ;
	    RECT 263.6000 76.3000 264.4000 76.4000 ;
	    RECT 278.0000 76.3000 278.8000 76.4000 ;
	    RECT 263.6000 75.7000 278.8000 76.3000 ;
	    RECT 263.6000 75.6000 264.4000 75.7000 ;
	    RECT 278.0000 75.6000 278.8000 75.7000 ;
	    RECT 279.6000 76.3000 280.4000 76.4000 ;
	    RECT 290.8000 76.3000 291.6000 76.4000 ;
	    RECT 279.6000 75.7000 291.6000 76.3000 ;
	    RECT 279.6000 75.6000 280.4000 75.7000 ;
	    RECT 290.8000 75.6000 291.6000 75.7000 ;
	    RECT 292.4000 76.3000 293.2000 76.4000 ;
	    RECT 318.0000 76.3000 318.8000 76.4000 ;
	    RECT 498.8000 76.3000 499.6000 76.4000 ;
	    RECT 506.8000 76.3000 507.6000 76.4000 ;
	    RECT 292.4000 75.7000 318.8000 76.3000 ;
	    RECT 292.4000 75.6000 293.2000 75.7000 ;
	    RECT 318.0000 75.6000 318.8000 75.7000 ;
	    RECT 330.9000 75.7000 456.3000 76.3000 ;
	    RECT 4.4000 74.3000 5.2000 74.4000 ;
	    RECT 15.6000 74.3000 16.4000 74.4000 ;
	    RECT 39.6000 74.3000 40.4000 74.4000 ;
	    RECT 4.4000 73.7000 40.4000 74.3000 ;
	    RECT 4.4000 73.6000 5.2000 73.7000 ;
	    RECT 15.6000 73.6000 16.4000 73.7000 ;
	    RECT 39.6000 73.6000 40.4000 73.7000 ;
	    RECT 42.8000 74.3000 43.6000 74.4000 ;
	    RECT 50.8000 74.3000 51.6000 74.4000 ;
	    RECT 42.8000 73.7000 51.6000 74.3000 ;
	    RECT 42.8000 73.6000 43.6000 73.7000 ;
	    RECT 50.8000 73.6000 51.6000 73.7000 ;
	    RECT 63.6000 74.3000 64.4000 74.4000 ;
	    RECT 71.6000 74.3000 72.4000 74.4000 ;
	    RECT 63.6000 73.7000 72.4000 74.3000 ;
	    RECT 63.6000 73.6000 64.4000 73.7000 ;
	    RECT 71.6000 73.6000 72.4000 73.7000 ;
	    RECT 92.4000 74.3000 93.2000 74.4000 ;
	    RECT 105.2000 74.3000 106.0000 74.4000 ;
	    RECT 92.4000 73.7000 106.0000 74.3000 ;
	    RECT 92.4000 73.6000 93.2000 73.7000 ;
	    RECT 105.2000 73.6000 106.0000 73.7000 ;
	    RECT 106.8000 74.3000 107.6000 74.4000 ;
	    RECT 122.8000 74.3000 123.6000 74.4000 ;
	    RECT 106.8000 73.7000 123.6000 74.3000 ;
	    RECT 106.8000 73.6000 107.6000 73.7000 ;
	    RECT 122.8000 73.6000 123.6000 73.7000 ;
	    RECT 130.8000 74.3000 131.6000 74.4000 ;
	    RECT 140.4000 74.3000 141.2000 74.4000 ;
	    RECT 330.9000 74.3000 331.5000 75.7000 ;
	    RECT 455.7000 74.4000 456.3000 75.7000 ;
	    RECT 498.8000 75.7000 507.6000 76.3000 ;
	    RECT 498.8000 75.6000 499.6000 75.7000 ;
	    RECT 506.8000 75.6000 507.6000 75.7000 ;
	    RECT 130.8000 73.7000 331.5000 74.3000 ;
	    RECT 334.0000 74.3000 334.8000 74.4000 ;
	    RECT 348.4000 74.3000 349.2000 74.4000 ;
	    RECT 394.8000 74.3000 395.6000 74.4000 ;
	    RECT 414.0000 74.3000 414.8000 74.4000 ;
	    RECT 334.0000 73.7000 414.8000 74.3000 ;
	    RECT 130.8000 73.6000 131.6000 73.7000 ;
	    RECT 140.4000 73.6000 141.2000 73.7000 ;
	    RECT 334.0000 73.6000 334.8000 73.7000 ;
	    RECT 348.4000 73.6000 349.2000 73.7000 ;
	    RECT 394.8000 73.6000 395.6000 73.7000 ;
	    RECT 414.0000 73.6000 414.8000 73.7000 ;
	    RECT 455.6000 74.3000 456.4000 74.4000 ;
	    RECT 474.8000 74.3000 475.6000 74.4000 ;
	    RECT 455.6000 73.7000 475.6000 74.3000 ;
	    RECT 455.6000 73.6000 456.4000 73.7000 ;
	    RECT 474.8000 73.6000 475.6000 73.7000 ;
	    RECT 482.8000 74.3000 483.6000 74.4000 ;
	    RECT 503.6000 74.3000 504.4000 74.4000 ;
	    RECT 482.8000 73.7000 504.4000 74.3000 ;
	    RECT 482.8000 73.6000 483.6000 73.7000 ;
	    RECT 503.6000 73.6000 504.4000 73.7000 ;
	    RECT 34.8000 72.3000 35.6000 72.4000 ;
	    RECT 46.0000 72.3000 46.8000 72.4000 ;
	    RECT 34.8000 71.7000 46.8000 72.3000 ;
	    RECT 34.8000 71.6000 35.6000 71.7000 ;
	    RECT 46.0000 71.6000 46.8000 71.7000 ;
	    RECT 81.2000 72.3000 82.0000 72.4000 ;
	    RECT 94.0000 72.3000 94.8000 72.4000 ;
	    RECT 81.2000 71.7000 94.8000 72.3000 ;
	    RECT 81.2000 71.6000 82.0000 71.7000 ;
	    RECT 94.0000 71.6000 94.8000 71.7000 ;
	    RECT 103.6000 72.3000 104.4000 72.4000 ;
	    RECT 113.2000 72.3000 114.0000 72.4000 ;
	    RECT 103.6000 71.7000 114.0000 72.3000 ;
	    RECT 103.6000 71.6000 104.4000 71.7000 ;
	    RECT 113.2000 71.6000 114.0000 71.7000 ;
	    RECT 129.2000 72.3000 130.0000 72.4000 ;
	    RECT 134.0000 72.3000 134.8000 72.4000 ;
	    RECT 129.2000 71.7000 134.8000 72.3000 ;
	    RECT 129.2000 71.6000 130.0000 71.7000 ;
	    RECT 134.0000 71.6000 134.8000 71.7000 ;
	    RECT 158.0000 72.3000 158.8000 72.4000 ;
	    RECT 166.0000 72.3000 166.8000 72.4000 ;
	    RECT 158.0000 71.7000 166.8000 72.3000 ;
	    RECT 158.0000 71.6000 158.8000 71.7000 ;
	    RECT 166.0000 71.6000 166.8000 71.7000 ;
	    RECT 196.4000 72.3000 197.2000 72.4000 ;
	    RECT 210.8000 72.3000 211.6000 72.4000 ;
	    RECT 196.4000 71.7000 211.6000 72.3000 ;
	    RECT 196.4000 71.6000 197.2000 71.7000 ;
	    RECT 210.8000 71.6000 211.6000 71.7000 ;
	    RECT 215.6000 72.3000 216.4000 72.4000 ;
	    RECT 223.6000 72.3000 224.4000 72.4000 ;
	    RECT 234.8000 72.3000 235.6000 72.4000 ;
	    RECT 215.6000 71.7000 235.6000 72.3000 ;
	    RECT 215.6000 71.6000 216.4000 71.7000 ;
	    RECT 223.6000 71.6000 224.4000 71.7000 ;
	    RECT 234.8000 71.6000 235.6000 71.7000 ;
	    RECT 239.6000 72.3000 240.4000 72.4000 ;
	    RECT 257.2000 72.3000 258.0000 72.4000 ;
	    RECT 263.6000 72.3000 264.4000 72.4000 ;
	    RECT 239.6000 71.7000 253.1000 72.3000 ;
	    RECT 239.6000 71.6000 240.4000 71.7000 ;
	    RECT 28.4000 70.3000 29.2000 70.4000 ;
	    RECT 52.4000 70.3000 53.2000 70.4000 ;
	    RECT 28.4000 69.7000 53.2000 70.3000 ;
	    RECT 28.4000 69.6000 29.2000 69.7000 ;
	    RECT 52.4000 69.6000 53.2000 69.7000 ;
	    RECT 127.6000 70.3000 128.4000 70.4000 ;
	    RECT 132.4000 70.3000 133.2000 70.4000 ;
	    RECT 127.6000 69.7000 133.2000 70.3000 ;
	    RECT 127.6000 69.6000 128.4000 69.7000 ;
	    RECT 132.4000 69.6000 133.2000 69.7000 ;
	    RECT 134.0000 70.3000 134.8000 70.4000 ;
	    RECT 145.2000 70.3000 146.0000 70.4000 ;
	    RECT 134.0000 69.7000 146.0000 70.3000 ;
	    RECT 134.0000 69.6000 134.8000 69.7000 ;
	    RECT 145.2000 69.6000 146.0000 69.7000 ;
	    RECT 146.8000 70.3000 147.6000 70.4000 ;
	    RECT 151.6000 70.3000 152.4000 70.4000 ;
	    RECT 159.6000 70.3000 160.4000 70.4000 ;
	    RECT 146.8000 69.7000 152.4000 70.3000 ;
	    RECT 146.8000 69.6000 147.6000 69.7000 ;
	    RECT 151.6000 69.6000 152.4000 69.7000 ;
	    RECT 153.3000 69.7000 160.4000 70.3000 ;
	    RECT 100.4000 68.3000 101.2000 68.4000 ;
	    RECT 102.0000 68.3000 102.8000 68.4000 ;
	    RECT 100.4000 67.7000 102.8000 68.3000 ;
	    RECT 100.4000 67.6000 101.2000 67.7000 ;
	    RECT 102.0000 67.6000 102.8000 67.7000 ;
	    RECT 126.0000 68.3000 126.8000 68.4000 ;
	    RECT 135.6000 68.3000 136.4000 68.4000 ;
	    RECT 142.0000 68.3000 142.8000 68.4000 ;
	    RECT 126.0000 67.7000 142.8000 68.3000 ;
	    RECT 126.0000 67.6000 126.8000 67.7000 ;
	    RECT 135.6000 67.6000 136.4000 67.7000 ;
	    RECT 142.0000 67.6000 142.8000 67.7000 ;
	    RECT 148.4000 68.3000 149.2000 68.4000 ;
	    RECT 153.3000 68.3000 153.9000 69.7000 ;
	    RECT 159.6000 69.6000 160.4000 69.7000 ;
	    RECT 162.8000 70.3000 163.6000 70.4000 ;
	    RECT 178.8000 70.3000 179.6000 70.4000 ;
	    RECT 162.8000 69.7000 179.6000 70.3000 ;
	    RECT 162.8000 69.6000 163.6000 69.7000 ;
	    RECT 178.8000 69.6000 179.6000 69.7000 ;
	    RECT 198.0000 70.3000 198.8000 70.4000 ;
	    RECT 206.0000 70.3000 206.8000 70.4000 ;
	    RECT 198.0000 69.7000 206.8000 70.3000 ;
	    RECT 198.0000 69.6000 198.8000 69.7000 ;
	    RECT 206.0000 69.6000 206.8000 69.7000 ;
	    RECT 207.6000 70.3000 208.4000 70.4000 ;
	    RECT 209.2000 70.3000 210.0000 70.4000 ;
	    RECT 207.6000 69.7000 210.0000 70.3000 ;
	    RECT 207.6000 69.6000 208.4000 69.7000 ;
	    RECT 209.2000 69.6000 210.0000 69.7000 ;
	    RECT 212.4000 70.3000 213.2000 70.4000 ;
	    RECT 231.6000 70.3000 232.4000 70.4000 ;
	    RECT 212.4000 69.7000 232.4000 70.3000 ;
	    RECT 212.4000 69.6000 213.2000 69.7000 ;
	    RECT 231.6000 69.6000 232.4000 69.7000 ;
	    RECT 233.2000 70.3000 234.0000 70.4000 ;
	    RECT 238.0000 70.3000 238.8000 70.4000 ;
	    RECT 233.2000 69.7000 238.8000 70.3000 ;
	    RECT 233.2000 69.6000 234.0000 69.7000 ;
	    RECT 238.0000 69.6000 238.8000 69.7000 ;
	    RECT 244.4000 69.6000 245.2000 70.4000 ;
	    RECT 247.6000 70.3000 248.4000 70.4000 ;
	    RECT 250.8000 70.3000 251.6000 70.4000 ;
	    RECT 247.6000 69.7000 251.6000 70.3000 ;
	    RECT 252.5000 70.3000 253.1000 71.7000 ;
	    RECT 257.2000 71.7000 264.4000 72.3000 ;
	    RECT 257.2000 71.6000 258.0000 71.7000 ;
	    RECT 263.6000 71.6000 264.4000 71.7000 ;
	    RECT 268.4000 72.3000 269.2000 72.4000 ;
	    RECT 274.8000 72.3000 275.6000 72.4000 ;
	    RECT 268.4000 71.7000 275.6000 72.3000 ;
	    RECT 268.4000 71.6000 269.2000 71.7000 ;
	    RECT 274.8000 71.6000 275.6000 71.7000 ;
	    RECT 276.4000 72.3000 277.2000 72.4000 ;
	    RECT 292.4000 72.3000 293.2000 72.4000 ;
	    RECT 276.4000 71.7000 293.2000 72.3000 ;
	    RECT 276.4000 71.6000 277.2000 71.7000 ;
	    RECT 292.4000 71.6000 293.2000 71.7000 ;
	    RECT 294.0000 72.3000 294.8000 72.4000 ;
	    RECT 305.2000 72.3000 306.0000 72.4000 ;
	    RECT 294.0000 71.7000 306.0000 72.3000 ;
	    RECT 294.0000 71.6000 294.8000 71.7000 ;
	    RECT 305.2000 71.6000 306.0000 71.7000 ;
	    RECT 306.8000 72.3000 307.6000 72.4000 ;
	    RECT 314.8000 72.3000 315.6000 72.4000 ;
	    RECT 306.8000 71.7000 315.6000 72.3000 ;
	    RECT 306.8000 71.6000 307.6000 71.7000 ;
	    RECT 314.8000 71.6000 315.6000 71.7000 ;
	    RECT 316.4000 72.3000 317.2000 72.4000 ;
	    RECT 321.2000 72.3000 322.0000 72.4000 ;
	    RECT 335.6000 72.3000 336.4000 72.4000 ;
	    RECT 316.4000 71.7000 336.4000 72.3000 ;
	    RECT 316.4000 71.6000 317.2000 71.7000 ;
	    RECT 321.2000 71.6000 322.0000 71.7000 ;
	    RECT 335.6000 71.6000 336.4000 71.7000 ;
	    RECT 359.6000 72.3000 360.4000 72.4000 ;
	    RECT 362.8000 72.3000 363.6000 72.4000 ;
	    RECT 359.6000 71.7000 363.6000 72.3000 ;
	    RECT 359.6000 71.6000 360.4000 71.7000 ;
	    RECT 362.8000 71.6000 363.6000 71.7000 ;
	    RECT 377.2000 72.3000 378.0000 72.4000 ;
	    RECT 385.2000 72.3000 386.0000 72.4000 ;
	    RECT 377.2000 71.7000 386.0000 72.3000 ;
	    RECT 377.2000 71.6000 378.0000 71.7000 ;
	    RECT 385.2000 71.6000 386.0000 71.7000 ;
	    RECT 407.6000 72.3000 408.4000 72.4000 ;
	    RECT 425.2000 72.3000 426.0000 72.4000 ;
	    RECT 407.6000 71.7000 426.0000 72.3000 ;
	    RECT 407.6000 71.6000 408.4000 71.7000 ;
	    RECT 425.2000 71.6000 426.0000 71.7000 ;
	    RECT 454.0000 72.3000 454.8000 72.4000 ;
	    RECT 455.6000 72.3000 456.4000 72.4000 ;
	    RECT 454.0000 71.7000 456.4000 72.3000 ;
	    RECT 454.0000 71.6000 454.8000 71.7000 ;
	    RECT 455.6000 71.6000 456.4000 71.7000 ;
	    RECT 468.4000 72.3000 469.2000 72.4000 ;
	    RECT 479.6000 72.3000 480.4000 72.4000 ;
	    RECT 468.4000 71.7000 480.4000 72.3000 ;
	    RECT 468.4000 71.6000 469.2000 71.7000 ;
	    RECT 479.6000 71.6000 480.4000 71.7000 ;
	    RECT 487.6000 72.3000 488.4000 72.4000 ;
	    RECT 506.8000 72.3000 507.6000 72.4000 ;
	    RECT 487.6000 71.7000 507.6000 72.3000 ;
	    RECT 487.6000 71.6000 488.4000 71.7000 ;
	    RECT 506.8000 71.6000 507.6000 71.7000 ;
	    RECT 258.8000 70.3000 259.6000 70.4000 ;
	    RECT 252.5000 69.7000 259.6000 70.3000 ;
	    RECT 247.6000 69.6000 248.4000 69.7000 ;
	    RECT 250.8000 69.6000 251.6000 69.7000 ;
	    RECT 258.8000 69.6000 259.6000 69.7000 ;
	    RECT 262.0000 70.3000 262.8000 70.4000 ;
	    RECT 271.6000 70.3000 272.4000 70.4000 ;
	    RECT 322.8000 70.3000 323.6000 70.4000 ;
	    RECT 332.4000 70.3000 333.2000 70.4000 ;
	    RECT 262.0000 69.7000 272.4000 70.3000 ;
	    RECT 262.0000 69.6000 262.8000 69.7000 ;
	    RECT 271.6000 69.6000 272.4000 69.7000 ;
	    RECT 273.3000 69.7000 321.9000 70.3000 ;
	    RECT 148.4000 67.7000 153.9000 68.3000 ;
	    RECT 154.8000 68.3000 155.6000 68.4000 ;
	    RECT 166.0000 68.3000 166.8000 68.4000 ;
	    RECT 154.8000 67.7000 166.8000 68.3000 ;
	    RECT 148.4000 67.6000 149.2000 67.7000 ;
	    RECT 154.8000 67.6000 155.6000 67.7000 ;
	    RECT 166.0000 67.6000 166.8000 67.7000 ;
	    RECT 167.6000 68.3000 168.4000 68.4000 ;
	    RECT 175.6000 68.3000 176.4000 68.4000 ;
	    RECT 167.6000 67.7000 176.4000 68.3000 ;
	    RECT 167.6000 67.6000 168.4000 67.7000 ;
	    RECT 175.6000 67.6000 176.4000 67.7000 ;
	    RECT 217.2000 68.3000 218.0000 68.4000 ;
	    RECT 218.8000 68.3000 219.6000 68.4000 ;
	    RECT 217.2000 67.7000 219.6000 68.3000 ;
	    RECT 217.2000 67.6000 218.0000 67.7000 ;
	    RECT 218.8000 67.6000 219.6000 67.7000 ;
	    RECT 226.8000 68.3000 227.6000 68.4000 ;
	    RECT 238.0000 68.3000 238.8000 68.4000 ;
	    RECT 226.8000 67.7000 238.8000 68.3000 ;
	    RECT 226.8000 67.6000 227.6000 67.7000 ;
	    RECT 238.0000 67.6000 238.8000 67.7000 ;
	    RECT 241.2000 68.3000 242.0000 68.4000 ;
	    RECT 249.2000 68.3000 250.0000 68.4000 ;
	    RECT 241.2000 67.7000 250.0000 68.3000 ;
	    RECT 241.2000 67.6000 242.0000 67.7000 ;
	    RECT 249.2000 67.6000 250.0000 67.7000 ;
	    RECT 263.6000 68.3000 264.4000 68.4000 ;
	    RECT 266.8000 68.3000 267.6000 68.4000 ;
	    RECT 263.6000 67.7000 267.6000 68.3000 ;
	    RECT 263.6000 67.6000 264.4000 67.7000 ;
	    RECT 266.8000 67.6000 267.6000 67.7000 ;
	    RECT 270.0000 67.6000 270.8000 68.4000 ;
	    RECT 271.6000 68.3000 272.4000 68.4000 ;
	    RECT 273.3000 68.3000 273.9000 69.7000 ;
	    RECT 321.3000 68.4000 321.9000 69.7000 ;
	    RECT 322.8000 69.7000 333.2000 70.3000 ;
	    RECT 322.8000 69.6000 323.6000 69.7000 ;
	    RECT 332.4000 69.6000 333.2000 69.7000 ;
	    RECT 354.8000 70.3000 355.6000 70.4000 ;
	    RECT 393.2000 70.3000 394.0000 70.4000 ;
	    RECT 394.8000 70.3000 395.6000 70.4000 ;
	    RECT 354.8000 69.7000 395.6000 70.3000 ;
	    RECT 354.8000 69.6000 355.6000 69.7000 ;
	    RECT 393.2000 69.6000 394.0000 69.7000 ;
	    RECT 394.8000 69.6000 395.6000 69.7000 ;
	    RECT 423.6000 70.3000 424.4000 70.4000 ;
	    RECT 428.4000 70.3000 429.2000 70.4000 ;
	    RECT 430.0000 70.3000 430.8000 70.4000 ;
	    RECT 423.6000 69.7000 430.8000 70.3000 ;
	    RECT 423.6000 69.6000 424.4000 69.7000 ;
	    RECT 428.4000 69.6000 429.2000 69.7000 ;
	    RECT 430.0000 69.6000 430.8000 69.7000 ;
	    RECT 271.6000 67.7000 273.9000 68.3000 ;
	    RECT 278.0000 68.3000 278.8000 68.4000 ;
	    RECT 287.6000 68.3000 288.4000 68.4000 ;
	    RECT 303.6000 68.3000 304.4000 68.4000 ;
	    RECT 278.0000 67.7000 304.4000 68.3000 ;
	    RECT 271.6000 67.6000 272.4000 67.7000 ;
	    RECT 278.0000 67.6000 278.8000 67.7000 ;
	    RECT 287.6000 67.6000 288.4000 67.7000 ;
	    RECT 303.6000 67.6000 304.4000 67.7000 ;
	    RECT 311.6000 68.3000 312.4000 68.4000 ;
	    RECT 316.4000 68.3000 317.2000 68.4000 ;
	    RECT 311.6000 67.7000 317.2000 68.3000 ;
	    RECT 311.6000 67.6000 312.4000 67.7000 ;
	    RECT 316.4000 67.6000 317.2000 67.7000 ;
	    RECT 321.2000 68.3000 322.0000 68.4000 ;
	    RECT 324.4000 68.3000 325.2000 68.4000 ;
	    RECT 321.2000 67.7000 325.2000 68.3000 ;
	    RECT 321.2000 67.6000 322.0000 67.7000 ;
	    RECT 324.4000 67.6000 325.2000 67.7000 ;
	    RECT 326.0000 68.3000 326.8000 68.4000 ;
	    RECT 330.8000 68.3000 331.6000 68.4000 ;
	    RECT 326.0000 67.7000 331.6000 68.3000 ;
	    RECT 326.0000 67.6000 326.8000 67.7000 ;
	    RECT 330.8000 67.6000 331.6000 67.7000 ;
	    RECT 332.4000 68.3000 333.2000 68.4000 ;
	    RECT 343.6000 68.3000 344.4000 68.4000 ;
	    RECT 332.4000 67.7000 344.4000 68.3000 ;
	    RECT 332.4000 67.6000 333.2000 67.7000 ;
	    RECT 343.6000 67.6000 344.4000 67.7000 ;
	    RECT 362.8000 68.3000 363.6000 68.4000 ;
	    RECT 383.6000 68.3000 384.4000 68.4000 ;
	    RECT 362.8000 67.7000 384.4000 68.3000 ;
	    RECT 362.8000 67.6000 363.6000 67.7000 ;
	    RECT 383.6000 67.6000 384.4000 67.7000 ;
	    RECT 388.4000 68.3000 389.2000 68.4000 ;
	    RECT 398.0000 68.3000 398.8000 68.4000 ;
	    RECT 388.4000 67.7000 398.8000 68.3000 ;
	    RECT 388.4000 67.6000 389.2000 67.7000 ;
	    RECT 398.0000 67.6000 398.8000 67.7000 ;
	    RECT 450.8000 68.3000 451.6000 68.4000 ;
	    RECT 495.6000 68.3000 496.4000 68.4000 ;
	    RECT 450.8000 67.7000 496.4000 68.3000 ;
	    RECT 450.8000 67.6000 451.6000 67.7000 ;
	    RECT 495.6000 67.6000 496.4000 67.7000 ;
	    RECT 38.0000 66.3000 38.8000 66.4000 ;
	    RECT 42.8000 66.3000 43.6000 66.4000 ;
	    RECT 54.0000 66.3000 54.8000 66.4000 ;
	    RECT 74.8000 66.3000 75.6000 66.4000 ;
	    RECT 38.0000 65.7000 75.6000 66.3000 ;
	    RECT 38.0000 65.6000 38.8000 65.7000 ;
	    RECT 42.8000 65.6000 43.6000 65.7000 ;
	    RECT 54.0000 65.6000 54.8000 65.7000 ;
	    RECT 74.8000 65.6000 75.6000 65.7000 ;
	    RECT 81.2000 66.3000 82.0000 66.4000 ;
	    RECT 84.4000 66.3000 85.2000 66.4000 ;
	    RECT 81.2000 65.7000 85.2000 66.3000 ;
	    RECT 81.2000 65.6000 82.0000 65.7000 ;
	    RECT 84.4000 65.6000 85.2000 65.7000 ;
	    RECT 132.4000 66.3000 133.2000 66.4000 ;
	    RECT 170.8000 66.3000 171.6000 66.4000 ;
	    RECT 183.6000 66.3000 184.4000 66.4000 ;
	    RECT 132.4000 65.7000 184.4000 66.3000 ;
	    RECT 132.4000 65.6000 133.2000 65.7000 ;
	    RECT 170.8000 65.6000 171.6000 65.7000 ;
	    RECT 183.6000 65.6000 184.4000 65.7000 ;
	    RECT 188.4000 66.3000 189.2000 66.4000 ;
	    RECT 217.2000 66.3000 218.0000 66.4000 ;
	    RECT 268.4000 66.3000 269.2000 66.4000 ;
	    RECT 188.4000 65.7000 218.0000 66.3000 ;
	    RECT 188.4000 65.6000 189.2000 65.7000 ;
	    RECT 217.2000 65.6000 218.0000 65.7000 ;
	    RECT 218.9000 65.7000 269.2000 66.3000 ;
	    RECT 9.2000 64.3000 10.0000 64.4000 ;
	    RECT 44.4000 64.3000 45.2000 64.4000 ;
	    RECT 9.2000 63.7000 45.2000 64.3000 ;
	    RECT 9.2000 63.6000 10.0000 63.7000 ;
	    RECT 44.4000 63.6000 45.2000 63.7000 ;
	    RECT 58.8000 64.3000 59.6000 64.4000 ;
	    RECT 154.8000 64.3000 155.6000 64.4000 ;
	    RECT 58.8000 63.7000 155.6000 64.3000 ;
	    RECT 58.8000 63.6000 59.6000 63.7000 ;
	    RECT 154.8000 63.6000 155.6000 63.7000 ;
	    RECT 158.0000 64.3000 158.8000 64.4000 ;
	    RECT 159.6000 64.3000 160.4000 64.4000 ;
	    RECT 158.0000 63.7000 160.4000 64.3000 ;
	    RECT 158.0000 63.6000 158.8000 63.7000 ;
	    RECT 159.6000 63.6000 160.4000 63.7000 ;
	    RECT 166.0000 64.3000 166.8000 64.4000 ;
	    RECT 177.2000 64.3000 178.0000 64.4000 ;
	    RECT 166.0000 63.7000 178.0000 64.3000 ;
	    RECT 166.0000 63.6000 166.8000 63.7000 ;
	    RECT 177.2000 63.6000 178.0000 63.7000 ;
	    RECT 178.8000 64.3000 179.6000 64.4000 ;
	    RECT 196.4000 64.3000 197.2000 64.4000 ;
	    RECT 178.8000 63.7000 197.2000 64.3000 ;
	    RECT 178.8000 63.6000 179.6000 63.7000 ;
	    RECT 196.4000 63.6000 197.2000 63.7000 ;
	    RECT 202.8000 64.3000 203.6000 64.4000 ;
	    RECT 218.9000 64.3000 219.5000 65.7000 ;
	    RECT 268.4000 65.6000 269.2000 65.7000 ;
	    RECT 274.8000 66.3000 275.6000 66.4000 ;
	    RECT 278.0000 66.3000 278.8000 66.4000 ;
	    RECT 274.8000 65.7000 278.8000 66.3000 ;
	    RECT 274.8000 65.6000 275.6000 65.7000 ;
	    RECT 278.0000 65.6000 278.8000 65.7000 ;
	    RECT 284.4000 66.3000 285.2000 66.4000 ;
	    RECT 295.6000 66.3000 296.4000 66.4000 ;
	    RECT 284.4000 65.7000 296.4000 66.3000 ;
	    RECT 284.4000 65.6000 285.2000 65.7000 ;
	    RECT 295.6000 65.6000 296.4000 65.7000 ;
	    RECT 311.6000 66.3000 312.4000 66.4000 ;
	    RECT 359.6000 66.3000 360.4000 66.4000 ;
	    RECT 364.4000 66.3000 365.2000 66.4000 ;
	    RECT 311.6000 65.7000 365.2000 66.3000 ;
	    RECT 311.6000 65.6000 312.4000 65.7000 ;
	    RECT 359.6000 65.6000 360.4000 65.7000 ;
	    RECT 364.4000 65.6000 365.2000 65.7000 ;
	    RECT 202.8000 63.7000 219.5000 64.3000 ;
	    RECT 236.4000 64.3000 237.2000 64.4000 ;
	    RECT 281.2000 64.3000 282.0000 64.4000 ;
	    RECT 446.0000 64.3000 446.8000 64.4000 ;
	    RECT 236.4000 63.7000 277.1000 64.3000 ;
	    RECT 202.8000 63.6000 203.6000 63.7000 ;
	    RECT 236.4000 63.6000 237.2000 63.7000 ;
	    RECT 276.5000 62.4000 277.1000 63.7000 ;
	    RECT 281.2000 63.7000 446.8000 64.3000 ;
	    RECT 281.2000 63.6000 282.0000 63.7000 ;
	    RECT 446.0000 63.6000 446.8000 63.7000 ;
	    RECT 14.0000 62.3000 14.8000 62.4000 ;
	    RECT 76.4000 62.3000 77.2000 62.4000 ;
	    RECT 134.0000 62.3000 134.8000 62.4000 ;
	    RECT 14.0000 61.7000 134.8000 62.3000 ;
	    RECT 14.0000 61.6000 14.8000 61.7000 ;
	    RECT 76.4000 61.6000 77.2000 61.7000 ;
	    RECT 134.0000 61.6000 134.8000 61.7000 ;
	    RECT 158.0000 62.3000 158.8000 62.4000 ;
	    RECT 177.2000 62.3000 178.0000 62.4000 ;
	    RECT 199.6000 62.3000 200.4000 62.4000 ;
	    RECT 207.6000 62.3000 208.4000 62.4000 ;
	    RECT 158.0000 61.7000 208.4000 62.3000 ;
	    RECT 158.0000 61.6000 158.8000 61.7000 ;
	    RECT 177.2000 61.6000 178.0000 61.7000 ;
	    RECT 199.6000 61.6000 200.4000 61.7000 ;
	    RECT 207.6000 61.6000 208.4000 61.7000 ;
	    RECT 209.2000 61.6000 210.0000 62.4000 ;
	    RECT 210.8000 62.3000 211.6000 62.4000 ;
	    RECT 234.8000 62.3000 235.6000 62.4000 ;
	    RECT 210.8000 61.7000 235.6000 62.3000 ;
	    RECT 210.8000 61.6000 211.6000 61.7000 ;
	    RECT 234.8000 61.6000 235.6000 61.7000 ;
	    RECT 276.4000 62.3000 277.2000 62.4000 ;
	    RECT 289.2000 62.3000 290.0000 62.4000 ;
	    RECT 276.4000 61.7000 290.0000 62.3000 ;
	    RECT 276.4000 61.6000 277.2000 61.7000 ;
	    RECT 289.2000 61.6000 290.0000 61.7000 ;
	    RECT 300.4000 62.3000 301.2000 62.4000 ;
	    RECT 337.2000 62.3000 338.0000 62.4000 ;
	    RECT 300.4000 61.7000 338.0000 62.3000 ;
	    RECT 300.4000 61.6000 301.2000 61.7000 ;
	    RECT 337.2000 61.6000 338.0000 61.7000 ;
	    RECT 338.8000 62.3000 339.6000 62.4000 ;
	    RECT 370.8000 62.3000 371.6000 62.4000 ;
	    RECT 338.8000 61.7000 371.6000 62.3000 ;
	    RECT 338.8000 61.6000 339.6000 61.7000 ;
	    RECT 370.8000 61.6000 371.6000 61.7000 ;
	    RECT 430.0000 62.3000 430.8000 62.4000 ;
	    RECT 462.0000 62.3000 462.8000 62.4000 ;
	    RECT 463.6000 62.3000 464.4000 62.4000 ;
	    RECT 430.0000 61.7000 464.4000 62.3000 ;
	    RECT 430.0000 61.6000 430.8000 61.7000 ;
	    RECT 462.0000 61.6000 462.8000 61.7000 ;
	    RECT 463.6000 61.6000 464.4000 61.7000 ;
	    RECT 116.4000 60.3000 117.2000 60.4000 ;
	    RECT 167.6000 60.3000 168.4000 60.4000 ;
	    RECT 116.4000 59.7000 168.4000 60.3000 ;
	    RECT 116.4000 59.6000 117.2000 59.7000 ;
	    RECT 167.6000 59.6000 168.4000 59.7000 ;
	    RECT 174.0000 60.3000 174.8000 60.4000 ;
	    RECT 220.4000 60.3000 221.2000 60.4000 ;
	    RECT 174.0000 59.7000 221.2000 60.3000 ;
	    RECT 174.0000 59.6000 174.8000 59.7000 ;
	    RECT 220.4000 59.6000 221.2000 59.7000 ;
	    RECT 265.2000 60.3000 266.0000 60.4000 ;
	    RECT 281.2000 60.3000 282.0000 60.4000 ;
	    RECT 265.2000 59.7000 282.0000 60.3000 ;
	    RECT 265.2000 59.6000 266.0000 59.7000 ;
	    RECT 281.2000 59.6000 282.0000 59.7000 ;
	    RECT 295.6000 60.3000 296.4000 60.4000 ;
	    RECT 306.8000 60.3000 307.6000 60.4000 ;
	    RECT 295.6000 59.7000 307.6000 60.3000 ;
	    RECT 295.6000 59.6000 296.4000 59.7000 ;
	    RECT 306.8000 59.6000 307.6000 59.7000 ;
	    RECT 308.4000 60.3000 309.2000 60.4000 ;
	    RECT 332.4000 60.3000 333.2000 60.4000 ;
	    RECT 390.0000 60.3000 390.8000 60.4000 ;
	    RECT 394.8000 60.3000 395.6000 60.4000 ;
	    RECT 308.4000 59.7000 389.1000 60.3000 ;
	    RECT 308.4000 59.6000 309.2000 59.7000 ;
	    RECT 332.4000 59.6000 333.2000 59.7000 ;
	    RECT 55.6000 58.3000 56.4000 58.4000 ;
	    RECT 89.2000 58.3000 90.0000 58.4000 ;
	    RECT 55.6000 57.7000 90.0000 58.3000 ;
	    RECT 55.6000 57.6000 56.4000 57.7000 ;
	    RECT 89.2000 57.6000 90.0000 57.7000 ;
	    RECT 100.4000 58.3000 101.2000 58.4000 ;
	    RECT 119.6000 58.3000 120.4000 58.4000 ;
	    RECT 100.4000 57.7000 120.4000 58.3000 ;
	    RECT 100.4000 57.6000 101.2000 57.7000 ;
	    RECT 119.6000 57.6000 120.4000 57.7000 ;
	    RECT 122.8000 58.3000 123.6000 58.4000 ;
	    RECT 159.6000 58.3000 160.4000 58.4000 ;
	    RECT 172.4000 58.3000 173.2000 58.4000 ;
	    RECT 204.4000 58.3000 205.2000 58.4000 ;
	    RECT 217.2000 58.3000 218.0000 58.4000 ;
	    RECT 223.6000 58.3000 224.4000 58.4000 ;
	    RECT 122.8000 57.7000 224.4000 58.3000 ;
	    RECT 122.8000 57.6000 123.6000 57.7000 ;
	    RECT 159.6000 57.6000 160.4000 57.7000 ;
	    RECT 172.4000 57.6000 173.2000 57.7000 ;
	    RECT 204.4000 57.6000 205.2000 57.7000 ;
	    RECT 217.2000 57.6000 218.0000 57.7000 ;
	    RECT 223.6000 57.6000 224.4000 57.7000 ;
	    RECT 230.0000 58.3000 230.8000 58.4000 ;
	    RECT 239.6000 58.3000 240.4000 58.4000 ;
	    RECT 241.2000 58.3000 242.0000 58.4000 ;
	    RECT 230.0000 57.7000 242.0000 58.3000 ;
	    RECT 230.0000 57.6000 230.8000 57.7000 ;
	    RECT 239.6000 57.6000 240.4000 57.7000 ;
	    RECT 241.2000 57.6000 242.0000 57.7000 ;
	    RECT 247.6000 57.6000 248.4000 58.4000 ;
	    RECT 262.0000 58.3000 262.8000 58.4000 ;
	    RECT 258.9000 57.7000 262.8000 58.3000 ;
	    RECT 33.2000 56.3000 34.0000 56.4000 ;
	    RECT 52.4000 56.3000 53.2000 56.4000 ;
	    RECT 33.2000 55.7000 53.2000 56.3000 ;
	    RECT 33.2000 55.6000 34.0000 55.7000 ;
	    RECT 52.4000 55.6000 53.2000 55.7000 ;
	    RECT 73.2000 56.3000 74.0000 56.4000 ;
	    RECT 84.4000 56.3000 85.2000 56.4000 ;
	    RECT 89.2000 56.3000 90.0000 56.4000 ;
	    RECT 73.2000 55.7000 90.0000 56.3000 ;
	    RECT 73.2000 55.6000 74.0000 55.7000 ;
	    RECT 84.4000 55.6000 85.2000 55.7000 ;
	    RECT 89.2000 55.6000 90.0000 55.7000 ;
	    RECT 90.8000 56.3000 91.6000 56.4000 ;
	    RECT 174.0000 56.3000 174.8000 56.4000 ;
	    RECT 90.8000 55.7000 174.8000 56.3000 ;
	    RECT 90.8000 55.6000 91.6000 55.7000 ;
	    RECT 174.0000 55.6000 174.8000 55.7000 ;
	    RECT 185.2000 56.3000 186.0000 56.4000 ;
	    RECT 190.0000 56.3000 190.8000 56.4000 ;
	    RECT 193.2000 56.3000 194.0000 56.4000 ;
	    RECT 185.2000 55.7000 194.0000 56.3000 ;
	    RECT 185.2000 55.6000 186.0000 55.7000 ;
	    RECT 190.0000 55.6000 190.8000 55.7000 ;
	    RECT 193.2000 55.6000 194.0000 55.7000 ;
	    RECT 196.4000 56.3000 197.2000 56.4000 ;
	    RECT 198.0000 56.3000 198.8000 56.4000 ;
	    RECT 212.4000 56.3000 213.2000 56.4000 ;
	    RECT 196.4000 55.7000 198.8000 56.3000 ;
	    RECT 196.4000 55.6000 197.2000 55.7000 ;
	    RECT 198.0000 55.6000 198.8000 55.7000 ;
	    RECT 199.7000 55.7000 213.2000 56.3000 ;
	    RECT 50.8000 54.3000 51.6000 54.4000 ;
	    RECT 52.4000 54.3000 53.2000 54.4000 ;
	    RECT 50.8000 53.7000 53.2000 54.3000 ;
	    RECT 50.8000 53.6000 51.6000 53.7000 ;
	    RECT 52.4000 53.6000 53.2000 53.7000 ;
	    RECT 57.2000 54.3000 58.0000 54.4000 ;
	    RECT 62.0000 54.3000 62.8000 54.4000 ;
	    RECT 57.2000 53.7000 62.8000 54.3000 ;
	    RECT 57.2000 53.6000 58.0000 53.7000 ;
	    RECT 62.0000 53.6000 62.8000 53.7000 ;
	    RECT 65.2000 54.3000 66.0000 54.4000 ;
	    RECT 87.6000 54.3000 88.4000 54.4000 ;
	    RECT 105.2000 54.3000 106.0000 54.4000 ;
	    RECT 154.8000 54.3000 155.6000 54.4000 ;
	    RECT 65.2000 53.7000 155.6000 54.3000 ;
	    RECT 65.2000 53.6000 66.0000 53.7000 ;
	    RECT 87.6000 53.6000 88.4000 53.7000 ;
	    RECT 105.2000 53.6000 106.0000 53.7000 ;
	    RECT 154.8000 53.6000 155.6000 53.7000 ;
	    RECT 162.8000 54.3000 163.6000 54.4000 ;
	    RECT 186.8000 54.3000 187.6000 54.4000 ;
	    RECT 162.8000 53.7000 187.6000 54.3000 ;
	    RECT 162.8000 53.6000 163.6000 53.7000 ;
	    RECT 186.8000 53.6000 187.6000 53.7000 ;
	    RECT 196.4000 54.3000 197.2000 54.4000 ;
	    RECT 199.7000 54.3000 200.3000 55.7000 ;
	    RECT 212.4000 55.6000 213.2000 55.7000 ;
	    RECT 222.0000 56.3000 222.8000 56.4000 ;
	    RECT 226.8000 56.3000 227.6000 56.4000 ;
	    RECT 222.0000 55.7000 227.6000 56.3000 ;
	    RECT 222.0000 55.6000 222.8000 55.7000 ;
	    RECT 226.8000 55.6000 227.6000 55.7000 ;
	    RECT 231.6000 56.3000 232.4000 56.4000 ;
	    RECT 258.9000 56.3000 259.5000 57.7000 ;
	    RECT 262.0000 57.6000 262.8000 57.7000 ;
	    RECT 273.2000 58.3000 274.0000 58.4000 ;
	    RECT 282.8000 58.3000 283.6000 58.4000 ;
	    RECT 302.0000 58.3000 302.8000 58.4000 ;
	    RECT 273.2000 57.7000 302.8000 58.3000 ;
	    RECT 273.2000 57.6000 274.0000 57.7000 ;
	    RECT 282.8000 57.6000 283.6000 57.7000 ;
	    RECT 302.0000 57.6000 302.8000 57.7000 ;
	    RECT 321.2000 58.3000 322.0000 58.4000 ;
	    RECT 334.0000 58.3000 334.8000 58.4000 ;
	    RECT 321.2000 57.7000 334.8000 58.3000 ;
	    RECT 321.2000 57.6000 322.0000 57.7000 ;
	    RECT 334.0000 57.6000 334.8000 57.7000 ;
	    RECT 335.6000 58.3000 336.4000 58.4000 ;
	    RECT 350.0000 58.3000 350.8000 58.4000 ;
	    RECT 388.5000 58.3000 389.1000 59.7000 ;
	    RECT 390.0000 59.7000 395.6000 60.3000 ;
	    RECT 390.0000 59.6000 390.8000 59.7000 ;
	    RECT 394.8000 59.6000 395.6000 59.7000 ;
	    RECT 410.8000 60.3000 411.6000 60.4000 ;
	    RECT 425.2000 60.3000 426.0000 60.4000 ;
	    RECT 433.2000 60.3000 434.0000 60.4000 ;
	    RECT 490.8000 60.3000 491.6000 60.4000 ;
	    RECT 410.8000 59.7000 434.0000 60.3000 ;
	    RECT 410.8000 59.6000 411.6000 59.7000 ;
	    RECT 425.2000 59.6000 426.0000 59.7000 ;
	    RECT 433.2000 59.6000 434.0000 59.7000 ;
	    RECT 434.9000 59.7000 491.6000 60.3000 ;
	    RECT 434.9000 58.3000 435.5000 59.7000 ;
	    RECT 490.8000 59.6000 491.6000 59.7000 ;
	    RECT 335.6000 57.7000 381.1000 58.3000 ;
	    RECT 388.5000 57.7000 435.5000 58.3000 ;
	    RECT 438.0000 58.3000 438.8000 58.4000 ;
	    RECT 482.8000 58.3000 483.6000 58.4000 ;
	    RECT 438.0000 57.7000 483.6000 58.3000 ;
	    RECT 335.6000 57.6000 336.4000 57.7000 ;
	    RECT 350.0000 57.6000 350.8000 57.7000 ;
	    RECT 231.6000 55.7000 259.5000 56.3000 ;
	    RECT 260.4000 56.3000 261.2000 56.4000 ;
	    RECT 263.6000 56.3000 264.4000 56.4000 ;
	    RECT 260.4000 55.7000 264.4000 56.3000 ;
	    RECT 231.6000 55.6000 232.4000 55.7000 ;
	    RECT 260.4000 55.6000 261.2000 55.7000 ;
	    RECT 263.6000 55.6000 264.4000 55.7000 ;
	    RECT 266.8000 56.3000 267.6000 56.4000 ;
	    RECT 290.8000 56.3000 291.6000 56.4000 ;
	    RECT 266.8000 55.7000 291.6000 56.3000 ;
	    RECT 266.8000 55.6000 267.6000 55.7000 ;
	    RECT 290.8000 55.6000 291.6000 55.7000 ;
	    RECT 295.6000 56.3000 296.4000 56.4000 ;
	    RECT 303.6000 56.3000 304.4000 56.4000 ;
	    RECT 295.6000 55.7000 304.4000 56.3000 ;
	    RECT 295.6000 55.6000 296.4000 55.7000 ;
	    RECT 303.6000 55.6000 304.4000 55.7000 ;
	    RECT 305.2000 56.3000 306.0000 56.4000 ;
	    RECT 314.8000 56.3000 315.6000 56.4000 ;
	    RECT 305.2000 55.7000 315.6000 56.3000 ;
	    RECT 305.2000 55.6000 306.0000 55.7000 ;
	    RECT 314.8000 55.6000 315.6000 55.7000 ;
	    RECT 318.0000 56.3000 318.8000 56.4000 ;
	    RECT 326.0000 56.3000 326.8000 56.4000 ;
	    RECT 318.0000 55.7000 326.8000 56.3000 ;
	    RECT 318.0000 55.6000 318.8000 55.7000 ;
	    RECT 326.0000 55.6000 326.8000 55.7000 ;
	    RECT 327.6000 56.3000 328.4000 56.4000 ;
	    RECT 343.6000 56.3000 344.4000 56.4000 ;
	    RECT 351.6000 56.3000 352.4000 56.4000 ;
	    RECT 327.6000 55.7000 352.4000 56.3000 ;
	    RECT 380.5000 56.3000 381.1000 57.7000 ;
	    RECT 438.0000 57.6000 438.8000 57.7000 ;
	    RECT 482.8000 57.6000 483.6000 57.7000 ;
	    RECT 409.2000 56.3000 410.0000 56.4000 ;
	    RECT 380.5000 55.7000 410.0000 56.3000 ;
	    RECT 327.6000 55.6000 328.4000 55.7000 ;
	    RECT 343.6000 55.6000 344.4000 55.7000 ;
	    RECT 351.6000 55.6000 352.4000 55.7000 ;
	    RECT 409.2000 55.6000 410.0000 55.7000 ;
	    RECT 422.0000 56.3000 422.8000 56.4000 ;
	    RECT 433.2000 56.3000 434.0000 56.4000 ;
	    RECT 422.0000 55.7000 434.0000 56.3000 ;
	    RECT 422.0000 55.6000 422.8000 55.7000 ;
	    RECT 433.2000 55.6000 434.0000 55.7000 ;
	    RECT 436.4000 56.3000 437.2000 56.4000 ;
	    RECT 473.2000 56.3000 474.0000 56.4000 ;
	    RECT 436.4000 55.7000 474.0000 56.3000 ;
	    RECT 436.4000 55.6000 437.2000 55.7000 ;
	    RECT 473.2000 55.6000 474.0000 55.7000 ;
	    RECT 196.4000 53.7000 200.3000 54.3000 ;
	    RECT 252.4000 54.3000 253.2000 54.4000 ;
	    RECT 282.8000 54.3000 283.6000 54.4000 ;
	    RECT 294.0000 54.3000 294.8000 54.4000 ;
	    RECT 252.4000 53.7000 294.8000 54.3000 ;
	    RECT 196.4000 53.6000 197.2000 53.7000 ;
	    RECT 252.4000 53.6000 253.2000 53.7000 ;
	    RECT 282.8000 53.6000 283.6000 53.7000 ;
	    RECT 294.0000 53.6000 294.8000 53.7000 ;
	    RECT 302.0000 54.3000 302.8000 54.4000 ;
	    RECT 334.0000 54.3000 334.8000 54.4000 ;
	    RECT 302.0000 53.7000 334.8000 54.3000 ;
	    RECT 302.0000 53.6000 302.8000 53.7000 ;
	    RECT 334.0000 53.6000 334.8000 53.7000 ;
	    RECT 337.2000 54.3000 338.0000 54.4000 ;
	    RECT 342.0000 54.3000 342.8000 54.4000 ;
	    RECT 337.2000 53.7000 342.8000 54.3000 ;
	    RECT 337.2000 53.6000 338.0000 53.7000 ;
	    RECT 342.0000 53.6000 342.8000 53.7000 ;
	    RECT 359.6000 54.3000 360.4000 54.4000 ;
	    RECT 375.6000 54.3000 376.4000 54.4000 ;
	    RECT 359.6000 53.7000 376.4000 54.3000 ;
	    RECT 359.6000 53.6000 360.4000 53.7000 ;
	    RECT 375.6000 53.6000 376.4000 53.7000 ;
	    RECT 390.0000 54.3000 390.8000 54.4000 ;
	    RECT 438.0000 54.3000 438.8000 54.4000 ;
	    RECT 390.0000 53.7000 438.8000 54.3000 ;
	    RECT 390.0000 53.6000 390.8000 53.7000 ;
	    RECT 438.0000 53.6000 438.8000 53.7000 ;
	    RECT 28.4000 52.3000 29.2000 52.4000 ;
	    RECT 46.0000 52.3000 46.8000 52.4000 ;
	    RECT 28.4000 51.7000 46.8000 52.3000 ;
	    RECT 28.4000 51.6000 29.2000 51.7000 ;
	    RECT 46.0000 51.6000 46.8000 51.7000 ;
	    RECT 50.8000 52.3000 51.6000 52.4000 ;
	    RECT 68.4000 52.3000 69.2000 52.4000 ;
	    RECT 126.0000 52.3000 126.8000 52.4000 ;
	    RECT 142.0000 52.3000 142.8000 52.4000 ;
	    RECT 50.8000 51.7000 54.7000 52.3000 ;
	    RECT 50.8000 51.6000 51.6000 51.7000 ;
	    RECT 42.8000 50.3000 43.6000 50.4000 ;
	    RECT 52.4000 50.3000 53.2000 50.4000 ;
	    RECT 42.8000 49.7000 53.2000 50.3000 ;
	    RECT 54.1000 50.3000 54.7000 51.7000 ;
	    RECT 68.4000 51.7000 142.8000 52.3000 ;
	    RECT 68.4000 51.6000 69.2000 51.7000 ;
	    RECT 126.0000 51.6000 126.8000 51.7000 ;
	    RECT 142.0000 51.6000 142.8000 51.7000 ;
	    RECT 151.6000 52.3000 152.4000 52.4000 ;
	    RECT 161.2000 52.3000 162.0000 52.4000 ;
	    RECT 151.6000 51.7000 162.0000 52.3000 ;
	    RECT 151.6000 51.6000 152.4000 51.7000 ;
	    RECT 161.2000 51.6000 162.0000 51.7000 ;
	    RECT 170.8000 52.3000 171.6000 52.4000 ;
	    RECT 188.4000 52.3000 189.2000 52.4000 ;
	    RECT 170.8000 51.7000 189.2000 52.3000 ;
	    RECT 170.8000 51.6000 171.6000 51.7000 ;
	    RECT 188.4000 51.6000 189.2000 51.7000 ;
	    RECT 191.6000 52.3000 192.4000 52.4000 ;
	    RECT 206.0000 52.3000 206.8000 52.4000 ;
	    RECT 191.6000 51.7000 206.8000 52.3000 ;
	    RECT 191.6000 51.6000 192.4000 51.7000 ;
	    RECT 206.0000 51.6000 206.8000 51.7000 ;
	    RECT 210.8000 52.3000 211.6000 52.4000 ;
	    RECT 218.8000 52.3000 219.6000 52.4000 ;
	    RECT 210.8000 51.7000 219.6000 52.3000 ;
	    RECT 210.8000 51.6000 211.6000 51.7000 ;
	    RECT 218.8000 51.6000 219.6000 51.7000 ;
	    RECT 226.8000 52.3000 227.6000 52.4000 ;
	    RECT 231.6000 52.3000 232.4000 52.4000 ;
	    RECT 226.8000 51.7000 232.4000 52.3000 ;
	    RECT 226.8000 51.6000 227.6000 51.7000 ;
	    RECT 231.6000 51.6000 232.4000 51.7000 ;
	    RECT 233.2000 52.3000 234.0000 52.4000 ;
	    RECT 239.6000 52.3000 240.4000 52.4000 ;
	    RECT 233.2000 51.7000 240.4000 52.3000 ;
	    RECT 233.2000 51.6000 234.0000 51.7000 ;
	    RECT 239.6000 51.6000 240.4000 51.7000 ;
	    RECT 250.8000 52.3000 251.6000 52.4000 ;
	    RECT 276.4000 52.3000 277.2000 52.4000 ;
	    RECT 310.0000 52.3000 310.8000 52.4000 ;
	    RECT 318.0000 52.3000 318.8000 52.4000 ;
	    RECT 351.6000 52.3000 352.4000 52.4000 ;
	    RECT 250.8000 51.7000 352.4000 52.3000 ;
	    RECT 250.8000 51.6000 251.6000 51.7000 ;
	    RECT 276.4000 51.6000 277.2000 51.7000 ;
	    RECT 310.0000 51.6000 310.8000 51.7000 ;
	    RECT 318.0000 51.6000 318.8000 51.7000 ;
	    RECT 351.6000 51.6000 352.4000 51.7000 ;
	    RECT 361.2000 52.3000 362.0000 52.4000 ;
	    RECT 369.2000 52.3000 370.0000 52.4000 ;
	    RECT 361.2000 51.7000 370.0000 52.3000 ;
	    RECT 361.2000 51.6000 362.0000 51.7000 ;
	    RECT 369.2000 51.6000 370.0000 51.7000 ;
	    RECT 378.8000 52.3000 379.6000 52.4000 ;
	    RECT 385.2000 52.3000 386.0000 52.4000 ;
	    RECT 378.8000 51.7000 386.0000 52.3000 ;
	    RECT 378.8000 51.6000 379.6000 51.7000 ;
	    RECT 385.2000 51.6000 386.0000 51.7000 ;
	    RECT 388.4000 51.6000 389.2000 52.4000 ;
	    RECT 409.2000 52.3000 410.0000 52.4000 ;
	    RECT 428.4000 52.3000 429.2000 52.4000 ;
	    RECT 409.2000 51.7000 429.2000 52.3000 ;
	    RECT 409.2000 51.6000 410.0000 51.7000 ;
	    RECT 428.4000 51.6000 429.2000 51.7000 ;
	    RECT 431.6000 52.3000 432.4000 52.4000 ;
	    RECT 436.4000 52.3000 437.2000 52.4000 ;
	    RECT 442.8000 52.3000 443.6000 52.4000 ;
	    RECT 446.0000 52.3000 446.8000 52.4000 ;
	    RECT 431.6000 51.7000 446.8000 52.3000 ;
	    RECT 431.6000 51.6000 432.4000 51.7000 ;
	    RECT 436.4000 51.6000 437.2000 51.7000 ;
	    RECT 442.8000 51.6000 443.6000 51.7000 ;
	    RECT 446.0000 51.6000 446.8000 51.7000 ;
	    RECT 470.0000 52.3000 470.8000 52.4000 ;
	    RECT 478.0000 52.3000 478.8000 52.4000 ;
	    RECT 487.6000 52.3000 488.4000 52.4000 ;
	    RECT 489.2000 52.3000 490.0000 52.4000 ;
	    RECT 470.0000 51.7000 490.0000 52.3000 ;
	    RECT 470.0000 51.6000 470.8000 51.7000 ;
	    RECT 478.0000 51.6000 478.8000 51.7000 ;
	    RECT 487.6000 51.6000 488.4000 51.7000 ;
	    RECT 489.2000 51.6000 490.0000 51.7000 ;
	    RECT 90.8000 50.3000 91.6000 50.4000 ;
	    RECT 54.1000 49.7000 91.6000 50.3000 ;
	    RECT 42.8000 49.6000 43.6000 49.7000 ;
	    RECT 52.4000 49.6000 53.2000 49.7000 ;
	    RECT 90.8000 49.6000 91.6000 49.7000 ;
	    RECT 92.4000 50.3000 93.2000 50.4000 ;
	    RECT 95.6000 50.3000 96.4000 50.4000 ;
	    RECT 92.4000 49.7000 96.4000 50.3000 ;
	    RECT 92.4000 49.6000 93.2000 49.7000 ;
	    RECT 95.6000 49.6000 96.4000 49.7000 ;
	    RECT 98.8000 50.3000 99.6000 50.4000 ;
	    RECT 106.8000 50.3000 107.6000 50.4000 ;
	    RECT 98.8000 49.7000 107.6000 50.3000 ;
	    RECT 98.8000 49.6000 99.6000 49.7000 ;
	    RECT 106.8000 49.6000 107.6000 49.7000 ;
	    RECT 166.0000 50.3000 166.8000 50.4000 ;
	    RECT 193.2000 50.3000 194.0000 50.4000 ;
	    RECT 166.0000 49.7000 194.0000 50.3000 ;
	    RECT 166.0000 49.6000 166.8000 49.7000 ;
	    RECT 193.2000 49.6000 194.0000 49.7000 ;
	    RECT 207.6000 50.3000 208.4000 50.4000 ;
	    RECT 212.4000 50.3000 213.2000 50.4000 ;
	    RECT 218.8000 50.3000 219.6000 50.4000 ;
	    RECT 207.6000 49.7000 219.6000 50.3000 ;
	    RECT 207.6000 49.6000 208.4000 49.7000 ;
	    RECT 212.4000 49.6000 213.2000 49.7000 ;
	    RECT 218.8000 49.6000 219.6000 49.7000 ;
	    RECT 220.4000 50.3000 221.2000 50.4000 ;
	    RECT 268.4000 50.3000 269.2000 50.4000 ;
	    RECT 220.4000 49.7000 269.2000 50.3000 ;
	    RECT 220.4000 49.6000 221.2000 49.7000 ;
	    RECT 268.4000 49.6000 269.2000 49.7000 ;
	    RECT 270.0000 50.3000 270.8000 50.4000 ;
	    RECT 278.0000 50.3000 278.8000 50.4000 ;
	    RECT 270.0000 49.7000 278.8000 50.3000 ;
	    RECT 270.0000 49.6000 270.8000 49.7000 ;
	    RECT 278.0000 49.6000 278.8000 49.7000 ;
	    RECT 279.6000 50.3000 280.4000 50.4000 ;
	    RECT 290.8000 50.3000 291.6000 50.4000 ;
	    RECT 297.2000 50.3000 298.0000 50.4000 ;
	    RECT 318.0000 50.3000 318.8000 50.4000 ;
	    RECT 279.6000 49.7000 298.0000 50.3000 ;
	    RECT 279.6000 49.6000 280.4000 49.7000 ;
	    RECT 290.8000 49.6000 291.6000 49.7000 ;
	    RECT 297.2000 49.6000 298.0000 49.7000 ;
	    RECT 298.9000 49.7000 318.8000 50.3000 ;
	    RECT 4.4000 48.3000 5.2000 48.4000 ;
	    RECT 20.4000 48.3000 21.2000 48.4000 ;
	    RECT 39.6000 48.3000 40.4000 48.4000 ;
	    RECT 4.4000 47.7000 40.4000 48.3000 ;
	    RECT 4.4000 47.6000 5.2000 47.7000 ;
	    RECT 20.4000 47.6000 21.2000 47.7000 ;
	    RECT 39.6000 47.6000 40.4000 47.7000 ;
	    RECT 42.8000 48.3000 43.6000 48.4000 ;
	    RECT 46.0000 48.3000 46.8000 48.4000 ;
	    RECT 42.8000 47.7000 46.8000 48.3000 ;
	    RECT 42.8000 47.6000 43.6000 47.7000 ;
	    RECT 46.0000 47.6000 46.8000 47.7000 ;
	    RECT 62.0000 48.3000 62.8000 48.4000 ;
	    RECT 158.0000 48.3000 158.8000 48.4000 ;
	    RECT 62.0000 47.7000 158.8000 48.3000 ;
	    RECT 62.0000 47.6000 62.8000 47.7000 ;
	    RECT 158.0000 47.6000 158.8000 47.7000 ;
	    RECT 174.0000 48.3000 174.8000 48.4000 ;
	    RECT 202.8000 48.3000 203.6000 48.4000 ;
	    RECT 174.0000 47.7000 203.6000 48.3000 ;
	    RECT 174.0000 47.6000 174.8000 47.7000 ;
	    RECT 202.8000 47.6000 203.6000 47.7000 ;
	    RECT 218.8000 48.3000 219.6000 48.4000 ;
	    RECT 246.0000 48.3000 246.8000 48.4000 ;
	    RECT 218.8000 47.7000 246.8000 48.3000 ;
	    RECT 218.8000 47.6000 219.6000 47.7000 ;
	    RECT 246.0000 47.6000 246.8000 47.7000 ;
	    RECT 257.2000 48.3000 258.0000 48.4000 ;
	    RECT 265.2000 48.3000 266.0000 48.4000 ;
	    RECT 271.6000 48.3000 272.4000 48.4000 ;
	    RECT 273.2000 48.3000 274.0000 48.4000 ;
	    RECT 257.2000 47.7000 274.0000 48.3000 ;
	    RECT 257.2000 47.6000 258.0000 47.7000 ;
	    RECT 265.2000 47.6000 266.0000 47.7000 ;
	    RECT 271.6000 47.6000 272.4000 47.7000 ;
	    RECT 273.2000 47.6000 274.0000 47.7000 ;
	    RECT 276.4000 48.3000 277.2000 48.4000 ;
	    RECT 298.9000 48.3000 299.5000 49.7000 ;
	    RECT 318.0000 49.6000 318.8000 49.7000 ;
	    RECT 329.2000 50.3000 330.0000 50.4000 ;
	    RECT 330.8000 50.3000 331.6000 50.4000 ;
	    RECT 329.2000 49.7000 331.6000 50.3000 ;
	    RECT 329.2000 49.6000 330.0000 49.7000 ;
	    RECT 330.8000 49.6000 331.6000 49.7000 ;
	    RECT 345.2000 50.3000 346.0000 50.4000 ;
	    RECT 364.4000 50.3000 365.2000 50.4000 ;
	    RECT 345.2000 49.7000 365.2000 50.3000 ;
	    RECT 345.2000 49.6000 346.0000 49.7000 ;
	    RECT 364.4000 49.6000 365.2000 49.7000 ;
	    RECT 393.2000 50.3000 394.0000 50.4000 ;
	    RECT 401.2000 50.3000 402.0000 50.4000 ;
	    RECT 393.2000 49.7000 402.0000 50.3000 ;
	    RECT 393.2000 49.6000 394.0000 49.7000 ;
	    RECT 401.2000 49.6000 402.0000 49.7000 ;
	    RECT 276.4000 47.7000 299.5000 48.3000 ;
	    RECT 302.0000 48.3000 302.8000 48.4000 ;
	    RECT 311.6000 48.3000 312.4000 48.4000 ;
	    RECT 302.0000 47.7000 312.4000 48.3000 ;
	    RECT 276.4000 47.6000 277.2000 47.7000 ;
	    RECT 302.0000 47.6000 302.8000 47.7000 ;
	    RECT 311.6000 47.6000 312.4000 47.7000 ;
	    RECT 324.4000 48.3000 325.2000 48.4000 ;
	    RECT 358.0000 48.3000 358.8000 48.4000 ;
	    RECT 324.4000 47.7000 358.8000 48.3000 ;
	    RECT 324.4000 47.6000 325.2000 47.7000 ;
	    RECT 358.0000 47.6000 358.8000 47.7000 ;
	    RECT 361.2000 48.3000 362.0000 48.4000 ;
	    RECT 385.2000 48.3000 386.0000 48.4000 ;
	    RECT 361.2000 47.7000 386.0000 48.3000 ;
	    RECT 361.2000 47.6000 362.0000 47.7000 ;
	    RECT 385.2000 47.6000 386.0000 47.7000 ;
	    RECT 468.4000 48.3000 469.2000 48.4000 ;
	    RECT 479.6000 48.3000 480.4000 48.4000 ;
	    RECT 486.0000 48.3000 486.8000 48.4000 ;
	    RECT 468.4000 47.7000 486.8000 48.3000 ;
	    RECT 468.4000 47.6000 469.2000 47.7000 ;
	    RECT 479.6000 47.6000 480.4000 47.7000 ;
	    RECT 486.0000 47.6000 486.8000 47.7000 ;
	    RECT 47.6000 46.3000 48.4000 46.4000 ;
	    RECT 58.8000 46.3000 59.6000 46.4000 ;
	    RECT 47.6000 45.7000 59.6000 46.3000 ;
	    RECT 47.6000 45.6000 48.4000 45.7000 ;
	    RECT 58.8000 45.6000 59.6000 45.7000 ;
	    RECT 82.8000 46.3000 83.6000 46.4000 ;
	    RECT 97.2000 46.3000 98.0000 46.4000 ;
	    RECT 82.8000 45.7000 98.0000 46.3000 ;
	    RECT 82.8000 45.6000 83.6000 45.7000 ;
	    RECT 97.2000 45.6000 98.0000 45.7000 ;
	    RECT 102.0000 46.3000 102.8000 46.4000 ;
	    RECT 113.2000 46.3000 114.0000 46.4000 ;
	    RECT 154.8000 46.3000 155.6000 46.4000 ;
	    RECT 167.6000 46.3000 168.4000 46.4000 ;
	    RECT 180.4000 46.3000 181.2000 46.4000 ;
	    RECT 102.0000 45.7000 181.2000 46.3000 ;
	    RECT 102.0000 45.6000 102.8000 45.7000 ;
	    RECT 113.2000 45.6000 114.0000 45.7000 ;
	    RECT 154.8000 45.6000 155.6000 45.7000 ;
	    RECT 167.6000 45.6000 168.4000 45.7000 ;
	    RECT 180.4000 45.6000 181.2000 45.7000 ;
	    RECT 222.0000 46.3000 222.8000 46.4000 ;
	    RECT 225.2000 46.3000 226.0000 46.4000 ;
	    RECT 233.2000 46.3000 234.0000 46.4000 ;
	    RECT 222.0000 45.7000 234.0000 46.3000 ;
	    RECT 222.0000 45.6000 222.8000 45.7000 ;
	    RECT 225.2000 45.6000 226.0000 45.7000 ;
	    RECT 233.2000 45.6000 234.0000 45.7000 ;
	    RECT 249.2000 46.3000 250.0000 46.4000 ;
	    RECT 263.6000 46.3000 264.4000 46.4000 ;
	    RECT 270.0000 46.3000 270.8000 46.4000 ;
	    RECT 281.2000 46.3000 282.0000 46.4000 ;
	    RECT 249.2000 45.7000 282.0000 46.3000 ;
	    RECT 249.2000 45.6000 250.0000 45.7000 ;
	    RECT 263.6000 45.6000 264.4000 45.7000 ;
	    RECT 270.0000 45.6000 270.8000 45.7000 ;
	    RECT 281.2000 45.6000 282.0000 45.7000 ;
	    RECT 290.8000 46.3000 291.6000 46.4000 ;
	    RECT 313.2000 46.3000 314.0000 46.4000 ;
	    RECT 346.8000 46.3000 347.6000 46.4000 ;
	    RECT 290.8000 45.7000 347.6000 46.3000 ;
	    RECT 290.8000 45.6000 291.6000 45.7000 ;
	    RECT 313.2000 45.6000 314.0000 45.7000 ;
	    RECT 346.8000 45.6000 347.6000 45.7000 ;
	    RECT 382.0000 46.3000 382.8000 46.4000 ;
	    RECT 385.2000 46.3000 386.0000 46.4000 ;
	    RECT 382.0000 45.7000 386.0000 46.3000 ;
	    RECT 382.0000 45.6000 382.8000 45.7000 ;
	    RECT 385.2000 45.6000 386.0000 45.7000 ;
	    RECT 111.6000 44.3000 112.4000 44.4000 ;
	    RECT 129.2000 44.3000 130.0000 44.4000 ;
	    RECT 111.6000 43.7000 130.0000 44.3000 ;
	    RECT 111.6000 43.6000 112.4000 43.7000 ;
	    RECT 129.2000 43.6000 130.0000 43.7000 ;
	    RECT 132.4000 44.3000 133.2000 44.4000 ;
	    RECT 174.0000 44.3000 174.8000 44.4000 ;
	    RECT 132.4000 43.7000 174.8000 44.3000 ;
	    RECT 132.4000 43.6000 133.2000 43.7000 ;
	    RECT 174.0000 43.6000 174.8000 43.7000 ;
	    RECT 217.2000 44.3000 218.0000 44.4000 ;
	    RECT 266.8000 44.3000 267.6000 44.4000 ;
	    RECT 298.8000 44.3000 299.6000 44.4000 ;
	    RECT 338.8000 44.3000 339.6000 44.4000 ;
	    RECT 217.2000 43.7000 339.6000 44.3000 ;
	    RECT 217.2000 43.6000 218.0000 43.7000 ;
	    RECT 266.8000 43.6000 267.6000 43.7000 ;
	    RECT 298.8000 43.6000 299.6000 43.7000 ;
	    RECT 338.8000 43.6000 339.6000 43.7000 ;
	    RECT 254.0000 42.3000 254.8000 42.4000 ;
	    RECT 262.0000 42.3000 262.8000 42.4000 ;
	    RECT 254.0000 41.7000 262.8000 42.3000 ;
	    RECT 254.0000 41.6000 254.8000 41.7000 ;
	    RECT 262.0000 41.6000 262.8000 41.7000 ;
	    RECT 263.6000 42.3000 264.4000 42.4000 ;
	    RECT 337.2000 42.3000 338.0000 42.4000 ;
	    RECT 263.6000 41.7000 338.0000 42.3000 ;
	    RECT 263.6000 41.6000 264.4000 41.7000 ;
	    RECT 337.2000 41.6000 338.0000 41.7000 ;
	    RECT 124.4000 40.3000 125.2000 40.4000 ;
	    RECT 172.4000 40.3000 173.2000 40.4000 ;
	    RECT 124.4000 39.7000 173.2000 40.3000 ;
	    RECT 124.4000 39.6000 125.2000 39.7000 ;
	    RECT 172.4000 39.6000 173.2000 39.7000 ;
	    RECT 177.2000 40.3000 178.0000 40.4000 ;
	    RECT 204.4000 40.3000 205.2000 40.4000 ;
	    RECT 177.2000 39.7000 205.2000 40.3000 ;
	    RECT 177.2000 39.6000 178.0000 39.7000 ;
	    RECT 204.4000 39.6000 205.2000 39.7000 ;
	    RECT 215.6000 40.3000 216.4000 40.4000 ;
	    RECT 292.4000 40.3000 293.2000 40.4000 ;
	    RECT 215.6000 39.7000 293.2000 40.3000 ;
	    RECT 215.6000 39.6000 216.4000 39.7000 ;
	    RECT 292.4000 39.6000 293.2000 39.7000 ;
	    RECT 294.0000 40.3000 294.8000 40.4000 ;
	    RECT 308.4000 40.3000 309.2000 40.4000 ;
	    RECT 294.0000 39.7000 309.2000 40.3000 ;
	    RECT 294.0000 39.6000 294.8000 39.7000 ;
	    RECT 308.4000 39.6000 309.2000 39.7000 ;
	    RECT 314.8000 40.3000 315.6000 40.4000 ;
	    RECT 401.2000 40.3000 402.0000 40.4000 ;
	    RECT 314.8000 39.7000 402.0000 40.3000 ;
	    RECT 314.8000 39.6000 315.6000 39.7000 ;
	    RECT 401.2000 39.6000 402.0000 39.7000 ;
	    RECT 49.2000 38.3000 50.0000 38.4000 ;
	    RECT 94.0000 38.3000 94.8000 38.4000 ;
	    RECT 49.2000 37.7000 94.8000 38.3000 ;
	    RECT 49.2000 37.6000 50.0000 37.7000 ;
	    RECT 94.0000 37.6000 94.8000 37.7000 ;
	    RECT 95.6000 38.3000 96.4000 38.4000 ;
	    RECT 134.0000 38.3000 134.8000 38.4000 ;
	    RECT 148.4000 38.3000 149.2000 38.4000 ;
	    RECT 95.6000 37.7000 104.3000 38.3000 ;
	    RECT 95.6000 37.6000 96.4000 37.7000 ;
	    RECT 14.0000 36.3000 14.8000 36.4000 ;
	    RECT 57.2000 36.3000 58.0000 36.4000 ;
	    RECT 14.0000 35.7000 58.0000 36.3000 ;
	    RECT 14.0000 35.6000 14.8000 35.7000 ;
	    RECT 57.2000 35.6000 58.0000 35.7000 ;
	    RECT 95.6000 36.3000 96.4000 36.4000 ;
	    RECT 102.0000 36.3000 102.8000 36.4000 ;
	    RECT 95.6000 35.7000 102.8000 36.3000 ;
	    RECT 103.7000 36.3000 104.3000 37.7000 ;
	    RECT 134.0000 37.7000 149.2000 38.3000 ;
	    RECT 134.0000 37.6000 134.8000 37.7000 ;
	    RECT 148.4000 37.6000 149.2000 37.7000 ;
	    RECT 188.4000 38.3000 189.2000 38.4000 ;
	    RECT 191.6000 38.3000 192.4000 38.4000 ;
	    RECT 188.4000 37.7000 192.4000 38.3000 ;
	    RECT 188.4000 37.6000 189.2000 37.7000 ;
	    RECT 191.6000 37.6000 192.4000 37.7000 ;
	    RECT 238.0000 38.3000 238.8000 38.4000 ;
	    RECT 382.0000 38.3000 382.8000 38.4000 ;
	    RECT 391.6000 38.3000 392.4000 38.4000 ;
	    RECT 238.0000 37.7000 392.4000 38.3000 ;
	    RECT 238.0000 37.6000 238.8000 37.7000 ;
	    RECT 382.0000 37.6000 382.8000 37.7000 ;
	    RECT 391.6000 37.6000 392.4000 37.7000 ;
	    RECT 401.2000 38.3000 402.0000 38.4000 ;
	    RECT 418.8000 38.3000 419.6000 38.4000 ;
	    RECT 401.2000 37.7000 419.6000 38.3000 ;
	    RECT 401.2000 37.6000 402.0000 37.7000 ;
	    RECT 418.8000 37.6000 419.6000 37.7000 ;
	    RECT 476.4000 38.3000 477.2000 38.4000 ;
	    RECT 486.0000 38.3000 486.8000 38.4000 ;
	    RECT 495.6000 38.3000 496.4000 38.4000 ;
	    RECT 476.4000 37.7000 496.4000 38.3000 ;
	    RECT 476.4000 37.6000 477.2000 37.7000 ;
	    RECT 486.0000 37.6000 486.8000 37.7000 ;
	    RECT 495.6000 37.6000 496.4000 37.7000 ;
	    RECT 260.4000 36.3000 261.2000 36.4000 ;
	    RECT 103.7000 35.7000 261.2000 36.3000 ;
	    RECT 95.6000 35.6000 96.4000 35.7000 ;
	    RECT 102.0000 35.6000 102.8000 35.7000 ;
	    RECT 260.4000 35.6000 261.2000 35.7000 ;
	    RECT 266.8000 36.3000 267.6000 36.4000 ;
	    RECT 300.4000 36.3000 301.2000 36.4000 ;
	    RECT 266.8000 35.7000 301.2000 36.3000 ;
	    RECT 266.8000 35.6000 267.6000 35.7000 ;
	    RECT 300.4000 35.6000 301.2000 35.7000 ;
	    RECT 311.6000 36.3000 312.4000 36.4000 ;
	    RECT 343.6000 36.3000 344.4000 36.4000 ;
	    RECT 353.2000 36.3000 354.0000 36.4000 ;
	    RECT 311.6000 35.7000 354.0000 36.3000 ;
	    RECT 311.6000 35.6000 312.4000 35.7000 ;
	    RECT 343.6000 35.6000 344.4000 35.7000 ;
	    RECT 353.2000 35.6000 354.0000 35.7000 ;
	    RECT 356.4000 36.3000 357.2000 36.4000 ;
	    RECT 362.8000 36.3000 363.6000 36.4000 ;
	    RECT 356.4000 35.7000 363.6000 36.3000 ;
	    RECT 356.4000 35.6000 357.2000 35.7000 ;
	    RECT 362.8000 35.6000 363.6000 35.7000 ;
	    RECT 415.6000 36.3000 416.4000 36.4000 ;
	    RECT 457.2000 36.3000 458.0000 36.4000 ;
	    RECT 415.6000 35.7000 458.0000 36.3000 ;
	    RECT 415.6000 35.6000 416.4000 35.7000 ;
	    RECT 457.2000 35.6000 458.0000 35.7000 ;
	    RECT 1.2000 34.3000 2.0000 34.4000 ;
	    RECT 46.0000 34.3000 46.8000 34.4000 ;
	    RECT 1.2000 33.7000 46.8000 34.3000 ;
	    RECT 1.2000 33.6000 2.0000 33.7000 ;
	    RECT 46.0000 33.6000 46.8000 33.7000 ;
	    RECT 62.0000 34.3000 62.8000 34.4000 ;
	    RECT 98.8000 34.3000 99.6000 34.4000 ;
	    RECT 62.0000 33.7000 99.6000 34.3000 ;
	    RECT 62.0000 33.6000 62.8000 33.7000 ;
	    RECT 98.8000 33.6000 99.6000 33.7000 ;
	    RECT 185.2000 34.3000 186.0000 34.4000 ;
	    RECT 233.2000 34.3000 234.0000 34.4000 ;
	    RECT 257.2000 34.3000 258.0000 34.4000 ;
	    RECT 185.2000 33.7000 224.3000 34.3000 ;
	    RECT 185.2000 33.6000 186.0000 33.7000 ;
	    RECT 94.0000 32.3000 94.8000 32.4000 ;
	    RECT 132.4000 32.3000 133.2000 32.4000 ;
	    RECT 134.0000 32.3000 134.8000 32.4000 ;
	    RECT 161.2000 32.3000 162.0000 32.4000 ;
	    RECT 186.8000 32.3000 187.6000 32.4000 ;
	    RECT 94.0000 31.7000 187.6000 32.3000 ;
	    RECT 94.0000 31.6000 94.8000 31.7000 ;
	    RECT 132.4000 31.6000 133.2000 31.7000 ;
	    RECT 134.0000 31.6000 134.8000 31.7000 ;
	    RECT 161.2000 31.6000 162.0000 31.7000 ;
	    RECT 186.8000 31.6000 187.6000 31.7000 ;
	    RECT 191.6000 32.3000 192.4000 32.4000 ;
	    RECT 201.2000 32.3000 202.0000 32.4000 ;
	    RECT 191.6000 31.7000 202.0000 32.3000 ;
	    RECT 191.6000 31.6000 192.4000 31.7000 ;
	    RECT 201.2000 31.6000 202.0000 31.7000 ;
	    RECT 214.0000 32.3000 214.8000 32.4000 ;
	    RECT 222.0000 32.3000 222.8000 32.4000 ;
	    RECT 214.0000 31.7000 222.8000 32.3000 ;
	    RECT 223.7000 32.3000 224.3000 33.7000 ;
	    RECT 233.2000 33.7000 258.0000 34.3000 ;
	    RECT 233.2000 33.6000 234.0000 33.7000 ;
	    RECT 257.2000 33.6000 258.0000 33.7000 ;
	    RECT 260.4000 34.3000 261.2000 34.4000 ;
	    RECT 263.6000 34.3000 264.4000 34.4000 ;
	    RECT 260.4000 33.7000 264.4000 34.3000 ;
	    RECT 260.4000 33.6000 261.2000 33.7000 ;
	    RECT 263.6000 33.6000 264.4000 33.7000 ;
	    RECT 265.2000 34.3000 266.0000 34.4000 ;
	    RECT 270.0000 34.3000 270.8000 34.4000 ;
	    RECT 265.2000 33.7000 270.8000 34.3000 ;
	    RECT 265.2000 33.6000 266.0000 33.7000 ;
	    RECT 270.0000 33.6000 270.8000 33.7000 ;
	    RECT 279.6000 34.3000 280.4000 34.4000 ;
	    RECT 287.6000 34.3000 288.4000 34.4000 ;
	    RECT 279.6000 33.7000 288.4000 34.3000 ;
	    RECT 279.6000 33.6000 280.4000 33.7000 ;
	    RECT 287.6000 33.6000 288.4000 33.7000 ;
	    RECT 289.2000 34.3000 290.0000 34.4000 ;
	    RECT 322.8000 34.3000 323.6000 34.4000 ;
	    RECT 481.2000 34.3000 482.0000 34.4000 ;
	    RECT 490.8000 34.3000 491.6000 34.4000 ;
	    RECT 289.2000 33.7000 491.6000 34.3000 ;
	    RECT 289.2000 33.6000 290.0000 33.7000 ;
	    RECT 322.8000 33.6000 323.6000 33.7000 ;
	    RECT 481.2000 33.6000 482.0000 33.7000 ;
	    RECT 490.8000 33.6000 491.6000 33.7000 ;
	    RECT 276.4000 32.3000 277.2000 32.4000 ;
	    RECT 223.7000 31.7000 277.2000 32.3000 ;
	    RECT 214.0000 31.6000 214.8000 31.7000 ;
	    RECT 222.0000 31.6000 222.8000 31.7000 ;
	    RECT 276.4000 31.6000 277.2000 31.7000 ;
	    RECT 281.2000 32.3000 282.0000 32.4000 ;
	    RECT 289.2000 32.3000 290.0000 32.4000 ;
	    RECT 300.4000 32.3000 301.2000 32.4000 ;
	    RECT 281.2000 31.7000 290.0000 32.3000 ;
	    RECT 281.2000 31.6000 282.0000 31.7000 ;
	    RECT 289.2000 31.6000 290.0000 31.7000 ;
	    RECT 297.3000 31.7000 301.2000 32.3000 ;
	    RECT 42.8000 30.3000 43.6000 30.4000 ;
	    RECT 54.0000 30.3000 54.8000 30.4000 ;
	    RECT 42.8000 29.7000 54.8000 30.3000 ;
	    RECT 42.8000 29.6000 43.6000 29.7000 ;
	    RECT 54.0000 29.6000 54.8000 29.7000 ;
	    RECT 63.6000 30.3000 64.4000 30.4000 ;
	    RECT 129.2000 30.3000 130.0000 30.4000 ;
	    RECT 63.6000 29.7000 130.0000 30.3000 ;
	    RECT 63.6000 29.6000 64.4000 29.7000 ;
	    RECT 129.2000 29.6000 130.0000 29.7000 ;
	    RECT 135.6000 30.3000 136.4000 30.4000 ;
	    RECT 162.8000 30.3000 163.6000 30.4000 ;
	    RECT 135.6000 29.7000 163.6000 30.3000 ;
	    RECT 135.6000 29.6000 136.4000 29.7000 ;
	    RECT 162.8000 29.6000 163.6000 29.7000 ;
	    RECT 180.4000 30.3000 181.2000 30.4000 ;
	    RECT 194.8000 30.3000 195.6000 30.4000 ;
	    RECT 180.4000 29.7000 195.6000 30.3000 ;
	    RECT 180.4000 29.6000 181.2000 29.7000 ;
	    RECT 194.8000 29.6000 195.6000 29.7000 ;
	    RECT 198.0000 30.3000 198.8000 30.4000 ;
	    RECT 225.2000 30.3000 226.0000 30.4000 ;
	    RECT 236.4000 30.3000 237.2000 30.4000 ;
	    RECT 198.0000 29.7000 237.2000 30.3000 ;
	    RECT 198.0000 29.6000 198.8000 29.7000 ;
	    RECT 225.2000 29.6000 226.0000 29.7000 ;
	    RECT 236.4000 29.6000 237.2000 29.7000 ;
	    RECT 263.6000 30.3000 264.4000 30.4000 ;
	    RECT 268.4000 30.3000 269.2000 30.4000 ;
	    RECT 263.6000 29.7000 269.2000 30.3000 ;
	    RECT 263.6000 29.6000 264.4000 29.7000 ;
	    RECT 268.4000 29.6000 269.2000 29.7000 ;
	    RECT 273.2000 30.3000 274.0000 30.4000 ;
	    RECT 274.8000 30.3000 275.6000 30.4000 ;
	    RECT 273.2000 29.7000 275.6000 30.3000 ;
	    RECT 273.2000 29.6000 274.0000 29.7000 ;
	    RECT 274.8000 29.6000 275.6000 29.7000 ;
	    RECT 276.4000 30.3000 277.2000 30.4000 ;
	    RECT 286.0000 30.3000 286.8000 30.4000 ;
	    RECT 276.4000 29.7000 286.8000 30.3000 ;
	    RECT 276.4000 29.6000 277.2000 29.7000 ;
	    RECT 286.0000 29.6000 286.8000 29.7000 ;
	    RECT 289.2000 30.3000 290.0000 30.4000 ;
	    RECT 297.3000 30.3000 297.9000 31.7000 ;
	    RECT 300.4000 31.6000 301.2000 31.7000 ;
	    RECT 306.8000 32.3000 307.6000 32.4000 ;
	    RECT 308.4000 32.3000 309.2000 32.4000 ;
	    RECT 306.8000 31.7000 309.2000 32.3000 ;
	    RECT 306.8000 31.6000 307.6000 31.7000 ;
	    RECT 308.4000 31.6000 309.2000 31.7000 ;
	    RECT 311.6000 32.3000 312.4000 32.4000 ;
	    RECT 316.4000 32.3000 317.2000 32.4000 ;
	    RECT 311.6000 31.7000 317.2000 32.3000 ;
	    RECT 311.6000 31.6000 312.4000 31.7000 ;
	    RECT 316.4000 31.6000 317.2000 31.7000 ;
	    RECT 318.0000 32.3000 318.8000 32.4000 ;
	    RECT 334.0000 32.3000 334.8000 32.4000 ;
	    RECT 318.0000 31.7000 334.8000 32.3000 ;
	    RECT 318.0000 31.6000 318.8000 31.7000 ;
	    RECT 334.0000 31.6000 334.8000 31.7000 ;
	    RECT 356.4000 32.3000 357.2000 32.4000 ;
	    RECT 364.4000 32.3000 365.2000 32.4000 ;
	    RECT 356.4000 31.7000 365.2000 32.3000 ;
	    RECT 356.4000 31.6000 357.2000 31.7000 ;
	    RECT 364.4000 31.6000 365.2000 31.7000 ;
	    RECT 394.8000 32.3000 395.6000 32.4000 ;
	    RECT 404.4000 32.3000 405.2000 32.4000 ;
	    RECT 415.6000 32.3000 416.4000 32.4000 ;
	    RECT 394.8000 31.7000 416.4000 32.3000 ;
	    RECT 394.8000 31.6000 395.6000 31.7000 ;
	    RECT 404.4000 31.6000 405.2000 31.7000 ;
	    RECT 415.6000 31.6000 416.4000 31.7000 ;
	    RECT 449.2000 32.3000 450.0000 32.4000 ;
	    RECT 466.8000 32.3000 467.6000 32.4000 ;
	    RECT 449.2000 31.7000 467.6000 32.3000 ;
	    RECT 449.2000 31.6000 450.0000 31.7000 ;
	    RECT 466.8000 31.6000 467.6000 31.7000 ;
	    RECT 289.2000 29.7000 297.9000 30.3000 ;
	    RECT 298.8000 30.3000 299.6000 30.4000 ;
	    RECT 366.0000 30.3000 366.8000 30.4000 ;
	    RECT 378.8000 30.3000 379.6000 30.4000 ;
	    RECT 388.4000 30.3000 389.2000 30.4000 ;
	    RECT 298.8000 29.7000 389.2000 30.3000 ;
	    RECT 289.2000 29.6000 290.0000 29.7000 ;
	    RECT 298.8000 29.6000 299.6000 29.7000 ;
	    RECT 366.0000 29.6000 366.8000 29.7000 ;
	    RECT 378.8000 29.6000 379.6000 29.7000 ;
	    RECT 388.4000 29.6000 389.2000 29.7000 ;
	    RECT 394.8000 30.3000 395.6000 30.4000 ;
	    RECT 398.0000 30.3000 398.8000 30.4000 ;
	    RECT 394.8000 29.7000 398.8000 30.3000 ;
	    RECT 394.8000 29.6000 395.6000 29.7000 ;
	    RECT 398.0000 29.6000 398.8000 29.7000 ;
	    RECT 414.0000 30.3000 414.8000 30.4000 ;
	    RECT 426.8000 30.3000 427.6000 30.4000 ;
	    RECT 414.0000 29.7000 427.6000 30.3000 ;
	    RECT 414.0000 29.6000 414.8000 29.7000 ;
	    RECT 426.8000 29.6000 427.6000 29.7000 ;
	    RECT 466.8000 30.3000 467.6000 30.4000 ;
	    RECT 476.4000 30.3000 477.2000 30.4000 ;
	    RECT 466.8000 29.7000 477.2000 30.3000 ;
	    RECT 466.8000 29.6000 467.6000 29.7000 ;
	    RECT 476.4000 29.6000 477.2000 29.7000 ;
	    RECT 489.2000 30.3000 490.0000 30.4000 ;
	    RECT 500.4000 30.3000 501.2000 30.4000 ;
	    RECT 489.2000 29.7000 501.2000 30.3000 ;
	    RECT 489.2000 29.6000 490.0000 29.7000 ;
	    RECT 500.4000 29.6000 501.2000 29.7000 ;
	    RECT 34.8000 28.3000 35.6000 28.4000 ;
	    RECT 44.4000 28.3000 45.2000 28.4000 ;
	    RECT 50.8000 28.3000 51.6000 28.4000 ;
	    RECT 71.6000 28.3000 72.4000 28.4000 ;
	    RECT 34.8000 27.7000 72.4000 28.3000 ;
	    RECT 34.8000 27.6000 35.6000 27.7000 ;
	    RECT 44.4000 27.6000 45.2000 27.7000 ;
	    RECT 50.8000 27.6000 51.6000 27.7000 ;
	    RECT 71.6000 27.6000 72.4000 27.7000 ;
	    RECT 76.4000 28.3000 77.2000 28.4000 ;
	    RECT 94.0000 28.3000 94.8000 28.4000 ;
	    RECT 76.4000 27.7000 94.8000 28.3000 ;
	    RECT 76.4000 27.6000 77.2000 27.7000 ;
	    RECT 94.0000 27.6000 94.8000 27.7000 ;
	    RECT 132.4000 28.3000 133.2000 28.4000 ;
	    RECT 135.6000 28.3000 136.4000 28.4000 ;
	    RECT 132.4000 27.7000 136.4000 28.3000 ;
	    RECT 132.4000 27.6000 133.2000 27.7000 ;
	    RECT 135.6000 27.6000 136.4000 27.7000 ;
	    RECT 154.8000 28.3000 155.6000 28.4000 ;
	    RECT 172.4000 28.3000 173.2000 28.4000 ;
	    RECT 154.8000 27.7000 173.2000 28.3000 ;
	    RECT 154.8000 27.6000 155.6000 27.7000 ;
	    RECT 172.4000 27.6000 173.2000 27.7000 ;
	    RECT 194.8000 28.3000 195.6000 28.4000 ;
	    RECT 215.6000 28.3000 216.4000 28.4000 ;
	    RECT 194.8000 27.7000 216.4000 28.3000 ;
	    RECT 194.8000 27.6000 195.6000 27.7000 ;
	    RECT 215.6000 27.6000 216.4000 27.7000 ;
	    RECT 230.0000 28.3000 230.8000 28.4000 ;
	    RECT 244.4000 28.3000 245.2000 28.4000 ;
	    RECT 278.0000 28.3000 278.8000 28.4000 ;
	    RECT 303.6000 28.3000 304.4000 28.4000 ;
	    RECT 230.0000 27.7000 304.4000 28.3000 ;
	    RECT 230.0000 27.6000 230.8000 27.7000 ;
	    RECT 244.4000 27.6000 245.2000 27.7000 ;
	    RECT 278.0000 27.6000 278.8000 27.7000 ;
	    RECT 303.6000 27.6000 304.4000 27.7000 ;
	    RECT 318.0000 28.3000 318.8000 28.4000 ;
	    RECT 319.6000 28.3000 320.4000 28.4000 ;
	    RECT 330.8000 28.3000 331.6000 28.4000 ;
	    RECT 318.0000 27.7000 331.6000 28.3000 ;
	    RECT 318.0000 27.6000 318.8000 27.7000 ;
	    RECT 319.6000 27.6000 320.4000 27.7000 ;
	    RECT 330.8000 27.6000 331.6000 27.7000 ;
	    RECT 334.0000 28.3000 334.8000 28.4000 ;
	    RECT 340.4000 28.3000 341.2000 28.4000 ;
	    RECT 369.2000 28.3000 370.0000 28.4000 ;
	    RECT 375.6000 28.3000 376.4000 28.4000 ;
	    RECT 334.0000 27.7000 339.5000 28.3000 ;
	    RECT 334.0000 27.6000 334.8000 27.7000 ;
	    RECT 140.4000 26.3000 141.2000 26.4000 ;
	    RECT 158.0000 26.3000 158.8000 26.4000 ;
	    RECT 140.4000 25.7000 158.8000 26.3000 ;
	    RECT 140.4000 25.6000 141.2000 25.7000 ;
	    RECT 158.0000 25.6000 158.8000 25.7000 ;
	    RECT 190.0000 26.3000 190.8000 26.4000 ;
	    RECT 196.4000 26.3000 197.2000 26.4000 ;
	    RECT 206.0000 26.3000 206.8000 26.4000 ;
	    RECT 209.2000 26.3000 210.0000 26.4000 ;
	    RECT 190.0000 25.7000 210.0000 26.3000 ;
	    RECT 190.0000 25.6000 190.8000 25.7000 ;
	    RECT 196.4000 25.6000 197.2000 25.7000 ;
	    RECT 206.0000 25.6000 206.8000 25.7000 ;
	    RECT 209.2000 25.6000 210.0000 25.7000 ;
	    RECT 220.4000 26.3000 221.2000 26.4000 ;
	    RECT 228.4000 26.3000 229.2000 26.4000 ;
	    RECT 263.6000 26.3000 264.4000 26.4000 ;
	    RECT 314.8000 26.3000 315.6000 26.4000 ;
	    RECT 324.4000 26.3000 325.2000 26.4000 ;
	    RECT 332.4000 26.3000 333.2000 26.4000 ;
	    RECT 220.4000 25.7000 333.2000 26.3000 ;
	    RECT 220.4000 25.6000 221.2000 25.7000 ;
	    RECT 228.4000 25.6000 229.2000 25.7000 ;
	    RECT 263.6000 25.6000 264.4000 25.7000 ;
	    RECT 314.8000 25.6000 315.6000 25.7000 ;
	    RECT 324.4000 25.6000 325.2000 25.7000 ;
	    RECT 332.4000 25.6000 333.2000 25.7000 ;
	    RECT 335.6000 26.3000 336.4000 26.4000 ;
	    RECT 337.2000 26.3000 338.0000 26.4000 ;
	    RECT 335.6000 25.7000 338.0000 26.3000 ;
	    RECT 338.9000 26.3000 339.5000 27.7000 ;
	    RECT 340.4000 27.7000 376.4000 28.3000 ;
	    RECT 340.4000 27.6000 341.2000 27.7000 ;
	    RECT 369.2000 27.6000 370.0000 27.7000 ;
	    RECT 375.6000 27.6000 376.4000 27.7000 ;
	    RECT 398.0000 28.3000 398.8000 28.4000 ;
	    RECT 425.2000 28.3000 426.0000 28.4000 ;
	    RECT 398.0000 27.7000 426.0000 28.3000 ;
	    RECT 398.0000 27.6000 398.8000 27.7000 ;
	    RECT 425.2000 27.6000 426.0000 27.7000 ;
	    RECT 454.0000 28.3000 454.8000 28.4000 ;
	    RECT 468.4000 28.3000 469.2000 28.4000 ;
	    RECT 454.0000 27.7000 469.2000 28.3000 ;
	    RECT 454.0000 27.6000 454.8000 27.7000 ;
	    RECT 468.4000 27.6000 469.2000 27.7000 ;
	    RECT 353.2000 26.3000 354.0000 26.4000 ;
	    RECT 374.0000 26.3000 374.8000 26.4000 ;
	    RECT 338.9000 25.7000 354.0000 26.3000 ;
	    RECT 335.6000 25.6000 336.4000 25.7000 ;
	    RECT 337.2000 25.6000 338.0000 25.7000 ;
	    RECT 353.2000 25.6000 354.0000 25.7000 ;
	    RECT 366.1000 25.7000 374.8000 26.3000 ;
	    RECT 366.1000 24.4000 366.7000 25.7000 ;
	    RECT 374.0000 25.6000 374.8000 25.7000 ;
	    RECT 438.0000 26.3000 438.8000 26.4000 ;
	    RECT 462.0000 26.3000 462.8000 26.4000 ;
	    RECT 438.0000 25.7000 462.8000 26.3000 ;
	    RECT 438.0000 25.6000 438.8000 25.7000 ;
	    RECT 462.0000 25.6000 462.8000 25.7000 ;
	    RECT 70.0000 24.3000 70.8000 24.4000 ;
	    RECT 79.6000 24.3000 80.4000 24.4000 ;
	    RECT 89.2000 24.3000 90.0000 24.4000 ;
	    RECT 70.0000 23.7000 90.0000 24.3000 ;
	    RECT 70.0000 23.6000 70.8000 23.7000 ;
	    RECT 79.6000 23.6000 80.4000 23.7000 ;
	    RECT 89.2000 23.6000 90.0000 23.7000 ;
	    RECT 100.4000 24.3000 101.2000 24.4000 ;
	    RECT 119.6000 24.3000 120.4000 24.4000 ;
	    RECT 124.4000 24.3000 125.2000 24.4000 ;
	    RECT 130.8000 24.3000 131.6000 24.4000 ;
	    RECT 100.4000 23.7000 131.6000 24.3000 ;
	    RECT 100.4000 23.6000 101.2000 23.7000 ;
	    RECT 119.6000 23.6000 120.4000 23.7000 ;
	    RECT 124.4000 23.6000 125.2000 23.7000 ;
	    RECT 130.8000 23.6000 131.6000 23.7000 ;
	    RECT 159.6000 24.3000 160.4000 24.4000 ;
	    RECT 215.6000 24.3000 216.4000 24.4000 ;
	    RECT 159.6000 23.7000 216.4000 24.3000 ;
	    RECT 159.6000 23.6000 160.4000 23.7000 ;
	    RECT 215.6000 23.6000 216.4000 23.7000 ;
	    RECT 218.8000 24.3000 219.6000 24.4000 ;
	    RECT 239.6000 24.3000 240.4000 24.4000 ;
	    RECT 308.4000 24.3000 309.2000 24.4000 ;
	    RECT 340.4000 24.3000 341.2000 24.4000 ;
	    RECT 218.8000 23.7000 240.4000 24.3000 ;
	    RECT 218.8000 23.6000 219.6000 23.7000 ;
	    RECT 239.6000 23.6000 240.4000 23.7000 ;
	    RECT 241.3000 23.7000 288.3000 24.3000 ;
	    RECT 98.8000 22.3000 99.6000 22.4000 ;
	    RECT 241.3000 22.3000 241.9000 23.7000 ;
	    RECT 98.8000 21.7000 241.9000 22.3000 ;
	    RECT 262.0000 22.3000 262.8000 22.4000 ;
	    RECT 286.0000 22.3000 286.8000 22.4000 ;
	    RECT 262.0000 21.7000 286.8000 22.3000 ;
	    RECT 287.7000 22.3000 288.3000 23.7000 ;
	    RECT 308.4000 23.7000 341.2000 24.3000 ;
	    RECT 308.4000 23.6000 309.2000 23.7000 ;
	    RECT 340.4000 23.6000 341.2000 23.7000 ;
	    RECT 342.0000 24.3000 342.8000 24.4000 ;
	    RECT 366.0000 24.3000 366.8000 24.4000 ;
	    RECT 342.0000 23.7000 366.8000 24.3000 ;
	    RECT 342.0000 23.6000 342.8000 23.7000 ;
	    RECT 366.0000 23.6000 366.8000 23.7000 ;
	    RECT 367.6000 24.3000 368.4000 24.4000 ;
	    RECT 417.2000 24.3000 418.0000 24.4000 ;
	    RECT 444.4000 24.3000 445.2000 24.4000 ;
	    RECT 367.6000 23.7000 445.2000 24.3000 ;
	    RECT 367.6000 23.6000 368.4000 23.7000 ;
	    RECT 417.2000 23.6000 418.0000 23.7000 ;
	    RECT 444.4000 23.6000 445.2000 23.7000 ;
	    RECT 311.6000 22.3000 312.4000 22.4000 ;
	    RECT 287.7000 21.7000 312.4000 22.3000 ;
	    RECT 98.8000 21.6000 99.6000 21.7000 ;
	    RECT 262.0000 21.6000 262.8000 21.7000 ;
	    RECT 286.0000 21.6000 286.8000 21.7000 ;
	    RECT 311.6000 21.6000 312.4000 21.7000 ;
	    RECT 314.8000 22.3000 315.6000 22.4000 ;
	    RECT 321.2000 22.3000 322.0000 22.4000 ;
	    RECT 314.8000 21.7000 322.0000 22.3000 ;
	    RECT 314.8000 21.6000 315.6000 21.7000 ;
	    RECT 321.2000 21.6000 322.0000 21.7000 ;
	    RECT 322.8000 22.3000 323.6000 22.4000 ;
	    RECT 327.6000 22.3000 328.4000 22.4000 ;
	    RECT 322.8000 21.7000 328.4000 22.3000 ;
	    RECT 322.8000 21.6000 323.6000 21.7000 ;
	    RECT 327.6000 21.6000 328.4000 21.7000 ;
	    RECT 329.2000 22.3000 330.0000 22.4000 ;
	    RECT 334.0000 22.3000 334.8000 22.4000 ;
	    RECT 329.2000 21.7000 334.8000 22.3000 ;
	    RECT 329.2000 21.6000 330.0000 21.7000 ;
	    RECT 334.0000 21.6000 334.8000 21.7000 ;
	    RECT 335.6000 22.3000 336.4000 22.4000 ;
	    RECT 346.8000 22.3000 347.6000 22.4000 ;
	    RECT 335.6000 21.7000 347.6000 22.3000 ;
	    RECT 335.6000 21.6000 336.4000 21.7000 ;
	    RECT 346.8000 21.6000 347.6000 21.7000 ;
	    RECT 348.4000 22.3000 349.2000 22.4000 ;
	    RECT 438.0000 22.3000 438.8000 22.4000 ;
	    RECT 348.4000 21.7000 438.8000 22.3000 ;
	    RECT 348.4000 21.6000 349.2000 21.7000 ;
	    RECT 438.0000 21.6000 438.8000 21.7000 ;
	    RECT 33.2000 20.3000 34.0000 20.4000 ;
	    RECT 42.8000 20.3000 43.6000 20.4000 ;
	    RECT 33.2000 19.7000 43.6000 20.3000 ;
	    RECT 33.2000 19.6000 34.0000 19.7000 ;
	    RECT 42.8000 19.6000 43.6000 19.7000 ;
	    RECT 113.2000 20.3000 114.0000 20.4000 ;
	    RECT 119.6000 20.3000 120.4000 20.4000 ;
	    RECT 113.2000 19.7000 120.4000 20.3000 ;
	    RECT 113.2000 19.6000 114.0000 19.7000 ;
	    RECT 119.6000 19.6000 120.4000 19.7000 ;
	    RECT 209.2000 20.3000 210.0000 20.4000 ;
	    RECT 218.8000 20.3000 219.6000 20.4000 ;
	    RECT 209.2000 19.7000 219.6000 20.3000 ;
	    RECT 209.2000 19.6000 210.0000 19.7000 ;
	    RECT 218.8000 19.6000 219.6000 19.7000 ;
	    RECT 236.4000 20.3000 237.2000 20.4000 ;
	    RECT 250.8000 20.3000 251.6000 20.4000 ;
	    RECT 236.4000 19.7000 251.6000 20.3000 ;
	    RECT 236.4000 19.6000 237.2000 19.7000 ;
	    RECT 250.8000 19.6000 251.6000 19.7000 ;
	    RECT 270.0000 20.3000 270.8000 20.4000 ;
	    RECT 348.4000 20.3000 349.2000 20.4000 ;
	    RECT 270.0000 19.7000 349.2000 20.3000 ;
	    RECT 270.0000 19.6000 270.8000 19.7000 ;
	    RECT 348.4000 19.6000 349.2000 19.7000 ;
	    RECT 359.6000 20.3000 360.4000 20.4000 ;
	    RECT 385.2000 20.3000 386.0000 20.4000 ;
	    RECT 359.6000 19.7000 386.0000 20.3000 ;
	    RECT 359.6000 19.6000 360.4000 19.7000 ;
	    RECT 385.2000 19.6000 386.0000 19.7000 ;
	    RECT 423.6000 20.3000 424.4000 20.4000 ;
	    RECT 455.6000 20.3000 456.4000 20.4000 ;
	    RECT 463.6000 20.3000 464.4000 20.4000 ;
	    RECT 423.6000 19.7000 464.4000 20.3000 ;
	    RECT 423.6000 19.6000 424.4000 19.7000 ;
	    RECT 455.6000 19.6000 456.4000 19.7000 ;
	    RECT 463.6000 19.6000 464.4000 19.7000 ;
	    RECT 479.6000 20.3000 480.4000 20.4000 ;
	    RECT 492.4000 20.3000 493.2000 20.4000 ;
	    RECT 479.6000 19.7000 493.2000 20.3000 ;
	    RECT 479.6000 19.6000 480.4000 19.7000 ;
	    RECT 492.4000 19.6000 493.2000 19.7000 ;
	    RECT 44.4000 18.3000 45.2000 18.4000 ;
	    RECT 126.0000 18.3000 126.8000 18.4000 ;
	    RECT 44.4000 17.7000 126.8000 18.3000 ;
	    RECT 44.4000 17.6000 45.2000 17.7000 ;
	    RECT 126.0000 17.6000 126.8000 17.7000 ;
	    RECT 135.6000 18.3000 136.4000 18.4000 ;
	    RECT 137.2000 18.3000 138.0000 18.4000 ;
	    RECT 142.0000 18.3000 142.8000 18.4000 ;
	    RECT 135.6000 17.7000 142.8000 18.3000 ;
	    RECT 135.6000 17.6000 136.4000 17.7000 ;
	    RECT 137.2000 17.6000 138.0000 17.7000 ;
	    RECT 142.0000 17.6000 142.8000 17.7000 ;
	    RECT 166.0000 18.3000 166.8000 18.4000 ;
	    RECT 169.2000 18.3000 170.0000 18.4000 ;
	    RECT 166.0000 17.7000 170.0000 18.3000 ;
	    RECT 166.0000 17.6000 166.8000 17.7000 ;
	    RECT 169.2000 17.6000 170.0000 17.7000 ;
	    RECT 207.6000 18.3000 208.4000 18.4000 ;
	    RECT 236.4000 18.3000 237.2000 18.4000 ;
	    RECT 207.6000 17.7000 237.2000 18.3000 ;
	    RECT 207.6000 17.6000 208.4000 17.7000 ;
	    RECT 236.4000 17.6000 237.2000 17.7000 ;
	    RECT 238.0000 18.3000 238.8000 18.4000 ;
	    RECT 471.6000 18.3000 472.4000 18.4000 ;
	    RECT 481.2000 18.3000 482.0000 18.4000 ;
	    RECT 238.0000 17.7000 482.0000 18.3000 ;
	    RECT 238.0000 17.6000 238.8000 17.7000 ;
	    RECT 471.6000 17.6000 472.4000 17.7000 ;
	    RECT 481.2000 17.6000 482.0000 17.7000 ;
	    RECT 46.0000 16.3000 46.8000 16.4000 ;
	    RECT 114.8000 16.3000 115.6000 16.4000 ;
	    RECT 46.0000 15.7000 115.6000 16.3000 ;
	    RECT 46.0000 15.6000 46.8000 15.7000 ;
	    RECT 114.8000 15.6000 115.6000 15.7000 ;
	    RECT 129.2000 16.3000 130.0000 16.4000 ;
	    RECT 222.0000 16.3000 222.8000 16.4000 ;
	    RECT 129.2000 15.7000 222.8000 16.3000 ;
	    RECT 129.2000 15.6000 130.0000 15.7000 ;
	    RECT 222.0000 15.6000 222.8000 15.7000 ;
	    RECT 234.8000 16.3000 235.6000 16.4000 ;
	    RECT 249.2000 16.3000 250.0000 16.4000 ;
	    RECT 270.0000 16.3000 270.8000 16.4000 ;
	    RECT 234.8000 15.7000 270.8000 16.3000 ;
	    RECT 234.8000 15.6000 235.6000 15.7000 ;
	    RECT 249.2000 15.6000 250.0000 15.7000 ;
	    RECT 270.0000 15.6000 270.8000 15.7000 ;
	    RECT 278.0000 16.3000 278.8000 16.4000 ;
	    RECT 282.8000 16.3000 283.6000 16.4000 ;
	    RECT 278.0000 15.7000 283.6000 16.3000 ;
	    RECT 278.0000 15.6000 278.8000 15.7000 ;
	    RECT 282.8000 15.6000 283.6000 15.7000 ;
	    RECT 286.0000 16.3000 286.8000 16.4000 ;
	    RECT 302.0000 16.3000 302.8000 16.4000 ;
	    RECT 353.2000 16.3000 354.0000 16.4000 ;
	    RECT 286.0000 15.7000 302.8000 16.3000 ;
	    RECT 286.0000 15.6000 286.8000 15.7000 ;
	    RECT 302.0000 15.6000 302.8000 15.7000 ;
	    RECT 305.3000 15.7000 354.0000 16.3000 ;
	    RECT 22.0000 14.3000 22.8000 14.4000 ;
	    RECT 58.8000 14.3000 59.6000 14.4000 ;
	    RECT 81.2000 14.3000 82.0000 14.4000 ;
	    RECT 84.4000 14.3000 85.2000 14.4000 ;
	    RECT 22.0000 13.7000 85.2000 14.3000 ;
	    RECT 22.0000 13.6000 22.8000 13.7000 ;
	    RECT 58.8000 13.6000 59.6000 13.7000 ;
	    RECT 81.2000 13.6000 82.0000 13.7000 ;
	    RECT 84.4000 13.6000 85.2000 13.7000 ;
	    RECT 92.4000 14.3000 93.2000 14.4000 ;
	    RECT 113.2000 14.3000 114.0000 14.4000 ;
	    RECT 92.4000 13.7000 114.0000 14.3000 ;
	    RECT 92.4000 13.6000 93.2000 13.7000 ;
	    RECT 113.2000 13.6000 114.0000 13.7000 ;
	    RECT 118.0000 14.3000 118.8000 14.4000 ;
	    RECT 121.2000 14.3000 122.0000 14.4000 ;
	    RECT 118.0000 13.7000 122.0000 14.3000 ;
	    RECT 118.0000 13.6000 118.8000 13.7000 ;
	    RECT 121.2000 13.6000 122.0000 13.7000 ;
	    RECT 154.8000 14.3000 155.6000 14.4000 ;
	    RECT 158.0000 14.3000 158.8000 14.4000 ;
	    RECT 154.8000 13.7000 158.8000 14.3000 ;
	    RECT 154.8000 13.6000 155.6000 13.7000 ;
	    RECT 158.0000 13.6000 158.8000 13.7000 ;
	    RECT 202.8000 14.3000 203.6000 14.4000 ;
	    RECT 214.0000 14.3000 214.8000 14.4000 ;
	    RECT 202.8000 13.7000 214.8000 14.3000 ;
	    RECT 202.8000 13.6000 203.6000 13.7000 ;
	    RECT 214.0000 13.6000 214.8000 13.7000 ;
	    RECT 233.2000 14.3000 234.0000 14.4000 ;
	    RECT 238.0000 14.3000 238.8000 14.4000 ;
	    RECT 233.2000 13.7000 238.8000 14.3000 ;
	    RECT 270.1000 14.3000 270.7000 15.6000 ;
	    RECT 289.2000 14.3000 290.0000 14.4000 ;
	    RECT 294.0000 14.3000 294.8000 14.4000 ;
	    RECT 270.1000 13.7000 290.0000 14.3000 ;
	    RECT 233.2000 13.6000 234.0000 13.7000 ;
	    RECT 238.0000 13.6000 238.8000 13.7000 ;
	    RECT 289.2000 13.6000 290.0000 13.7000 ;
	    RECT 290.9000 13.7000 294.8000 14.3000 ;
	    RECT 23.6000 12.3000 24.4000 12.4000 ;
	    RECT 41.2000 12.3000 42.0000 12.4000 ;
	    RECT 23.6000 11.7000 42.0000 12.3000 ;
	    RECT 23.6000 11.6000 24.4000 11.7000 ;
	    RECT 41.2000 11.6000 42.0000 11.7000 ;
	    RECT 54.0000 12.3000 54.8000 12.4000 ;
	    RECT 73.2000 12.3000 74.0000 12.4000 ;
	    RECT 54.0000 11.7000 74.0000 12.3000 ;
	    RECT 54.0000 11.6000 54.8000 11.7000 ;
	    RECT 73.2000 11.6000 74.0000 11.7000 ;
	    RECT 76.4000 12.3000 77.2000 12.4000 ;
	    RECT 113.2000 12.3000 114.0000 12.4000 ;
	    RECT 76.4000 11.7000 114.0000 12.3000 ;
	    RECT 76.4000 11.6000 77.2000 11.7000 ;
	    RECT 113.2000 11.6000 114.0000 11.7000 ;
	    RECT 178.8000 12.3000 179.6000 12.4000 ;
	    RECT 180.4000 12.3000 181.2000 12.4000 ;
	    RECT 178.8000 11.7000 181.2000 12.3000 ;
	    RECT 178.8000 11.6000 179.6000 11.7000 ;
	    RECT 180.4000 11.6000 181.2000 11.7000 ;
	    RECT 182.0000 12.3000 182.8000 12.4000 ;
	    RECT 196.4000 12.3000 197.2000 12.4000 ;
	    RECT 182.0000 11.7000 197.2000 12.3000 ;
	    RECT 182.0000 11.6000 182.8000 11.7000 ;
	    RECT 196.4000 11.6000 197.2000 11.7000 ;
	    RECT 212.4000 12.3000 213.2000 12.4000 ;
	    RECT 217.2000 12.3000 218.0000 12.4000 ;
	    RECT 212.4000 11.7000 218.0000 12.3000 ;
	    RECT 212.4000 11.6000 213.2000 11.7000 ;
	    RECT 217.2000 11.6000 218.0000 11.7000 ;
	    RECT 226.8000 12.3000 227.6000 12.4000 ;
	    RECT 231.6000 12.3000 232.4000 12.4000 ;
	    RECT 286.0000 12.3000 286.8000 12.4000 ;
	    RECT 290.9000 12.3000 291.5000 13.7000 ;
	    RECT 294.0000 13.6000 294.8000 13.7000 ;
	    RECT 298.8000 14.3000 299.6000 14.4000 ;
	    RECT 305.3000 14.3000 305.9000 15.7000 ;
	    RECT 353.2000 15.6000 354.0000 15.7000 ;
	    RECT 366.0000 16.3000 366.8000 16.4000 ;
	    RECT 369.2000 16.3000 370.0000 16.4000 ;
	    RECT 366.0000 15.7000 370.0000 16.3000 ;
	    RECT 366.0000 15.6000 366.8000 15.7000 ;
	    RECT 369.2000 15.6000 370.0000 15.7000 ;
	    RECT 401.2000 16.3000 402.0000 16.4000 ;
	    RECT 418.8000 16.3000 419.6000 16.4000 ;
	    RECT 401.2000 15.7000 419.6000 16.3000 ;
	    RECT 401.2000 15.6000 402.0000 15.7000 ;
	    RECT 418.8000 15.6000 419.6000 15.7000 ;
	    RECT 298.8000 13.7000 305.9000 14.3000 ;
	    RECT 318.0000 14.3000 318.8000 14.4000 ;
	    RECT 324.4000 14.3000 325.2000 14.4000 ;
	    RECT 318.0000 13.7000 325.2000 14.3000 ;
	    RECT 298.8000 13.6000 299.6000 13.7000 ;
	    RECT 318.0000 13.6000 318.8000 13.7000 ;
	    RECT 324.4000 13.6000 325.2000 13.7000 ;
	    RECT 329.2000 14.3000 330.0000 14.4000 ;
	    RECT 330.8000 14.3000 331.6000 14.4000 ;
	    RECT 329.2000 13.7000 331.6000 14.3000 ;
	    RECT 329.2000 13.6000 330.0000 13.7000 ;
	    RECT 330.8000 13.6000 331.6000 13.7000 ;
	    RECT 332.4000 14.3000 333.2000 14.4000 ;
	    RECT 337.2000 14.3000 338.0000 14.4000 ;
	    RECT 332.4000 13.7000 338.0000 14.3000 ;
	    RECT 332.4000 13.6000 333.2000 13.7000 ;
	    RECT 337.2000 13.6000 338.0000 13.7000 ;
	    RECT 343.6000 13.6000 344.4000 14.4000 ;
	    RECT 380.4000 14.3000 381.2000 14.4000 ;
	    RECT 423.6000 14.3000 424.4000 14.4000 ;
	    RECT 380.4000 13.7000 424.4000 14.3000 ;
	    RECT 380.4000 13.6000 381.2000 13.7000 ;
	    RECT 423.6000 13.6000 424.4000 13.7000 ;
	    RECT 425.2000 14.3000 426.0000 14.4000 ;
	    RECT 454.0000 14.3000 454.8000 14.4000 ;
	    RECT 425.2000 13.7000 454.8000 14.3000 ;
	    RECT 425.2000 13.6000 426.0000 13.7000 ;
	    RECT 454.0000 13.6000 454.8000 13.7000 ;
	    RECT 460.4000 14.3000 461.2000 14.4000 ;
	    RECT 470.0000 14.3000 470.8000 14.4000 ;
	    RECT 460.4000 13.7000 470.8000 14.3000 ;
	    RECT 460.4000 13.6000 461.2000 13.7000 ;
	    RECT 470.0000 13.6000 470.8000 13.7000 ;
	    RECT 478.0000 14.3000 478.8000 14.4000 ;
	    RECT 487.6000 14.3000 488.4000 14.4000 ;
	    RECT 478.0000 13.7000 488.4000 14.3000 ;
	    RECT 478.0000 13.6000 478.8000 13.7000 ;
	    RECT 487.6000 13.6000 488.4000 13.7000 ;
	    RECT 226.8000 11.7000 285.1000 12.3000 ;
	    RECT 226.8000 11.6000 227.6000 11.7000 ;
	    RECT 231.6000 11.6000 232.4000 11.7000 ;
	    RECT 10.8000 10.3000 11.6000 10.4000 ;
	    RECT 30.0000 10.3000 30.8000 10.4000 ;
	    RECT 10.8000 9.7000 30.8000 10.3000 ;
	    RECT 10.8000 9.6000 11.6000 9.7000 ;
	    RECT 30.0000 9.6000 30.8000 9.7000 ;
	    RECT 33.2000 10.3000 34.0000 10.4000 ;
	    RECT 41.2000 10.3000 42.0000 10.4000 ;
	    RECT 33.2000 9.7000 42.0000 10.3000 ;
	    RECT 33.2000 9.6000 34.0000 9.7000 ;
	    RECT 41.2000 9.6000 42.0000 9.7000 ;
	    RECT 76.4000 10.3000 77.2000 10.4000 ;
	    RECT 100.4000 10.3000 101.2000 10.4000 ;
	    RECT 76.4000 9.7000 101.2000 10.3000 ;
	    RECT 76.4000 9.6000 77.2000 9.7000 ;
	    RECT 100.4000 9.6000 101.2000 9.7000 ;
	    RECT 119.6000 10.3000 120.4000 10.4000 ;
	    RECT 126.0000 10.3000 126.8000 10.4000 ;
	    RECT 119.6000 9.7000 126.8000 10.3000 ;
	    RECT 119.6000 9.6000 120.4000 9.7000 ;
	    RECT 126.0000 9.6000 126.8000 9.7000 ;
	    RECT 201.2000 10.3000 202.0000 10.4000 ;
	    RECT 222.0000 10.3000 222.8000 10.4000 ;
	    RECT 201.2000 9.7000 222.8000 10.3000 ;
	    RECT 201.2000 9.6000 202.0000 9.7000 ;
	    RECT 222.0000 9.6000 222.8000 9.7000 ;
	    RECT 225.2000 10.3000 226.0000 10.4000 ;
	    RECT 234.8000 10.3000 235.6000 10.4000 ;
	    RECT 225.2000 9.7000 235.6000 10.3000 ;
	    RECT 225.2000 9.6000 226.0000 9.7000 ;
	    RECT 234.8000 9.6000 235.6000 9.7000 ;
	    RECT 244.4000 10.3000 245.2000 10.4000 ;
	    RECT 266.8000 10.3000 267.6000 10.4000 ;
	    RECT 279.6000 10.3000 280.4000 10.4000 ;
	    RECT 244.4000 9.7000 280.4000 10.3000 ;
	    RECT 284.5000 10.3000 285.1000 11.7000 ;
	    RECT 286.0000 11.7000 291.5000 12.3000 ;
	    RECT 292.4000 12.3000 293.2000 12.4000 ;
	    RECT 297.2000 12.3000 298.0000 12.4000 ;
	    RECT 298.8000 12.3000 299.6000 12.4000 ;
	    RECT 292.4000 11.7000 299.6000 12.3000 ;
	    RECT 286.0000 11.6000 286.8000 11.7000 ;
	    RECT 292.4000 11.6000 293.2000 11.7000 ;
	    RECT 297.2000 11.6000 298.0000 11.7000 ;
	    RECT 298.8000 11.6000 299.6000 11.7000 ;
	    RECT 300.4000 12.3000 301.2000 12.4000 ;
	    RECT 319.6000 12.3000 320.4000 12.4000 ;
	    RECT 300.4000 11.7000 320.4000 12.3000 ;
	    RECT 300.4000 11.6000 301.2000 11.7000 ;
	    RECT 319.6000 11.6000 320.4000 11.7000 ;
	    RECT 322.8000 12.3000 323.6000 12.4000 ;
	    RECT 324.4000 12.3000 325.2000 12.4000 ;
	    RECT 327.6000 12.3000 328.4000 12.4000 ;
	    RECT 322.8000 11.7000 328.4000 12.3000 ;
	    RECT 322.8000 11.6000 323.6000 11.7000 ;
	    RECT 324.4000 11.6000 325.2000 11.7000 ;
	    RECT 327.6000 11.6000 328.4000 11.7000 ;
	    RECT 330.8000 12.3000 331.6000 12.4000 ;
	    RECT 358.0000 12.3000 358.8000 12.4000 ;
	    RECT 330.8000 11.7000 358.8000 12.3000 ;
	    RECT 330.8000 11.6000 331.6000 11.7000 ;
	    RECT 358.0000 11.6000 358.8000 11.7000 ;
	    RECT 417.2000 12.3000 418.0000 12.4000 ;
	    RECT 422.0000 12.3000 422.8000 12.4000 ;
	    RECT 446.0000 12.3000 446.8000 12.4000 ;
	    RECT 450.8000 12.3000 451.6000 12.4000 ;
	    RECT 417.2000 11.7000 451.6000 12.3000 ;
	    RECT 417.2000 11.6000 418.0000 11.7000 ;
	    RECT 422.0000 11.6000 422.8000 11.7000 ;
	    RECT 446.0000 11.6000 446.8000 11.7000 ;
	    RECT 450.8000 11.6000 451.6000 11.7000 ;
	    RECT 289.2000 10.3000 290.0000 10.4000 ;
	    RECT 322.8000 10.3000 323.6000 10.4000 ;
	    RECT 284.5000 9.7000 288.3000 10.3000 ;
	    RECT 244.4000 9.6000 245.2000 9.7000 ;
	    RECT 266.8000 9.6000 267.6000 9.7000 ;
	    RECT 279.6000 9.6000 280.4000 9.7000 ;
	    RECT 196.4000 8.3000 197.2000 8.4000 ;
	    RECT 241.2000 8.3000 242.0000 8.4000 ;
	    RECT 278.0000 8.3000 278.8000 8.4000 ;
	    RECT 196.4000 7.7000 278.8000 8.3000 ;
	    RECT 196.4000 7.6000 197.2000 7.7000 ;
	    RECT 241.2000 7.6000 242.0000 7.7000 ;
	    RECT 278.0000 7.6000 278.8000 7.7000 ;
	    RECT 282.8000 8.3000 283.6000 8.4000 ;
	    RECT 286.0000 8.3000 286.8000 8.4000 ;
	    RECT 282.8000 7.7000 286.8000 8.3000 ;
	    RECT 287.7000 8.3000 288.3000 9.7000 ;
	    RECT 289.2000 9.7000 323.6000 10.3000 ;
	    RECT 289.2000 9.6000 290.0000 9.7000 ;
	    RECT 322.8000 9.6000 323.6000 9.7000 ;
	    RECT 337.2000 10.3000 338.0000 10.4000 ;
	    RECT 361.2000 10.3000 362.0000 10.4000 ;
	    RECT 388.4000 10.3000 389.2000 10.4000 ;
	    RECT 414.0000 10.3000 414.8000 10.4000 ;
	    RECT 337.2000 9.7000 414.8000 10.3000 ;
	    RECT 337.2000 9.6000 338.0000 9.7000 ;
	    RECT 361.2000 9.6000 362.0000 9.7000 ;
	    RECT 388.4000 9.6000 389.2000 9.7000 ;
	    RECT 414.0000 9.6000 414.8000 9.7000 ;
	    RECT 438.0000 10.3000 438.8000 10.4000 ;
	    RECT 447.6000 10.3000 448.4000 10.4000 ;
	    RECT 438.0000 9.7000 448.4000 10.3000 ;
	    RECT 438.0000 9.6000 438.8000 9.7000 ;
	    RECT 447.6000 9.6000 448.4000 9.7000 ;
	    RECT 300.4000 8.3000 301.2000 8.4000 ;
	    RECT 287.7000 7.7000 301.2000 8.3000 ;
	    RECT 282.8000 7.6000 283.6000 7.7000 ;
	    RECT 286.0000 7.6000 286.8000 7.7000 ;
	    RECT 300.4000 7.6000 301.2000 7.7000 ;
	    RECT 313.2000 8.3000 314.0000 8.4000 ;
	    RECT 314.8000 8.3000 315.6000 8.4000 ;
	    RECT 313.2000 7.7000 315.6000 8.3000 ;
	    RECT 313.2000 7.6000 314.0000 7.7000 ;
	    RECT 314.8000 7.6000 315.6000 7.7000 ;
	    RECT 316.4000 8.3000 317.2000 8.4000 ;
	    RECT 356.4000 8.3000 357.2000 8.4000 ;
	    RECT 425.2000 8.3000 426.0000 8.4000 ;
	    RECT 316.4000 7.7000 426.0000 8.3000 ;
	    RECT 316.4000 7.6000 317.2000 7.7000 ;
	    RECT 356.4000 7.6000 357.2000 7.7000 ;
	    RECT 425.2000 7.6000 426.0000 7.7000 ;
	    RECT 338.8000 6.3000 339.6000 6.4000 ;
	    RECT 362.8000 6.3000 363.6000 6.4000 ;
	    RECT 338.8000 5.7000 363.6000 6.3000 ;
	    RECT 338.8000 5.6000 339.6000 5.7000 ;
	    RECT 362.8000 5.6000 363.6000 5.7000 ;
	    RECT 124.4000 4.3000 125.2000 4.4000 ;
	    RECT 338.8000 4.3000 339.6000 4.4000 ;
	    RECT 462.0000 4.3000 462.8000 4.4000 ;
	    RECT 124.4000 3.7000 339.6000 4.3000 ;
	    RECT 124.4000 3.6000 125.2000 3.7000 ;
	    RECT 338.8000 3.6000 339.6000 3.7000 ;
	    RECT 393.3000 3.7000 462.8000 4.3000 ;
	    RECT 276.4000 2.3000 277.2000 2.4000 ;
	    RECT 332.4000 2.3000 333.2000 2.4000 ;
	    RECT 393.3000 2.3000 393.9000 3.7000 ;
	    RECT 462.0000 3.6000 462.8000 3.7000 ;
	    RECT 276.4000 1.7000 393.9000 2.3000 ;
	    RECT 276.4000 1.6000 277.2000 1.7000 ;
	    RECT 332.4000 1.6000 333.2000 1.7000 ;
         LAYER metal4 ;
	    RECT 61.8000 259.4000 63.0000 296.6000 ;
	    RECT 71.4000 255.4000 72.6000 318.6000 ;
	    RECT 116.2000 307.4000 117.4000 312.6000 ;
	    RECT 74.6000 225.4000 75.8000 256.6000 ;
	    RECT 61.8000 213.4000 63.0000 224.6000 ;
	    RECT 84.2000 221.4000 85.4000 292.6000 ;
	    RECT 87.4000 285.4000 88.6000 294.6000 ;
	    RECT 97.0000 251.4000 98.2000 288.6000 ;
	    RECT 100.2000 267.4000 101.4000 280.6000 ;
	    RECT 93.8000 211.4000 95.0000 228.6000 ;
	    RECT 119.4000 215.4000 120.6000 310.6000 ;
	    RECT 129.0000 287.4000 130.2000 332.6000 ;
	    RECT 138.6000 303.4000 139.8000 312.6000 ;
	    RECT 129.0000 259.4000 130.2000 268.6000 ;
	    RECT 132.2000 261.4000 133.4000 292.6000 ;
	    RECT 148.2000 275.4000 149.4000 312.6000 ;
	    RECT 151.4000 291.4000 152.6000 338.6000 ;
	    RECT 135.4000 211.4000 136.6000 230.6000 ;
	    RECT 141.8000 225.4000 143.0000 266.6000 ;
	    RECT 161.0000 255.4000 162.2000 310.6000 ;
	    RECT 164.2000 293.4000 165.4000 336.6000 ;
	    RECT 218.6000 332.6000 219.8000 334.6000 ;
	    RECT 36.2000 125.4000 37.4000 192.6000 ;
	    RECT 113.0000 181.4000 114.2000 198.6000 ;
	    RECT 145.0000 185.4000 146.2000 242.6000 ;
	    RECT 148.2000 229.4000 149.4000 250.6000 ;
	    RECT 52.2000 53.4000 53.4000 104.6000 ;
	    RECT 74.6000 101.4000 75.8000 136.6000 ;
	    RECT 68.2000 91.4000 69.4000 100.6000 ;
	    RECT 81.0000 87.4000 82.2000 166.6000 ;
	    RECT 87.4000 139.4000 88.6000 144.6000 ;
	    RECT 97.0000 81.4000 98.2000 98.6000 ;
	    RECT 116.2000 91.4000 117.4000 146.6000 ;
	    RECT 119.4000 93.4000 120.6000 124.6000 ;
	    RECT 132.2000 95.4000 133.4000 164.6000 ;
	    RECT 151.4000 163.4000 152.6000 220.6000 ;
	    RECT 154.6000 171.4000 155.8000 222.6000 ;
	    RECT 141.8000 115.4000 143.0000 128.6000 ;
	    RECT 135.4000 103.4000 136.6000 112.6000 ;
	    RECT 100.2000 67.4000 101.4000 86.6000 ;
	    RECT 119.4000 57.4000 120.6000 78.6000 ;
	    RECT 122.6000 73.4000 123.8000 92.6000 ;
	    RECT 129.0000 29.4000 130.2000 72.6000 ;
	    RECT 145.0000 69.4000 146.2000 136.6000 ;
	    RECT 154.6000 131.4000 155.8000 138.6000 ;
	    RECT 154.6000 105.4000 155.8000 112.6000 ;
	    RECT 157.8000 111.4000 159.0000 168.6000 ;
	    RECT 161.0000 147.4000 162.2000 250.6000 ;
	    RECT 164.2000 247.4000 165.4000 290.6000 ;
	    RECT 170.6000 289.4000 171.8000 298.6000 ;
	    RECT 170.6000 227.4000 171.8000 280.6000 ;
	    RECT 186.6000 277.4000 187.8000 294.6000 ;
	    RECT 183.4000 265.4000 184.6000 276.6000 ;
	    RECT 177.0000 229.4000 178.2000 262.6000 ;
	    RECT 186.6000 251.4000 187.8000 272.6000 ;
	    RECT 189.8000 269.4000 191.0000 332.6000 ;
	    RECT 215.4000 331.4000 219.8000 332.6000 ;
	    RECT 263.4000 331.4000 264.6000 336.6000 ;
	    RECT 215.4000 328.6000 216.6000 331.4000 ;
	    RECT 212.2000 327.4000 216.6000 328.6000 ;
	    RECT 193.0000 249.4000 194.2000 280.6000 ;
	    RECT 199.4000 279.4000 200.6000 310.6000 ;
	    RECT 202.6000 293.4000 203.8000 308.6000 ;
	    RECT 202.6000 265.4000 203.8000 288.6000 ;
	    RECT 205.8000 269.4000 207.0000 310.6000 ;
	    RECT 215.4000 293.4000 216.6000 320.6000 ;
	    RECT 228.2000 307.4000 229.4000 322.6000 ;
	    RECT 263.4000 305.4000 264.6000 312.6000 ;
	    RECT 164.2000 205.4000 165.4000 218.6000 ;
	    RECT 164.2000 131.4000 165.4000 150.6000 ;
	    RECT 170.6000 149.4000 171.8000 182.6000 ;
	    RECT 173.8000 159.4000 175.0000 206.6000 ;
	    RECT 173.8000 141.4000 175.0000 156.6000 ;
	    RECT 177.0000 137.4000 178.2000 224.6000 ;
	    RECT 186.6000 219.4000 187.8000 248.6000 ;
	    RECT 189.8000 227.4000 191.0000 246.6000 ;
	    RECT 196.2000 245.4000 197.4000 252.6000 ;
	    RECT 183.4000 208.6000 184.6000 216.6000 ;
	    RECT 193.0000 208.6000 194.2000 216.6000 ;
	    RECT 183.4000 207.4000 186.2000 208.6000 ;
	    RECT 188.2000 207.4000 194.2000 208.6000 ;
	    RECT 180.2000 145.4000 181.4000 184.6000 ;
	    RECT 183.4000 105.4000 184.6000 188.6000 ;
	    RECT 193.0000 171.4000 194.2000 202.6000 ;
	    RECT 196.2000 185.4000 197.4000 230.6000 ;
	    RECT 199.4000 209.4000 200.6000 246.6000 ;
	    RECT 202.6000 241.4000 203.8000 246.6000 ;
	    RECT 202.6000 212.6000 203.8000 216.6000 ;
	    RECT 205.8000 215.4000 207.0000 264.6000 ;
	    RECT 209.0000 239.4000 210.2000 264.6000 ;
	    RECT 212.2000 251.4000 213.4000 278.6000 ;
	    RECT 215.4000 265.4000 216.6000 272.6000 ;
	    RECT 218.6000 249.4000 219.8000 286.6000 ;
	    RECT 215.4000 235.4000 219.8000 236.6000 ;
	    RECT 209.0000 212.6000 210.2000 218.6000 ;
	    RECT 202.6000 211.4000 210.2000 212.6000 ;
	    RECT 199.4000 187.4000 200.6000 196.6000 ;
	    RECT 199.4000 149.4000 200.6000 180.6000 ;
	    RECT 205.8000 167.4000 207.0000 200.6000 ;
	    RECT 212.2000 197.4000 213.4000 230.6000 ;
	    RECT 218.6000 219.4000 219.8000 235.4000 ;
	    RECT 221.8000 213.4000 223.0000 294.6000 ;
	    RECT 225.0000 217.4000 226.2000 224.6000 ;
	    RECT 228.2000 215.4000 229.4000 270.6000 ;
	    RECT 234.6000 265.4000 235.8000 272.6000 ;
	    RECT 244.2000 269.4000 245.4000 290.6000 ;
	    RECT 250.6000 277.4000 251.8000 286.6000 ;
	    RECT 234.6000 225.4000 235.8000 258.6000 ;
	    RECT 244.2000 225.4000 245.4000 244.6000 ;
	    RECT 250.6000 235.4000 251.8000 264.6000 ;
	    RECT 266.6000 259.4000 267.8000 296.6000 ;
	    RECT 266.6000 251.4000 269.4000 252.6000 ;
	    RECT 266.6000 244.6000 267.8000 251.4000 ;
	    RECT 263.4000 243.4000 267.8000 244.6000 ;
	    RECT 231.4000 211.4000 232.6000 220.6000 ;
	    RECT 202.6000 143.4000 203.8000 160.6000 ;
	    RECT 205.8000 108.6000 207.0000 156.6000 ;
	    RECT 209.0000 151.4000 210.2000 190.6000 ;
	    RECT 221.8000 185.4000 223.0000 200.6000 ;
	    RECT 215.4000 175.4000 216.6000 184.6000 ;
	    RECT 161.0000 87.4000 162.2000 92.6000 ;
	    RECT 173.8000 83.4000 175.0000 92.6000 ;
	    RECT 148.2000 37.4000 149.4000 68.6000 ;
	    RECT 154.6000 63.4000 155.8000 68.6000 ;
	    RECT 157.8000 13.4000 159.0000 64.6000 ;
	    RECT 167.4000 59.4000 168.6000 68.6000 ;
	    RECT 177.0000 63.4000 178.2000 84.6000 ;
	    RECT 173.8000 47.4000 175.0000 56.6000 ;
	    RECT 193.0000 55.4000 194.2000 90.6000 ;
	    RECT 196.2000 55.4000 197.4000 108.6000 ;
	    RECT 202.6000 107.4000 207.0000 108.6000 ;
	    RECT 202.6000 91.4000 203.8000 107.4000 ;
	    RECT 205.8000 79.4000 207.0000 104.6000 ;
	    RECT 209.0000 69.4000 210.2000 148.6000 ;
	    RECT 215.4000 131.4000 216.6000 150.6000 ;
	    RECT 212.2000 69.4000 213.4000 104.6000 ;
	    RECT 215.4000 87.4000 216.6000 114.6000 ;
	    RECT 218.6000 107.4000 219.8000 164.6000 ;
	    RECT 221.8000 121.4000 223.0000 160.6000 ;
	    RECT 225.0000 133.4000 226.2000 198.6000 ;
	    RECT 228.2000 169.4000 229.4000 206.6000 ;
	    RECT 234.6000 171.4000 235.8000 214.6000 ;
	    RECT 250.6000 213.4000 251.8000 224.6000 ;
	    RECT 263.4000 219.4000 264.6000 230.6000 ;
	    RECT 237.8000 165.4000 239.0000 210.6000 ;
	    RECT 241.0000 191.4000 242.2000 208.6000 ;
	    RECT 244.2000 199.4000 245.4000 210.6000 ;
	    RECT 266.6000 205.4000 267.8000 232.6000 ;
	    RECT 269.8000 197.4000 271.0000 212.6000 ;
	    RECT 273.0000 211.4000 274.2000 332.6000 ;
	    RECT 298.6000 329.4000 299.8000 334.6000 ;
	    RECT 289.0000 289.4000 290.2000 324.6000 ;
	    RECT 276.2000 283.4000 277.4000 288.6000 ;
	    RECT 279.4000 275.4000 280.6000 288.6000 ;
	    RECT 292.2000 271.4000 293.4000 318.6000 ;
	    RECT 298.6000 263.4000 299.8000 310.6000 ;
	    RECT 308.2000 285.4000 309.4000 296.6000 ;
	    RECT 327.4000 271.4000 328.6000 284.6000 ;
	    RECT 305.0000 264.6000 306.2000 266.6000 ;
	    RECT 305.0000 263.4000 315.8000 264.6000 ;
	    RECT 276.2000 195.4000 277.4000 260.6000 ;
	    RECT 301.8000 241.4000 303.0000 260.6000 ;
	    RECT 282.6000 227.4000 283.8000 232.6000 ;
	    RECT 228.2000 139.4000 229.4000 156.6000 ;
	    RECT 234.6000 111.4000 235.8000 146.6000 ;
	    RECT 237.8000 127.4000 239.0000 156.6000 ;
	    RECT 241.0000 137.4000 242.2000 186.6000 ;
	    RECT 244.2000 129.4000 245.4000 160.6000 ;
	    RECT 263.4000 133.4000 264.6000 162.6000 ;
	    RECT 266.6000 141.4000 267.8000 152.6000 ;
	    RECT 279.4000 149.4000 280.6000 186.6000 ;
	    RECT 180.2000 11.4000 181.4000 30.6000 ;
	    RECT 209.0000 19.4000 210.2000 62.6000 ;
	    RECT 218.6000 47.4000 219.8000 68.6000 ;
	    RECT 234.6000 61.4000 235.8000 78.6000 ;
	    RECT 237.8000 13.4000 239.0000 76.6000 ;
	    RECT 241.0000 57.4000 242.2000 98.6000 ;
	    RECT 244.2000 69.4000 245.4000 124.6000 ;
	    RECT 282.6000 121.4000 283.8000 200.6000 ;
	    RECT 285.8000 179.4000 287.0000 224.6000 ;
	    RECT 289.0000 221.4000 290.2000 240.6000 ;
	    RECT 308.2000 201.4000 309.4000 220.6000 ;
	    RECT 333.8000 219.4000 335.0000 286.6000 ;
	    RECT 353.0000 268.6000 354.2000 270.6000 ;
	    RECT 372.2000 269.4000 373.4000 314.6000 ;
	    RECT 353.0000 267.4000 357.4000 268.6000 ;
	    RECT 356.2000 263.4000 357.4000 267.4000 ;
	    RECT 285.8000 121.4000 287.0000 166.6000 ;
	    RECT 295.4000 149.4000 296.6000 182.6000 ;
	    RECT 247.4000 91.4000 248.6000 102.6000 ;
	    RECT 263.4000 91.4000 264.6000 106.6000 ;
	    RECT 276.2000 93.4000 277.4000 114.6000 ;
	    RECT 282.6000 85.4000 283.8000 100.6000 ;
	    RECT 247.4000 57.4000 248.6000 82.6000 ;
	    RECT 263.4000 55.4000 264.6000 76.6000 ;
	    RECT 266.6000 43.4000 267.8000 80.6000 ;
	    RECT 269.8000 45.4000 271.0000 68.6000 ;
	    RECT 273.0000 29.4000 274.2000 58.6000 ;
	    RECT 276.2000 51.4000 277.4000 80.6000 ;
	    RECT 276.2000 31.4000 277.4000 48.6000 ;
	    RECT 282.6000 15.4000 283.8000 54.6000 ;
	    RECT 285.8000 21.4000 287.0000 100.6000 ;
	    RECT 289.0000 61.4000 290.2000 112.6000 ;
	    RECT 292.2000 93.4000 293.4000 136.6000 ;
	    RECT 295.4000 119.4000 296.6000 136.6000 ;
	    RECT 301.8000 129.4000 303.0000 140.6000 ;
	    RECT 311.4000 139.4000 312.6000 152.6000 ;
	    RECT 317.8000 143.4000 319.0000 162.6000 ;
	    RECT 308.2000 133.4000 309.4000 138.6000 ;
	    RECT 330.6000 131.4000 331.8000 194.6000 ;
	    RECT 343.4000 193.4000 344.6000 252.6000 ;
	    RECT 346.6000 213.4000 347.8000 240.6000 ;
	    RECT 298.6000 103.4000 299.8000 108.6000 ;
	    RECT 317.8000 95.4000 319.0000 126.6000 ;
	    RECT 292.2000 71.4000 293.4000 76.6000 ;
	    RECT 295.4000 55.4000 296.6000 94.6000 ;
	    RECT 289.0000 9.4000 290.2000 32.6000 ;
	    RECT 298.6000 11.4000 299.8000 44.6000 ;
	    RECT 308.2000 31.4000 309.4000 82.6000 ;
	    RECT 321.0000 67.4000 322.2000 120.6000 ;
	    RECT 343.4000 109.4000 344.6000 186.6000 ;
	    RECT 356.2000 167.4000 357.4000 206.6000 ;
	    RECT 346.6000 107.4000 347.8000 158.6000 ;
	    RECT 362.6000 147.4000 363.8000 254.6000 ;
	    RECT 349.8000 121.4000 351.0000 126.6000 ;
	    RECT 333.8000 56.6000 335.0000 58.6000 ;
	    RECT 311.4000 21.4000 312.6000 32.6000 ;
	    RECT 314.6000 21.4000 315.8000 56.6000 ;
	    RECT 333.8000 55.4000 338.2000 56.6000 ;
	    RECT 337.0000 53.4000 338.2000 55.4000 ;
	    RECT 317.8000 27.4000 319.0000 52.6000 ;
	    RECT 317.8000 12.6000 319.0000 14.6000 ;
	    RECT 314.6000 11.4000 319.0000 12.6000 ;
	    RECT 324.2000 11.4000 325.4000 48.6000 ;
	    RECT 330.6000 13.4000 331.8000 50.6000 ;
	    RECT 333.8000 21.4000 335.0000 28.6000 ;
	    RECT 314.6000 7.4000 315.8000 11.4000 ;
	    RECT 337.0000 9.4000 338.2000 26.6000 ;
	    RECT 340.2000 23.4000 341.4000 28.6000 ;
	    RECT 343.4000 13.4000 344.6000 56.6000 ;
	    RECT 353.0000 15.4000 354.2000 100.6000 ;
	    RECT 359.4000 93.4000 360.6000 130.6000 ;
	    RECT 381.8000 83.4000 383.0000 260.6000 ;
	    RECT 391.4000 229.4000 392.6000 332.6000 ;
	    RECT 417.0000 271.4000 418.2000 298.6000 ;
	    RECT 429.8000 257.4000 431.0000 298.6000 ;
	    RECT 420.2000 249.4000 421.4000 256.6000 ;
	    RECT 413.8000 233.4000 415.0000 238.6000 ;
	    RECT 385.0000 143.4000 386.2000 194.6000 ;
	    RECT 388.2000 51.4000 389.4000 86.6000 ;
	    RECT 394.6000 69.4000 395.8000 210.6000 ;
	    RECT 413.8000 141.4000 415.0000 214.6000 ;
	    RECT 449.0000 213.4000 450.2000 262.6000 ;
	    RECT 474.6000 229.4000 475.8000 272.6000 ;
	    RECT 452.2000 165.4000 453.4000 184.6000 ;
	    RECT 477.8000 173.4000 479.0000 268.6000 ;
	    RECT 481.0000 243.4000 482.2000 254.6000 ;
	    RECT 487.4000 243.4000 488.6000 296.6000 ;
	    RECT 493.8000 175.4000 495.0000 190.6000 ;
	    RECT 397.8000 67.4000 399.0000 134.6000 ;
	    RECT 503.4000 133.4000 504.6000 260.6000 ;
	    RECT 506.6000 253.4000 507.8000 286.6000 ;
	    RECT 506.6000 193.4000 507.8000 250.6000 ;
	    RECT 506.6000 169.4000 507.8000 188.6000 ;
	    RECT 429.8000 69.4000 431.0000 130.6000 ;
	    RECT 455.4000 71.4000 456.6000 106.6000 ;
	    RECT 461.8000 61.4000 463.0000 100.6000 ;
	    RECT 465.0000 79.4000 466.2000 114.6000 ;
	    RECT 487.4000 51.4000 488.6000 124.6000 ;
	    RECT 506.6000 75.4000 507.8000 136.6000 ;
	    RECT 509.8000 123.4000 511.0000 290.6000 ;
   END
END internal_register
