magic
tech scmos
magscale 1 2
timestamp 1588175369
<< metal1 >>
rect 1914 1814 1926 1816
rect 1899 1806 1901 1814
rect 1909 1806 1911 1814
rect 1919 1806 1921 1814
rect 1929 1806 1931 1814
rect 1939 1806 1941 1814
rect 1914 1804 1926 1806
rect 1901 1777 1964 1783
rect 1805 1757 1843 1763
rect 2068 1757 2083 1763
rect 2557 1737 2604 1743
rect 1741 1717 1763 1723
rect 2013 1717 2028 1723
rect 682 1614 694 1616
rect 667 1606 669 1614
rect 677 1606 679 1614
rect 687 1606 689 1614
rect 697 1606 699 1614
rect 707 1606 709 1614
rect 682 1604 694 1606
rect 532 1576 534 1584
rect 365 1517 380 1523
rect 45 1497 60 1503
rect 644 1497 739 1503
rect 749 1497 771 1503
rect 1565 1497 1603 1503
rect 1748 1497 1763 1503
rect 1956 1497 2019 1503
rect 2148 1497 2163 1503
rect 493 1477 515 1483
rect 1588 1477 1603 1483
rect 2221 1477 2236 1483
rect 637 1457 700 1463
rect 781 1457 796 1463
rect 1517 1457 1555 1463
rect 1914 1414 1926 1416
rect 1899 1406 1901 1414
rect 1909 1406 1911 1414
rect 1919 1406 1921 1414
rect 1929 1406 1931 1414
rect 1939 1406 1941 1414
rect 1914 1404 1926 1406
rect 77 1337 115 1343
rect 1613 1343 1619 1363
rect 1677 1357 1699 1363
rect 2493 1357 2508 1363
rect 1508 1337 1523 1343
rect 1613 1337 1628 1343
rect 1748 1337 1756 1343
rect 1764 1337 1842 1343
rect 45 1317 60 1323
rect 1485 1317 1523 1323
rect 2494 1317 2531 1323
rect 2557 1277 2604 1283
rect 682 1214 694 1216
rect 667 1206 669 1214
rect 677 1206 679 1214
rect 687 1206 689 1214
rect 697 1206 699 1214
rect 707 1206 709 1214
rect 682 1204 694 1206
rect 500 1176 502 1184
rect 954 1176 956 1184
rect 2548 1176 2550 1184
rect 778 1136 780 1144
rect 157 1117 172 1123
rect 205 1103 211 1116
rect 205 1097 243 1103
rect 365 1097 396 1103
rect 532 1097 563 1103
rect 644 1097 659 1103
rect 781 1097 819 1103
rect 884 1097 899 1103
rect 1660 1103 1668 1104
rect 1629 1097 1668 1103
rect 1757 1097 1772 1103
rect 1876 1097 1955 1103
rect 2477 1097 2492 1103
rect 301 1077 339 1083
rect 1588 1077 1603 1083
rect 1981 1077 1996 1083
rect 2420 1077 2435 1083
rect 2445 1077 2483 1083
rect 36 1056 44 1064
rect 77 1057 92 1063
rect 621 1057 643 1063
rect 2397 1057 2419 1063
rect 452 1036 454 1044
rect 1914 1014 1926 1016
rect 1899 1006 1901 1014
rect 1909 1006 1911 1014
rect 1919 1006 1921 1014
rect 1929 1006 1931 1014
rect 1939 1006 1941 1014
rect 1914 1004 1926 1006
rect 637 957 739 963
rect 1709 957 1731 963
rect 157 923 163 943
rect 877 937 892 943
rect 1640 937 1660 943
rect 1789 943 1795 963
rect 1780 937 1795 943
rect 1853 943 1859 963
rect 1917 957 1980 963
rect 1828 937 1843 943
rect 1853 937 1868 943
rect 2052 937 2067 943
rect 2589 937 2604 943
rect 140 917 163 923
rect 173 917 188 923
rect 140 912 148 917
rect 285 917 300 923
rect 1588 917 1604 923
rect 1596 912 1604 917
rect 1821 917 1852 923
rect 1956 917 2003 923
rect 2452 917 2467 923
rect 2493 923 2499 936
rect 2493 917 2515 923
rect 61 897 76 903
rect 132 897 147 903
rect 797 897 835 903
rect 1917 897 1964 903
rect 2436 897 2451 903
rect 109 877 140 883
rect 900 877 915 883
rect 1812 836 1814 844
rect 682 814 694 816
rect 667 806 669 814
rect 677 806 679 814
rect 687 806 689 814
rect 697 806 699 814
rect 707 806 709 814
rect 682 804 694 806
rect 746 776 748 784
rect 1594 776 1596 784
rect 1549 737 1572 743
rect 1976 736 1980 744
rect 237 703 243 723
rect 676 717 700 723
rect 205 697 243 703
rect 381 697 467 703
rect 509 697 540 703
rect 125 677 163 683
rect 125 657 131 677
rect 301 683 307 696
rect 285 677 307 683
rect 509 677 515 697
rect 637 697 684 703
rect 1037 697 1075 703
rect 1085 697 1100 703
rect 1597 697 1628 703
rect 573 677 588 683
rect 781 683 787 696
rect 765 677 787 683
rect 820 677 835 683
rect 925 677 940 683
rect 1357 677 1372 683
rect 1661 683 1667 703
rect 2036 697 2051 703
rect 2132 697 2163 703
rect 1661 677 1692 683
rect 1876 677 1923 683
rect 2173 683 2179 703
rect 2077 677 2115 683
rect 2173 677 2204 683
rect 1645 657 1660 663
rect 954 636 956 644
rect 1914 614 1926 616
rect 1899 606 1901 614
rect 1909 606 1911 614
rect 1919 606 1921 614
rect 1929 606 1931 614
rect 1939 606 1941 614
rect 1914 604 1926 606
rect 2116 576 2120 584
rect 1053 557 1068 563
rect 1140 557 1171 563
rect 1549 557 1571 563
rect 781 537 812 543
rect 845 537 892 543
rect 964 537 979 543
rect 1060 537 1091 543
rect 2189 543 2195 556
rect 2173 537 2195 543
rect 205 517 259 523
rect 852 517 867 523
rect 989 517 1004 523
rect 964 477 995 483
rect 1082 436 1084 444
rect 1988 437 2051 443
rect 682 414 694 416
rect 667 406 669 414
rect 677 406 679 414
rect 687 406 689 414
rect 697 406 699 414
rect 707 406 709 414
rect 682 404 694 406
rect 1908 377 1971 383
rect 45 297 82 303
rect 493 297 547 303
rect 676 297 755 303
rect 1028 297 1043 303
rect 1053 297 1068 303
rect 820 277 883 283
rect 909 277 963 283
rect 1021 277 1059 283
rect 828 276 836 277
rect 429 257 444 263
rect 973 257 1004 263
rect 884 236 886 244
rect 1914 214 1926 216
rect 1899 206 1901 214
rect 1909 206 1911 214
rect 1919 206 1921 214
rect 1929 206 1931 214
rect 1939 206 1941 214
rect 1914 204 1926 206
rect 1844 137 1859 143
rect 2477 137 2492 143
rect 525 117 540 123
rect 909 117 946 123
rect 1309 117 1348 123
rect 1340 116 1348 117
rect 1726 117 1763 123
rect 1821 117 1859 123
rect 1917 117 1964 123
rect 2493 117 2515 123
rect 2532 117 2547 123
rect 396 112 404 116
rect 381 97 403 103
rect 653 37 716 43
rect 682 14 694 16
rect 667 6 669 14
rect 677 6 679 14
rect 687 6 689 14
rect 697 6 699 14
rect 707 6 709 14
rect 682 4 694 6
<< m2contact >>
rect 1891 1806 1899 1814
rect 1901 1806 1909 1814
rect 1911 1806 1919 1814
rect 1921 1806 1929 1814
rect 1931 1806 1939 1814
rect 1941 1806 1949 1814
rect 1660 1776 1668 1784
rect 1708 1776 1716 1784
rect 1788 1776 1796 1784
rect 1964 1776 1972 1784
rect 1980 1776 1988 1784
rect 188 1756 196 1764
rect 540 1756 548 1764
rect 1100 1756 1108 1764
rect 1436 1756 1444 1764
rect 1724 1756 1732 1764
rect 1852 1756 1860 1764
rect 2028 1756 2036 1764
rect 2060 1756 2068 1764
rect 2236 1756 2244 1764
rect 2476 1756 2484 1764
rect 2508 1756 2516 1764
rect 220 1736 228 1744
rect 572 1736 580 1744
rect 780 1736 788 1744
rect 908 1736 916 1744
rect 1132 1736 1140 1744
rect 1404 1736 1412 1744
rect 1598 1736 1606 1744
rect 1772 1736 1780 1744
rect 2268 1736 2276 1744
rect 2604 1736 2612 1744
rect 316 1716 324 1724
rect 460 1716 468 1724
rect 1132 1716 1140 1724
rect 1324 1716 1332 1724
rect 1628 1716 1636 1724
rect 1676 1716 1684 1724
rect 1820 1716 1828 1724
rect 1868 1716 1876 1724
rect 2028 1716 2036 1724
rect 2268 1716 2276 1724
rect 2412 1716 2420 1724
rect 2524 1716 2532 1724
rect 316 1696 324 1704
rect 636 1700 644 1708
rect 1196 1700 1204 1708
rect 1308 1696 1316 1704
rect 2364 1696 2372 1704
rect 2444 1676 2452 1684
rect 28 1636 36 1644
rect 316 1636 324 1644
rect 380 1636 388 1644
rect 636 1636 644 1644
rect 940 1636 948 1644
rect 1196 1636 1204 1644
rect 1308 1636 1316 1644
rect 2044 1636 2052 1644
rect 2364 1636 2372 1644
rect 2460 1636 2468 1644
rect 2492 1636 2500 1644
rect 659 1606 667 1614
rect 669 1606 677 1614
rect 679 1606 687 1614
rect 689 1606 697 1614
rect 699 1606 707 1614
rect 709 1606 717 1614
rect 524 1576 532 1584
rect 572 1576 580 1584
rect 1228 1576 1236 1584
rect 1516 1576 1524 1584
rect 1708 1576 1716 1584
rect 1788 1576 1796 1584
rect 2108 1576 2116 1584
rect 2572 1576 2580 1584
rect 268 1556 276 1564
rect 1068 1558 1076 1566
rect 2316 1558 2324 1566
rect 332 1512 340 1520
rect 380 1516 388 1524
rect 556 1516 564 1524
rect 620 1516 628 1524
rect 1068 1512 1076 1520
rect 1228 1516 1236 1524
rect 2316 1512 2324 1520
rect 60 1496 68 1504
rect 268 1496 276 1504
rect 412 1496 420 1504
rect 444 1496 452 1504
rect 524 1496 532 1504
rect 604 1496 612 1504
rect 636 1496 644 1504
rect 892 1496 900 1504
rect 1100 1496 1108 1504
rect 1180 1496 1188 1504
rect 1260 1496 1268 1504
rect 1324 1496 1332 1504
rect 1644 1496 1652 1504
rect 1660 1496 1668 1504
rect 1676 1496 1684 1504
rect 1740 1496 1748 1504
rect 1948 1496 1956 1504
rect 2060 1496 2068 1504
rect 2076 1496 2084 1504
rect 2124 1496 2132 1504
rect 2140 1496 2148 1504
rect 2172 1496 2180 1504
rect 2220 1496 2228 1504
rect 2268 1496 2276 1504
rect 2284 1496 2292 1504
rect 12 1476 20 1484
rect 268 1476 276 1484
rect 460 1476 468 1484
rect 1004 1476 1012 1484
rect 1148 1476 1156 1484
rect 1324 1476 1332 1484
rect 1580 1476 1588 1484
rect 1804 1476 1812 1484
rect 2236 1476 2244 1484
rect 2380 1476 2388 1484
rect 236 1456 244 1464
rect 476 1456 484 1464
rect 700 1456 708 1464
rect 716 1456 724 1464
rect 796 1456 804 1464
rect 812 1456 820 1464
rect 972 1456 980 1464
rect 1356 1456 1364 1464
rect 1740 1456 1748 1464
rect 2412 1456 2420 1464
rect 76 1436 84 1444
rect 1724 1436 1732 1444
rect 1916 1436 1924 1444
rect 2044 1436 2052 1444
rect 1891 1406 1899 1414
rect 1901 1406 1909 1414
rect 1911 1406 1919 1414
rect 1921 1406 1929 1414
rect 1931 1406 1939 1414
rect 1941 1406 1949 1414
rect 124 1376 132 1384
rect 60 1356 68 1364
rect 140 1356 148 1364
rect 316 1356 324 1364
rect 732 1356 740 1364
rect 1228 1356 1236 1364
rect 1388 1356 1396 1364
rect 1468 1356 1476 1364
rect 284 1336 292 1344
rect 700 1336 708 1344
rect 924 1336 932 1344
rect 1052 1336 1060 1344
rect 1196 1336 1204 1344
rect 1500 1336 1508 1344
rect 1996 1356 2004 1364
rect 2332 1356 2340 1364
rect 2508 1356 2516 1364
rect 1628 1336 1636 1344
rect 1708 1336 1716 1344
rect 1724 1336 1732 1344
rect 1740 1336 1748 1344
rect 1756 1336 1764 1344
rect 2028 1336 2036 1344
rect 2300 1336 2308 1344
rect 60 1316 68 1324
rect 92 1316 100 1324
rect 396 1316 404 1324
rect 588 1316 596 1324
rect 812 1316 820 1324
rect 1196 1316 1204 1324
rect 1308 1316 1316 1324
rect 1452 1316 1460 1324
rect 1564 1316 1572 1324
rect 1580 1316 1588 1324
rect 1596 1316 1604 1324
rect 1644 1316 1652 1324
rect 1740 1316 1748 1324
rect 2108 1316 2116 1324
rect 2204 1316 2212 1324
rect 188 1296 196 1304
rect 636 1300 644 1308
rect 1132 1300 1140 1308
rect 1676 1296 1684 1304
rect 2092 1300 2100 1308
rect 2236 1300 2244 1308
rect 12 1276 20 1284
rect 2604 1276 2612 1284
rect 1132 1254 1140 1262
rect 2236 1254 2244 1262
rect 188 1236 196 1244
rect 476 1236 484 1244
rect 636 1236 644 1244
rect 892 1236 900 1244
rect 1420 1236 1428 1244
rect 2092 1236 2100 1244
rect 659 1206 667 1214
rect 669 1206 677 1214
rect 679 1206 687 1214
rect 689 1206 697 1214
rect 699 1206 707 1214
rect 709 1206 717 1214
rect 492 1176 500 1184
rect 956 1176 964 1184
rect 1052 1176 1060 1184
rect 1436 1176 1444 1184
rect 2012 1176 2020 1184
rect 2540 1176 2548 1184
rect 2268 1158 2276 1166
rect 268 1136 276 1144
rect 780 1136 788 1144
rect 988 1136 996 1144
rect 1068 1136 1076 1144
rect 1148 1136 1156 1144
rect 1516 1136 1524 1144
rect 44 1116 52 1124
rect 172 1116 180 1124
rect 204 1116 212 1124
rect 380 1116 388 1124
rect 460 1116 468 1124
rect 524 1116 532 1124
rect 540 1116 548 1124
rect 748 1116 756 1124
rect 924 1116 932 1124
rect 1036 1116 1044 1124
rect 1100 1116 1108 1124
rect 1436 1116 1444 1124
rect 1580 1116 1588 1124
rect 1724 1116 1732 1124
rect 92 1096 100 1104
rect 2268 1112 2276 1120
rect 2396 1116 2404 1124
rect 284 1096 292 1104
rect 348 1096 356 1104
rect 396 1096 404 1104
rect 492 1096 500 1104
rect 524 1096 532 1104
rect 572 1096 580 1104
rect 636 1096 644 1104
rect 668 1096 676 1104
rect 876 1096 884 1104
rect 908 1096 916 1104
rect 956 1096 964 1104
rect 1020 1096 1028 1104
rect 1052 1096 1060 1104
rect 1420 1096 1428 1104
rect 1484 1096 1492 1104
rect 1532 1096 1540 1104
rect 1692 1096 1700 1104
rect 1772 1096 1780 1104
rect 1820 1096 1828 1104
rect 1868 1096 1876 1104
rect 2204 1096 2212 1104
rect 2316 1096 2324 1104
rect 2364 1096 2372 1104
rect 2460 1096 2468 1104
rect 2492 1096 2500 1104
rect 2508 1096 2516 1104
rect 2524 1096 2532 1104
rect 2572 1096 2580 1104
rect 12 1076 20 1084
rect 172 1076 180 1084
rect 220 1076 228 1084
rect 412 1076 420 1084
rect 428 1076 436 1084
rect 476 1076 484 1084
rect 588 1076 596 1084
rect 796 1076 804 1084
rect 844 1080 852 1088
rect 860 1076 868 1084
rect 972 1076 980 1084
rect 1340 1076 1348 1084
rect 1548 1076 1556 1084
rect 1580 1076 1588 1084
rect 1644 1076 1652 1084
rect 1772 1076 1780 1084
rect 1788 1076 1796 1084
rect 1996 1076 2004 1084
rect 2204 1076 2212 1084
rect 2348 1076 2356 1084
rect 2412 1076 2420 1084
rect 44 1056 52 1064
rect 60 1056 68 1064
rect 92 1056 100 1064
rect 108 1056 116 1064
rect 140 1056 148 1064
rect 316 1056 324 1064
rect 396 1056 404 1064
rect 604 1056 612 1064
rect 876 1056 884 1064
rect 1116 1056 1124 1064
rect 1308 1056 1316 1064
rect 1580 1056 1588 1064
rect 2172 1056 2180 1064
rect 2492 1056 2500 1064
rect 124 1036 132 1044
rect 204 1036 212 1044
rect 268 1036 276 1044
rect 444 1036 452 1044
rect 1724 1036 1732 1044
rect 1836 1036 1844 1044
rect 1891 1006 1899 1014
rect 1901 1006 1909 1014
rect 1911 1006 1919 1014
rect 1921 1006 1929 1014
rect 1931 1006 1939 1014
rect 1941 1006 1949 1014
rect 636 976 644 984
rect 2412 976 2420 984
rect 76 956 84 964
rect 476 956 484 964
rect 1068 956 1076 964
rect 1404 956 1412 964
rect 1692 956 1700 964
rect 44 916 52 924
rect 124 916 132 924
rect 300 936 308 944
rect 444 936 452 944
rect 812 936 820 944
rect 844 936 852 944
rect 892 936 900 944
rect 1100 936 1108 944
rect 1372 936 1380 944
rect 1660 936 1668 944
rect 1676 936 1684 944
rect 1772 936 1780 944
rect 1820 936 1828 944
rect 1980 956 1988 964
rect 2044 956 2052 964
rect 2076 956 2084 964
rect 2252 956 2260 964
rect 1868 936 1876 944
rect 2012 936 2020 944
rect 2044 936 2052 944
rect 2220 936 2228 944
rect 2492 936 2500 944
rect 2604 936 2612 944
rect 188 916 196 924
rect 236 916 244 924
rect 300 916 308 924
rect 556 916 564 924
rect 764 916 772 924
rect 860 916 868 924
rect 1196 916 1204 924
rect 1276 916 1284 924
rect 1580 916 1588 924
rect 1612 916 1620 924
rect 1660 916 1668 924
rect 1756 916 1764 924
rect 1852 916 1860 924
rect 1884 916 1892 924
rect 1948 916 1956 924
rect 2332 916 2340 924
rect 2444 916 2452 924
rect 2476 916 2484 924
rect 2556 916 2564 924
rect 76 896 84 904
rect 124 896 132 904
rect 188 896 196 904
rect 252 896 260 904
rect 268 896 276 904
rect 380 900 388 908
rect 780 896 788 904
rect 1164 900 1172 908
rect 1276 896 1284 904
rect 1724 896 1732 904
rect 1964 896 1972 904
rect 2156 900 2164 908
rect 2428 896 2436 904
rect 12 876 20 884
rect 140 876 148 884
rect 220 876 228 884
rect 892 876 900 884
rect 1628 876 1636 884
rect 2540 876 2548 884
rect 380 854 388 862
rect 2156 854 2164 862
rect 124 836 132 844
rect 236 836 244 844
rect 764 836 772 844
rect 1164 836 1172 844
rect 1276 836 1284 844
rect 1564 836 1572 844
rect 1804 836 1812 844
rect 2044 836 2052 844
rect 659 806 667 814
rect 669 806 677 814
rect 679 806 687 814
rect 689 806 697 814
rect 699 806 707 814
rect 709 806 717 814
rect 748 776 756 784
rect 844 776 852 784
rect 1548 776 1556 784
rect 1596 776 1604 784
rect 2572 776 2580 784
rect 2316 758 2324 766
rect 1980 736 1988 744
rect 220 716 228 724
rect 76 696 84 704
rect 188 696 196 704
rect 348 716 356 724
rect 572 716 580 724
rect 668 716 676 724
rect 700 716 708 724
rect 716 716 724 724
rect 940 716 948 724
rect 1100 716 1108 724
rect 1164 716 1172 724
rect 1740 716 1748 724
rect 1836 716 1844 724
rect 2028 716 2036 724
rect 2316 712 2324 720
rect 268 696 276 704
rect 300 696 308 704
rect 28 676 36 684
rect 92 676 100 684
rect 12 656 20 664
rect 172 676 180 684
rect 252 676 260 684
rect 396 676 404 684
rect 412 676 420 684
rect 540 696 548 704
rect 684 696 692 704
rect 748 696 756 704
rect 780 696 788 704
rect 876 696 884 704
rect 908 696 916 704
rect 988 696 996 704
rect 1100 696 1108 704
rect 1132 696 1140 704
rect 1212 696 1220 704
rect 1516 696 1524 704
rect 1628 696 1636 704
rect 524 676 532 684
rect 588 676 596 684
rect 604 676 612 684
rect 812 676 820 684
rect 940 676 948 684
rect 972 676 980 684
rect 1004 676 1012 684
rect 1052 676 1060 684
rect 1116 676 1124 684
rect 1180 676 1188 684
rect 1372 676 1380 684
rect 1612 676 1620 684
rect 1676 696 1684 704
rect 1804 696 1812 704
rect 2028 696 2036 704
rect 2060 696 2068 704
rect 2092 696 2100 704
rect 2124 696 2132 704
rect 1692 676 1700 684
rect 1772 676 1780 684
rect 1788 676 1796 684
rect 1820 676 1828 684
rect 1868 676 1876 684
rect 2012 676 2020 684
rect 2188 696 2196 704
rect 2284 696 2292 704
rect 2204 676 2212 684
rect 2380 676 2388 684
rect 140 656 148 664
rect 332 656 340 664
rect 588 656 596 664
rect 812 656 820 664
rect 1036 656 1044 664
rect 1628 656 1636 664
rect 1660 656 1668 664
rect 1724 656 1732 664
rect 2124 656 2132 664
rect 2140 656 2148 664
rect 2236 656 2244 664
rect 2412 656 2420 664
rect 60 636 68 644
rect 108 636 116 644
rect 316 636 324 644
rect 348 636 356 644
rect 796 636 804 644
rect 956 636 964 644
rect 1164 636 1172 644
rect 1244 636 1252 644
rect 1484 636 1492 644
rect 1548 636 1556 644
rect 1708 636 1716 644
rect 1740 636 1748 644
rect 2220 636 2228 644
rect 1891 606 1899 614
rect 1901 606 1909 614
rect 1911 606 1919 614
rect 1921 606 1929 614
rect 1931 606 1939 614
rect 1941 606 1949 614
rect 1116 576 1124 584
rect 2108 576 2116 584
rect 2204 576 2212 584
rect 2540 576 2548 584
rect 12 556 20 564
rect 476 556 484 564
rect 892 556 900 564
rect 1068 556 1076 564
rect 1100 556 1108 564
rect 1132 556 1140 564
rect 1324 556 1332 564
rect 1788 556 1796 564
rect 1948 556 1956 564
rect 2060 556 2068 564
rect 2188 556 2196 564
rect 2380 556 2388 564
rect 124 536 132 544
rect 172 536 180 544
rect 236 536 244 544
rect 300 536 308 544
rect 444 536 452 544
rect 748 536 756 544
rect 812 536 820 544
rect 828 536 836 544
rect 892 536 900 544
rect 956 536 964 544
rect 1052 536 1060 544
rect 1356 536 1364 544
rect 1500 536 1508 544
rect 1596 536 1604 544
rect 1756 536 1764 544
rect 2076 536 2084 544
rect 2348 536 2356 544
rect 44 516 52 524
rect 92 516 100 524
rect 156 516 164 524
rect 188 516 196 524
rect 284 516 292 524
rect 348 516 356 524
rect 556 516 564 524
rect 638 516 646 524
rect 732 516 740 524
rect 796 516 804 524
rect 844 516 852 524
rect 940 516 948 524
rect 1004 516 1012 524
rect 1020 516 1028 524
rect 1068 516 1076 524
rect 1420 516 1428 524
rect 1516 516 1524 524
rect 1612 516 1620 524
rect 1868 516 1876 524
rect 2252 516 2260 524
rect 108 496 116 504
rect 220 496 228 504
rect 380 500 388 508
rect 748 496 756 504
rect 812 496 820 504
rect 1004 496 1012 504
rect 1036 496 1044 504
rect 1452 496 1460 504
rect 1548 496 1556 504
rect 1660 496 1668 504
rect 2284 500 2292 508
rect 44 476 52 484
rect 76 476 84 484
rect 956 476 964 484
rect 380 454 388 462
rect 2284 454 2292 462
rect 92 436 100 444
rect 268 436 276 444
rect 908 436 916 444
rect 1084 436 1092 444
rect 1452 436 1460 444
rect 1564 436 1572 444
rect 1660 436 1668 444
rect 1980 436 1988 444
rect 2204 436 2212 444
rect 659 406 667 414
rect 669 406 677 414
rect 679 406 687 414
rect 689 406 697 414
rect 699 406 707 414
rect 709 406 717 414
rect 76 376 84 384
rect 364 376 372 384
rect 940 376 948 384
rect 1468 376 1476 384
rect 1900 376 1908 384
rect 2268 376 2276 384
rect 1212 358 1220 366
rect 1564 358 1572 366
rect 828 336 836 344
rect 364 316 372 324
rect 508 316 516 324
rect 732 316 740 324
rect 796 316 804 324
rect 988 316 996 324
rect 1212 312 1220 320
rect 1564 312 1572 320
rect 2124 316 2132 324
rect 2268 316 2276 324
rect 348 296 356 304
rect 444 296 452 304
rect 476 296 484 304
rect 572 296 580 304
rect 604 296 612 304
rect 636 296 644 304
rect 668 296 676 304
rect 764 296 772 304
rect 812 296 820 304
rect 860 296 868 304
rect 924 296 932 304
rect 940 296 948 304
rect 1020 296 1028 304
rect 1068 296 1076 304
rect 1100 296 1108 304
rect 1132 296 1140 304
rect 1196 296 1204 304
rect 1388 296 1396 304
rect 1740 296 1748 304
rect 1852 296 1860 304
rect 1996 296 2004 304
rect 2012 296 2020 304
rect 2092 296 2100 304
rect 2140 296 2148 304
rect 2156 296 2164 304
rect 2204 296 2212 304
rect 2284 296 2292 304
rect 12 276 20 284
rect 268 276 276 284
rect 460 276 468 284
rect 524 276 532 284
rect 588 276 596 284
rect 652 276 660 284
rect 780 276 788 284
rect 812 276 820 284
rect 1084 276 1092 284
rect 1276 276 1284 284
rect 1628 276 1636 284
rect 2364 276 2372 284
rect 236 256 244 264
rect 412 256 420 264
rect 444 256 452 264
rect 1068 256 1076 264
rect 1308 256 1316 264
rect 1660 256 1668 264
rect 2060 256 2068 264
rect 2108 256 2116 264
rect 2396 256 2404 264
rect 572 236 580 244
rect 876 236 884 244
rect 1820 236 1828 244
rect 1884 236 1892 244
rect 2044 236 2052 244
rect 2076 236 2084 244
rect 2188 236 2196 244
rect 2556 236 2564 244
rect 1891 206 1899 214
rect 1901 206 1909 214
rect 1911 206 1919 214
rect 1921 206 1929 214
rect 1931 206 1939 214
rect 1941 206 1949 214
rect 28 176 36 184
rect 812 176 820 184
rect 940 176 948 184
rect 1372 176 1380 184
rect 2108 176 2116 184
rect 2460 176 2468 184
rect 188 156 196 164
rect 364 156 372 164
rect 476 156 484 164
rect 796 156 804 164
rect 1100 156 1108 164
rect 1564 156 1572 164
rect 1724 156 1732 164
rect 1804 156 1812 164
rect 2268 156 2276 164
rect 2444 156 2452 164
rect 2524 156 2532 164
rect 220 136 228 144
rect 492 136 500 144
rect 748 136 756 144
rect 780 136 788 144
rect 1132 136 1140 144
rect 1276 136 1284 144
rect 1324 136 1332 144
rect 1532 136 1540 144
rect 1836 136 1844 144
rect 2300 136 2308 144
rect 2492 136 2500 144
rect 316 116 324 124
rect 396 116 404 124
rect 412 116 420 124
rect 460 116 468 124
rect 508 116 516 124
rect 540 116 548 124
rect 588 116 596 124
rect 620 116 628 124
rect 764 116 772 124
rect 860 116 868 124
rect 1196 116 1204 124
rect 1228 116 1236 124
rect 1644 116 1652 124
rect 1900 116 1908 124
rect 1964 116 1972 124
rect 1996 116 2004 124
rect 2044 116 2052 124
rect 2188 116 2196 124
rect 2524 116 2532 124
rect 316 96 324 104
rect 604 96 612 104
rect 732 96 740 104
rect 1228 96 1236 104
rect 1468 100 1476 108
rect 2364 100 2372 108
rect 428 76 436 84
rect 444 76 452 84
rect 540 76 548 84
rect 572 76 580 84
rect 588 56 596 64
rect 316 36 324 44
rect 716 36 724 44
rect 828 36 836 44
rect 876 36 884 44
rect 1228 36 1236 44
rect 1468 36 1476 44
rect 1788 36 1796 44
rect 2028 36 2036 44
rect 2076 36 2084 44
rect 2364 36 2372 44
rect 2572 36 2580 44
rect 659 6 667 14
rect 669 6 677 14
rect 679 6 687 14
rect 689 6 697 14
rect 699 6 707 14
rect 709 6 717 14
<< metal2 >>
rect 589 1824 595 1863
rect 29 1544 35 1636
rect 61 1504 67 1536
rect 13 1484 19 1496
rect 61 1364 67 1496
rect 125 1384 131 1616
rect 189 1604 195 1756
rect 221 1624 227 1736
rect 324 1717 332 1723
rect 317 1644 323 1696
rect 237 1464 243 1596
rect 269 1504 275 1556
rect 333 1520 339 1716
rect 573 1644 579 1736
rect 637 1644 643 1700
rect 381 1584 387 1636
rect 525 1584 531 1636
rect 573 1584 579 1616
rect 682 1614 694 1616
rect 667 1606 669 1614
rect 677 1606 679 1614
rect 687 1606 689 1614
rect 697 1606 699 1614
rect 707 1606 709 1614
rect 682 1604 694 1606
rect 388 1517 403 1523
rect 141 1364 147 1436
rect 237 1404 243 1456
rect 317 1364 323 1396
rect 13 1284 19 1296
rect 45 1124 51 1176
rect 61 1164 67 1316
rect 93 1264 99 1316
rect 141 1224 147 1356
rect 285 1304 291 1336
rect 397 1324 403 1517
rect 445 1504 451 1576
rect 413 1484 419 1496
rect 445 1484 451 1496
rect 461 1484 467 1496
rect 477 1464 483 1476
rect 189 1244 195 1296
rect 93 1104 99 1136
rect 100 1097 115 1103
rect 13 1084 19 1096
rect 61 1064 67 1076
rect 109 1064 115 1097
rect 68 1057 83 1063
rect 77 964 83 1057
rect 13 884 19 896
rect 45 824 51 916
rect 93 723 99 1056
rect 125 924 131 1036
rect 141 904 147 1056
rect 141 884 147 896
rect 205 883 211 1036
rect 253 984 259 1216
rect 477 1184 483 1236
rect 493 1184 499 1296
rect 605 1184 611 1496
rect 701 1364 707 1456
rect 733 1444 739 1756
rect 781 1744 787 1756
rect 909 1744 915 1863
rect 1085 1824 1091 1863
rect 1645 1857 1667 1863
rect 909 1604 915 1736
rect 1005 1504 1011 1636
rect 1101 1624 1107 1756
rect 1133 1744 1139 1816
rect 1661 1784 1667 1857
rect 1405 1744 1411 1776
rect 1693 1763 1699 1863
rect 1709 1857 1731 1863
rect 1709 1784 1715 1857
rect 1693 1757 1715 1763
rect 1069 1520 1075 1558
rect 1133 1504 1139 1716
rect 1197 1644 1203 1700
rect 1309 1644 1315 1696
rect 1229 1524 1235 1576
rect 1325 1504 1331 1716
rect 1437 1624 1443 1756
rect 1677 1724 1683 1736
rect 797 1464 803 1496
rect 733 1364 739 1436
rect 637 1244 643 1300
rect 701 1284 707 1336
rect 893 1324 899 1496
rect 1005 1484 1011 1496
rect 1149 1484 1155 1496
rect 973 1444 979 1456
rect 1261 1424 1267 1496
rect 1325 1464 1331 1476
rect 1357 1464 1363 1616
rect 1517 1584 1523 1716
rect 1661 1504 1667 1636
rect 1709 1584 1715 1757
rect 1773 1763 1779 1863
rect 1837 1857 1859 1863
rect 1853 1764 1859 1857
rect 1965 1857 1987 1863
rect 1914 1814 1926 1816
rect 1899 1806 1901 1814
rect 1909 1806 1911 1814
rect 1919 1806 1921 1814
rect 1929 1806 1931 1814
rect 1939 1806 1941 1814
rect 1914 1804 1926 1806
rect 1965 1784 1971 1857
rect 2013 1824 2019 1863
rect 1981 1784 1987 1816
rect 1773 1757 1795 1763
rect 1725 1744 1731 1756
rect 1773 1644 1779 1736
rect 1789 1584 1795 1757
rect 2029 1724 2035 1756
rect 1821 1644 1827 1716
rect 682 1214 694 1216
rect 667 1206 669 1214
rect 677 1206 679 1214
rect 687 1206 689 1214
rect 697 1206 699 1214
rect 707 1206 709 1214
rect 682 1204 694 1206
rect 285 1104 291 1176
rect 525 1124 531 1136
rect 349 1104 355 1116
rect 317 1064 323 1096
rect 253 904 259 976
rect 269 904 275 1036
rect 381 984 387 1116
rect 461 1104 467 1116
rect 429 1084 435 1096
rect 477 1084 483 1116
rect 493 1084 499 1096
rect 445 944 451 1036
rect 285 937 300 943
rect 205 877 220 883
rect 125 724 131 836
rect 77 717 99 723
rect 77 704 83 717
rect 141 704 147 876
rect 237 724 243 836
rect 189 704 195 716
rect 13 664 19 676
rect 29 664 35 676
rect 13 564 19 656
rect 45 524 51 656
rect 77 523 83 696
rect 93 684 99 696
rect 93 543 99 676
rect 141 664 147 676
rect 109 564 115 636
rect 173 544 179 676
rect 93 537 115 543
rect 77 517 92 523
rect 109 504 115 537
rect 125 504 131 536
rect 189 524 195 696
rect 221 664 227 716
rect 253 703 259 896
rect 285 704 291 937
rect 381 862 387 900
rect 477 844 483 956
rect 237 697 259 703
rect 237 604 243 697
rect 269 644 275 696
rect 333 644 339 656
rect 221 504 227 596
rect 237 544 243 556
rect 301 544 307 596
rect 285 504 291 516
rect 93 304 99 436
rect 13 284 19 296
rect 237 264 243 476
rect 269 284 275 436
rect 317 404 323 636
rect 349 544 355 636
rect 397 604 403 676
rect 413 664 419 676
rect 525 664 531 676
rect 541 644 547 696
rect 349 304 355 516
rect 381 462 387 500
rect 477 484 483 556
rect 557 524 563 916
rect 573 724 579 816
rect 589 764 595 1076
rect 605 1064 611 1156
rect 765 1084 771 1176
rect 797 1084 803 1096
rect 637 984 643 1056
rect 765 924 771 1076
rect 893 1063 899 1236
rect 957 1184 963 1276
rect 1037 1144 1043 1356
rect 1053 1344 1059 1356
rect 1309 1324 1315 1416
rect 1357 1364 1363 1456
rect 1133 1262 1139 1300
rect 1053 1184 1059 1256
rect 925 1124 931 1136
rect 1037 1124 1043 1136
rect 1069 1124 1075 1136
rect 909 1084 915 1096
rect 893 1057 915 1063
rect 845 944 851 956
rect 893 924 899 936
rect 682 814 694 816
rect 667 806 669 814
rect 677 806 679 814
rect 687 806 689 814
rect 697 806 699 814
rect 707 806 709 814
rect 682 804 694 806
rect 749 784 755 896
rect 765 744 771 836
rect 573 623 579 716
rect 589 684 595 716
rect 669 704 675 716
rect 701 703 707 716
rect 733 703 739 716
rect 877 704 883 756
rect 701 697 739 703
rect 605 664 611 676
rect 589 624 595 656
rect 573 617 588 623
rect 557 464 563 516
rect 365 324 371 376
rect 445 304 451 396
rect 589 324 595 596
rect 605 524 611 656
rect 749 644 755 696
rect 797 644 803 656
rect 733 524 739 596
rect 749 564 755 636
rect 682 414 694 416
rect 667 406 669 414
rect 677 406 679 414
rect 687 406 689 414
rect 697 406 699 414
rect 707 406 709 414
rect 682 404 694 406
rect 733 384 739 516
rect 237 204 243 256
rect 189 164 195 196
rect 349 124 355 296
rect 445 283 451 296
rect 429 277 451 283
rect 397 257 412 263
rect 397 124 403 257
rect 317 44 323 96
rect 429 84 435 277
rect 461 164 467 276
rect 477 104 483 156
rect 493 144 499 156
rect 493 24 499 136
rect 509 124 515 296
rect 589 284 595 316
rect 525 264 531 276
rect 573 144 579 236
rect 589 143 595 276
rect 621 184 627 316
rect 733 204 739 316
rect 765 304 771 356
rect 781 284 787 556
rect 797 524 803 636
rect 813 604 819 656
rect 813 504 819 536
rect 877 504 883 696
rect 893 624 899 876
rect 909 704 915 1057
rect 909 684 915 696
rect 893 564 899 616
rect 797 263 803 316
rect 813 304 819 496
rect 925 483 931 1096
rect 973 1084 979 1096
rect 1021 1084 1027 1096
rect 1117 1044 1123 1056
rect 1069 964 1075 976
rect 1101 944 1107 956
rect 1197 924 1203 1316
rect 1309 1244 1315 1316
rect 1357 1184 1363 1356
rect 1453 1324 1459 1496
rect 1581 1464 1587 1476
rect 1645 1444 1651 1496
rect 1661 1344 1667 1496
rect 1677 1364 1683 1496
rect 1741 1464 1747 1496
rect 1725 1444 1731 1456
rect 1725 1344 1731 1436
rect 1741 1344 1747 1456
rect 1581 1324 1587 1336
rect 1549 1317 1564 1323
rect 941 724 947 736
rect 1101 724 1107 916
rect 1165 844 1171 900
rect 1213 784 1219 1076
rect 1309 1064 1315 1176
rect 1309 984 1315 1056
rect 1341 1044 1347 1076
rect 1405 964 1411 1176
rect 1421 1104 1427 1236
rect 1437 1124 1443 1176
rect 1517 1124 1523 1136
rect 1485 1084 1491 1096
rect 1549 1084 1555 1317
rect 1629 1184 1635 1336
rect 1588 1117 1603 1123
rect 1581 1084 1587 1096
rect 1597 1084 1603 1117
rect 1373 944 1379 956
rect 1277 844 1283 896
rect 1108 717 1123 723
rect 941 684 947 716
rect 941 624 947 676
rect 957 564 963 636
rect 973 544 979 676
rect 989 664 995 696
rect 1005 684 1011 696
rect 1117 684 1123 717
rect 1133 704 1139 716
rect 1165 704 1171 716
rect 1213 704 1219 776
rect 1373 684 1379 856
rect 1517 704 1523 1076
rect 1588 1057 1603 1063
rect 1581 924 1587 1036
rect 1549 784 1555 896
rect 941 504 947 516
rect 925 477 947 483
rect 909 344 915 436
rect 941 384 947 477
rect 957 364 963 476
rect 957 303 963 356
rect 973 304 979 536
rect 989 324 995 616
rect 1021 524 1027 596
rect 1053 544 1059 676
rect 1117 584 1123 656
rect 1165 584 1171 636
rect 1069 564 1075 576
rect 1133 564 1139 576
rect 1245 564 1251 636
rect 1485 584 1491 636
rect 1245 484 1251 556
rect 1021 304 1027 316
rect 948 297 963 303
rect 797 257 819 263
rect 589 137 604 143
rect 605 104 611 136
rect 621 124 627 176
rect 749 144 755 156
rect 765 124 771 216
rect 797 164 803 196
rect 813 184 819 257
rect 861 204 867 296
rect 1085 284 1091 436
rect 1197 304 1203 456
rect 1325 383 1331 556
rect 1357 544 1363 576
rect 1517 524 1523 676
rect 1565 644 1571 836
rect 1421 424 1427 516
rect 1453 444 1459 496
rect 1309 377 1331 383
rect 1213 320 1219 358
rect 1133 284 1139 296
rect 877 224 883 236
rect 1069 204 1075 256
rect 941 184 947 196
rect 1101 164 1107 176
rect 1133 144 1139 156
rect 1197 124 1203 296
rect 1309 264 1315 377
rect 1389 304 1395 416
rect 1469 384 1475 416
rect 1309 184 1315 256
rect 1517 244 1523 516
rect 1549 504 1555 636
rect 1565 404 1571 436
rect 1581 424 1587 916
rect 1597 784 1603 1057
rect 1613 904 1619 916
rect 1629 704 1635 876
rect 1629 644 1635 656
rect 1613 524 1619 596
rect 1645 544 1651 1076
rect 1661 944 1667 1336
rect 1677 1124 1683 1296
rect 1725 923 1731 1036
rect 1741 963 1747 1316
rect 1757 1083 1763 1336
rect 1780 1097 1795 1103
rect 1789 1084 1795 1097
rect 1757 1077 1772 1083
rect 1741 957 1756 963
rect 1757 924 1763 956
rect 1725 917 1747 923
rect 1661 884 1667 916
rect 1677 704 1683 876
rect 1741 743 1747 917
rect 1773 904 1779 936
rect 1789 884 1795 1076
rect 1837 964 1843 1036
rect 1853 924 1859 1476
rect 1869 1184 1875 1716
rect 2045 1524 2051 1636
rect 2061 1504 2067 1636
rect 2109 1584 2115 1736
rect 2237 1643 2243 1756
rect 2477 1724 2483 1756
rect 2237 1637 2259 1643
rect 2125 1504 2131 1516
rect 2221 1504 2227 1596
rect 2077 1484 2083 1496
rect 1914 1414 1926 1416
rect 1899 1406 1901 1414
rect 1909 1406 1911 1414
rect 1919 1406 1921 1414
rect 1929 1406 1931 1414
rect 1939 1406 1941 1414
rect 1914 1404 1926 1406
rect 1997 1364 2003 1436
rect 2045 1404 2051 1436
rect 2109 1324 2115 1396
rect 2093 1244 2099 1300
rect 2141 1204 2147 1496
rect 2173 1464 2179 1496
rect 2253 1444 2259 1637
rect 2269 1504 2275 1716
rect 2365 1644 2371 1696
rect 2413 1684 2419 1716
rect 2445 1684 2451 1696
rect 2461 1604 2467 1636
rect 2317 1520 2323 1558
rect 1914 1014 1926 1016
rect 1899 1006 1901 1014
rect 1909 1006 1911 1014
rect 1919 1006 1921 1014
rect 1929 1006 1931 1014
rect 1939 1006 1941 1014
rect 1914 1004 1926 1006
rect 1725 737 1747 743
rect 1661 444 1667 496
rect 1565 320 1571 358
rect 1629 284 1635 396
rect 1677 383 1683 576
rect 1693 444 1699 676
rect 1725 664 1731 737
rect 1741 704 1747 716
rect 1805 704 1811 836
rect 1869 684 1875 936
rect 1885 924 1891 956
rect 1949 924 1955 956
rect 1965 904 1971 1116
rect 1997 1084 2003 1096
rect 2173 1064 2179 1436
rect 2285 1404 2291 1496
rect 2413 1444 2419 1456
rect 2205 1324 2211 1396
rect 2333 1364 2339 1416
rect 2205 1104 2211 1316
rect 2237 1262 2243 1300
rect 2269 1120 2275 1158
rect 2493 1124 2499 1636
rect 2509 1364 2515 1756
rect 2573 1584 2579 1716
rect 2077 964 2083 1056
rect 2173 1004 2179 1056
rect 2013 684 2019 896
rect 2029 724 2035 736
rect 2045 684 2051 836
rect 1789 664 1795 676
rect 1869 644 1875 676
rect 1709 624 1715 636
rect 1741 604 1747 636
rect 1757 544 1763 616
rect 1914 614 1926 616
rect 1899 606 1901 614
rect 1909 606 1911 614
rect 1919 606 1921 614
rect 1929 606 1931 614
rect 1939 606 1941 614
rect 1914 604 1926 606
rect 1789 564 1795 576
rect 2013 564 2019 676
rect 1869 404 1875 516
rect 1661 377 1683 383
rect 1661 264 1667 377
rect 1741 304 1747 396
rect 1901 384 1907 396
rect 1661 164 1667 256
rect 1277 124 1283 136
rect 541 84 547 96
rect 541 24 547 76
rect 589 64 595 96
rect 1229 44 1235 96
rect 461 -23 467 16
rect 509 -23 515 16
rect 682 14 694 16
rect 667 6 669 14
rect 677 6 679 14
rect 687 6 689 14
rect 697 6 699 14
rect 707 6 709 14
rect 682 4 694 6
rect 749 -23 755 36
rect 829 -17 835 36
rect 877 -17 883 36
rect 1325 -17 1331 136
rect 1741 124 1747 296
rect 1869 237 1884 243
rect 1469 44 1475 100
rect 1789 -17 1795 36
rect 1869 24 1875 237
rect 1914 214 1926 216
rect 1899 206 1901 214
rect 1909 206 1911 214
rect 1919 206 1921 214
rect 1929 206 1931 214
rect 1939 206 1941 214
rect 1914 204 1926 206
rect 1965 124 1971 296
rect 1981 124 1987 436
rect 1997 304 2003 316
rect 2013 304 2019 556
rect 2077 544 2083 956
rect 2221 944 2227 1016
rect 2317 1003 2323 1096
rect 2349 1064 2355 1076
rect 2413 1024 2419 1076
rect 2317 997 2339 1003
rect 2253 964 2259 996
rect 2093 704 2099 936
rect 2333 924 2339 997
rect 2429 904 2435 1116
rect 2509 1104 2515 1196
rect 2541 1184 2547 1336
rect 2605 1284 2611 1296
rect 2573 1104 2579 1116
rect 2468 1097 2483 1103
rect 2477 924 2483 1097
rect 2493 984 2499 1056
rect 2493 944 2499 976
rect 2157 862 2163 900
rect 2445 824 2451 916
rect 2109 584 2115 716
rect 2189 704 2195 796
rect 2125 644 2131 656
rect 2141 550 2147 656
rect 2189 564 2195 636
rect 2205 584 2211 676
rect 2237 664 2243 816
rect 2477 804 2483 916
rect 2317 720 2323 758
rect 2221 544 2227 636
rect 2253 524 2259 696
rect 2381 584 2387 656
rect 2381 564 2387 576
rect 2157 304 2163 336
rect 2061 244 2067 256
rect 1997 124 2003 236
rect 2045 143 2051 236
rect 2077 164 2083 236
rect 2109 184 2115 256
rect 2045 137 2067 143
rect 829 -23 851 -17
rect 877 -23 899 -17
rect 1325 -23 1363 -17
rect 1773 -23 1795 -17
rect 1981 -23 1987 16
rect 2029 -17 2035 36
rect 2061 -17 2067 137
rect 2109 124 2115 176
rect 2173 123 2179 396
rect 2205 344 2211 436
rect 2253 404 2259 516
rect 2285 462 2291 500
rect 2269 324 2275 376
rect 2205 304 2211 316
rect 2285 304 2291 396
rect 2381 383 2387 556
rect 2509 503 2515 1096
rect 2557 924 2563 1056
rect 2541 884 2547 896
rect 2557 783 2563 916
rect 2557 777 2572 783
rect 2541 584 2547 636
rect 2493 497 2515 503
rect 2381 377 2403 383
rect 2189 144 2195 236
rect 2269 164 2275 236
rect 2365 224 2371 276
rect 2397 264 2403 377
rect 2493 304 2499 497
rect 2397 244 2403 256
rect 2461 184 2467 216
rect 2493 144 2499 296
rect 2525 164 2531 236
rect 2525 124 2531 156
rect 2173 117 2188 123
rect 2365 44 2371 100
rect 2013 -23 2035 -17
rect 2045 -23 2067 -17
rect 2077 -23 2083 36
rect 2573 -17 2579 36
rect 2557 -23 2579 -17
<< m3contact >>
rect 588 1816 596 1824
rect 188 1756 196 1764
rect 540 1756 548 1764
rect 732 1756 740 1764
rect 780 1756 788 1764
rect 124 1616 132 1624
rect 28 1536 36 1544
rect 60 1536 68 1544
rect 12 1496 20 1504
rect 76 1436 84 1444
rect 332 1716 340 1724
rect 460 1716 468 1724
rect 220 1616 228 1624
rect 188 1596 196 1604
rect 236 1596 244 1604
rect 524 1636 532 1644
rect 572 1636 580 1644
rect 572 1616 580 1624
rect 659 1606 667 1614
rect 669 1606 677 1614
rect 679 1606 687 1614
rect 689 1606 697 1614
rect 699 1606 707 1614
rect 709 1606 717 1614
rect 380 1576 388 1584
rect 444 1576 452 1584
rect 268 1476 276 1484
rect 140 1436 148 1444
rect 236 1396 244 1404
rect 316 1396 324 1404
rect 12 1296 20 1304
rect 44 1176 52 1184
rect 92 1256 100 1264
rect 556 1516 564 1524
rect 620 1516 628 1524
rect 460 1496 468 1504
rect 524 1496 532 1504
rect 636 1496 644 1504
rect 412 1476 420 1484
rect 444 1476 452 1484
rect 476 1476 484 1484
rect 396 1316 404 1324
rect 588 1316 596 1324
rect 284 1296 292 1304
rect 492 1296 500 1304
rect 140 1216 148 1224
rect 252 1216 260 1224
rect 60 1156 68 1164
rect 92 1136 100 1144
rect 172 1116 180 1124
rect 204 1116 212 1124
rect 12 1096 20 1104
rect 60 1076 68 1084
rect 172 1076 180 1084
rect 220 1076 228 1084
rect 44 1056 52 1064
rect 140 1056 148 1064
rect 12 896 20 904
rect 76 896 84 904
rect 44 816 52 824
rect 188 916 196 924
rect 124 896 132 904
rect 140 896 148 904
rect 188 896 196 904
rect 716 1456 724 1464
rect 1084 1816 1092 1824
rect 1132 1816 1140 1824
rect 940 1636 948 1644
rect 1004 1636 1012 1644
rect 908 1596 916 1604
rect 1404 1776 1412 1784
rect 1100 1616 1108 1624
rect 1596 1736 1598 1744
rect 1598 1736 1604 1744
rect 1676 1736 1684 1744
rect 1516 1716 1524 1724
rect 1628 1716 1636 1724
rect 1356 1616 1364 1624
rect 1436 1616 1444 1624
rect 796 1496 804 1504
rect 1004 1496 1012 1504
rect 1100 1496 1108 1504
rect 1132 1496 1140 1504
rect 1148 1496 1156 1504
rect 1180 1496 1188 1504
rect 812 1456 820 1464
rect 732 1436 740 1444
rect 700 1356 708 1364
rect 972 1436 980 1444
rect 1660 1636 1668 1644
rect 1788 1776 1796 1784
rect 1891 1806 1899 1814
rect 1901 1806 1909 1814
rect 1911 1806 1919 1814
rect 1921 1806 1929 1814
rect 1931 1806 1939 1814
rect 1941 1806 1949 1814
rect 1980 1816 1988 1824
rect 2012 1816 2020 1824
rect 1724 1736 1732 1744
rect 1772 1636 1780 1644
rect 2028 1756 2036 1764
rect 2060 1756 2068 1764
rect 2108 1736 2116 1744
rect 1820 1636 1828 1644
rect 1452 1496 1460 1504
rect 1324 1456 1332 1464
rect 1260 1416 1268 1424
rect 1308 1416 1316 1424
rect 1036 1356 1044 1364
rect 1052 1356 1060 1364
rect 1228 1356 1236 1364
rect 924 1336 932 1344
rect 812 1316 820 1324
rect 892 1316 900 1324
rect 700 1276 708 1284
rect 956 1276 964 1284
rect 659 1206 667 1214
rect 669 1206 677 1214
rect 679 1206 687 1214
rect 689 1206 697 1214
rect 699 1206 707 1214
rect 709 1206 717 1214
rect 284 1176 292 1184
rect 476 1176 484 1184
rect 604 1176 612 1184
rect 764 1176 772 1184
rect 268 1136 276 1144
rect 604 1156 612 1164
rect 524 1136 532 1144
rect 348 1116 356 1124
rect 476 1116 484 1124
rect 540 1116 548 1124
rect 316 1096 324 1104
rect 316 1056 324 1064
rect 252 976 260 984
rect 236 916 244 924
rect 396 1096 404 1104
rect 428 1096 436 1104
rect 460 1096 468 1104
rect 524 1096 532 1104
rect 572 1096 580 1104
rect 412 1076 420 1084
rect 492 1076 500 1084
rect 396 1056 404 1064
rect 380 976 388 984
rect 124 716 132 724
rect 188 716 196 724
rect 236 716 244 724
rect 92 696 100 704
rect 140 696 148 704
rect 188 696 196 704
rect 12 676 20 684
rect 28 656 36 664
rect 44 656 52 664
rect 12 556 20 564
rect 60 636 68 644
rect 140 676 148 684
rect 172 676 180 684
rect 108 556 116 564
rect 300 916 308 924
rect 476 836 484 844
rect 348 716 356 724
rect 220 656 228 664
rect 284 696 292 704
rect 300 696 308 704
rect 252 676 260 684
rect 396 676 404 684
rect 268 636 276 644
rect 332 636 340 644
rect 220 596 228 604
rect 236 596 244 604
rect 300 596 308 604
rect 156 516 164 524
rect 236 556 244 564
rect 124 496 132 504
rect 284 496 292 504
rect 44 476 52 484
rect 76 476 84 484
rect 236 476 244 484
rect 76 376 84 384
rect 12 296 20 304
rect 92 296 100 304
rect 412 656 420 664
rect 524 656 532 664
rect 540 636 548 644
rect 396 596 404 604
rect 348 536 356 544
rect 444 536 452 544
rect 316 396 324 404
rect 572 816 580 824
rect 748 1116 756 1124
rect 636 1096 644 1104
rect 668 1096 676 1104
rect 780 1136 788 1144
rect 796 1096 804 1104
rect 876 1096 884 1104
rect 764 1076 772 1084
rect 844 1080 852 1084
rect 844 1076 852 1080
rect 860 1076 868 1084
rect 604 1056 612 1064
rect 636 1056 644 1064
rect 876 1056 884 1064
rect 1196 1336 1204 1344
rect 1356 1356 1364 1364
rect 1388 1356 1396 1364
rect 1052 1256 1060 1264
rect 924 1136 932 1144
rect 988 1136 996 1144
rect 1036 1136 1044 1144
rect 1148 1136 1156 1144
rect 924 1116 932 1124
rect 1068 1116 1076 1124
rect 1100 1116 1108 1124
rect 924 1096 932 1104
rect 956 1096 964 1104
rect 972 1096 980 1104
rect 1052 1096 1060 1104
rect 908 1076 916 1084
rect 844 956 852 964
rect 812 936 820 944
rect 892 936 900 944
rect 860 916 868 924
rect 892 916 900 924
rect 748 896 756 904
rect 780 896 788 904
rect 659 806 667 814
rect 669 806 677 814
rect 679 806 687 814
rect 689 806 697 814
rect 699 806 707 814
rect 709 806 717 814
rect 588 756 596 764
rect 844 776 852 784
rect 876 756 884 764
rect 764 736 772 744
rect 588 716 596 724
rect 716 716 724 724
rect 732 716 740 724
rect 668 696 676 704
rect 684 696 692 704
rect 780 696 788 704
rect 876 696 884 704
rect 604 656 612 664
rect 588 616 596 624
rect 588 596 596 604
rect 476 476 484 484
rect 556 456 564 464
rect 444 396 452 404
rect 812 676 820 684
rect 796 656 804 664
rect 748 636 756 644
rect 732 596 740 604
rect 748 556 756 564
rect 780 556 788 564
rect 748 536 756 544
rect 604 516 612 524
rect 636 516 638 524
rect 638 516 644 524
rect 659 406 667 414
rect 669 406 677 414
rect 679 406 687 414
rect 689 406 697 414
rect 699 406 707 414
rect 709 406 717 414
rect 748 496 756 504
rect 732 376 740 384
rect 764 356 772 364
rect 508 316 516 324
rect 588 316 596 324
rect 620 316 628 324
rect 732 316 740 324
rect 476 296 484 304
rect 508 296 516 304
rect 572 296 580 304
rect 188 196 196 204
rect 236 196 244 204
rect 28 176 36 184
rect 220 136 228 144
rect 364 156 372 164
rect 316 116 324 124
rect 348 116 356 124
rect 412 116 420 124
rect 444 256 452 264
rect 460 156 468 164
rect 492 156 500 164
rect 460 116 468 124
rect 476 96 484 104
rect 444 76 452 84
rect 604 296 612 304
rect 524 256 532 264
rect 572 136 580 144
rect 636 296 644 304
rect 668 296 676 304
rect 652 276 660 284
rect 812 596 820 604
rect 828 536 836 544
rect 844 516 852 524
rect 908 676 916 684
rect 892 616 900 624
rect 892 536 900 544
rect 812 496 820 504
rect 876 496 884 504
rect 972 1076 980 1084
rect 1020 1076 1028 1084
rect 1116 1036 1124 1044
rect 1068 976 1076 984
rect 1100 956 1108 964
rect 1308 1236 1316 1244
rect 1580 1456 1588 1464
rect 1644 1436 1652 1444
rect 1468 1356 1476 1364
rect 1804 1476 1812 1484
rect 1852 1476 1860 1484
rect 1724 1456 1732 1464
rect 1676 1356 1684 1364
rect 1500 1336 1508 1344
rect 1580 1336 1588 1344
rect 1660 1336 1668 1344
rect 1708 1336 1716 1344
rect 1420 1236 1428 1244
rect 1308 1176 1316 1184
rect 1356 1176 1364 1184
rect 1404 1176 1412 1184
rect 1212 1076 1220 1084
rect 1100 916 1108 924
rect 1196 916 1204 924
rect 940 736 948 744
rect 1340 1036 1348 1044
rect 1308 976 1316 984
rect 1516 1116 1524 1124
rect 1532 1096 1540 1104
rect 1564 1316 1572 1324
rect 1596 1316 1604 1324
rect 1644 1316 1652 1324
rect 1628 1176 1636 1184
rect 1580 1096 1588 1104
rect 1484 1076 1492 1084
rect 1516 1076 1524 1084
rect 1596 1076 1604 1084
rect 1372 956 1380 964
rect 1276 916 1284 924
rect 1372 856 1380 864
rect 1212 776 1220 784
rect 1004 696 1012 704
rect 1100 696 1108 704
rect 972 676 980 684
rect 940 616 948 624
rect 956 556 964 564
rect 1132 716 1140 724
rect 1164 696 1172 704
rect 1580 1036 1588 1044
rect 1548 896 1556 904
rect 1116 676 1124 684
rect 1180 676 1188 684
rect 1516 676 1524 684
rect 988 656 996 664
rect 1036 656 1044 664
rect 988 616 996 624
rect 956 536 964 544
rect 972 536 980 544
rect 940 496 948 504
rect 956 356 964 364
rect 828 336 836 344
rect 908 336 916 344
rect 924 296 932 304
rect 1020 596 1028 604
rect 1116 656 1124 664
rect 1068 576 1076 584
rect 1132 576 1140 584
rect 1164 576 1172 584
rect 1356 576 1364 584
rect 1484 576 1492 584
rect 1100 556 1108 564
rect 1244 556 1252 564
rect 1324 556 1332 564
rect 1004 516 1012 524
rect 1068 516 1076 524
rect 1004 496 1012 504
rect 1036 496 1044 504
rect 1244 476 1252 484
rect 1196 456 1204 464
rect 1020 316 1028 324
rect 972 296 980 304
rect 1068 296 1076 304
rect 812 276 820 284
rect 764 216 772 224
rect 732 196 740 204
rect 620 176 628 184
rect 604 136 612 144
rect 540 116 548 124
rect 588 116 596 124
rect 748 156 756 164
rect 796 196 804 204
rect 1500 536 1508 544
rect 1564 636 1572 644
rect 1388 416 1396 424
rect 1420 416 1428 424
rect 1468 416 1476 424
rect 1100 296 1108 304
rect 1132 276 1140 284
rect 876 216 884 224
rect 860 196 868 204
rect 940 196 948 204
rect 1068 196 1076 204
rect 1100 176 1108 184
rect 1132 156 1140 164
rect 780 136 788 144
rect 1276 276 1284 284
rect 1612 896 1620 904
rect 1628 876 1636 884
rect 1612 676 1620 684
rect 1628 636 1636 644
rect 1612 596 1620 604
rect 1596 536 1604 544
rect 1740 1316 1748 1324
rect 1676 1116 1684 1124
rect 1724 1116 1732 1124
rect 1692 1096 1700 1104
rect 1692 956 1700 964
rect 1676 936 1684 944
rect 1820 1096 1828 1104
rect 1756 956 1764 964
rect 1724 896 1732 904
rect 1660 876 1668 884
rect 1676 876 1684 884
rect 1772 896 1780 904
rect 1836 956 1844 964
rect 1820 936 1828 944
rect 2060 1636 2068 1644
rect 2044 1516 2052 1524
rect 2268 1736 2276 1744
rect 2476 1716 2484 1724
rect 2220 1596 2228 1604
rect 2124 1516 2132 1524
rect 1948 1496 1956 1504
rect 2060 1496 2068 1504
rect 2140 1496 2148 1504
rect 2076 1476 2084 1484
rect 1916 1436 1924 1444
rect 1996 1436 2004 1444
rect 1891 1406 1899 1414
rect 1901 1406 1909 1414
rect 1911 1406 1919 1414
rect 1921 1406 1929 1414
rect 1931 1406 1939 1414
rect 1941 1406 1949 1414
rect 2044 1396 2052 1404
rect 2108 1396 2116 1404
rect 2028 1336 2036 1344
rect 2236 1476 2244 1484
rect 2172 1456 2180 1464
rect 2444 1696 2452 1704
rect 2412 1676 2420 1684
rect 2460 1596 2468 1604
rect 2172 1436 2180 1444
rect 2252 1436 2260 1444
rect 2140 1196 2148 1204
rect 1868 1176 1876 1184
rect 2012 1176 2020 1184
rect 1964 1116 1972 1124
rect 1868 1096 1876 1104
rect 1891 1006 1899 1014
rect 1901 1006 1909 1014
rect 1911 1006 1919 1014
rect 1921 1006 1929 1014
rect 1931 1006 1939 1014
rect 1941 1006 1949 1014
rect 1884 956 1892 964
rect 1948 956 1956 964
rect 1788 876 1796 884
rect 1660 656 1668 664
rect 1676 576 1684 584
rect 1644 536 1652 544
rect 1580 416 1588 424
rect 1564 396 1572 404
rect 1628 396 1636 404
rect 1836 716 1844 724
rect 1740 696 1748 704
rect 1996 1096 2004 1104
rect 2380 1476 2388 1484
rect 2412 1436 2420 1444
rect 2332 1416 2340 1424
rect 2204 1396 2212 1404
rect 2284 1396 2292 1404
rect 2300 1336 2308 1344
rect 2604 1736 2612 1744
rect 2524 1716 2532 1724
rect 2572 1716 2580 1724
rect 2540 1336 2548 1344
rect 2508 1196 2516 1204
rect 2396 1116 2404 1124
rect 2428 1116 2436 1124
rect 2492 1116 2500 1124
rect 2364 1096 2372 1104
rect 2204 1076 2212 1084
rect 2076 1056 2084 1064
rect 2220 1016 2228 1024
rect 2172 996 2180 1004
rect 1980 956 1988 964
rect 2044 956 2052 964
rect 2012 936 2020 944
rect 2044 936 2052 944
rect 2012 896 2020 904
rect 1980 736 1988 744
rect 2028 736 2036 744
rect 2028 696 2036 704
rect 2060 696 2068 704
rect 1772 676 1780 684
rect 1820 676 1828 684
rect 2044 676 2052 684
rect 1788 656 1796 664
rect 1868 636 1876 644
rect 1708 616 1716 624
rect 1756 616 1764 624
rect 1740 596 1748 604
rect 1891 606 1899 614
rect 1901 606 1909 614
rect 1911 606 1919 614
rect 1921 606 1929 614
rect 1931 606 1939 614
rect 1941 606 1949 614
rect 1788 576 1796 584
rect 1948 556 1956 564
rect 2012 556 2020 564
rect 2060 556 2068 564
rect 1692 436 1700 444
rect 1980 436 1988 444
rect 1740 396 1748 404
rect 1868 396 1876 404
rect 1900 396 1908 404
rect 1852 296 1860 304
rect 1964 296 1972 304
rect 1516 236 1524 244
rect 1308 176 1316 184
rect 1372 176 1380 184
rect 1564 156 1572 164
rect 1660 156 1668 164
rect 1724 156 1732 164
rect 1532 136 1540 144
rect 860 116 868 124
rect 1228 116 1236 124
rect 1276 116 1284 124
rect 540 96 548 104
rect 588 96 596 104
rect 732 96 740 104
rect 572 76 580 84
rect 716 36 724 44
rect 748 36 756 44
rect 460 16 468 24
rect 492 16 500 24
rect 508 16 516 24
rect 540 16 548 24
rect 659 6 667 14
rect 669 6 677 14
rect 679 6 687 14
rect 689 6 697 14
rect 699 6 707 14
rect 709 6 717 14
rect 1820 236 1828 244
rect 1804 156 1812 164
rect 1836 136 1844 144
rect 1644 116 1652 124
rect 1740 116 1748 124
rect 1891 206 1899 214
rect 1901 206 1909 214
rect 1911 206 1919 214
rect 1921 206 1929 214
rect 1931 206 1939 214
rect 1941 206 1949 214
rect 1996 316 2004 324
rect 2252 996 2260 1004
rect 2348 1056 2356 1064
rect 2412 1016 2420 1024
rect 2092 936 2100 944
rect 2412 976 2420 984
rect 2604 1296 2612 1304
rect 2572 1116 2580 1124
rect 2460 1096 2468 1104
rect 2492 1096 2500 1104
rect 2524 1096 2532 1104
rect 2492 976 2500 984
rect 2236 816 2244 824
rect 2444 816 2452 824
rect 2188 796 2196 804
rect 2108 716 2116 724
rect 2124 696 2132 704
rect 2124 636 2132 644
rect 2188 636 2196 644
rect 2476 796 2484 804
rect 2252 696 2260 704
rect 2284 696 2292 704
rect 2220 536 2228 544
rect 2380 676 2388 684
rect 2380 656 2388 664
rect 2412 656 2420 664
rect 2380 576 2388 584
rect 2348 536 2356 544
rect 2172 396 2180 404
rect 2156 336 2164 344
rect 2124 316 2132 324
rect 2092 296 2100 304
rect 2140 296 2148 304
rect 1996 236 2004 244
rect 2060 236 2068 244
rect 2076 156 2084 164
rect 1900 116 1908 124
rect 1980 116 1988 124
rect 2044 116 2052 124
rect 1868 16 1876 24
rect 1980 16 1988 24
rect 2108 116 2116 124
rect 2252 396 2260 404
rect 2284 396 2292 404
rect 2204 336 2212 344
rect 2204 316 2212 324
rect 2556 1056 2564 1064
rect 2604 936 2612 944
rect 2540 896 2548 904
rect 2540 636 2548 644
rect 2268 236 2276 244
rect 2492 296 2500 304
rect 2396 236 2404 244
rect 2364 216 2372 224
rect 2460 216 2468 224
rect 2444 156 2452 164
rect 2524 236 2532 244
rect 2556 236 2564 244
rect 2188 136 2196 144
rect 2300 136 2308 144
<< metal3 >>
rect 1092 1817 1132 1823
rect 1988 1817 2012 1823
rect 1890 1814 1950 1816
rect 1890 1806 1891 1814
rect 1900 1806 1901 1814
rect 1939 1806 1940 1814
rect 1949 1806 1950 1814
rect 1890 1804 1950 1806
rect 1412 1777 1788 1783
rect 196 1757 540 1763
rect 548 1757 732 1763
rect 740 1757 780 1763
rect 2036 1757 2060 1763
rect 1604 1737 1676 1743
rect 1684 1737 1724 1743
rect 2116 1737 2268 1743
rect 2612 1737 2643 1743
rect 340 1717 460 1723
rect 1524 1717 1628 1723
rect 2484 1717 2524 1723
rect 2532 1717 2572 1723
rect 2452 1697 2643 1703
rect 532 1637 572 1643
rect 948 1637 1004 1643
rect 1668 1637 1772 1643
rect 1780 1637 1820 1643
rect 1828 1637 2060 1643
rect 132 1617 220 1623
rect 580 1617 588 1623
rect 1108 1617 1356 1623
rect 1364 1617 1436 1623
rect 658 1614 718 1616
rect 658 1606 659 1614
rect 668 1606 669 1614
rect 707 1606 708 1614
rect 717 1606 718 1614
rect 658 1604 718 1606
rect 196 1597 236 1603
rect 2228 1597 2460 1603
rect 388 1577 444 1583
rect 36 1537 60 1543
rect 564 1517 620 1523
rect 2052 1517 2124 1523
rect -35 1497 12 1503
rect 468 1497 524 1503
rect 532 1497 636 1503
rect 804 1497 1004 1503
rect 1108 1497 1132 1503
rect 1140 1497 1148 1503
rect 1188 1497 1452 1503
rect 1460 1497 1948 1503
rect 1956 1497 1996 1503
rect 2068 1497 2140 1503
rect 276 1477 412 1483
rect 452 1477 476 1483
rect 916 1477 1388 1483
rect 1396 1477 1804 1483
rect 1860 1477 2076 1483
rect 2244 1477 2380 1483
rect 724 1457 812 1463
rect 1332 1457 1580 1463
rect 1732 1457 2172 1463
rect 84 1437 140 1443
rect 740 1437 972 1443
rect 1652 1437 1836 1443
rect 1924 1437 1996 1443
rect 2004 1437 2172 1443
rect 2180 1437 2252 1443
rect 2260 1437 2412 1443
rect 2333 1424 2339 1437
rect 1268 1417 1308 1423
rect 1890 1414 1950 1416
rect 1890 1406 1891 1414
rect 1900 1406 1901 1414
rect 1939 1406 1940 1414
rect 1949 1406 1950 1414
rect 1890 1404 1950 1406
rect 244 1397 316 1403
rect 2052 1397 2108 1403
rect 2116 1397 2204 1403
rect 2212 1397 2284 1403
rect 708 1357 1036 1363
rect 1060 1357 1228 1363
rect 1236 1357 1356 1363
rect 1396 1357 1468 1363
rect 1476 1357 1676 1363
rect 916 1337 924 1343
rect 1204 1337 1500 1343
rect 1588 1337 1660 1343
rect 1716 1337 2028 1343
rect 2308 1337 2540 1343
rect 404 1317 588 1323
rect 820 1317 892 1323
rect 1572 1317 1596 1323
rect 1652 1317 1740 1323
rect -35 1297 12 1303
rect 292 1297 492 1303
rect 2612 1297 2643 1303
rect 708 1277 956 1283
rect 100 1257 1052 1263
rect 1316 1237 1420 1243
rect 148 1217 252 1223
rect 658 1214 718 1216
rect 658 1206 659 1214
rect 668 1206 669 1214
rect 707 1206 708 1214
rect 717 1206 718 1214
rect 658 1204 718 1206
rect 2148 1197 2508 1203
rect -35 1177 44 1183
rect 52 1177 284 1183
rect 484 1177 604 1183
rect 612 1177 764 1183
rect 1316 1177 1356 1183
rect 1364 1177 1404 1183
rect 1636 1177 1868 1183
rect 1876 1177 2012 1183
rect 68 1157 604 1163
rect -35 1137 92 1143
rect 100 1137 268 1143
rect 532 1137 780 1143
rect 932 1137 988 1143
rect 1044 1137 1148 1143
rect 180 1117 204 1123
rect 212 1117 348 1123
rect 484 1117 540 1123
rect 548 1117 748 1123
rect 756 1117 924 1123
rect 1076 1117 1100 1123
rect 1524 1117 1676 1123
rect 1684 1117 1724 1123
rect 1732 1117 1964 1123
rect 1972 1117 2396 1123
rect 2404 1117 2428 1123
rect 2500 1117 2572 1123
rect -35 1097 12 1103
rect 20 1097 316 1103
rect 404 1097 428 1103
rect 468 1097 524 1103
rect 580 1097 636 1103
rect 676 1097 796 1103
rect 804 1097 876 1103
rect 932 1097 956 1103
rect 980 1097 1052 1103
rect 1060 1097 1532 1103
rect 1540 1097 1580 1103
rect 1700 1097 1820 1103
rect 1828 1097 1868 1103
rect 2004 1097 2364 1103
rect 2372 1097 2460 1103
rect 2500 1097 2524 1103
rect -35 1077 60 1083
rect -35 1057 -29 1077
rect 68 1077 172 1083
rect 180 1077 220 1083
rect 420 1077 492 1083
rect 772 1077 844 1083
rect 868 1077 908 1083
rect 916 1077 972 1083
rect 1028 1077 1212 1083
rect 1220 1077 1484 1083
rect 1492 1077 1516 1083
rect 1604 1077 2204 1083
rect 52 1057 140 1063
rect 324 1057 396 1063
rect 612 1057 636 1063
rect 845 1063 851 1076
rect 845 1057 876 1063
rect 2084 1057 2348 1063
rect 2356 1057 2556 1063
rect 1124 1037 1340 1043
rect 1348 1037 1580 1043
rect 2228 1017 2412 1023
rect 1890 1014 1950 1016
rect 1890 1006 1891 1014
rect 1900 1006 1901 1014
rect 1939 1006 1940 1014
rect 1949 1006 1950 1014
rect 1890 1004 1950 1006
rect 2180 997 2252 1003
rect 260 977 380 983
rect 1076 977 1308 983
rect 2420 977 2492 983
rect 852 957 1100 963
rect 1380 957 1692 963
rect 1764 957 1836 963
rect 1844 957 1884 963
rect 1892 957 1948 963
rect 1988 957 2044 963
rect 820 937 892 943
rect 1684 937 1820 943
rect 1844 937 2012 943
rect 2020 937 2044 943
rect 2052 937 2092 943
rect 2612 937 2643 943
rect 196 917 236 923
rect 308 917 860 923
rect 900 917 1100 923
rect 1204 917 1276 923
rect -35 897 12 903
rect 84 897 124 903
rect 148 897 188 903
rect 756 897 780 903
rect 1556 897 1612 903
rect 1620 897 1724 903
rect 1780 897 2012 903
rect 2548 897 2643 903
rect 1636 877 1660 883
rect 1668 877 1676 883
rect 1684 877 1788 883
rect 1380 857 1388 863
rect 484 837 492 843
rect 52 817 572 823
rect 2244 817 2444 823
rect 658 814 718 816
rect 658 806 659 814
rect 668 806 669 814
rect 707 806 708 814
rect 717 806 718 814
rect 658 804 718 806
rect 2196 797 2476 803
rect 852 777 1212 783
rect 596 757 876 763
rect 772 737 940 743
rect 1988 737 2028 743
rect 132 717 188 723
rect 244 717 348 723
rect 596 717 716 723
rect 740 717 1132 723
rect 1844 717 2108 723
rect 100 697 140 703
rect 196 697 284 703
rect 292 697 300 703
rect 381 697 668 703
rect -35 663 -29 683
rect 20 677 140 683
rect 148 677 172 683
rect 381 683 387 697
rect 692 697 780 703
rect 884 697 1004 703
rect 1108 697 1164 703
rect 1748 697 2028 703
rect 2068 697 2124 703
rect 2260 697 2284 703
rect 260 677 387 683
rect 404 677 812 683
rect 916 677 972 683
rect 1124 677 1180 683
rect 1524 677 1612 683
rect 1780 677 1820 683
rect 2052 677 2380 683
rect -35 657 28 663
rect 36 657 44 663
rect 52 657 220 663
rect 420 657 524 663
rect 532 657 604 663
rect 804 657 988 663
rect 1044 657 1116 663
rect 1668 657 1788 663
rect 2388 657 2412 663
rect 68 637 268 643
rect 276 637 332 643
rect 548 637 748 643
rect 1572 637 1628 643
rect 1636 637 1804 643
rect 1812 637 1868 643
rect 2132 637 2188 643
rect 2196 637 2412 643
rect 2420 637 2540 643
rect 596 617 892 623
rect 948 617 988 623
rect 1716 617 1756 623
rect 1890 614 1950 616
rect 1890 606 1891 614
rect 1900 606 1901 614
rect 1939 606 1940 614
rect 1949 606 1950 614
rect 1890 604 1950 606
rect 228 597 236 603
rect 244 597 300 603
rect 308 597 396 603
rect 404 597 588 603
rect 740 597 812 603
rect 820 597 1020 603
rect 1620 597 1740 603
rect 884 577 1068 583
rect 1076 577 1132 583
rect 1172 577 1356 583
rect 1492 577 1676 583
rect 1684 577 1788 583
rect 1796 577 2380 583
rect -35 557 12 563
rect 116 557 236 563
rect 756 557 780 563
rect 788 557 956 563
rect 964 557 1100 563
rect 1252 557 1324 563
rect 1956 557 2012 563
rect 2020 557 2060 563
rect 356 537 444 543
rect 756 537 828 543
rect 900 537 956 543
rect 980 537 1500 543
rect 1508 537 1596 543
rect 1604 537 1644 543
rect 2228 537 2348 543
rect 164 517 604 523
rect 612 517 636 523
rect 644 517 844 523
rect 1012 517 1068 523
rect -35 497 124 503
rect 292 497 748 503
rect 820 497 876 503
rect 948 497 1004 503
rect 1012 497 1036 503
rect 52 477 76 483
rect 244 477 476 483
rect 484 477 492 483
rect 500 477 1244 483
rect 564 457 1196 463
rect 1700 437 1980 443
rect 1396 417 1420 423
rect 1476 417 1580 423
rect 658 414 718 416
rect 658 406 659 414
rect 668 406 669 414
rect 707 406 708 414
rect 717 406 718 414
rect 658 404 718 406
rect 324 397 444 403
rect 1572 397 1628 403
rect 1748 397 1868 403
rect 1876 397 1900 403
rect 1908 397 2172 403
rect 2180 397 2252 403
rect 2260 397 2284 403
rect 84 377 732 383
rect 772 357 956 363
rect 836 337 908 343
rect 2164 337 2204 343
rect 516 317 588 323
rect 628 317 732 323
rect 740 317 1020 323
rect 1396 317 1996 323
rect 2132 317 2204 323
rect -35 297 12 303
rect 100 297 476 303
rect 484 297 508 303
rect 580 297 604 303
rect 644 297 668 303
rect 932 297 972 303
rect 1076 297 1100 303
rect 1812 297 1852 303
rect 1972 297 2092 303
rect 2100 297 2140 303
rect 2148 297 2492 303
rect 660 277 812 283
rect 1140 277 1276 283
rect 452 257 524 263
rect 1524 237 1820 243
rect 1828 237 1996 243
rect 2004 237 2060 243
rect 2276 237 2396 243
rect 2532 237 2556 243
rect 772 217 876 223
rect 2372 217 2460 223
rect 1890 214 1950 216
rect 1890 206 1891 214
rect 1900 206 1901 214
rect 1939 206 1940 214
rect 1949 206 1950 214
rect 1890 204 1950 206
rect 196 197 236 203
rect 740 197 796 203
rect 868 197 940 203
rect 948 197 1068 203
rect 36 177 620 183
rect 1108 177 1308 183
rect 1380 177 1388 183
rect 372 157 460 163
rect 468 157 492 163
rect 756 157 1132 163
rect 1572 157 1660 163
rect 1732 157 1804 163
rect 2084 157 2444 163
rect 228 137 572 143
rect 612 137 780 143
rect 1540 137 1836 143
rect 2196 137 2300 143
rect 324 117 348 123
rect 420 117 460 123
rect 548 117 588 123
rect 868 117 876 123
rect 1236 117 1276 123
rect 1652 117 1740 123
rect 1908 117 1980 123
rect 2052 117 2108 123
rect 484 97 540 103
rect 596 97 732 103
rect 452 77 572 83
rect 724 37 748 43
rect 468 17 492 23
rect 516 17 540 23
rect 1876 17 1980 23
rect 658 14 718 16
rect 658 6 659 14
rect 668 6 669 14
rect 707 6 708 14
rect 717 6 718 14
rect 658 4 718 6
<< m4contact >>
rect 588 1816 596 1824
rect 1892 1806 1899 1814
rect 1899 1806 1900 1814
rect 1904 1806 1909 1814
rect 1909 1806 1911 1814
rect 1911 1806 1912 1814
rect 1916 1806 1919 1814
rect 1919 1806 1921 1814
rect 1921 1806 1924 1814
rect 1928 1806 1929 1814
rect 1929 1806 1931 1814
rect 1931 1806 1936 1814
rect 1940 1806 1941 1814
rect 1941 1806 1948 1814
rect 2412 1676 2420 1684
rect 588 1616 596 1624
rect 660 1606 667 1614
rect 667 1606 668 1614
rect 672 1606 677 1614
rect 677 1606 679 1614
rect 679 1606 680 1614
rect 684 1606 687 1614
rect 687 1606 689 1614
rect 689 1606 692 1614
rect 696 1606 697 1614
rect 697 1606 699 1614
rect 699 1606 704 1614
rect 708 1606 709 1614
rect 709 1606 716 1614
rect 908 1596 916 1604
rect 1996 1496 2004 1504
rect 908 1476 916 1484
rect 1388 1476 1396 1484
rect 1836 1436 1844 1444
rect 1892 1406 1899 1414
rect 1899 1406 1900 1414
rect 1904 1406 1909 1414
rect 1909 1406 1911 1414
rect 1911 1406 1912 1414
rect 1916 1406 1919 1414
rect 1919 1406 1921 1414
rect 1921 1406 1924 1414
rect 1928 1406 1929 1414
rect 1929 1406 1931 1414
rect 1931 1406 1936 1414
rect 1940 1406 1941 1414
rect 1941 1406 1948 1414
rect 908 1336 916 1344
rect 660 1206 667 1214
rect 667 1206 668 1214
rect 672 1206 677 1214
rect 677 1206 679 1214
rect 679 1206 680 1214
rect 684 1206 687 1214
rect 687 1206 689 1214
rect 689 1206 692 1214
rect 696 1206 697 1214
rect 697 1206 699 1214
rect 699 1206 704 1214
rect 708 1206 709 1214
rect 709 1206 716 1214
rect 1892 1006 1899 1014
rect 1899 1006 1900 1014
rect 1904 1006 1909 1014
rect 1909 1006 1911 1014
rect 1911 1006 1912 1014
rect 1916 1006 1919 1014
rect 1919 1006 1921 1014
rect 1921 1006 1924 1014
rect 1928 1006 1929 1014
rect 1929 1006 1931 1014
rect 1931 1006 1936 1014
rect 1940 1006 1941 1014
rect 1941 1006 1948 1014
rect 1836 936 1844 944
rect 1388 856 1396 864
rect 492 836 500 844
rect 660 806 667 814
rect 667 806 668 814
rect 672 806 677 814
rect 677 806 679 814
rect 679 806 680 814
rect 684 806 687 814
rect 687 806 689 814
rect 689 806 692 814
rect 696 806 697 814
rect 697 806 699 814
rect 699 806 704 814
rect 708 806 709 814
rect 709 806 716 814
rect 1804 636 1812 644
rect 2412 636 2420 644
rect 1892 606 1899 614
rect 1899 606 1900 614
rect 1904 606 1909 614
rect 1909 606 1911 614
rect 1911 606 1912 614
rect 1916 606 1919 614
rect 1919 606 1921 614
rect 1921 606 1924 614
rect 1928 606 1929 614
rect 1929 606 1931 614
rect 1931 606 1936 614
rect 1940 606 1941 614
rect 1941 606 1948 614
rect 876 576 884 584
rect 492 476 500 484
rect 660 406 667 414
rect 667 406 668 414
rect 672 406 677 414
rect 677 406 679 414
rect 679 406 680 414
rect 684 406 687 414
rect 687 406 689 414
rect 689 406 692 414
rect 696 406 697 414
rect 697 406 699 414
rect 699 406 704 414
rect 708 406 709 414
rect 709 406 716 414
rect 1388 316 1396 324
rect 1996 316 2004 324
rect 1804 296 1812 304
rect 1892 206 1899 214
rect 1899 206 1900 214
rect 1904 206 1909 214
rect 1909 206 1911 214
rect 1911 206 1912 214
rect 1916 206 1919 214
rect 1919 206 1921 214
rect 1921 206 1924 214
rect 1928 206 1929 214
rect 1929 206 1931 214
rect 1931 206 1936 214
rect 1940 206 1941 214
rect 1941 206 1948 214
rect 1388 176 1396 184
rect 876 116 884 124
rect 660 6 667 14
rect 667 6 668 14
rect 672 6 677 14
rect 677 6 679 14
rect 679 6 680 14
rect 684 6 687 14
rect 687 6 689 14
rect 689 6 692 14
rect 696 6 697 14
rect 697 6 699 14
rect 699 6 704 14
rect 708 6 709 14
rect 709 6 716 14
<< metal4 >>
rect 586 1824 598 1826
rect 586 1816 588 1824
rect 596 1816 598 1824
rect 586 1624 598 1816
rect 586 1616 588 1624
rect 596 1616 598 1624
rect 586 1614 598 1616
rect 656 1614 720 1816
rect 656 1606 660 1614
rect 668 1606 672 1614
rect 680 1606 684 1614
rect 692 1606 696 1614
rect 704 1606 708 1614
rect 716 1606 720 1614
rect 1888 1814 1952 1816
rect 1888 1806 1892 1814
rect 1900 1806 1904 1814
rect 1912 1806 1916 1814
rect 1924 1806 1928 1814
rect 1936 1806 1940 1814
rect 1948 1806 1952 1814
rect 656 1214 720 1606
rect 906 1604 918 1606
rect 906 1596 908 1604
rect 916 1596 918 1604
rect 906 1484 918 1596
rect 906 1476 908 1484
rect 916 1476 918 1484
rect 906 1344 918 1476
rect 906 1336 908 1344
rect 916 1336 918 1344
rect 906 1334 918 1336
rect 1386 1484 1398 1486
rect 1386 1476 1388 1484
rect 1396 1476 1398 1484
rect 656 1206 660 1214
rect 668 1206 672 1214
rect 680 1206 684 1214
rect 692 1206 696 1214
rect 704 1206 708 1214
rect 716 1206 720 1214
rect 490 844 502 846
rect 490 836 492 844
rect 500 836 502 844
rect 490 484 502 836
rect 490 476 492 484
rect 500 476 502 484
rect 490 474 502 476
rect 656 814 720 1206
rect 1386 864 1398 1476
rect 1834 1444 1846 1446
rect 1834 1436 1836 1444
rect 1844 1436 1846 1444
rect 1834 944 1846 1436
rect 1834 936 1836 944
rect 1844 936 1846 944
rect 1834 934 1846 936
rect 1888 1414 1952 1806
rect 2410 1684 2422 1686
rect 2410 1676 2412 1684
rect 2420 1676 2422 1684
rect 1888 1406 1892 1414
rect 1900 1406 1904 1414
rect 1912 1406 1916 1414
rect 1924 1406 1928 1414
rect 1936 1406 1940 1414
rect 1948 1406 1952 1414
rect 1888 1014 1952 1406
rect 1888 1006 1892 1014
rect 1900 1006 1904 1014
rect 1912 1006 1916 1014
rect 1924 1006 1928 1014
rect 1936 1006 1940 1014
rect 1948 1006 1952 1014
rect 1386 856 1388 864
rect 1396 856 1398 864
rect 1386 854 1398 856
rect 656 806 660 814
rect 668 806 672 814
rect 680 806 684 814
rect 692 806 696 814
rect 704 806 708 814
rect 716 806 720 814
rect 656 414 720 806
rect 1802 644 1814 646
rect 1802 636 1804 644
rect 1812 636 1814 644
rect 656 406 660 414
rect 668 406 672 414
rect 680 406 684 414
rect 692 406 696 414
rect 704 406 708 414
rect 716 406 720 414
rect 656 14 720 406
rect 874 584 886 586
rect 874 576 876 584
rect 884 576 886 584
rect 874 124 886 576
rect 1386 324 1398 326
rect 1386 316 1388 324
rect 1396 316 1398 324
rect 1386 184 1398 316
rect 1802 304 1814 636
rect 1802 296 1804 304
rect 1812 296 1814 304
rect 1802 294 1814 296
rect 1888 614 1952 1006
rect 1888 606 1892 614
rect 1900 606 1904 614
rect 1912 606 1916 614
rect 1924 606 1928 614
rect 1936 606 1940 614
rect 1948 606 1952 614
rect 1386 176 1388 184
rect 1396 176 1398 184
rect 1386 174 1398 176
rect 1888 214 1952 606
rect 1994 1504 2006 1506
rect 1994 1496 1996 1504
rect 2004 1496 2006 1504
rect 1994 324 2006 1496
rect 2410 644 2422 1676
rect 2410 636 2412 644
rect 2420 636 2422 644
rect 2410 634 2422 636
rect 1994 316 1996 324
rect 2004 316 2006 324
rect 1994 314 2006 316
rect 1888 206 1892 214
rect 1900 206 1904 214
rect 1912 206 1916 214
rect 1924 206 1928 214
rect 1936 206 1940 214
rect 1948 206 1952 214
rect 874 116 876 124
rect 884 116 886 124
rect 874 114 886 116
rect 656 6 660 14
rect 668 6 672 14
rect 680 6 684 14
rect 692 6 696 14
rect 704 6 708 14
rect 716 6 720 14
rect 656 -10 720 6
rect 1888 -10 1952 206
use DFFSR  _307_
timestamp 1588175369
transform -1 0 360 0 -1 210
box -4 -6 356 206
use INVX1  _233_
timestamp 1588175369
transform 1 0 360 0 -1 210
box -4 -6 36 206
use BUFX2  _264_
timestamp 1588175369
transform -1 0 56 0 1 210
box -4 -6 52 206
use DFFSR  _305_
timestamp 1588175369
transform -1 0 408 0 1 210
box -4 -6 356 206
use OAI21X1  _238_
timestamp 1588175369
transform 1 0 456 0 1 210
box -4 -6 68 206
use NOR2X1  _235_
timestamp 1588175369
transform 1 0 408 0 1 210
box -4 -6 52 206
use INVX1  _246_
timestamp 1588175369
transform -1 0 488 0 -1 210
box -4 -6 36 206
use NAND3X1  _247_
timestamp 1588175369
transform 1 0 392 0 -1 210
box -4 -6 68 206
use OAI22X1  _244_
timestamp 1588175369
transform 1 0 520 0 1 210
box -4 -6 84 206
use OAI21X1  _245_
timestamp 1588175369
transform 1 0 488 0 -1 210
box -4 -6 68 206
use AND2X2  _243_
timestamp 1588175369
transform -1 0 664 0 1 210
box -4 -6 68 206
use BUFX2  _266_
timestamp 1588175369
transform 1 0 616 0 -1 210
box -4 -6 52 206
use NAND3X1  _248_
timestamp 1588175369
transform -1 0 616 0 -1 210
box -4 -6 68 206
use FILL  SFILL7120x2100
timestamp 1588175369
transform 1 0 712 0 1 210
box -4 -6 20 206
use FILL  SFILL6960x2100
timestamp 1588175369
transform 1 0 696 0 1 210
box -4 -6 20 206
use FILL  SFILL6800x2100
timestamp 1588175369
transform 1 0 680 0 1 210
box -4 -6 20 206
use FILL  SFILL6640x2100
timestamp 1588175369
transform 1 0 664 0 1 210
box -4 -6 20 206
use FILL  SFILL7120x100
timestamp 1588175369
transform -1 0 728 0 -1 210
box -4 -6 20 206
use FILL  SFILL6960x100
timestamp 1588175369
transform -1 0 712 0 -1 210
box -4 -6 20 206
use FILL  SFILL6800x100
timestamp 1588175369
transform -1 0 696 0 -1 210
box -4 -6 20 206
use FILL  SFILL6640x100
timestamp 1588175369
transform -1 0 680 0 -1 210
box -4 -6 20 206
use OAI21X1  _242_
timestamp 1588175369
transform -1 0 792 0 1 210
box -4 -6 68 206
use OAI21X1  _250_
timestamp 1588175369
transform -1 0 792 0 -1 210
box -4 -6 68 206
use AOI22X1  _249_
timestamp 1588175369
transform -1 0 936 0 1 210
box -4 -6 84 206
use NAND3X1  _241_
timestamp 1588175369
transform 1 0 792 0 1 210
box -4 -6 68 206
use BUFX2  _267_
timestamp 1588175369
transform -1 0 920 0 -1 210
box -4 -6 52 206
use BUFX2  _265_
timestamp 1588175369
transform -1 0 872 0 -1 210
box -4 -6 52 206
use INVX1  _239_
timestamp 1588175369
transform 1 0 792 0 -1 210
box -4 -6 36 206
use AND2X2  _258_
timestamp 1588175369
transform 1 0 1080 0 1 210
box -4 -6 68 206
use NOR2X1  _126_
timestamp 1588175369
transform -1 0 1080 0 1 210
box -4 -6 52 206
use NAND2X1  _128_
timestamp 1588175369
transform -1 0 1032 0 1 210
box -4 -6 52 206
use NOR2X1  _129_
timestamp 1588175369
transform -1 0 984 0 1 210
box -4 -6 52 206
use DFFSR  _308_
timestamp 1588175369
transform -1 0 1272 0 -1 210
box -4 -6 356 206
use BUFX2  BUFX2_insert9
timestamp 1588175369
transform -1 0 1320 0 -1 210
box -4 -6 52 206
use INVX8  _259_
timestamp 1588175369
transform 1 0 1320 0 -1 210
box -4 -6 84 206
use DFFSR  _295_
timestamp 1588175369
transform 1 0 1400 0 -1 210
box -4 -6 356 206
use DFFSR  _288_
timestamp 1588175369
transform 1 0 1144 0 1 210
box -4 -6 356 206
use BUFX2  _273_
timestamp 1588175369
transform 1 0 1752 0 -1 210
box -4 -6 52 206
use INVX1  _146_
timestamp 1588175369
transform 1 0 1800 0 -1 210
box -4 -6 36 206
use DFFSR  _309_
timestamp 1588175369
transform 1 0 1496 0 1 210
box -4 -6 356 206
use BUFX2  _282_
timestamp 1588175369
transform 1 0 1848 0 1 210
box -4 -6 52 206
use FILL  SFILL18960x2100
timestamp 1588175369
transform 1 0 1896 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_insert11
timestamp 1588175369
transform -1 0 2008 0 1 210
box -4 -6 52 206
use FILL  SFILL19280x100
timestamp 1588175369
transform -1 0 1944 0 -1 210
box -4 -6 20 206
use FILL  SFILL19440x100
timestamp 1588175369
transform -1 0 1960 0 -1 210
box -4 -6 20 206
use FILL  SFILL19600x100
timestamp 1588175369
transform -1 0 1976 0 -1 210
box -4 -6 20 206
use FILL  SFILL19760x100
timestamp 1588175369
transform -1 0 1992 0 -1 210
box -4 -6 20 206
use FILL  SFILL19120x2100
timestamp 1588175369
transform 1 0 1912 0 1 210
box -4 -6 20 206
use FILL  SFILL19280x2100
timestamp 1588175369
transform 1 0 1928 0 1 210
box -4 -6 20 206
use FILL  SFILL19440x2100
timestamp 1588175369
transform 1 0 1944 0 1 210
box -4 -6 20 206
use MUX2X1  _148_
timestamp 1588175369
transform -1 0 1928 0 -1 210
box -4 -6 100 206
use MUX2X1  _160_
timestamp 1588175369
transform 1 0 2136 0 1 210
box -4 -6 100 206
use INVX1  _158_
timestamp 1588175369
transform 1 0 2104 0 1 210
box -4 -6 36 206
use NOR2X1  _138_
timestamp 1588175369
transform 1 0 2056 0 1 210
box -4 -6 52 206
use BUFX2  _281_
timestamp 1588175369
transform 1 0 2008 0 1 210
box -4 -6 52 206
use BUFX2  _277_
timestamp 1588175369
transform 1 0 2040 0 -1 210
box -4 -6 52 206
use BUFX2  _278_
timestamp 1588175369
transform 1 0 1992 0 -1 210
box -4 -6 52 206
use DFFSR  _299_
timestamp 1588175369
transform -1 0 2440 0 -1 210
box -4 -6 356 206
use AOI21X1  _139_
timestamp 1588175369
transform -1 0 2504 0 -1 210
box -4 -6 68 206
use INVX1  _136_
timestamp 1588175369
transform -1 0 2536 0 -1 210
box -4 -6 36 206
use DFFSR  _292_
timestamp 1588175369
transform 1 0 2232 0 1 210
box -4 -6 356 206
use BUFX2  _270_
timestamp 1588175369
transform 1 0 2536 0 -1 210
box -4 -6 52 206
use FILL  FILL24560x100
timestamp 1588175369
transform -1 0 2600 0 -1 210
box -4 -6 20 206
use FILL  FILL24560x2100
timestamp 1588175369
transform 1 0 2584 0 1 210
box -4 -6 20 206
use NOR2X1  _236_
timestamp 1588175369
transform 1 0 8 0 -1 610
box -4 -6 52 206
use NAND3X1  _237_
timestamp 1588175369
transform -1 0 120 0 -1 610
box -4 -6 68 206
use BUFX2  _262_
timestamp 1588175369
transform -1 0 168 0 -1 610
box -4 -6 52 206
use OAI21X1  _220_
timestamp 1588175369
transform 1 0 168 0 -1 610
box -4 -6 68 206
use OAI22X1  _224_
timestamp 1588175369
transform 1 0 232 0 -1 610
box -4 -6 84 206
use DFFSR  _303_
timestamp 1588175369
transform 1 0 312 0 -1 610
box -4 -6 356 206
use AOI22X1  _223_
timestamp 1588175369
transform -1 0 808 0 -1 610
box -4 -6 84 206
use FILL  SFILL6640x4100
timestamp 1588175369
transform -1 0 680 0 -1 610
box -4 -6 20 206
use FILL  SFILL6800x4100
timestamp 1588175369
transform -1 0 696 0 -1 610
box -4 -6 20 206
use FILL  SFILL6960x4100
timestamp 1588175369
transform -1 0 712 0 -1 610
box -4 -6 20 206
use FILL  SFILL7120x4100
timestamp 1588175369
transform -1 0 728 0 -1 610
box -4 -6 20 206
use NAND2X1  _222_
timestamp 1588175369
transform -1 0 856 0 -1 610
box -4 -6 52 206
use NOR2X1  _123_
timestamp 1588175369
transform -1 0 904 0 -1 610
box -4 -6 52 206
use AND2X2  _240_
timestamp 1588175369
transform -1 0 968 0 -1 610
box -4 -6 68 206
use NAND2X1  _125_
timestamp 1588175369
transform 1 0 968 0 -1 610
box -4 -6 52 206
use NOR2X1  _124_
timestamp 1588175369
transform -1 0 1064 0 -1 610
box -4 -6 52 206
use NOR2X1  _228_
timestamp 1588175369
transform -1 0 1112 0 -1 610
box -4 -6 52 206
use INVX1  _229_
timestamp 1588175369
transform -1 0 1144 0 -1 610
box -4 -6 36 206
use DFFSR  _306_
timestamp 1588175369
transform -1 0 1496 0 -1 610
box -4 -6 356 206
use OAI21X1  _173_
timestamp 1588175369
transform 1 0 1496 0 -1 610
box -4 -6 68 206
use AOI21X1  _174_
timestamp 1588175369
transform -1 0 1624 0 -1 610
box -4 -6 68 206
use DFFSR  _312_
timestamp 1588175369
transform 1 0 1624 0 -1 610
box -4 -6 356 206
use INVX1  _147_
timestamp 1588175369
transform -1 0 2072 0 -1 610
box -4 -6 36 206
use XNOR2X1  _164_
timestamp 1588175369
transform 1 0 2072 0 -1 610
box -4 -6 116 206
use FILL  SFILL19760x4100
timestamp 1588175369
transform -1 0 1992 0 -1 610
box -4 -6 20 206
use FILL  SFILL19920x4100
timestamp 1588175369
transform -1 0 2008 0 -1 610
box -4 -6 20 206
use FILL  SFILL20080x4100
timestamp 1588175369
transform -1 0 2024 0 -1 610
box -4 -6 20 206
use FILL  SFILL20240x4100
timestamp 1588175369
transform -1 0 2040 0 -1 610
box -4 -6 20 206
use INVX1  _159_
timestamp 1588175369
transform 1 0 2184 0 -1 610
box -4 -6 36 206
use DFFSR  _316_
timestamp 1588175369
transform 1 0 2216 0 -1 610
box -4 -6 356 206
use FILL  FILL24400x4100
timestamp 1588175369
transform -1 0 2584 0 -1 610
box -4 -6 20 206
use FILL  FILL24560x4100
timestamp 1588175369
transform -1 0 2600 0 -1 610
box -4 -6 20 206
use OR2X2  _226_
timestamp 1588175369
transform 1 0 8 0 1 610
box -4 -6 68 206
use AOI21X1  _219_
timestamp 1588175369
transform 1 0 72 0 1 610
box -4 -6 68 206
use INVX1  _217_
timestamp 1588175369
transform 1 0 136 0 1 610
box -4 -6 36 206
use OAI21X1  _225_
timestamp 1588175369
transform 1 0 168 0 1 610
box -4 -6 68 206
use OAI21X1  _227_
timestamp 1588175369
transform -1 0 296 0 1 610
box -4 -6 68 206
use NOR2X1  _234_
timestamp 1588175369
transform -1 0 344 0 1 610
box -4 -6 52 206
use OAI21X1  _207_
timestamp 1588175369
transform -1 0 408 0 1 610
box -4 -6 68 206
use XOR2X1  _202_
timestamp 1588175369
transform -1 0 520 0 1 610
box -4 -6 116 206
use OAI21X1  _213_
timestamp 1588175369
transform 1 0 520 0 1 610
box -4 -6 68 206
use OR2X2  _212_
timestamp 1588175369
transform 1 0 584 0 1 610
box -4 -6 68 206
use OAI21X1  _214_
timestamp 1588175369
transform -1 0 776 0 1 610
box -4 -6 68 206
use FILL  SFILL6480x6100
timestamp 1588175369
transform 1 0 648 0 1 610
box -4 -6 20 206
use FILL  SFILL6640x6100
timestamp 1588175369
transform 1 0 664 0 1 610
box -4 -6 20 206
use FILL  SFILL6800x6100
timestamp 1588175369
transform 1 0 680 0 1 610
box -4 -6 20 206
use FILL  SFILL6960x6100
timestamp 1588175369
transform 1 0 696 0 1 610
box -4 -6 20 206
use NOR2X1  _221_
timestamp 1588175369
transform -1 0 824 0 1 610
box -4 -6 52 206
use INVX4  _121_
timestamp 1588175369
transform 1 0 824 0 1 610
box -4 -6 52 206
use AND2X2  _196_
timestamp 1588175369
transform -1 0 936 0 1 610
box -4 -6 68 206
use NAND2X1  _201_
timestamp 1588175369
transform -1 0 984 0 1 610
box -4 -6 52 206
use AOI21X1  _230_
timestamp 1588175369
transform 1 0 984 0 1 610
box -4 -6 68 206
use OAI21X1  _231_
timestamp 1588175369
transform 1 0 1048 0 1 610
box -4 -6 68 206
use OAI21X1  _232_
timestamp 1588175369
transform 1 0 1112 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert6
timestamp 1588175369
transform -1 0 1224 0 1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert0
timestamp 1588175369
transform -1 0 1368 0 1 610
box -4 -6 148 206
use CLKBUF1  CLKBUF1_insert2
timestamp 1588175369
transform 1 0 1368 0 1 610
box -4 -6 148 206
use BUFX2  BUFX2_insert7
timestamp 1588175369
transform 1 0 1512 0 1 610
box -4 -6 52 206
use OAI21X1  _255_
timestamp 1588175369
transform -1 0 1624 0 1 610
box -4 -6 68 206
use NOR2X1  _165_
timestamp 1588175369
transform 1 0 1624 0 1 610
box -4 -6 52 206
use AOI21X1  _178_
timestamp 1588175369
transform 1 0 1672 0 1 610
box -4 -6 68 206
use NAND2X1  _172_
timestamp 1588175369
transform -1 0 1784 0 1 610
box -4 -6 52 206
use OAI21X1  _167_
timestamp 1588175369
transform 1 0 1784 0 1 610
box -4 -6 68 206
use XNOR2X1  _170_
timestamp 1588175369
transform -1 0 2024 0 1 610
box -4 -6 116 206
use OAI21X1  _171_
timestamp 1588175369
transform -1 0 2088 0 1 610
box -4 -6 68 206
use NOR2X1  _168_
timestamp 1588175369
transform -1 0 2136 0 1 610
box -4 -6 52 206
use NOR2X1  _169_
timestamp 1588175369
transform 1 0 2136 0 1 610
box -4 -6 52 206
use FILL  SFILL18480x6100
timestamp 1588175369
transform 1 0 1848 0 1 610
box -4 -6 20 206
use FILL  SFILL18640x6100
timestamp 1588175369
transform 1 0 1864 0 1 610
box -4 -6 20 206
use FILL  SFILL18800x6100
timestamp 1588175369
transform 1 0 1880 0 1 610
box -4 -6 20 206
use FILL  SFILL18960x6100
timestamp 1588175369
transform 1 0 1896 0 1 610
box -4 -6 20 206
use AOI21X1  _186_
timestamp 1588175369
transform 1 0 2184 0 1 610
box -4 -6 68 206
use DFFSR  _314_
timestamp 1588175369
transform 1 0 2248 0 1 610
box -4 -6 356 206
use BUFX2  _263_
timestamp 1588175369
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use INVX1  _203_
timestamp 1588175369
transform -1 0 88 0 -1 1010
box -4 -6 36 206
use NAND3X1  _210_
timestamp 1588175369
transform -1 0 152 0 -1 1010
box -4 -6 68 206
use NAND2X1  _204_
timestamp 1588175369
transform 1 0 152 0 -1 1010
box -4 -6 52 206
use NAND3X1  _206_
timestamp 1588175369
transform -1 0 264 0 -1 1010
box -4 -6 68 206
use NAND2X1  _211_
timestamp 1588175369
transform -1 0 312 0 -1 1010
box -4 -6 52 206
use DFFSR  _302_
timestamp 1588175369
transform 1 0 312 0 -1 1010
box -4 -6 356 206
use NOR2X1  _127_
timestamp 1588175369
transform 1 0 728 0 -1 1010
box -4 -6 52 206
use FILL  SFILL6640x8100
timestamp 1588175369
transform -1 0 680 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6800x8100
timestamp 1588175369
transform -1 0 696 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6960x8100
timestamp 1588175369
transform -1 0 712 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7120x8100
timestamp 1588175369
transform -1 0 728 0 -1 1010
box -4 -6 20 206
use NAND2X1  _215_
timestamp 1588175369
transform -1 0 824 0 -1 1010
box -4 -6 52 206
use OAI21X1  _216_
timestamp 1588175369
transform -1 0 888 0 -1 1010
box -4 -6 68 206
use DFFSR  _304_
timestamp 1588175369
transform -1 0 1240 0 -1 1010
box -4 -6 356 206
use DFFSR  _313_
timestamp 1588175369
transform 1 0 1240 0 -1 1010
box -4 -6 356 206
use NAND3X1  _137_
timestamp 1588175369
transform 1 0 1592 0 -1 1010
box -4 -6 68 206
use AOI21X1  _180_
timestamp 1588175369
transform 1 0 1656 0 -1 1010
box -4 -6 68 206
use OAI21X1  _179_
timestamp 1588175369
transform -1 0 1784 0 -1 1010
box -4 -6 68 206
use NOR2X1  _166_
timestamp 1588175369
transform 1 0 1784 0 -1 1010
box -4 -6 52 206
use INVX1  _150_
timestamp 1588175369
transform -1 0 1864 0 -1 1010
box -4 -6 36 206
use OAI21X1  _181_
timestamp 1588175369
transform 1 0 1864 0 -1 1010
box -4 -6 68 206
use AOI21X1  _182_
timestamp 1588175369
transform 1 0 1992 0 -1 1010
box -4 -6 68 206
use INVX1  _153_
timestamp 1588175369
transform -1 0 2088 0 -1 1010
box -4 -6 36 206
use DFFSR  _315_
timestamp 1588175369
transform 1 0 2088 0 -1 1010
box -4 -6 356 206
use FILL  SFILL19280x8100
timestamp 1588175369
transform -1 0 1944 0 -1 1010
box -4 -6 20 206
use FILL  SFILL19440x8100
timestamp 1588175369
transform -1 0 1960 0 -1 1010
box -4 -6 20 206
use FILL  SFILL19600x8100
timestamp 1588175369
transform -1 0 1976 0 -1 1010
box -4 -6 20 206
use FILL  SFILL19760x8100
timestamp 1588175369
transform -1 0 1992 0 -1 1010
box -4 -6 20 206
use OAI21X1  _185_
timestamp 1588175369
transform -1 0 2504 0 -1 1010
box -4 -6 68 206
use BUFX2  _284_
timestamp 1588175369
transform 1 0 2504 0 -1 1010
box -4 -6 52 206
use BUFX2  _283_
timestamp 1588175369
transform 1 0 2552 0 -1 1010
box -4 -6 52 206
use NAND2X1  _193_
timestamp 1588175369
transform 1 0 8 0 1 1010
box -4 -6 52 206
use NOR2X1  _218_
timestamp 1588175369
transform 1 0 56 0 1 1010
box -4 -6 52 206
use INVX1  _209_
timestamp 1588175369
transform 1 0 104 0 1 1010
box -4 -6 36 206
use INVX1  _194_
timestamp 1588175369
transform 1 0 136 0 1 1010
box -4 -6 36 206
use NAND2X1  _205_
timestamp 1588175369
transform 1 0 168 0 1 1010
box -4 -6 52 206
use OAI21X1  _208_
timestamp 1588175369
transform 1 0 216 0 1 1010
box -4 -6 68 206
use NOR2X1  _192_
timestamp 1588175369
transform -1 0 328 0 1 1010
box -4 -6 52 206
use OAI21X1  _195_
timestamp 1588175369
transform 1 0 328 0 1 1010
box -4 -6 68 206
use NAND2X1  _200_
timestamp 1588175369
transform 1 0 424 0 1 1010
box -4 -6 52 206
use INVX1  _187_
timestamp 1588175369
transform 1 0 392 0 1 1010
box -4 -6 36 206
use OAI21X1  _191_
timestamp 1588175369
transform 1 0 472 0 1 1010
box -4 -6 68 206
use OAI21X1  _199_
timestamp 1588175369
transform -1 0 600 0 1 1010
box -4 -6 68 206
use NOR2X1  _198_
timestamp 1588175369
transform 1 0 632 0 1 1010
box -4 -6 52 206
use INVX1  _197_
timestamp 1588175369
transform 1 0 600 0 1 1010
box -4 -6 36 206
use FILL  SFILL7280x10100
timestamp 1588175369
transform 1 0 728 0 1 1010
box -4 -6 20 206
use FILL  SFILL7120x10100
timestamp 1588175369
transform 1 0 712 0 1 1010
box -4 -6 20 206
use FILL  SFILL6960x10100
timestamp 1588175369
transform 1 0 696 0 1 1010
box -4 -6 20 206
use FILL  SFILL6800x10100
timestamp 1588175369
transform 1 0 680 0 1 1010
box -4 -6 20 206
use OAI21X1  _190_
timestamp 1588175369
transform -1 0 808 0 1 1010
box -4 -6 68 206
use AND2X2  _189_
timestamp 1588175369
transform -1 0 872 0 1 1010
box -4 -6 68 206
use NOR2X1  _188_
timestamp 1588175369
transform 1 0 872 0 1 1010
box -4 -6 52 206
use OAI21X1  _130_
timestamp 1588175369
transform -1 0 984 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert8
timestamp 1588175369
transform -1 0 1032 0 1 1010
box -4 -6 52 206
use NAND3X1  _253_
timestamp 1588175369
transform 1 0 1032 0 1 1010
box -4 -6 68 206
use INVX1  _252_
timestamp 1588175369
transform -1 0 1128 0 1 1010
box -4 -6 36 206
use DFFSR  _290_
timestamp 1588175369
transform -1 0 1480 0 1 1010
box -4 -6 356 206
use BUFX2  BUFX2_insert5
timestamp 1588175369
transform 1 0 1480 0 1 1010
box -4 -6 52 206
use AOI21X1  _256_
timestamp 1588175369
transform 1 0 1528 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert15
timestamp 1588175369
transform -1 0 1640 0 1 1010
box -4 -6 52 206
use INVX8  _122_
timestamp 1588175369
transform 1 0 1640 0 1 1010
box -4 -6 84 206
use OAI21X1  _177_
timestamp 1588175369
transform -1 0 1784 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert14
timestamp 1588175369
transform -1 0 1832 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert16
timestamp 1588175369
transform -1 0 1880 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert17
timestamp 1588175369
transform 1 0 1944 0 1 1010
box -4 -6 52 206
use DFFSR  _310_
timestamp 1588175369
transform -1 0 2344 0 1 1010
box -4 -6 356 206
use FILL  SFILL18800x10100
timestamp 1588175369
transform 1 0 1880 0 1 1010
box -4 -6 20 206
use FILL  SFILL18960x10100
timestamp 1588175369
transform 1 0 1896 0 1 1010
box -4 -6 20 206
use FILL  SFILL19120x10100
timestamp 1588175369
transform 1 0 1912 0 1 1010
box -4 -6 20 206
use FILL  SFILL19280x10100
timestamp 1588175369
transform 1 0 1928 0 1 1010
box -4 -6 20 206
use OAI21X1  _183_
timestamp 1588175369
transform 1 0 2344 0 1 1010
box -4 -6 68 206
use AOI21X1  _184_
timestamp 1588175369
transform -1 0 2472 0 1 1010
box -4 -6 68 206
use INVX1  _156_
timestamp 1588175369
transform -1 0 2504 0 1 1010
box -4 -6 36 206
use MUX2X1  _157_
timestamp 1588175369
transform 1 0 2504 0 1 1010
box -4 -6 100 206
use BUFX2  _261_
timestamp 1588175369
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use INVX1  _251_
timestamp 1588175369
transform 1 0 56 0 -1 1410
box -4 -6 36 206
use AOI21X1  _254_
timestamp 1588175369
transform 1 0 88 0 -1 1410
box -4 -6 68 206
use DFFSR  _301_
timestamp 1588175369
transform 1 0 152 0 -1 1410
box -4 -6 356 206
use DFFSR  _289_
timestamp 1588175369
transform 1 0 568 0 -1 1410
box -4 -6 356 206
use FILL  SFILL5040x12100
timestamp 1588175369
transform -1 0 520 0 -1 1410
box -4 -6 20 206
use FILL  SFILL5200x12100
timestamp 1588175369
transform -1 0 536 0 -1 1410
box -4 -6 20 206
use FILL  SFILL5360x12100
timestamp 1588175369
transform -1 0 552 0 -1 1410
box -4 -6 20 206
use FILL  SFILL5520x12100
timestamp 1588175369
transform -1 0 568 0 -1 1410
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert1
timestamp 1588175369
transform 1 0 920 0 -1 1410
box -4 -6 148 206
use DFFSR  _293_
timestamp 1588175369
transform 1 0 1064 0 -1 1410
box -4 -6 356 206
use BUFX2  BUFX2_insert12
timestamp 1588175369
transform -1 0 1464 0 -1 1410
box -4 -6 52 206
use INVX1  _140_
timestamp 1588175369
transform 1 0 1464 0 -1 1410
box -4 -6 36 206
use MUX2X1  _142_
timestamp 1588175369
transform -1 0 1592 0 -1 1410
box -4 -6 100 206
use INVX1  _141_
timestamp 1588175369
transform -1 0 1624 0 -1 1410
box -4 -6 36 206
use OAI21X1  _175_
timestamp 1588175369
transform 1 0 1624 0 -1 1410
box -4 -6 68 206
use AOI21X1  _176_
timestamp 1588175369
transform -1 0 1752 0 -1 1410
box -4 -6 68 206
use FILL  SFILL17520x12100
timestamp 1588175369
transform -1 0 1768 0 -1 1410
box -4 -6 20 206
use FILL  SFILL17680x12100
timestamp 1588175369
transform -1 0 1784 0 -1 1410
box -4 -6 20 206
use FILL  SFILL17840x12100
timestamp 1588175369
transform -1 0 1800 0 -1 1410
box -4 -6 20 206
use FILL  SFILL18000x12100
timestamp 1588175369
transform -1 0 1816 0 -1 1410
box -4 -6 20 206
use DFFSR  _311_
timestamp 1588175369
transform -1 0 2168 0 -1 1410
box -4 -6 356 206
use DFFSR  _298_
timestamp 1588175369
transform 1 0 2168 0 -1 1410
box -4 -6 356 206
use BUFX2  _276_
timestamp 1588175369
transform 1 0 2520 0 -1 1410
box -4 -6 52 206
use FILL  FILL24400x12100
timestamp 1588175369
transform -1 0 2584 0 -1 1410
box -4 -6 20 206
use FILL  FILL24560x12100
timestamp 1588175369
transform -1 0 2600 0 -1 1410
box -4 -6 20 206
use BUFX2  _268_
timestamp 1588175369
transform -1 0 56 0 1 1410
box -4 -6 52 206
use DFFSR  _286_
timestamp 1588175369
transform -1 0 408 0 1 1410
box -4 -6 356 206
use AND2X2  _257_
timestamp 1588175369
transform -1 0 472 0 1 1410
box -4 -6 68 206
use OAI21X1  _135_
timestamp 1588175369
transform 1 0 504 0 1 1410
box -4 -6 68 206
use INVX1  _132_
timestamp 1588175369
transform 1 0 472 0 1 1410
box -4 -6 36 206
use BUFX2  _260_
timestamp 1588175369
transform -1 0 616 0 1 1410
box -4 -6 52 206
use FILL  SFILL6480x14100
timestamp 1588175369
transform 1 0 648 0 1 1410
box -4 -6 20 206
use INVX1  _131_
timestamp 1588175369
transform -1 0 648 0 1 1410
box -4 -6 36 206
use FILL  SFILL6960x14100
timestamp 1588175369
transform 1 0 696 0 1 1410
box -4 -6 20 206
use FILL  SFILL6800x14100
timestamp 1588175369
transform 1 0 680 0 1 1410
box -4 -6 20 206
use FILL  SFILL6640x14100
timestamp 1588175369
transform 1 0 664 0 1 1410
box -4 -6 20 206
use NOR2X1  _134_
timestamp 1588175369
transform 1 0 712 0 1 1410
box -4 -6 52 206
use INVX1  _133_
timestamp 1588175369
transform -1 0 792 0 1 1410
box -4 -6 36 206
use DFFSR  _318_
timestamp 1588175369
transform -1 0 1144 0 1 1410
box -4 -6 356 206
use BUFX2  BUFX2_insert10
timestamp 1588175369
transform -1 0 1192 0 1 1410
box -4 -6 52 206
use DFFSR  _297_
timestamp 1588175369
transform 1 0 1192 0 1 1410
box -4 -6 356 206
use INVX1  _152_
timestamp 1588175369
transform 1 0 1544 0 1 1410
box -4 -6 36 206
use MUX2X1  _154_
timestamp 1588175369
transform -1 0 1672 0 1 1410
box -4 -6 100 206
use BUFX2  _271_
timestamp 1588175369
transform 1 0 1672 0 1 1410
box -4 -6 52 206
use INVX1  _144_
timestamp 1588175369
transform -1 0 1752 0 1 1410
box -4 -6 36 206
use BUFX2  _280_
timestamp 1588175369
transform 1 0 1752 0 1 1410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert3
timestamp 1588175369
transform 1 0 1800 0 1 1410
box -4 -6 148 206
use BUFX2  BUFX2_insert13
timestamp 1588175369
transform 1 0 2008 0 1 1410
box -4 -6 52 206
use MUX2X1  _151_
timestamp 1588175369
transform 1 0 2056 0 1 1410
box -4 -6 100 206
use MUX2X1  _145_
timestamp 1588175369
transform 1 0 2152 0 1 1410
box -4 -6 100 206
use FILL  SFILL19440x14100
timestamp 1588175369
transform 1 0 1944 0 1 1410
box -4 -6 20 206
use FILL  SFILL19600x14100
timestamp 1588175369
transform 1 0 1960 0 1 1410
box -4 -6 20 206
use FILL  SFILL19760x14100
timestamp 1588175369
transform 1 0 1976 0 1 1410
box -4 -6 20 206
use FILL  SFILL19920x14100
timestamp 1588175369
transform 1 0 1992 0 1 1410
box -4 -6 20 206
use DFFSR  _294_
timestamp 1588175369
transform 1 0 2248 0 1 1410
box -4 -6 356 206
use DFFSR  _300_
timestamp 1588175369
transform -1 0 360 0 -1 1810
box -4 -6 356 206
use DFFSR  _287_
timestamp 1588175369
transform -1 0 712 0 -1 1810
box -4 -6 356 206
use FILL  SFILL7120x16100
timestamp 1588175369
transform -1 0 728 0 -1 1810
box -4 -6 20 206
use FILL  SFILL7280x16100
timestamp 1588175369
transform -1 0 744 0 -1 1810
box -4 -6 20 206
use CLKBUF1  CLKBUF1_insert4
timestamp 1588175369
transform -1 0 920 0 -1 1810
box -4 -6 148 206
use DFFSR  _317_
timestamp 1588175369
transform -1 0 1272 0 -1 1810
box -4 -6 356 206
use FILL  SFILL7440x16100
timestamp 1588175369
transform -1 0 760 0 -1 1810
box -4 -6 20 206
use FILL  SFILL7600x16100
timestamp 1588175369
transform -1 0 776 0 -1 1810
box -4 -6 20 206
use DFFSR  _291_
timestamp 1588175369
transform 1 0 1272 0 -1 1810
box -4 -6 356 206
use BUFX2  _275_
timestamp 1588175369
transform 1 0 1624 0 -1 1810
box -4 -6 52 206
use BUFX2  _269_
timestamp 1588175369
transform 1 0 1672 0 -1 1810
box -4 -6 52 206
use INVX1  _161_
timestamp 1588175369
transform 1 0 1720 0 -1 1810
box -4 -6 36 206
use AOI21X1  _163_
timestamp 1588175369
transform 1 0 1752 0 -1 1810
box -4 -6 68 206
use NOR2X1  _162_
timestamp 1588175369
transform -1 0 1864 0 -1 1810
box -4 -6 52 206
use BUFX2  _279_
timestamp 1588175369
transform 1 0 1864 0 -1 1810
box -4 -6 52 206
use BUFX2  _274_
timestamp 1588175369
transform -1 0 2024 0 -1 1810
box -4 -6 52 206
use INVX1  _149_
timestamp 1588175369
transform 1 0 2024 0 -1 1810
box -4 -6 36 206
use DFFSR  _296_
timestamp 1588175369
transform -1 0 2408 0 -1 1810
box -4 -6 356 206
use FILL  SFILL19120x16100
timestamp 1588175369
transform -1 0 1928 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19280x16100
timestamp 1588175369
transform -1 0 1944 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19440x16100
timestamp 1588175369
transform -1 0 1960 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19600x16100
timestamp 1588175369
transform -1 0 1976 0 -1 1810
box -4 -6 20 206
use BUFX2  _285_
timestamp 1588175369
transform 1 0 2408 0 -1 1810
box -4 -6 52 206
use INVX1  _143_
timestamp 1588175369
transform -1 0 2488 0 -1 1810
box -4 -6 36 206
use INVX1  _155_
timestamp 1588175369
transform -1 0 2520 0 -1 1810
box -4 -6 36 206
use BUFX2  _272_
timestamp 1588175369
transform 1 0 2520 0 -1 1810
box -4 -6 52 206
use FILL  FILL24400x16100
timestamp 1588175369
transform -1 0 2584 0 -1 1810
box -4 -6 20 206
use FILL  FILL24560x16100
timestamp 1588175369
transform -1 0 2600 0 -1 1810
box -4 -6 20 206
<< labels >>
flabel metal4 s 1888 -10 1952 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 656 -10 720 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 509 -23 515 -17 7 FreeSans 24 270 0 0 N[8]
port 2 nsew
flabel metal2 s 461 -23 467 -17 7 FreeSans 24 270 0 0 N[7]
port 3 nsew
flabel metal3 s -35 677 -29 683 7 FreeSans 24 0 0 0 N[6]
port 4 nsew
flabel metal3 s -35 557 -29 563 7 FreeSans 24 0 0 0 N[5]
port 5 nsew
flabel metal3 s -35 1137 -29 1143 7 FreeSans 24 0 0 0 N[4]
port 6 nsew
flabel metal3 s -35 1057 -29 1063 7 FreeSans 24 0 0 0 N[3]
port 7 nsew
flabel metal3 s -35 1177 -29 1183 7 FreeSans 24 0 0 0 N[2]
port 8 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 N[1]
port 9 nsew
flabel metal2 s 1837 1857 1843 1863 3 FreeSans 24 90 0 0 N[0]
port 10 nsew
flabel metal2 s 909 1857 915 1863 3 FreeSans 24 90 0 0 clock
port 11 nsew
flabel metal2 s 893 -23 899 -17 7 FreeSans 24 270 0 0 counter[7]
port 12 nsew
flabel metal2 s 749 -23 755 -17 7 FreeSans 24 270 0 0 counter[6]
port 13 nsew
flabel metal2 s 845 -23 851 -17 7 FreeSans 24 270 0 0 counter[5]
port 14 nsew
flabel metal3 s -35 297 -29 303 7 FreeSans 24 0 0 0 counter[4]
port 15 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 counter[3]
port 16 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 counter[2]
port 17 nsew
flabel metal3 s -35 1297 -29 1303 7 FreeSans 24 0 0 0 counter[1]
port 18 nsew
flabel metal2 s 589 1857 595 1863 3 FreeSans 24 90 0 0 counter[0]
port 19 nsew
flabel metal3 s -35 1497 -29 1503 7 FreeSans 24 0 0 0 done
port 20 nsew
flabel metal2 s 2077 -23 2083 -17 7 FreeSans 24 270 0 0 dp[8]
port 21 nsew
flabel metal3 s 2637 1297 2643 1303 3 FreeSans 24 0 0 0 dp[7]
port 22 nsew
flabel metal2 s 1645 1857 1651 1863 3 FreeSans 24 90 0 0 dp[6]
port 23 nsew
flabel metal2 s 2013 1857 2019 1863 3 FreeSans 24 90 0 0 dp[5]
port 24 nsew
flabel metal2 s 1773 -23 1779 -17 7 FreeSans 24 270 0 0 dp[4]
port 25 nsew
flabel metal3 s 2637 1737 2643 1743 3 FreeSans 24 0 0 0 dp[3]
port 26 nsew
flabel metal2 s 1693 1857 1699 1863 3 FreeSans 24 90 0 0 dp[2]
port 27 nsew
flabel metal2 s 2557 -23 2563 -17 7 FreeSans 24 270 0 0 dp[1]
port 28 nsew
flabel metal2 s 1725 1857 1731 1863 3 FreeSans 24 90 0 0 dp[0]
port 29 nsew
flabel metal2 s 1357 -23 1363 -17 7 FreeSans 24 270 0 0 reset
port 30 nsew
flabel metal3 s 2637 1697 2643 1703 3 FreeSans 24 0 0 0 sr[7]
port 31 nsew
flabel metal3 s 2637 897 2643 903 3 FreeSans 24 0 0 0 sr[6]
port 32 nsew
flabel metal3 s 2637 937 2643 943 3 FreeSans 24 0 0 0 sr[5]
port 33 nsew
flabel metal2 s 1981 -23 1987 -17 7 FreeSans 24 270 0 0 sr[4]
port 34 nsew
flabel metal2 s 2045 -23 2051 -17 7 FreeSans 24 270 0 0 sr[3]
port 35 nsew
flabel metal2 s 1773 1857 1779 1863 3 FreeSans 24 90 0 0 sr[2]
port 36 nsew
flabel metal2 s 1981 1857 1987 1863 3 FreeSans 24 90 0 0 sr[1]
port 37 nsew
flabel metal2 s 2013 -23 2019 -17 7 FreeSans 24 270 0 0 sr[0]
port 38 nsew
flabel metal2 s 1085 1857 1091 1863 3 FreeSans 24 90 0 0 start
port 39 nsew
<< end >>
